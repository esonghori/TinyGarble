
module MUX_N512_0 ( A, B, S, O );
  input [511:0] A;
  input [511:0] B;
  output [511:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024;

  XOR U1 ( .A(A[9]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U4 ( .A(A[99]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U7 ( .A(A[98]), .B(n5), .Z(O[98]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[98]), .B(A[98]), .Z(n6) );
  XOR U10 ( .A(A[97]), .B(n7), .Z(O[97]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[97]), .B(A[97]), .Z(n8) );
  XOR U13 ( .A(A[96]), .B(n9), .Z(O[96]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[96]), .B(A[96]), .Z(n10) );
  XOR U16 ( .A(A[95]), .B(n11), .Z(O[95]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[95]), .B(A[95]), .Z(n12) );
  XOR U19 ( .A(A[94]), .B(n13), .Z(O[94]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[94]), .B(A[94]), .Z(n14) );
  XOR U22 ( .A(A[93]), .B(n15), .Z(O[93]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[93]), .B(A[93]), .Z(n16) );
  XOR U25 ( .A(A[92]), .B(n17), .Z(O[92]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[92]), .B(A[92]), .Z(n18) );
  XOR U28 ( .A(A[91]), .B(n19), .Z(O[91]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[91]), .B(A[91]), .Z(n20) );
  XOR U31 ( .A(A[90]), .B(n21), .Z(O[90]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[90]), .B(A[90]), .Z(n22) );
  XOR U34 ( .A(A[8]), .B(n23), .Z(O[8]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR U37 ( .A(A[89]), .B(n25), .Z(O[89]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[89]), .B(A[89]), .Z(n26) );
  XOR U40 ( .A(A[88]), .B(n27), .Z(O[88]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[88]), .B(A[88]), .Z(n28) );
  XOR U43 ( .A(A[87]), .B(n29), .Z(O[87]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[87]), .B(A[87]), .Z(n30) );
  XOR U46 ( .A(A[86]), .B(n31), .Z(O[86]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[86]), .B(A[86]), .Z(n32) );
  XOR U49 ( .A(A[85]), .B(n33), .Z(O[85]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[85]), .B(A[85]), .Z(n34) );
  XOR U52 ( .A(A[84]), .B(n35), .Z(O[84]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[84]), .B(A[84]), .Z(n36) );
  XOR U55 ( .A(A[83]), .B(n37), .Z(O[83]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[83]), .B(A[83]), .Z(n38) );
  XOR U58 ( .A(A[82]), .B(n39), .Z(O[82]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[82]), .B(A[82]), .Z(n40) );
  XOR U61 ( .A(A[81]), .B(n41), .Z(O[81]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[81]), .B(A[81]), .Z(n42) );
  XOR U64 ( .A(A[80]), .B(n43), .Z(O[80]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[80]), .B(A[80]), .Z(n44) );
  XOR U67 ( .A(A[7]), .B(n45), .Z(O[7]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[7]), .B(A[7]), .Z(n46) );
  XOR U70 ( .A(A[79]), .B(n47), .Z(O[79]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[79]), .B(A[79]), .Z(n48) );
  XOR U73 ( .A(A[78]), .B(n49), .Z(O[78]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[78]), .B(A[78]), .Z(n50) );
  XOR U76 ( .A(A[77]), .B(n51), .Z(O[77]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[77]), .B(A[77]), .Z(n52) );
  XOR U79 ( .A(A[76]), .B(n53), .Z(O[76]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[76]), .B(A[76]), .Z(n54) );
  XOR U82 ( .A(A[75]), .B(n55), .Z(O[75]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[75]), .B(A[75]), .Z(n56) );
  XOR U85 ( .A(A[74]), .B(n57), .Z(O[74]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[74]), .B(A[74]), .Z(n58) );
  XOR U88 ( .A(A[73]), .B(n59), .Z(O[73]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[73]), .B(A[73]), .Z(n60) );
  XOR U91 ( .A(A[72]), .B(n61), .Z(O[72]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[72]), .B(A[72]), .Z(n62) );
  XOR U94 ( .A(A[71]), .B(n63), .Z(O[71]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[71]), .B(A[71]), .Z(n64) );
  XOR U97 ( .A(A[70]), .B(n65), .Z(O[70]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[70]), .B(A[70]), .Z(n66) );
  XOR U100 ( .A(A[6]), .B(n67), .Z(O[6]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[6]), .B(A[6]), .Z(n68) );
  XOR U103 ( .A(A[69]), .B(n69), .Z(O[69]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[69]), .B(A[69]), .Z(n70) );
  XOR U106 ( .A(A[68]), .B(n71), .Z(O[68]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[68]), .B(A[68]), .Z(n72) );
  XOR U109 ( .A(A[67]), .B(n73), .Z(O[67]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[67]), .B(A[67]), .Z(n74) );
  XOR U112 ( .A(A[66]), .B(n75), .Z(O[66]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[66]), .B(A[66]), .Z(n76) );
  XOR U115 ( .A(A[65]), .B(n77), .Z(O[65]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[65]), .B(A[65]), .Z(n78) );
  XOR U118 ( .A(A[64]), .B(n79), .Z(O[64]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[64]), .B(A[64]), .Z(n80) );
  XOR U121 ( .A(A[63]), .B(n81), .Z(O[63]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[63]), .B(A[63]), .Z(n82) );
  XOR U124 ( .A(A[62]), .B(n83), .Z(O[62]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[62]), .B(A[62]), .Z(n84) );
  XOR U127 ( .A(A[61]), .B(n85), .Z(O[61]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[61]), .B(A[61]), .Z(n86) );
  XOR U130 ( .A(A[60]), .B(n87), .Z(O[60]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[60]), .B(A[60]), .Z(n88) );
  XOR U133 ( .A(A[5]), .B(n89), .Z(O[5]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[5]), .B(A[5]), .Z(n90) );
  XOR U136 ( .A(A[59]), .B(n91), .Z(O[59]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[59]), .B(A[59]), .Z(n92) );
  XOR U139 ( .A(A[58]), .B(n93), .Z(O[58]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[58]), .B(A[58]), .Z(n94) );
  XOR U142 ( .A(A[57]), .B(n95), .Z(O[57]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[57]), .B(A[57]), .Z(n96) );
  XOR U145 ( .A(A[56]), .B(n97), .Z(O[56]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[56]), .B(A[56]), .Z(n98) );
  XOR U148 ( .A(A[55]), .B(n99), .Z(O[55]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[55]), .B(A[55]), .Z(n100) );
  XOR U151 ( .A(A[54]), .B(n101), .Z(O[54]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[54]), .B(A[54]), .Z(n102) );
  XOR U154 ( .A(A[53]), .B(n103), .Z(O[53]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[53]), .B(A[53]), .Z(n104) );
  XOR U157 ( .A(A[52]), .B(n105), .Z(O[52]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[52]), .B(A[52]), .Z(n106) );
  XOR U160 ( .A(A[51]), .B(n107), .Z(O[51]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[51]), .B(A[51]), .Z(n108) );
  XOR U163 ( .A(A[511]), .B(n109), .Z(O[511]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[511]), .B(A[511]), .Z(n110) );
  XOR U166 ( .A(A[510]), .B(n111), .Z(O[510]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[510]), .B(A[510]), .Z(n112) );
  XOR U169 ( .A(A[50]), .B(n113), .Z(O[50]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[50]), .B(A[50]), .Z(n114) );
  XOR U172 ( .A(A[509]), .B(n115), .Z(O[509]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[509]), .B(A[509]), .Z(n116) );
  XOR U175 ( .A(A[508]), .B(n117), .Z(O[508]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[508]), .B(A[508]), .Z(n118) );
  XOR U178 ( .A(A[507]), .B(n119), .Z(O[507]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[507]), .B(A[507]), .Z(n120) );
  XOR U181 ( .A(A[506]), .B(n121), .Z(O[506]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[506]), .B(A[506]), .Z(n122) );
  XOR U184 ( .A(A[505]), .B(n123), .Z(O[505]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[505]), .B(A[505]), .Z(n124) );
  XOR U187 ( .A(A[504]), .B(n125), .Z(O[504]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[504]), .B(A[504]), .Z(n126) );
  XOR U190 ( .A(A[503]), .B(n127), .Z(O[503]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[503]), .B(A[503]), .Z(n128) );
  XOR U193 ( .A(A[502]), .B(n129), .Z(O[502]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[502]), .B(A[502]), .Z(n130) );
  XOR U196 ( .A(A[501]), .B(n131), .Z(O[501]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[501]), .B(A[501]), .Z(n132) );
  XOR U199 ( .A(A[500]), .B(n133), .Z(O[500]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[500]), .B(A[500]), .Z(n134) );
  XOR U202 ( .A(A[4]), .B(n135), .Z(O[4]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[4]), .B(A[4]), .Z(n136) );
  XOR U205 ( .A(A[49]), .B(n137), .Z(O[49]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[49]), .B(A[49]), .Z(n138) );
  XOR U208 ( .A(A[499]), .B(n139), .Z(O[499]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[499]), .B(A[499]), .Z(n140) );
  XOR U211 ( .A(A[498]), .B(n141), .Z(O[498]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[498]), .B(A[498]), .Z(n142) );
  XOR U214 ( .A(A[497]), .B(n143), .Z(O[497]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[497]), .B(A[497]), .Z(n144) );
  XOR U217 ( .A(A[496]), .B(n145), .Z(O[496]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[496]), .B(A[496]), .Z(n146) );
  XOR U220 ( .A(A[495]), .B(n147), .Z(O[495]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[495]), .B(A[495]), .Z(n148) );
  XOR U223 ( .A(A[494]), .B(n149), .Z(O[494]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[494]), .B(A[494]), .Z(n150) );
  XOR U226 ( .A(A[493]), .B(n151), .Z(O[493]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[493]), .B(A[493]), .Z(n152) );
  XOR U229 ( .A(A[492]), .B(n153), .Z(O[492]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[492]), .B(A[492]), .Z(n154) );
  XOR U232 ( .A(A[491]), .B(n155), .Z(O[491]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[491]), .B(A[491]), .Z(n156) );
  XOR U235 ( .A(A[490]), .B(n157), .Z(O[490]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[490]), .B(A[490]), .Z(n158) );
  XOR U238 ( .A(A[48]), .B(n159), .Z(O[48]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[48]), .B(A[48]), .Z(n160) );
  XOR U241 ( .A(A[489]), .B(n161), .Z(O[489]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[489]), .B(A[489]), .Z(n162) );
  XOR U244 ( .A(A[488]), .B(n163), .Z(O[488]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[488]), .B(A[488]), .Z(n164) );
  XOR U247 ( .A(A[487]), .B(n165), .Z(O[487]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[487]), .B(A[487]), .Z(n166) );
  XOR U250 ( .A(A[486]), .B(n167), .Z(O[486]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[486]), .B(A[486]), .Z(n168) );
  XOR U253 ( .A(A[485]), .B(n169), .Z(O[485]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[485]), .B(A[485]), .Z(n170) );
  XOR U256 ( .A(A[484]), .B(n171), .Z(O[484]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[484]), .B(A[484]), .Z(n172) );
  XOR U259 ( .A(A[483]), .B(n173), .Z(O[483]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[483]), .B(A[483]), .Z(n174) );
  XOR U262 ( .A(A[482]), .B(n175), .Z(O[482]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[482]), .B(A[482]), .Z(n176) );
  XOR U265 ( .A(A[481]), .B(n177), .Z(O[481]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[481]), .B(A[481]), .Z(n178) );
  XOR U268 ( .A(A[480]), .B(n179), .Z(O[480]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[480]), .B(A[480]), .Z(n180) );
  XOR U271 ( .A(A[47]), .B(n181), .Z(O[47]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[47]), .B(A[47]), .Z(n182) );
  XOR U274 ( .A(A[479]), .B(n183), .Z(O[479]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[479]), .B(A[479]), .Z(n184) );
  XOR U277 ( .A(A[478]), .B(n185), .Z(O[478]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[478]), .B(A[478]), .Z(n186) );
  XOR U280 ( .A(A[477]), .B(n187), .Z(O[477]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[477]), .B(A[477]), .Z(n188) );
  XOR U283 ( .A(A[476]), .B(n189), .Z(O[476]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[476]), .B(A[476]), .Z(n190) );
  XOR U286 ( .A(A[475]), .B(n191), .Z(O[475]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[475]), .B(A[475]), .Z(n192) );
  XOR U289 ( .A(A[474]), .B(n193), .Z(O[474]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[474]), .B(A[474]), .Z(n194) );
  XOR U292 ( .A(A[473]), .B(n195), .Z(O[473]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[473]), .B(A[473]), .Z(n196) );
  XOR U295 ( .A(A[472]), .B(n197), .Z(O[472]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[472]), .B(A[472]), .Z(n198) );
  XOR U298 ( .A(A[471]), .B(n199), .Z(O[471]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[471]), .B(A[471]), .Z(n200) );
  XOR U301 ( .A(A[470]), .B(n201), .Z(O[470]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[470]), .B(A[470]), .Z(n202) );
  XOR U304 ( .A(A[46]), .B(n203), .Z(O[46]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[46]), .B(A[46]), .Z(n204) );
  XOR U307 ( .A(A[469]), .B(n205), .Z(O[469]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[469]), .B(A[469]), .Z(n206) );
  XOR U310 ( .A(A[468]), .B(n207), .Z(O[468]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[468]), .B(A[468]), .Z(n208) );
  XOR U313 ( .A(A[467]), .B(n209), .Z(O[467]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[467]), .B(A[467]), .Z(n210) );
  XOR U316 ( .A(A[466]), .B(n211), .Z(O[466]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[466]), .B(A[466]), .Z(n212) );
  XOR U319 ( .A(A[465]), .B(n213), .Z(O[465]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[465]), .B(A[465]), .Z(n214) );
  XOR U322 ( .A(A[464]), .B(n215), .Z(O[464]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[464]), .B(A[464]), .Z(n216) );
  XOR U325 ( .A(A[463]), .B(n217), .Z(O[463]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[463]), .B(A[463]), .Z(n218) );
  XOR U328 ( .A(A[462]), .B(n219), .Z(O[462]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[462]), .B(A[462]), .Z(n220) );
  XOR U331 ( .A(A[461]), .B(n221), .Z(O[461]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[461]), .B(A[461]), .Z(n222) );
  XOR U334 ( .A(A[460]), .B(n223), .Z(O[460]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[460]), .B(A[460]), .Z(n224) );
  XOR U337 ( .A(A[45]), .B(n225), .Z(O[45]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[45]), .B(A[45]), .Z(n226) );
  XOR U340 ( .A(A[459]), .B(n227), .Z(O[459]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[459]), .B(A[459]), .Z(n228) );
  XOR U343 ( .A(A[458]), .B(n229), .Z(O[458]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[458]), .B(A[458]), .Z(n230) );
  XOR U346 ( .A(A[457]), .B(n231), .Z(O[457]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[457]), .B(A[457]), .Z(n232) );
  XOR U349 ( .A(A[456]), .B(n233), .Z(O[456]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[456]), .B(A[456]), .Z(n234) );
  XOR U352 ( .A(A[455]), .B(n235), .Z(O[455]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[455]), .B(A[455]), .Z(n236) );
  XOR U355 ( .A(A[454]), .B(n237), .Z(O[454]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[454]), .B(A[454]), .Z(n238) );
  XOR U358 ( .A(A[453]), .B(n239), .Z(O[453]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[453]), .B(A[453]), .Z(n240) );
  XOR U361 ( .A(A[452]), .B(n241), .Z(O[452]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[452]), .B(A[452]), .Z(n242) );
  XOR U364 ( .A(A[451]), .B(n243), .Z(O[451]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[451]), .B(A[451]), .Z(n244) );
  XOR U367 ( .A(A[450]), .B(n245), .Z(O[450]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[450]), .B(A[450]), .Z(n246) );
  XOR U370 ( .A(A[44]), .B(n247), .Z(O[44]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[44]), .B(A[44]), .Z(n248) );
  XOR U373 ( .A(A[449]), .B(n249), .Z(O[449]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[449]), .B(A[449]), .Z(n250) );
  XOR U376 ( .A(A[448]), .B(n251), .Z(O[448]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[448]), .B(A[448]), .Z(n252) );
  XOR U379 ( .A(A[447]), .B(n253), .Z(O[447]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[447]), .B(A[447]), .Z(n254) );
  XOR U382 ( .A(A[446]), .B(n255), .Z(O[446]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[446]), .B(A[446]), .Z(n256) );
  XOR U385 ( .A(A[445]), .B(n257), .Z(O[445]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[445]), .B(A[445]), .Z(n258) );
  XOR U388 ( .A(A[444]), .B(n259), .Z(O[444]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[444]), .B(A[444]), .Z(n260) );
  XOR U391 ( .A(A[443]), .B(n261), .Z(O[443]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[443]), .B(A[443]), .Z(n262) );
  XOR U394 ( .A(A[442]), .B(n263), .Z(O[442]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[442]), .B(A[442]), .Z(n264) );
  XOR U397 ( .A(A[441]), .B(n265), .Z(O[441]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[441]), .B(A[441]), .Z(n266) );
  XOR U400 ( .A(A[440]), .B(n267), .Z(O[440]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[440]), .B(A[440]), .Z(n268) );
  XOR U403 ( .A(A[43]), .B(n269), .Z(O[43]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[43]), .B(A[43]), .Z(n270) );
  XOR U406 ( .A(A[439]), .B(n271), .Z(O[439]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[439]), .B(A[439]), .Z(n272) );
  XOR U409 ( .A(A[438]), .B(n273), .Z(O[438]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[438]), .B(A[438]), .Z(n274) );
  XOR U412 ( .A(A[437]), .B(n275), .Z(O[437]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[437]), .B(A[437]), .Z(n276) );
  XOR U415 ( .A(A[436]), .B(n277), .Z(O[436]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[436]), .B(A[436]), .Z(n278) );
  XOR U418 ( .A(A[435]), .B(n279), .Z(O[435]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[435]), .B(A[435]), .Z(n280) );
  XOR U421 ( .A(A[434]), .B(n281), .Z(O[434]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[434]), .B(A[434]), .Z(n282) );
  XOR U424 ( .A(A[433]), .B(n283), .Z(O[433]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[433]), .B(A[433]), .Z(n284) );
  XOR U427 ( .A(A[432]), .B(n285), .Z(O[432]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[432]), .B(A[432]), .Z(n286) );
  XOR U430 ( .A(A[431]), .B(n287), .Z(O[431]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[431]), .B(A[431]), .Z(n288) );
  XOR U433 ( .A(A[430]), .B(n289), .Z(O[430]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[430]), .B(A[430]), .Z(n290) );
  XOR U436 ( .A(A[42]), .B(n291), .Z(O[42]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[42]), .B(A[42]), .Z(n292) );
  XOR U439 ( .A(A[429]), .B(n293), .Z(O[429]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[429]), .B(A[429]), .Z(n294) );
  XOR U442 ( .A(A[428]), .B(n295), .Z(O[428]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[428]), .B(A[428]), .Z(n296) );
  XOR U445 ( .A(A[427]), .B(n297), .Z(O[427]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[427]), .B(A[427]), .Z(n298) );
  XOR U448 ( .A(A[426]), .B(n299), .Z(O[426]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[426]), .B(A[426]), .Z(n300) );
  XOR U451 ( .A(A[425]), .B(n301), .Z(O[425]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[425]), .B(A[425]), .Z(n302) );
  XOR U454 ( .A(A[424]), .B(n303), .Z(O[424]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[424]), .B(A[424]), .Z(n304) );
  XOR U457 ( .A(A[423]), .B(n305), .Z(O[423]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[423]), .B(A[423]), .Z(n306) );
  XOR U460 ( .A(A[422]), .B(n307), .Z(O[422]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[422]), .B(A[422]), .Z(n308) );
  XOR U463 ( .A(A[421]), .B(n309), .Z(O[421]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[421]), .B(A[421]), .Z(n310) );
  XOR U466 ( .A(A[420]), .B(n311), .Z(O[420]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[420]), .B(A[420]), .Z(n312) );
  XOR U469 ( .A(A[41]), .B(n313), .Z(O[41]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[41]), .B(A[41]), .Z(n314) );
  XOR U472 ( .A(A[419]), .B(n315), .Z(O[419]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[419]), .B(A[419]), .Z(n316) );
  XOR U475 ( .A(A[418]), .B(n317), .Z(O[418]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[418]), .B(A[418]), .Z(n318) );
  XOR U478 ( .A(A[417]), .B(n319), .Z(O[417]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[417]), .B(A[417]), .Z(n320) );
  XOR U481 ( .A(A[416]), .B(n321), .Z(O[416]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[416]), .B(A[416]), .Z(n322) );
  XOR U484 ( .A(A[415]), .B(n323), .Z(O[415]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[415]), .B(A[415]), .Z(n324) );
  XOR U487 ( .A(A[414]), .B(n325), .Z(O[414]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[414]), .B(A[414]), .Z(n326) );
  XOR U490 ( .A(A[413]), .B(n327), .Z(O[413]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[413]), .B(A[413]), .Z(n328) );
  XOR U493 ( .A(A[412]), .B(n329), .Z(O[412]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[412]), .B(A[412]), .Z(n330) );
  XOR U496 ( .A(A[411]), .B(n331), .Z(O[411]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[411]), .B(A[411]), .Z(n332) );
  XOR U499 ( .A(A[410]), .B(n333), .Z(O[410]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[410]), .B(A[410]), .Z(n334) );
  XOR U502 ( .A(A[40]), .B(n335), .Z(O[40]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[40]), .B(A[40]), .Z(n336) );
  XOR U505 ( .A(A[409]), .B(n337), .Z(O[409]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[409]), .B(A[409]), .Z(n338) );
  XOR U508 ( .A(A[408]), .B(n339), .Z(O[408]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[408]), .B(A[408]), .Z(n340) );
  XOR U511 ( .A(A[407]), .B(n341), .Z(O[407]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[407]), .B(A[407]), .Z(n342) );
  XOR U514 ( .A(A[406]), .B(n343), .Z(O[406]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[406]), .B(A[406]), .Z(n344) );
  XOR U517 ( .A(A[405]), .B(n345), .Z(O[405]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[405]), .B(A[405]), .Z(n346) );
  XOR U520 ( .A(A[404]), .B(n347), .Z(O[404]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[404]), .B(A[404]), .Z(n348) );
  XOR U523 ( .A(A[403]), .B(n349), .Z(O[403]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[403]), .B(A[403]), .Z(n350) );
  XOR U526 ( .A(A[402]), .B(n351), .Z(O[402]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[402]), .B(A[402]), .Z(n352) );
  XOR U529 ( .A(A[401]), .B(n353), .Z(O[401]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[401]), .B(A[401]), .Z(n354) );
  XOR U532 ( .A(A[400]), .B(n355), .Z(O[400]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[400]), .B(A[400]), .Z(n356) );
  XOR U535 ( .A(A[3]), .B(n357), .Z(O[3]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[3]), .B(A[3]), .Z(n358) );
  XOR U538 ( .A(A[39]), .B(n359), .Z(O[39]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[39]), .B(A[39]), .Z(n360) );
  XOR U541 ( .A(A[399]), .B(n361), .Z(O[399]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[399]), .B(A[399]), .Z(n362) );
  XOR U544 ( .A(A[398]), .B(n363), .Z(O[398]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[398]), .B(A[398]), .Z(n364) );
  XOR U547 ( .A(A[397]), .B(n365), .Z(O[397]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[397]), .B(A[397]), .Z(n366) );
  XOR U550 ( .A(A[396]), .B(n367), .Z(O[396]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[396]), .B(A[396]), .Z(n368) );
  XOR U553 ( .A(A[395]), .B(n369), .Z(O[395]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[395]), .B(A[395]), .Z(n370) );
  XOR U556 ( .A(A[394]), .B(n371), .Z(O[394]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[394]), .B(A[394]), .Z(n372) );
  XOR U559 ( .A(A[393]), .B(n373), .Z(O[393]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[393]), .B(A[393]), .Z(n374) );
  XOR U562 ( .A(A[392]), .B(n375), .Z(O[392]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[392]), .B(A[392]), .Z(n376) );
  XOR U565 ( .A(A[391]), .B(n377), .Z(O[391]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[391]), .B(A[391]), .Z(n378) );
  XOR U568 ( .A(A[390]), .B(n379), .Z(O[390]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[390]), .B(A[390]), .Z(n380) );
  XOR U571 ( .A(A[38]), .B(n381), .Z(O[38]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[38]), .B(A[38]), .Z(n382) );
  XOR U574 ( .A(A[389]), .B(n383), .Z(O[389]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[389]), .B(A[389]), .Z(n384) );
  XOR U577 ( .A(A[388]), .B(n385), .Z(O[388]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[388]), .B(A[388]), .Z(n386) );
  XOR U580 ( .A(A[387]), .B(n387), .Z(O[387]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[387]), .B(A[387]), .Z(n388) );
  XOR U583 ( .A(A[386]), .B(n389), .Z(O[386]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[386]), .B(A[386]), .Z(n390) );
  XOR U586 ( .A(A[385]), .B(n391), .Z(O[385]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[385]), .B(A[385]), .Z(n392) );
  XOR U589 ( .A(A[384]), .B(n393), .Z(O[384]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[384]), .B(A[384]), .Z(n394) );
  XOR U592 ( .A(A[383]), .B(n395), .Z(O[383]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[383]), .B(A[383]), .Z(n396) );
  XOR U595 ( .A(A[382]), .B(n397), .Z(O[382]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[382]), .B(A[382]), .Z(n398) );
  XOR U598 ( .A(A[381]), .B(n399), .Z(O[381]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[381]), .B(A[381]), .Z(n400) );
  XOR U601 ( .A(A[380]), .B(n401), .Z(O[380]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[380]), .B(A[380]), .Z(n402) );
  XOR U604 ( .A(A[37]), .B(n403), .Z(O[37]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[37]), .B(A[37]), .Z(n404) );
  XOR U607 ( .A(A[379]), .B(n405), .Z(O[379]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[379]), .B(A[379]), .Z(n406) );
  XOR U610 ( .A(A[378]), .B(n407), .Z(O[378]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[378]), .B(A[378]), .Z(n408) );
  XOR U613 ( .A(A[377]), .B(n409), .Z(O[377]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[377]), .B(A[377]), .Z(n410) );
  XOR U616 ( .A(A[376]), .B(n411), .Z(O[376]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[376]), .B(A[376]), .Z(n412) );
  XOR U619 ( .A(A[375]), .B(n413), .Z(O[375]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[375]), .B(A[375]), .Z(n414) );
  XOR U622 ( .A(A[374]), .B(n415), .Z(O[374]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[374]), .B(A[374]), .Z(n416) );
  XOR U625 ( .A(A[373]), .B(n417), .Z(O[373]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[373]), .B(A[373]), .Z(n418) );
  XOR U628 ( .A(A[372]), .B(n419), .Z(O[372]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[372]), .B(A[372]), .Z(n420) );
  XOR U631 ( .A(A[371]), .B(n421), .Z(O[371]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[371]), .B(A[371]), .Z(n422) );
  XOR U634 ( .A(A[370]), .B(n423), .Z(O[370]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[370]), .B(A[370]), .Z(n424) );
  XOR U637 ( .A(A[36]), .B(n425), .Z(O[36]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[36]), .B(A[36]), .Z(n426) );
  XOR U640 ( .A(A[369]), .B(n427), .Z(O[369]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[369]), .B(A[369]), .Z(n428) );
  XOR U643 ( .A(A[368]), .B(n429), .Z(O[368]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[368]), .B(A[368]), .Z(n430) );
  XOR U646 ( .A(A[367]), .B(n431), .Z(O[367]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[367]), .B(A[367]), .Z(n432) );
  XOR U649 ( .A(A[366]), .B(n433), .Z(O[366]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[366]), .B(A[366]), .Z(n434) );
  XOR U652 ( .A(A[365]), .B(n435), .Z(O[365]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[365]), .B(A[365]), .Z(n436) );
  XOR U655 ( .A(A[364]), .B(n437), .Z(O[364]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[364]), .B(A[364]), .Z(n438) );
  XOR U658 ( .A(A[363]), .B(n439), .Z(O[363]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[363]), .B(A[363]), .Z(n440) );
  XOR U661 ( .A(A[362]), .B(n441), .Z(O[362]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[362]), .B(A[362]), .Z(n442) );
  XOR U664 ( .A(A[361]), .B(n443), .Z(O[361]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[361]), .B(A[361]), .Z(n444) );
  XOR U667 ( .A(A[360]), .B(n445), .Z(O[360]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[360]), .B(A[360]), .Z(n446) );
  XOR U670 ( .A(A[35]), .B(n447), .Z(O[35]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[35]), .B(A[35]), .Z(n448) );
  XOR U673 ( .A(A[359]), .B(n449), .Z(O[359]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[359]), .B(A[359]), .Z(n450) );
  XOR U676 ( .A(A[358]), .B(n451), .Z(O[358]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[358]), .B(A[358]), .Z(n452) );
  XOR U679 ( .A(A[357]), .B(n453), .Z(O[357]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[357]), .B(A[357]), .Z(n454) );
  XOR U682 ( .A(A[356]), .B(n455), .Z(O[356]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[356]), .B(A[356]), .Z(n456) );
  XOR U685 ( .A(A[355]), .B(n457), .Z(O[355]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[355]), .B(A[355]), .Z(n458) );
  XOR U688 ( .A(A[354]), .B(n459), .Z(O[354]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[354]), .B(A[354]), .Z(n460) );
  XOR U691 ( .A(A[353]), .B(n461), .Z(O[353]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[353]), .B(A[353]), .Z(n462) );
  XOR U694 ( .A(A[352]), .B(n463), .Z(O[352]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[352]), .B(A[352]), .Z(n464) );
  XOR U697 ( .A(A[351]), .B(n465), .Z(O[351]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[351]), .B(A[351]), .Z(n466) );
  XOR U700 ( .A(A[350]), .B(n467), .Z(O[350]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[350]), .B(A[350]), .Z(n468) );
  XOR U703 ( .A(A[34]), .B(n469), .Z(O[34]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[34]), .B(A[34]), .Z(n470) );
  XOR U706 ( .A(A[349]), .B(n471), .Z(O[349]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[349]), .B(A[349]), .Z(n472) );
  XOR U709 ( .A(A[348]), .B(n473), .Z(O[348]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[348]), .B(A[348]), .Z(n474) );
  XOR U712 ( .A(A[347]), .B(n475), .Z(O[347]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[347]), .B(A[347]), .Z(n476) );
  XOR U715 ( .A(A[346]), .B(n477), .Z(O[346]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[346]), .B(A[346]), .Z(n478) );
  XOR U718 ( .A(A[345]), .B(n479), .Z(O[345]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[345]), .B(A[345]), .Z(n480) );
  XOR U721 ( .A(A[344]), .B(n481), .Z(O[344]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[344]), .B(A[344]), .Z(n482) );
  XOR U724 ( .A(A[343]), .B(n483), .Z(O[343]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[343]), .B(A[343]), .Z(n484) );
  XOR U727 ( .A(A[342]), .B(n485), .Z(O[342]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[342]), .B(A[342]), .Z(n486) );
  XOR U730 ( .A(A[341]), .B(n487), .Z(O[341]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[341]), .B(A[341]), .Z(n488) );
  XOR U733 ( .A(A[340]), .B(n489), .Z(O[340]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[340]), .B(A[340]), .Z(n490) );
  XOR U736 ( .A(A[33]), .B(n491), .Z(O[33]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[33]), .B(A[33]), .Z(n492) );
  XOR U739 ( .A(A[339]), .B(n493), .Z(O[339]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[339]), .B(A[339]), .Z(n494) );
  XOR U742 ( .A(A[338]), .B(n495), .Z(O[338]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[338]), .B(A[338]), .Z(n496) );
  XOR U745 ( .A(A[337]), .B(n497), .Z(O[337]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[337]), .B(A[337]), .Z(n498) );
  XOR U748 ( .A(A[336]), .B(n499), .Z(O[336]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[336]), .B(A[336]), .Z(n500) );
  XOR U751 ( .A(A[335]), .B(n501), .Z(O[335]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[335]), .B(A[335]), .Z(n502) );
  XOR U754 ( .A(A[334]), .B(n503), .Z(O[334]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[334]), .B(A[334]), .Z(n504) );
  XOR U757 ( .A(A[333]), .B(n505), .Z(O[333]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[333]), .B(A[333]), .Z(n506) );
  XOR U760 ( .A(A[332]), .B(n507), .Z(O[332]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[332]), .B(A[332]), .Z(n508) );
  XOR U763 ( .A(A[331]), .B(n509), .Z(O[331]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[331]), .B(A[331]), .Z(n510) );
  XOR U766 ( .A(A[330]), .B(n511), .Z(O[330]) );
  AND U767 ( .A(S), .B(n512), .Z(n511) );
  XOR U768 ( .A(B[330]), .B(A[330]), .Z(n512) );
  XOR U769 ( .A(A[32]), .B(n513), .Z(O[32]) );
  AND U770 ( .A(S), .B(n514), .Z(n513) );
  XOR U771 ( .A(B[32]), .B(A[32]), .Z(n514) );
  XOR U772 ( .A(A[329]), .B(n515), .Z(O[329]) );
  AND U773 ( .A(S), .B(n516), .Z(n515) );
  XOR U774 ( .A(B[329]), .B(A[329]), .Z(n516) );
  XOR U775 ( .A(A[328]), .B(n517), .Z(O[328]) );
  AND U776 ( .A(S), .B(n518), .Z(n517) );
  XOR U777 ( .A(B[328]), .B(A[328]), .Z(n518) );
  XOR U778 ( .A(A[327]), .B(n519), .Z(O[327]) );
  AND U779 ( .A(S), .B(n520), .Z(n519) );
  XOR U780 ( .A(B[327]), .B(A[327]), .Z(n520) );
  XOR U781 ( .A(A[326]), .B(n521), .Z(O[326]) );
  AND U782 ( .A(S), .B(n522), .Z(n521) );
  XOR U783 ( .A(B[326]), .B(A[326]), .Z(n522) );
  XOR U784 ( .A(A[325]), .B(n523), .Z(O[325]) );
  AND U785 ( .A(S), .B(n524), .Z(n523) );
  XOR U786 ( .A(B[325]), .B(A[325]), .Z(n524) );
  XOR U787 ( .A(A[324]), .B(n525), .Z(O[324]) );
  AND U788 ( .A(S), .B(n526), .Z(n525) );
  XOR U789 ( .A(B[324]), .B(A[324]), .Z(n526) );
  XOR U790 ( .A(A[323]), .B(n527), .Z(O[323]) );
  AND U791 ( .A(S), .B(n528), .Z(n527) );
  XOR U792 ( .A(B[323]), .B(A[323]), .Z(n528) );
  XOR U793 ( .A(A[322]), .B(n529), .Z(O[322]) );
  AND U794 ( .A(S), .B(n530), .Z(n529) );
  XOR U795 ( .A(B[322]), .B(A[322]), .Z(n530) );
  XOR U796 ( .A(A[321]), .B(n531), .Z(O[321]) );
  AND U797 ( .A(S), .B(n532), .Z(n531) );
  XOR U798 ( .A(B[321]), .B(A[321]), .Z(n532) );
  XOR U799 ( .A(A[320]), .B(n533), .Z(O[320]) );
  AND U800 ( .A(S), .B(n534), .Z(n533) );
  XOR U801 ( .A(B[320]), .B(A[320]), .Z(n534) );
  XOR U802 ( .A(A[31]), .B(n535), .Z(O[31]) );
  AND U803 ( .A(S), .B(n536), .Z(n535) );
  XOR U804 ( .A(B[31]), .B(A[31]), .Z(n536) );
  XOR U805 ( .A(A[319]), .B(n537), .Z(O[319]) );
  AND U806 ( .A(S), .B(n538), .Z(n537) );
  XOR U807 ( .A(B[319]), .B(A[319]), .Z(n538) );
  XOR U808 ( .A(A[318]), .B(n539), .Z(O[318]) );
  AND U809 ( .A(S), .B(n540), .Z(n539) );
  XOR U810 ( .A(B[318]), .B(A[318]), .Z(n540) );
  XOR U811 ( .A(A[317]), .B(n541), .Z(O[317]) );
  AND U812 ( .A(S), .B(n542), .Z(n541) );
  XOR U813 ( .A(B[317]), .B(A[317]), .Z(n542) );
  XOR U814 ( .A(A[316]), .B(n543), .Z(O[316]) );
  AND U815 ( .A(S), .B(n544), .Z(n543) );
  XOR U816 ( .A(B[316]), .B(A[316]), .Z(n544) );
  XOR U817 ( .A(A[315]), .B(n545), .Z(O[315]) );
  AND U818 ( .A(S), .B(n546), .Z(n545) );
  XOR U819 ( .A(B[315]), .B(A[315]), .Z(n546) );
  XOR U820 ( .A(A[314]), .B(n547), .Z(O[314]) );
  AND U821 ( .A(S), .B(n548), .Z(n547) );
  XOR U822 ( .A(B[314]), .B(A[314]), .Z(n548) );
  XOR U823 ( .A(A[313]), .B(n549), .Z(O[313]) );
  AND U824 ( .A(S), .B(n550), .Z(n549) );
  XOR U825 ( .A(B[313]), .B(A[313]), .Z(n550) );
  XOR U826 ( .A(A[312]), .B(n551), .Z(O[312]) );
  AND U827 ( .A(S), .B(n552), .Z(n551) );
  XOR U828 ( .A(B[312]), .B(A[312]), .Z(n552) );
  XOR U829 ( .A(A[311]), .B(n553), .Z(O[311]) );
  AND U830 ( .A(S), .B(n554), .Z(n553) );
  XOR U831 ( .A(B[311]), .B(A[311]), .Z(n554) );
  XOR U832 ( .A(A[310]), .B(n555), .Z(O[310]) );
  AND U833 ( .A(S), .B(n556), .Z(n555) );
  XOR U834 ( .A(B[310]), .B(A[310]), .Z(n556) );
  XOR U835 ( .A(A[30]), .B(n557), .Z(O[30]) );
  AND U836 ( .A(S), .B(n558), .Z(n557) );
  XOR U837 ( .A(B[30]), .B(A[30]), .Z(n558) );
  XOR U838 ( .A(A[309]), .B(n559), .Z(O[309]) );
  AND U839 ( .A(S), .B(n560), .Z(n559) );
  XOR U840 ( .A(B[309]), .B(A[309]), .Z(n560) );
  XOR U841 ( .A(A[308]), .B(n561), .Z(O[308]) );
  AND U842 ( .A(S), .B(n562), .Z(n561) );
  XOR U843 ( .A(B[308]), .B(A[308]), .Z(n562) );
  XOR U844 ( .A(A[307]), .B(n563), .Z(O[307]) );
  AND U845 ( .A(S), .B(n564), .Z(n563) );
  XOR U846 ( .A(B[307]), .B(A[307]), .Z(n564) );
  XOR U847 ( .A(A[306]), .B(n565), .Z(O[306]) );
  AND U848 ( .A(S), .B(n566), .Z(n565) );
  XOR U849 ( .A(B[306]), .B(A[306]), .Z(n566) );
  XOR U850 ( .A(A[305]), .B(n567), .Z(O[305]) );
  AND U851 ( .A(S), .B(n568), .Z(n567) );
  XOR U852 ( .A(B[305]), .B(A[305]), .Z(n568) );
  XOR U853 ( .A(A[304]), .B(n569), .Z(O[304]) );
  AND U854 ( .A(S), .B(n570), .Z(n569) );
  XOR U855 ( .A(B[304]), .B(A[304]), .Z(n570) );
  XOR U856 ( .A(A[303]), .B(n571), .Z(O[303]) );
  AND U857 ( .A(S), .B(n572), .Z(n571) );
  XOR U858 ( .A(B[303]), .B(A[303]), .Z(n572) );
  XOR U859 ( .A(A[302]), .B(n573), .Z(O[302]) );
  AND U860 ( .A(S), .B(n574), .Z(n573) );
  XOR U861 ( .A(B[302]), .B(A[302]), .Z(n574) );
  XOR U862 ( .A(A[301]), .B(n575), .Z(O[301]) );
  AND U863 ( .A(S), .B(n576), .Z(n575) );
  XOR U864 ( .A(B[301]), .B(A[301]), .Z(n576) );
  XOR U865 ( .A(A[300]), .B(n577), .Z(O[300]) );
  AND U866 ( .A(S), .B(n578), .Z(n577) );
  XOR U867 ( .A(B[300]), .B(A[300]), .Z(n578) );
  XOR U868 ( .A(A[2]), .B(n579), .Z(O[2]) );
  AND U869 ( .A(S), .B(n580), .Z(n579) );
  XOR U870 ( .A(B[2]), .B(A[2]), .Z(n580) );
  XOR U871 ( .A(A[29]), .B(n581), .Z(O[29]) );
  AND U872 ( .A(S), .B(n582), .Z(n581) );
  XOR U873 ( .A(B[29]), .B(A[29]), .Z(n582) );
  XOR U874 ( .A(A[299]), .B(n583), .Z(O[299]) );
  AND U875 ( .A(S), .B(n584), .Z(n583) );
  XOR U876 ( .A(B[299]), .B(A[299]), .Z(n584) );
  XOR U877 ( .A(A[298]), .B(n585), .Z(O[298]) );
  AND U878 ( .A(S), .B(n586), .Z(n585) );
  XOR U879 ( .A(B[298]), .B(A[298]), .Z(n586) );
  XOR U880 ( .A(A[297]), .B(n587), .Z(O[297]) );
  AND U881 ( .A(S), .B(n588), .Z(n587) );
  XOR U882 ( .A(B[297]), .B(A[297]), .Z(n588) );
  XOR U883 ( .A(A[296]), .B(n589), .Z(O[296]) );
  AND U884 ( .A(S), .B(n590), .Z(n589) );
  XOR U885 ( .A(B[296]), .B(A[296]), .Z(n590) );
  XOR U886 ( .A(A[295]), .B(n591), .Z(O[295]) );
  AND U887 ( .A(S), .B(n592), .Z(n591) );
  XOR U888 ( .A(B[295]), .B(A[295]), .Z(n592) );
  XOR U889 ( .A(A[294]), .B(n593), .Z(O[294]) );
  AND U890 ( .A(S), .B(n594), .Z(n593) );
  XOR U891 ( .A(B[294]), .B(A[294]), .Z(n594) );
  XOR U892 ( .A(A[293]), .B(n595), .Z(O[293]) );
  AND U893 ( .A(S), .B(n596), .Z(n595) );
  XOR U894 ( .A(B[293]), .B(A[293]), .Z(n596) );
  XOR U895 ( .A(A[292]), .B(n597), .Z(O[292]) );
  AND U896 ( .A(S), .B(n598), .Z(n597) );
  XOR U897 ( .A(B[292]), .B(A[292]), .Z(n598) );
  XOR U898 ( .A(A[291]), .B(n599), .Z(O[291]) );
  AND U899 ( .A(S), .B(n600), .Z(n599) );
  XOR U900 ( .A(B[291]), .B(A[291]), .Z(n600) );
  XOR U901 ( .A(A[290]), .B(n601), .Z(O[290]) );
  AND U902 ( .A(S), .B(n602), .Z(n601) );
  XOR U903 ( .A(B[290]), .B(A[290]), .Z(n602) );
  XOR U904 ( .A(A[28]), .B(n603), .Z(O[28]) );
  AND U905 ( .A(S), .B(n604), .Z(n603) );
  XOR U906 ( .A(B[28]), .B(A[28]), .Z(n604) );
  XOR U907 ( .A(A[289]), .B(n605), .Z(O[289]) );
  AND U908 ( .A(S), .B(n606), .Z(n605) );
  XOR U909 ( .A(B[289]), .B(A[289]), .Z(n606) );
  XOR U910 ( .A(A[288]), .B(n607), .Z(O[288]) );
  AND U911 ( .A(S), .B(n608), .Z(n607) );
  XOR U912 ( .A(B[288]), .B(A[288]), .Z(n608) );
  XOR U913 ( .A(A[287]), .B(n609), .Z(O[287]) );
  AND U914 ( .A(S), .B(n610), .Z(n609) );
  XOR U915 ( .A(B[287]), .B(A[287]), .Z(n610) );
  XOR U916 ( .A(A[286]), .B(n611), .Z(O[286]) );
  AND U917 ( .A(S), .B(n612), .Z(n611) );
  XOR U918 ( .A(B[286]), .B(A[286]), .Z(n612) );
  XOR U919 ( .A(A[285]), .B(n613), .Z(O[285]) );
  AND U920 ( .A(S), .B(n614), .Z(n613) );
  XOR U921 ( .A(B[285]), .B(A[285]), .Z(n614) );
  XOR U922 ( .A(A[284]), .B(n615), .Z(O[284]) );
  AND U923 ( .A(S), .B(n616), .Z(n615) );
  XOR U924 ( .A(B[284]), .B(A[284]), .Z(n616) );
  XOR U925 ( .A(A[283]), .B(n617), .Z(O[283]) );
  AND U926 ( .A(S), .B(n618), .Z(n617) );
  XOR U927 ( .A(B[283]), .B(A[283]), .Z(n618) );
  XOR U928 ( .A(A[282]), .B(n619), .Z(O[282]) );
  AND U929 ( .A(S), .B(n620), .Z(n619) );
  XOR U930 ( .A(B[282]), .B(A[282]), .Z(n620) );
  XOR U931 ( .A(A[281]), .B(n621), .Z(O[281]) );
  AND U932 ( .A(S), .B(n622), .Z(n621) );
  XOR U933 ( .A(B[281]), .B(A[281]), .Z(n622) );
  XOR U934 ( .A(A[280]), .B(n623), .Z(O[280]) );
  AND U935 ( .A(S), .B(n624), .Z(n623) );
  XOR U936 ( .A(B[280]), .B(A[280]), .Z(n624) );
  XOR U937 ( .A(A[27]), .B(n625), .Z(O[27]) );
  AND U938 ( .A(S), .B(n626), .Z(n625) );
  XOR U939 ( .A(B[27]), .B(A[27]), .Z(n626) );
  XOR U940 ( .A(A[279]), .B(n627), .Z(O[279]) );
  AND U941 ( .A(S), .B(n628), .Z(n627) );
  XOR U942 ( .A(B[279]), .B(A[279]), .Z(n628) );
  XOR U943 ( .A(A[278]), .B(n629), .Z(O[278]) );
  AND U944 ( .A(S), .B(n630), .Z(n629) );
  XOR U945 ( .A(B[278]), .B(A[278]), .Z(n630) );
  XOR U946 ( .A(A[277]), .B(n631), .Z(O[277]) );
  AND U947 ( .A(S), .B(n632), .Z(n631) );
  XOR U948 ( .A(B[277]), .B(A[277]), .Z(n632) );
  XOR U949 ( .A(A[276]), .B(n633), .Z(O[276]) );
  AND U950 ( .A(S), .B(n634), .Z(n633) );
  XOR U951 ( .A(B[276]), .B(A[276]), .Z(n634) );
  XOR U952 ( .A(A[275]), .B(n635), .Z(O[275]) );
  AND U953 ( .A(S), .B(n636), .Z(n635) );
  XOR U954 ( .A(B[275]), .B(A[275]), .Z(n636) );
  XOR U955 ( .A(A[274]), .B(n637), .Z(O[274]) );
  AND U956 ( .A(S), .B(n638), .Z(n637) );
  XOR U957 ( .A(B[274]), .B(A[274]), .Z(n638) );
  XOR U958 ( .A(A[273]), .B(n639), .Z(O[273]) );
  AND U959 ( .A(S), .B(n640), .Z(n639) );
  XOR U960 ( .A(B[273]), .B(A[273]), .Z(n640) );
  XOR U961 ( .A(A[272]), .B(n641), .Z(O[272]) );
  AND U962 ( .A(S), .B(n642), .Z(n641) );
  XOR U963 ( .A(B[272]), .B(A[272]), .Z(n642) );
  XOR U964 ( .A(A[271]), .B(n643), .Z(O[271]) );
  AND U965 ( .A(S), .B(n644), .Z(n643) );
  XOR U966 ( .A(B[271]), .B(A[271]), .Z(n644) );
  XOR U967 ( .A(A[270]), .B(n645), .Z(O[270]) );
  AND U968 ( .A(S), .B(n646), .Z(n645) );
  XOR U969 ( .A(B[270]), .B(A[270]), .Z(n646) );
  XOR U970 ( .A(A[26]), .B(n647), .Z(O[26]) );
  AND U971 ( .A(S), .B(n648), .Z(n647) );
  XOR U972 ( .A(B[26]), .B(A[26]), .Z(n648) );
  XOR U973 ( .A(A[269]), .B(n649), .Z(O[269]) );
  AND U974 ( .A(S), .B(n650), .Z(n649) );
  XOR U975 ( .A(B[269]), .B(A[269]), .Z(n650) );
  XOR U976 ( .A(A[268]), .B(n651), .Z(O[268]) );
  AND U977 ( .A(S), .B(n652), .Z(n651) );
  XOR U978 ( .A(B[268]), .B(A[268]), .Z(n652) );
  XOR U979 ( .A(A[267]), .B(n653), .Z(O[267]) );
  AND U980 ( .A(S), .B(n654), .Z(n653) );
  XOR U981 ( .A(B[267]), .B(A[267]), .Z(n654) );
  XOR U982 ( .A(A[266]), .B(n655), .Z(O[266]) );
  AND U983 ( .A(S), .B(n656), .Z(n655) );
  XOR U984 ( .A(B[266]), .B(A[266]), .Z(n656) );
  XOR U985 ( .A(A[265]), .B(n657), .Z(O[265]) );
  AND U986 ( .A(S), .B(n658), .Z(n657) );
  XOR U987 ( .A(B[265]), .B(A[265]), .Z(n658) );
  XOR U988 ( .A(A[264]), .B(n659), .Z(O[264]) );
  AND U989 ( .A(S), .B(n660), .Z(n659) );
  XOR U990 ( .A(B[264]), .B(A[264]), .Z(n660) );
  XOR U991 ( .A(A[263]), .B(n661), .Z(O[263]) );
  AND U992 ( .A(S), .B(n662), .Z(n661) );
  XOR U993 ( .A(B[263]), .B(A[263]), .Z(n662) );
  XOR U994 ( .A(A[262]), .B(n663), .Z(O[262]) );
  AND U995 ( .A(S), .B(n664), .Z(n663) );
  XOR U996 ( .A(B[262]), .B(A[262]), .Z(n664) );
  XOR U997 ( .A(A[261]), .B(n665), .Z(O[261]) );
  AND U998 ( .A(S), .B(n666), .Z(n665) );
  XOR U999 ( .A(B[261]), .B(A[261]), .Z(n666) );
  XOR U1000 ( .A(A[260]), .B(n667), .Z(O[260]) );
  AND U1001 ( .A(S), .B(n668), .Z(n667) );
  XOR U1002 ( .A(B[260]), .B(A[260]), .Z(n668) );
  XOR U1003 ( .A(A[25]), .B(n669), .Z(O[25]) );
  AND U1004 ( .A(S), .B(n670), .Z(n669) );
  XOR U1005 ( .A(B[25]), .B(A[25]), .Z(n670) );
  XOR U1006 ( .A(A[259]), .B(n671), .Z(O[259]) );
  AND U1007 ( .A(S), .B(n672), .Z(n671) );
  XOR U1008 ( .A(B[259]), .B(A[259]), .Z(n672) );
  XOR U1009 ( .A(A[258]), .B(n673), .Z(O[258]) );
  AND U1010 ( .A(S), .B(n674), .Z(n673) );
  XOR U1011 ( .A(B[258]), .B(A[258]), .Z(n674) );
  XOR U1012 ( .A(A[257]), .B(n675), .Z(O[257]) );
  AND U1013 ( .A(S), .B(n676), .Z(n675) );
  XOR U1014 ( .A(B[257]), .B(A[257]), .Z(n676) );
  XOR U1015 ( .A(A[256]), .B(n677), .Z(O[256]) );
  AND U1016 ( .A(S), .B(n678), .Z(n677) );
  XOR U1017 ( .A(B[256]), .B(A[256]), .Z(n678) );
  XOR U1018 ( .A(A[255]), .B(n679), .Z(O[255]) );
  AND U1019 ( .A(S), .B(n680), .Z(n679) );
  XOR U1020 ( .A(B[255]), .B(A[255]), .Z(n680) );
  XOR U1021 ( .A(A[254]), .B(n681), .Z(O[254]) );
  AND U1022 ( .A(S), .B(n682), .Z(n681) );
  XOR U1023 ( .A(B[254]), .B(A[254]), .Z(n682) );
  XOR U1024 ( .A(A[253]), .B(n683), .Z(O[253]) );
  AND U1025 ( .A(S), .B(n684), .Z(n683) );
  XOR U1026 ( .A(B[253]), .B(A[253]), .Z(n684) );
  XOR U1027 ( .A(A[252]), .B(n685), .Z(O[252]) );
  AND U1028 ( .A(S), .B(n686), .Z(n685) );
  XOR U1029 ( .A(B[252]), .B(A[252]), .Z(n686) );
  XOR U1030 ( .A(A[251]), .B(n687), .Z(O[251]) );
  AND U1031 ( .A(S), .B(n688), .Z(n687) );
  XOR U1032 ( .A(B[251]), .B(A[251]), .Z(n688) );
  XOR U1033 ( .A(A[250]), .B(n689), .Z(O[250]) );
  AND U1034 ( .A(S), .B(n690), .Z(n689) );
  XOR U1035 ( .A(B[250]), .B(A[250]), .Z(n690) );
  XOR U1036 ( .A(A[24]), .B(n691), .Z(O[24]) );
  AND U1037 ( .A(S), .B(n692), .Z(n691) );
  XOR U1038 ( .A(B[24]), .B(A[24]), .Z(n692) );
  XOR U1039 ( .A(A[249]), .B(n693), .Z(O[249]) );
  AND U1040 ( .A(S), .B(n694), .Z(n693) );
  XOR U1041 ( .A(B[249]), .B(A[249]), .Z(n694) );
  XOR U1042 ( .A(A[248]), .B(n695), .Z(O[248]) );
  AND U1043 ( .A(S), .B(n696), .Z(n695) );
  XOR U1044 ( .A(B[248]), .B(A[248]), .Z(n696) );
  XOR U1045 ( .A(A[247]), .B(n697), .Z(O[247]) );
  AND U1046 ( .A(S), .B(n698), .Z(n697) );
  XOR U1047 ( .A(B[247]), .B(A[247]), .Z(n698) );
  XOR U1048 ( .A(A[246]), .B(n699), .Z(O[246]) );
  AND U1049 ( .A(S), .B(n700), .Z(n699) );
  XOR U1050 ( .A(B[246]), .B(A[246]), .Z(n700) );
  XOR U1051 ( .A(A[245]), .B(n701), .Z(O[245]) );
  AND U1052 ( .A(S), .B(n702), .Z(n701) );
  XOR U1053 ( .A(B[245]), .B(A[245]), .Z(n702) );
  XOR U1054 ( .A(A[244]), .B(n703), .Z(O[244]) );
  AND U1055 ( .A(S), .B(n704), .Z(n703) );
  XOR U1056 ( .A(B[244]), .B(A[244]), .Z(n704) );
  XOR U1057 ( .A(A[243]), .B(n705), .Z(O[243]) );
  AND U1058 ( .A(S), .B(n706), .Z(n705) );
  XOR U1059 ( .A(B[243]), .B(A[243]), .Z(n706) );
  XOR U1060 ( .A(A[242]), .B(n707), .Z(O[242]) );
  AND U1061 ( .A(S), .B(n708), .Z(n707) );
  XOR U1062 ( .A(B[242]), .B(A[242]), .Z(n708) );
  XOR U1063 ( .A(A[241]), .B(n709), .Z(O[241]) );
  AND U1064 ( .A(S), .B(n710), .Z(n709) );
  XOR U1065 ( .A(B[241]), .B(A[241]), .Z(n710) );
  XOR U1066 ( .A(A[240]), .B(n711), .Z(O[240]) );
  AND U1067 ( .A(S), .B(n712), .Z(n711) );
  XOR U1068 ( .A(B[240]), .B(A[240]), .Z(n712) );
  XOR U1069 ( .A(A[23]), .B(n713), .Z(O[23]) );
  AND U1070 ( .A(S), .B(n714), .Z(n713) );
  XOR U1071 ( .A(B[23]), .B(A[23]), .Z(n714) );
  XOR U1072 ( .A(A[239]), .B(n715), .Z(O[239]) );
  AND U1073 ( .A(S), .B(n716), .Z(n715) );
  XOR U1074 ( .A(B[239]), .B(A[239]), .Z(n716) );
  XOR U1075 ( .A(A[238]), .B(n717), .Z(O[238]) );
  AND U1076 ( .A(S), .B(n718), .Z(n717) );
  XOR U1077 ( .A(B[238]), .B(A[238]), .Z(n718) );
  XOR U1078 ( .A(A[237]), .B(n719), .Z(O[237]) );
  AND U1079 ( .A(S), .B(n720), .Z(n719) );
  XOR U1080 ( .A(B[237]), .B(A[237]), .Z(n720) );
  XOR U1081 ( .A(A[236]), .B(n721), .Z(O[236]) );
  AND U1082 ( .A(S), .B(n722), .Z(n721) );
  XOR U1083 ( .A(B[236]), .B(A[236]), .Z(n722) );
  XOR U1084 ( .A(A[235]), .B(n723), .Z(O[235]) );
  AND U1085 ( .A(S), .B(n724), .Z(n723) );
  XOR U1086 ( .A(B[235]), .B(A[235]), .Z(n724) );
  XOR U1087 ( .A(A[234]), .B(n725), .Z(O[234]) );
  AND U1088 ( .A(S), .B(n726), .Z(n725) );
  XOR U1089 ( .A(B[234]), .B(A[234]), .Z(n726) );
  XOR U1090 ( .A(A[233]), .B(n727), .Z(O[233]) );
  AND U1091 ( .A(S), .B(n728), .Z(n727) );
  XOR U1092 ( .A(B[233]), .B(A[233]), .Z(n728) );
  XOR U1093 ( .A(A[232]), .B(n729), .Z(O[232]) );
  AND U1094 ( .A(S), .B(n730), .Z(n729) );
  XOR U1095 ( .A(B[232]), .B(A[232]), .Z(n730) );
  XOR U1096 ( .A(A[231]), .B(n731), .Z(O[231]) );
  AND U1097 ( .A(S), .B(n732), .Z(n731) );
  XOR U1098 ( .A(B[231]), .B(A[231]), .Z(n732) );
  XOR U1099 ( .A(A[230]), .B(n733), .Z(O[230]) );
  AND U1100 ( .A(S), .B(n734), .Z(n733) );
  XOR U1101 ( .A(B[230]), .B(A[230]), .Z(n734) );
  XOR U1102 ( .A(A[22]), .B(n735), .Z(O[22]) );
  AND U1103 ( .A(S), .B(n736), .Z(n735) );
  XOR U1104 ( .A(B[22]), .B(A[22]), .Z(n736) );
  XOR U1105 ( .A(A[229]), .B(n737), .Z(O[229]) );
  AND U1106 ( .A(S), .B(n738), .Z(n737) );
  XOR U1107 ( .A(B[229]), .B(A[229]), .Z(n738) );
  XOR U1108 ( .A(A[228]), .B(n739), .Z(O[228]) );
  AND U1109 ( .A(S), .B(n740), .Z(n739) );
  XOR U1110 ( .A(B[228]), .B(A[228]), .Z(n740) );
  XOR U1111 ( .A(A[227]), .B(n741), .Z(O[227]) );
  AND U1112 ( .A(S), .B(n742), .Z(n741) );
  XOR U1113 ( .A(B[227]), .B(A[227]), .Z(n742) );
  XOR U1114 ( .A(A[226]), .B(n743), .Z(O[226]) );
  AND U1115 ( .A(S), .B(n744), .Z(n743) );
  XOR U1116 ( .A(B[226]), .B(A[226]), .Z(n744) );
  XOR U1117 ( .A(A[225]), .B(n745), .Z(O[225]) );
  AND U1118 ( .A(S), .B(n746), .Z(n745) );
  XOR U1119 ( .A(B[225]), .B(A[225]), .Z(n746) );
  XOR U1120 ( .A(A[224]), .B(n747), .Z(O[224]) );
  AND U1121 ( .A(S), .B(n748), .Z(n747) );
  XOR U1122 ( .A(B[224]), .B(A[224]), .Z(n748) );
  XOR U1123 ( .A(A[223]), .B(n749), .Z(O[223]) );
  AND U1124 ( .A(S), .B(n750), .Z(n749) );
  XOR U1125 ( .A(B[223]), .B(A[223]), .Z(n750) );
  XOR U1126 ( .A(A[222]), .B(n751), .Z(O[222]) );
  AND U1127 ( .A(S), .B(n752), .Z(n751) );
  XOR U1128 ( .A(B[222]), .B(A[222]), .Z(n752) );
  XOR U1129 ( .A(A[221]), .B(n753), .Z(O[221]) );
  AND U1130 ( .A(S), .B(n754), .Z(n753) );
  XOR U1131 ( .A(B[221]), .B(A[221]), .Z(n754) );
  XOR U1132 ( .A(A[220]), .B(n755), .Z(O[220]) );
  AND U1133 ( .A(S), .B(n756), .Z(n755) );
  XOR U1134 ( .A(B[220]), .B(A[220]), .Z(n756) );
  XOR U1135 ( .A(A[21]), .B(n757), .Z(O[21]) );
  AND U1136 ( .A(S), .B(n758), .Z(n757) );
  XOR U1137 ( .A(B[21]), .B(A[21]), .Z(n758) );
  XOR U1138 ( .A(A[219]), .B(n759), .Z(O[219]) );
  AND U1139 ( .A(S), .B(n760), .Z(n759) );
  XOR U1140 ( .A(B[219]), .B(A[219]), .Z(n760) );
  XOR U1141 ( .A(A[218]), .B(n761), .Z(O[218]) );
  AND U1142 ( .A(S), .B(n762), .Z(n761) );
  XOR U1143 ( .A(B[218]), .B(A[218]), .Z(n762) );
  XOR U1144 ( .A(A[217]), .B(n763), .Z(O[217]) );
  AND U1145 ( .A(S), .B(n764), .Z(n763) );
  XOR U1146 ( .A(B[217]), .B(A[217]), .Z(n764) );
  XOR U1147 ( .A(A[216]), .B(n765), .Z(O[216]) );
  AND U1148 ( .A(S), .B(n766), .Z(n765) );
  XOR U1149 ( .A(B[216]), .B(A[216]), .Z(n766) );
  XOR U1150 ( .A(A[215]), .B(n767), .Z(O[215]) );
  AND U1151 ( .A(S), .B(n768), .Z(n767) );
  XOR U1152 ( .A(B[215]), .B(A[215]), .Z(n768) );
  XOR U1153 ( .A(A[214]), .B(n769), .Z(O[214]) );
  AND U1154 ( .A(S), .B(n770), .Z(n769) );
  XOR U1155 ( .A(B[214]), .B(A[214]), .Z(n770) );
  XOR U1156 ( .A(A[213]), .B(n771), .Z(O[213]) );
  AND U1157 ( .A(S), .B(n772), .Z(n771) );
  XOR U1158 ( .A(B[213]), .B(A[213]), .Z(n772) );
  XOR U1159 ( .A(A[212]), .B(n773), .Z(O[212]) );
  AND U1160 ( .A(S), .B(n774), .Z(n773) );
  XOR U1161 ( .A(B[212]), .B(A[212]), .Z(n774) );
  XOR U1162 ( .A(A[211]), .B(n775), .Z(O[211]) );
  AND U1163 ( .A(S), .B(n776), .Z(n775) );
  XOR U1164 ( .A(B[211]), .B(A[211]), .Z(n776) );
  XOR U1165 ( .A(A[210]), .B(n777), .Z(O[210]) );
  AND U1166 ( .A(S), .B(n778), .Z(n777) );
  XOR U1167 ( .A(B[210]), .B(A[210]), .Z(n778) );
  XOR U1168 ( .A(A[20]), .B(n779), .Z(O[20]) );
  AND U1169 ( .A(S), .B(n780), .Z(n779) );
  XOR U1170 ( .A(B[20]), .B(A[20]), .Z(n780) );
  XOR U1171 ( .A(A[209]), .B(n781), .Z(O[209]) );
  AND U1172 ( .A(S), .B(n782), .Z(n781) );
  XOR U1173 ( .A(B[209]), .B(A[209]), .Z(n782) );
  XOR U1174 ( .A(A[208]), .B(n783), .Z(O[208]) );
  AND U1175 ( .A(S), .B(n784), .Z(n783) );
  XOR U1176 ( .A(B[208]), .B(A[208]), .Z(n784) );
  XOR U1177 ( .A(A[207]), .B(n785), .Z(O[207]) );
  AND U1178 ( .A(S), .B(n786), .Z(n785) );
  XOR U1179 ( .A(B[207]), .B(A[207]), .Z(n786) );
  XOR U1180 ( .A(A[206]), .B(n787), .Z(O[206]) );
  AND U1181 ( .A(S), .B(n788), .Z(n787) );
  XOR U1182 ( .A(B[206]), .B(A[206]), .Z(n788) );
  XOR U1183 ( .A(A[205]), .B(n789), .Z(O[205]) );
  AND U1184 ( .A(S), .B(n790), .Z(n789) );
  XOR U1185 ( .A(B[205]), .B(A[205]), .Z(n790) );
  XOR U1186 ( .A(A[204]), .B(n791), .Z(O[204]) );
  AND U1187 ( .A(S), .B(n792), .Z(n791) );
  XOR U1188 ( .A(B[204]), .B(A[204]), .Z(n792) );
  XOR U1189 ( .A(A[203]), .B(n793), .Z(O[203]) );
  AND U1190 ( .A(S), .B(n794), .Z(n793) );
  XOR U1191 ( .A(B[203]), .B(A[203]), .Z(n794) );
  XOR U1192 ( .A(A[202]), .B(n795), .Z(O[202]) );
  AND U1193 ( .A(S), .B(n796), .Z(n795) );
  XOR U1194 ( .A(B[202]), .B(A[202]), .Z(n796) );
  XOR U1195 ( .A(A[201]), .B(n797), .Z(O[201]) );
  AND U1196 ( .A(S), .B(n798), .Z(n797) );
  XOR U1197 ( .A(B[201]), .B(A[201]), .Z(n798) );
  XOR U1198 ( .A(A[200]), .B(n799), .Z(O[200]) );
  AND U1199 ( .A(S), .B(n800), .Z(n799) );
  XOR U1200 ( .A(B[200]), .B(A[200]), .Z(n800) );
  XOR U1201 ( .A(A[1]), .B(n801), .Z(O[1]) );
  AND U1202 ( .A(S), .B(n802), .Z(n801) );
  XOR U1203 ( .A(B[1]), .B(A[1]), .Z(n802) );
  XOR U1204 ( .A(A[19]), .B(n803), .Z(O[19]) );
  AND U1205 ( .A(S), .B(n804), .Z(n803) );
  XOR U1206 ( .A(B[19]), .B(A[19]), .Z(n804) );
  XOR U1207 ( .A(A[199]), .B(n805), .Z(O[199]) );
  AND U1208 ( .A(S), .B(n806), .Z(n805) );
  XOR U1209 ( .A(B[199]), .B(A[199]), .Z(n806) );
  XOR U1210 ( .A(A[198]), .B(n807), .Z(O[198]) );
  AND U1211 ( .A(S), .B(n808), .Z(n807) );
  XOR U1212 ( .A(B[198]), .B(A[198]), .Z(n808) );
  XOR U1213 ( .A(A[197]), .B(n809), .Z(O[197]) );
  AND U1214 ( .A(S), .B(n810), .Z(n809) );
  XOR U1215 ( .A(B[197]), .B(A[197]), .Z(n810) );
  XOR U1216 ( .A(A[196]), .B(n811), .Z(O[196]) );
  AND U1217 ( .A(S), .B(n812), .Z(n811) );
  XOR U1218 ( .A(B[196]), .B(A[196]), .Z(n812) );
  XOR U1219 ( .A(A[195]), .B(n813), .Z(O[195]) );
  AND U1220 ( .A(S), .B(n814), .Z(n813) );
  XOR U1221 ( .A(B[195]), .B(A[195]), .Z(n814) );
  XOR U1222 ( .A(A[194]), .B(n815), .Z(O[194]) );
  AND U1223 ( .A(S), .B(n816), .Z(n815) );
  XOR U1224 ( .A(B[194]), .B(A[194]), .Z(n816) );
  XOR U1225 ( .A(A[193]), .B(n817), .Z(O[193]) );
  AND U1226 ( .A(S), .B(n818), .Z(n817) );
  XOR U1227 ( .A(B[193]), .B(A[193]), .Z(n818) );
  XOR U1228 ( .A(A[192]), .B(n819), .Z(O[192]) );
  AND U1229 ( .A(S), .B(n820), .Z(n819) );
  XOR U1230 ( .A(B[192]), .B(A[192]), .Z(n820) );
  XOR U1231 ( .A(A[191]), .B(n821), .Z(O[191]) );
  AND U1232 ( .A(S), .B(n822), .Z(n821) );
  XOR U1233 ( .A(B[191]), .B(A[191]), .Z(n822) );
  XOR U1234 ( .A(A[190]), .B(n823), .Z(O[190]) );
  AND U1235 ( .A(S), .B(n824), .Z(n823) );
  XOR U1236 ( .A(B[190]), .B(A[190]), .Z(n824) );
  XOR U1237 ( .A(A[18]), .B(n825), .Z(O[18]) );
  AND U1238 ( .A(S), .B(n826), .Z(n825) );
  XOR U1239 ( .A(B[18]), .B(A[18]), .Z(n826) );
  XOR U1240 ( .A(A[189]), .B(n827), .Z(O[189]) );
  AND U1241 ( .A(S), .B(n828), .Z(n827) );
  XOR U1242 ( .A(B[189]), .B(A[189]), .Z(n828) );
  XOR U1243 ( .A(A[188]), .B(n829), .Z(O[188]) );
  AND U1244 ( .A(S), .B(n830), .Z(n829) );
  XOR U1245 ( .A(B[188]), .B(A[188]), .Z(n830) );
  XOR U1246 ( .A(A[187]), .B(n831), .Z(O[187]) );
  AND U1247 ( .A(S), .B(n832), .Z(n831) );
  XOR U1248 ( .A(B[187]), .B(A[187]), .Z(n832) );
  XOR U1249 ( .A(A[186]), .B(n833), .Z(O[186]) );
  AND U1250 ( .A(S), .B(n834), .Z(n833) );
  XOR U1251 ( .A(B[186]), .B(A[186]), .Z(n834) );
  XOR U1252 ( .A(A[185]), .B(n835), .Z(O[185]) );
  AND U1253 ( .A(S), .B(n836), .Z(n835) );
  XOR U1254 ( .A(B[185]), .B(A[185]), .Z(n836) );
  XOR U1255 ( .A(A[184]), .B(n837), .Z(O[184]) );
  AND U1256 ( .A(S), .B(n838), .Z(n837) );
  XOR U1257 ( .A(B[184]), .B(A[184]), .Z(n838) );
  XOR U1258 ( .A(A[183]), .B(n839), .Z(O[183]) );
  AND U1259 ( .A(S), .B(n840), .Z(n839) );
  XOR U1260 ( .A(B[183]), .B(A[183]), .Z(n840) );
  XOR U1261 ( .A(A[182]), .B(n841), .Z(O[182]) );
  AND U1262 ( .A(S), .B(n842), .Z(n841) );
  XOR U1263 ( .A(B[182]), .B(A[182]), .Z(n842) );
  XOR U1264 ( .A(A[181]), .B(n843), .Z(O[181]) );
  AND U1265 ( .A(S), .B(n844), .Z(n843) );
  XOR U1266 ( .A(B[181]), .B(A[181]), .Z(n844) );
  XOR U1267 ( .A(A[180]), .B(n845), .Z(O[180]) );
  AND U1268 ( .A(S), .B(n846), .Z(n845) );
  XOR U1269 ( .A(B[180]), .B(A[180]), .Z(n846) );
  XOR U1270 ( .A(A[17]), .B(n847), .Z(O[17]) );
  AND U1271 ( .A(S), .B(n848), .Z(n847) );
  XOR U1272 ( .A(B[17]), .B(A[17]), .Z(n848) );
  XOR U1273 ( .A(A[179]), .B(n849), .Z(O[179]) );
  AND U1274 ( .A(S), .B(n850), .Z(n849) );
  XOR U1275 ( .A(B[179]), .B(A[179]), .Z(n850) );
  XOR U1276 ( .A(A[178]), .B(n851), .Z(O[178]) );
  AND U1277 ( .A(S), .B(n852), .Z(n851) );
  XOR U1278 ( .A(B[178]), .B(A[178]), .Z(n852) );
  XOR U1279 ( .A(A[177]), .B(n853), .Z(O[177]) );
  AND U1280 ( .A(S), .B(n854), .Z(n853) );
  XOR U1281 ( .A(B[177]), .B(A[177]), .Z(n854) );
  XOR U1282 ( .A(A[176]), .B(n855), .Z(O[176]) );
  AND U1283 ( .A(S), .B(n856), .Z(n855) );
  XOR U1284 ( .A(B[176]), .B(A[176]), .Z(n856) );
  XOR U1285 ( .A(A[175]), .B(n857), .Z(O[175]) );
  AND U1286 ( .A(S), .B(n858), .Z(n857) );
  XOR U1287 ( .A(B[175]), .B(A[175]), .Z(n858) );
  XOR U1288 ( .A(A[174]), .B(n859), .Z(O[174]) );
  AND U1289 ( .A(S), .B(n860), .Z(n859) );
  XOR U1290 ( .A(B[174]), .B(A[174]), .Z(n860) );
  XOR U1291 ( .A(A[173]), .B(n861), .Z(O[173]) );
  AND U1292 ( .A(S), .B(n862), .Z(n861) );
  XOR U1293 ( .A(B[173]), .B(A[173]), .Z(n862) );
  XOR U1294 ( .A(A[172]), .B(n863), .Z(O[172]) );
  AND U1295 ( .A(S), .B(n864), .Z(n863) );
  XOR U1296 ( .A(B[172]), .B(A[172]), .Z(n864) );
  XOR U1297 ( .A(A[171]), .B(n865), .Z(O[171]) );
  AND U1298 ( .A(S), .B(n866), .Z(n865) );
  XOR U1299 ( .A(B[171]), .B(A[171]), .Z(n866) );
  XOR U1300 ( .A(A[170]), .B(n867), .Z(O[170]) );
  AND U1301 ( .A(S), .B(n868), .Z(n867) );
  XOR U1302 ( .A(B[170]), .B(A[170]), .Z(n868) );
  XOR U1303 ( .A(A[16]), .B(n869), .Z(O[16]) );
  AND U1304 ( .A(S), .B(n870), .Z(n869) );
  XOR U1305 ( .A(B[16]), .B(A[16]), .Z(n870) );
  XOR U1306 ( .A(A[169]), .B(n871), .Z(O[169]) );
  AND U1307 ( .A(S), .B(n872), .Z(n871) );
  XOR U1308 ( .A(B[169]), .B(A[169]), .Z(n872) );
  XOR U1309 ( .A(A[168]), .B(n873), .Z(O[168]) );
  AND U1310 ( .A(S), .B(n874), .Z(n873) );
  XOR U1311 ( .A(B[168]), .B(A[168]), .Z(n874) );
  XOR U1312 ( .A(A[167]), .B(n875), .Z(O[167]) );
  AND U1313 ( .A(S), .B(n876), .Z(n875) );
  XOR U1314 ( .A(B[167]), .B(A[167]), .Z(n876) );
  XOR U1315 ( .A(A[166]), .B(n877), .Z(O[166]) );
  AND U1316 ( .A(S), .B(n878), .Z(n877) );
  XOR U1317 ( .A(B[166]), .B(A[166]), .Z(n878) );
  XOR U1318 ( .A(A[165]), .B(n879), .Z(O[165]) );
  AND U1319 ( .A(S), .B(n880), .Z(n879) );
  XOR U1320 ( .A(B[165]), .B(A[165]), .Z(n880) );
  XOR U1321 ( .A(A[164]), .B(n881), .Z(O[164]) );
  AND U1322 ( .A(S), .B(n882), .Z(n881) );
  XOR U1323 ( .A(B[164]), .B(A[164]), .Z(n882) );
  XOR U1324 ( .A(A[163]), .B(n883), .Z(O[163]) );
  AND U1325 ( .A(S), .B(n884), .Z(n883) );
  XOR U1326 ( .A(B[163]), .B(A[163]), .Z(n884) );
  XOR U1327 ( .A(A[162]), .B(n885), .Z(O[162]) );
  AND U1328 ( .A(S), .B(n886), .Z(n885) );
  XOR U1329 ( .A(B[162]), .B(A[162]), .Z(n886) );
  XOR U1330 ( .A(A[161]), .B(n887), .Z(O[161]) );
  AND U1331 ( .A(S), .B(n888), .Z(n887) );
  XOR U1332 ( .A(B[161]), .B(A[161]), .Z(n888) );
  XOR U1333 ( .A(A[160]), .B(n889), .Z(O[160]) );
  AND U1334 ( .A(S), .B(n890), .Z(n889) );
  XOR U1335 ( .A(B[160]), .B(A[160]), .Z(n890) );
  XOR U1336 ( .A(A[15]), .B(n891), .Z(O[15]) );
  AND U1337 ( .A(S), .B(n892), .Z(n891) );
  XOR U1338 ( .A(B[15]), .B(A[15]), .Z(n892) );
  XOR U1339 ( .A(A[159]), .B(n893), .Z(O[159]) );
  AND U1340 ( .A(S), .B(n894), .Z(n893) );
  XOR U1341 ( .A(B[159]), .B(A[159]), .Z(n894) );
  XOR U1342 ( .A(A[158]), .B(n895), .Z(O[158]) );
  AND U1343 ( .A(S), .B(n896), .Z(n895) );
  XOR U1344 ( .A(B[158]), .B(A[158]), .Z(n896) );
  XOR U1345 ( .A(A[157]), .B(n897), .Z(O[157]) );
  AND U1346 ( .A(S), .B(n898), .Z(n897) );
  XOR U1347 ( .A(B[157]), .B(A[157]), .Z(n898) );
  XOR U1348 ( .A(A[156]), .B(n899), .Z(O[156]) );
  AND U1349 ( .A(S), .B(n900), .Z(n899) );
  XOR U1350 ( .A(B[156]), .B(A[156]), .Z(n900) );
  XOR U1351 ( .A(A[155]), .B(n901), .Z(O[155]) );
  AND U1352 ( .A(S), .B(n902), .Z(n901) );
  XOR U1353 ( .A(B[155]), .B(A[155]), .Z(n902) );
  XOR U1354 ( .A(A[154]), .B(n903), .Z(O[154]) );
  AND U1355 ( .A(S), .B(n904), .Z(n903) );
  XOR U1356 ( .A(B[154]), .B(A[154]), .Z(n904) );
  XOR U1357 ( .A(A[153]), .B(n905), .Z(O[153]) );
  AND U1358 ( .A(S), .B(n906), .Z(n905) );
  XOR U1359 ( .A(B[153]), .B(A[153]), .Z(n906) );
  XOR U1360 ( .A(A[152]), .B(n907), .Z(O[152]) );
  AND U1361 ( .A(S), .B(n908), .Z(n907) );
  XOR U1362 ( .A(B[152]), .B(A[152]), .Z(n908) );
  XOR U1363 ( .A(A[151]), .B(n909), .Z(O[151]) );
  AND U1364 ( .A(S), .B(n910), .Z(n909) );
  XOR U1365 ( .A(B[151]), .B(A[151]), .Z(n910) );
  XOR U1366 ( .A(A[150]), .B(n911), .Z(O[150]) );
  AND U1367 ( .A(S), .B(n912), .Z(n911) );
  XOR U1368 ( .A(B[150]), .B(A[150]), .Z(n912) );
  XOR U1369 ( .A(A[14]), .B(n913), .Z(O[14]) );
  AND U1370 ( .A(S), .B(n914), .Z(n913) );
  XOR U1371 ( .A(B[14]), .B(A[14]), .Z(n914) );
  XOR U1372 ( .A(A[149]), .B(n915), .Z(O[149]) );
  AND U1373 ( .A(S), .B(n916), .Z(n915) );
  XOR U1374 ( .A(B[149]), .B(A[149]), .Z(n916) );
  XOR U1375 ( .A(A[148]), .B(n917), .Z(O[148]) );
  AND U1376 ( .A(S), .B(n918), .Z(n917) );
  XOR U1377 ( .A(B[148]), .B(A[148]), .Z(n918) );
  XOR U1378 ( .A(A[147]), .B(n919), .Z(O[147]) );
  AND U1379 ( .A(S), .B(n920), .Z(n919) );
  XOR U1380 ( .A(B[147]), .B(A[147]), .Z(n920) );
  XOR U1381 ( .A(A[146]), .B(n921), .Z(O[146]) );
  AND U1382 ( .A(S), .B(n922), .Z(n921) );
  XOR U1383 ( .A(B[146]), .B(A[146]), .Z(n922) );
  XOR U1384 ( .A(A[145]), .B(n923), .Z(O[145]) );
  AND U1385 ( .A(S), .B(n924), .Z(n923) );
  XOR U1386 ( .A(B[145]), .B(A[145]), .Z(n924) );
  XOR U1387 ( .A(A[144]), .B(n925), .Z(O[144]) );
  AND U1388 ( .A(S), .B(n926), .Z(n925) );
  XOR U1389 ( .A(B[144]), .B(A[144]), .Z(n926) );
  XOR U1390 ( .A(A[143]), .B(n927), .Z(O[143]) );
  AND U1391 ( .A(S), .B(n928), .Z(n927) );
  XOR U1392 ( .A(B[143]), .B(A[143]), .Z(n928) );
  XOR U1393 ( .A(A[142]), .B(n929), .Z(O[142]) );
  AND U1394 ( .A(S), .B(n930), .Z(n929) );
  XOR U1395 ( .A(B[142]), .B(A[142]), .Z(n930) );
  XOR U1396 ( .A(A[141]), .B(n931), .Z(O[141]) );
  AND U1397 ( .A(S), .B(n932), .Z(n931) );
  XOR U1398 ( .A(B[141]), .B(A[141]), .Z(n932) );
  XOR U1399 ( .A(A[140]), .B(n933), .Z(O[140]) );
  AND U1400 ( .A(S), .B(n934), .Z(n933) );
  XOR U1401 ( .A(B[140]), .B(A[140]), .Z(n934) );
  XOR U1402 ( .A(A[13]), .B(n935), .Z(O[13]) );
  AND U1403 ( .A(S), .B(n936), .Z(n935) );
  XOR U1404 ( .A(B[13]), .B(A[13]), .Z(n936) );
  XOR U1405 ( .A(A[139]), .B(n937), .Z(O[139]) );
  AND U1406 ( .A(S), .B(n938), .Z(n937) );
  XOR U1407 ( .A(B[139]), .B(A[139]), .Z(n938) );
  XOR U1408 ( .A(A[138]), .B(n939), .Z(O[138]) );
  AND U1409 ( .A(S), .B(n940), .Z(n939) );
  XOR U1410 ( .A(B[138]), .B(A[138]), .Z(n940) );
  XOR U1411 ( .A(A[137]), .B(n941), .Z(O[137]) );
  AND U1412 ( .A(S), .B(n942), .Z(n941) );
  XOR U1413 ( .A(B[137]), .B(A[137]), .Z(n942) );
  XOR U1414 ( .A(A[136]), .B(n943), .Z(O[136]) );
  AND U1415 ( .A(S), .B(n944), .Z(n943) );
  XOR U1416 ( .A(B[136]), .B(A[136]), .Z(n944) );
  XOR U1417 ( .A(A[135]), .B(n945), .Z(O[135]) );
  AND U1418 ( .A(S), .B(n946), .Z(n945) );
  XOR U1419 ( .A(B[135]), .B(A[135]), .Z(n946) );
  XOR U1420 ( .A(A[134]), .B(n947), .Z(O[134]) );
  AND U1421 ( .A(S), .B(n948), .Z(n947) );
  XOR U1422 ( .A(B[134]), .B(A[134]), .Z(n948) );
  XOR U1423 ( .A(A[133]), .B(n949), .Z(O[133]) );
  AND U1424 ( .A(S), .B(n950), .Z(n949) );
  XOR U1425 ( .A(B[133]), .B(A[133]), .Z(n950) );
  XOR U1426 ( .A(A[132]), .B(n951), .Z(O[132]) );
  AND U1427 ( .A(S), .B(n952), .Z(n951) );
  XOR U1428 ( .A(B[132]), .B(A[132]), .Z(n952) );
  XOR U1429 ( .A(A[131]), .B(n953), .Z(O[131]) );
  AND U1430 ( .A(S), .B(n954), .Z(n953) );
  XOR U1431 ( .A(B[131]), .B(A[131]), .Z(n954) );
  XOR U1432 ( .A(A[130]), .B(n955), .Z(O[130]) );
  AND U1433 ( .A(S), .B(n956), .Z(n955) );
  XOR U1434 ( .A(B[130]), .B(A[130]), .Z(n956) );
  XOR U1435 ( .A(A[12]), .B(n957), .Z(O[12]) );
  AND U1436 ( .A(S), .B(n958), .Z(n957) );
  XOR U1437 ( .A(B[12]), .B(A[12]), .Z(n958) );
  XOR U1438 ( .A(A[129]), .B(n959), .Z(O[129]) );
  AND U1439 ( .A(S), .B(n960), .Z(n959) );
  XOR U1440 ( .A(B[129]), .B(A[129]), .Z(n960) );
  XOR U1441 ( .A(A[128]), .B(n961), .Z(O[128]) );
  AND U1442 ( .A(S), .B(n962), .Z(n961) );
  XOR U1443 ( .A(B[128]), .B(A[128]), .Z(n962) );
  XOR U1444 ( .A(A[127]), .B(n963), .Z(O[127]) );
  AND U1445 ( .A(S), .B(n964), .Z(n963) );
  XOR U1446 ( .A(B[127]), .B(A[127]), .Z(n964) );
  XOR U1447 ( .A(A[126]), .B(n965), .Z(O[126]) );
  AND U1448 ( .A(S), .B(n966), .Z(n965) );
  XOR U1449 ( .A(B[126]), .B(A[126]), .Z(n966) );
  XOR U1450 ( .A(A[125]), .B(n967), .Z(O[125]) );
  AND U1451 ( .A(S), .B(n968), .Z(n967) );
  XOR U1452 ( .A(B[125]), .B(A[125]), .Z(n968) );
  XOR U1453 ( .A(A[124]), .B(n969), .Z(O[124]) );
  AND U1454 ( .A(S), .B(n970), .Z(n969) );
  XOR U1455 ( .A(B[124]), .B(A[124]), .Z(n970) );
  XOR U1456 ( .A(A[123]), .B(n971), .Z(O[123]) );
  AND U1457 ( .A(S), .B(n972), .Z(n971) );
  XOR U1458 ( .A(B[123]), .B(A[123]), .Z(n972) );
  XOR U1459 ( .A(A[122]), .B(n973), .Z(O[122]) );
  AND U1460 ( .A(S), .B(n974), .Z(n973) );
  XOR U1461 ( .A(B[122]), .B(A[122]), .Z(n974) );
  XOR U1462 ( .A(A[121]), .B(n975), .Z(O[121]) );
  AND U1463 ( .A(S), .B(n976), .Z(n975) );
  XOR U1464 ( .A(B[121]), .B(A[121]), .Z(n976) );
  XOR U1465 ( .A(A[120]), .B(n977), .Z(O[120]) );
  AND U1466 ( .A(S), .B(n978), .Z(n977) );
  XOR U1467 ( .A(B[120]), .B(A[120]), .Z(n978) );
  XOR U1468 ( .A(A[11]), .B(n979), .Z(O[11]) );
  AND U1469 ( .A(S), .B(n980), .Z(n979) );
  XOR U1470 ( .A(B[11]), .B(A[11]), .Z(n980) );
  XOR U1471 ( .A(A[119]), .B(n981), .Z(O[119]) );
  AND U1472 ( .A(S), .B(n982), .Z(n981) );
  XOR U1473 ( .A(B[119]), .B(A[119]), .Z(n982) );
  XOR U1474 ( .A(A[118]), .B(n983), .Z(O[118]) );
  AND U1475 ( .A(S), .B(n984), .Z(n983) );
  XOR U1476 ( .A(B[118]), .B(A[118]), .Z(n984) );
  XOR U1477 ( .A(A[117]), .B(n985), .Z(O[117]) );
  AND U1478 ( .A(S), .B(n986), .Z(n985) );
  XOR U1479 ( .A(B[117]), .B(A[117]), .Z(n986) );
  XOR U1480 ( .A(A[116]), .B(n987), .Z(O[116]) );
  AND U1481 ( .A(S), .B(n988), .Z(n987) );
  XOR U1482 ( .A(B[116]), .B(A[116]), .Z(n988) );
  XOR U1483 ( .A(A[115]), .B(n989), .Z(O[115]) );
  AND U1484 ( .A(S), .B(n990), .Z(n989) );
  XOR U1485 ( .A(B[115]), .B(A[115]), .Z(n990) );
  XOR U1486 ( .A(A[114]), .B(n991), .Z(O[114]) );
  AND U1487 ( .A(S), .B(n992), .Z(n991) );
  XOR U1488 ( .A(B[114]), .B(A[114]), .Z(n992) );
  XOR U1489 ( .A(A[113]), .B(n993), .Z(O[113]) );
  AND U1490 ( .A(S), .B(n994), .Z(n993) );
  XOR U1491 ( .A(B[113]), .B(A[113]), .Z(n994) );
  XOR U1492 ( .A(A[112]), .B(n995), .Z(O[112]) );
  AND U1493 ( .A(S), .B(n996), .Z(n995) );
  XOR U1494 ( .A(B[112]), .B(A[112]), .Z(n996) );
  XOR U1495 ( .A(A[111]), .B(n997), .Z(O[111]) );
  AND U1496 ( .A(S), .B(n998), .Z(n997) );
  XOR U1497 ( .A(B[111]), .B(A[111]), .Z(n998) );
  XOR U1498 ( .A(A[110]), .B(n999), .Z(O[110]) );
  AND U1499 ( .A(S), .B(n1000), .Z(n999) );
  XOR U1500 ( .A(B[110]), .B(A[110]), .Z(n1000) );
  XOR U1501 ( .A(A[10]), .B(n1001), .Z(O[10]) );
  AND U1502 ( .A(S), .B(n1002), .Z(n1001) );
  XOR U1503 ( .A(B[10]), .B(A[10]), .Z(n1002) );
  XOR U1504 ( .A(A[109]), .B(n1003), .Z(O[109]) );
  AND U1505 ( .A(S), .B(n1004), .Z(n1003) );
  XOR U1506 ( .A(B[109]), .B(A[109]), .Z(n1004) );
  XOR U1507 ( .A(A[108]), .B(n1005), .Z(O[108]) );
  AND U1508 ( .A(S), .B(n1006), .Z(n1005) );
  XOR U1509 ( .A(B[108]), .B(A[108]), .Z(n1006) );
  XOR U1510 ( .A(A[107]), .B(n1007), .Z(O[107]) );
  AND U1511 ( .A(S), .B(n1008), .Z(n1007) );
  XOR U1512 ( .A(B[107]), .B(A[107]), .Z(n1008) );
  XOR U1513 ( .A(A[106]), .B(n1009), .Z(O[106]) );
  AND U1514 ( .A(S), .B(n1010), .Z(n1009) );
  XOR U1515 ( .A(B[106]), .B(A[106]), .Z(n1010) );
  XOR U1516 ( .A(A[105]), .B(n1011), .Z(O[105]) );
  AND U1517 ( .A(S), .B(n1012), .Z(n1011) );
  XOR U1518 ( .A(B[105]), .B(A[105]), .Z(n1012) );
  XOR U1519 ( .A(A[104]), .B(n1013), .Z(O[104]) );
  AND U1520 ( .A(S), .B(n1014), .Z(n1013) );
  XOR U1521 ( .A(B[104]), .B(A[104]), .Z(n1014) );
  XOR U1522 ( .A(A[103]), .B(n1015), .Z(O[103]) );
  AND U1523 ( .A(S), .B(n1016), .Z(n1015) );
  XOR U1524 ( .A(B[103]), .B(A[103]), .Z(n1016) );
  XOR U1525 ( .A(A[102]), .B(n1017), .Z(O[102]) );
  AND U1526 ( .A(S), .B(n1018), .Z(n1017) );
  XOR U1527 ( .A(B[102]), .B(A[102]), .Z(n1018) );
  XOR U1528 ( .A(A[101]), .B(n1019), .Z(O[101]) );
  AND U1529 ( .A(S), .B(n1020), .Z(n1019) );
  XOR U1530 ( .A(B[101]), .B(A[101]), .Z(n1020) );
  XOR U1531 ( .A(A[100]), .B(n1021), .Z(O[100]) );
  AND U1532 ( .A(S), .B(n1022), .Z(n1021) );
  XOR U1533 ( .A(B[100]), .B(A[100]), .Z(n1022) );
  XOR U1534 ( .A(A[0]), .B(n1023), .Z(O[0]) );
  AND U1535 ( .A(S), .B(n1024), .Z(n1023) );
  XOR U1536 ( .A(B[0]), .B(A[0]), .Z(n1024) );
endmodule


module MUX_N514_0 ( A, B, S, O );
  input [513:0] A;
  input [513:0] B;
  output [513:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[511]), .A(S), .Z(O[511]) );
  ANDN U56 ( .B(A[510]), .A(S), .Z(O[510]) );
  ANDN U57 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U58 ( .B(A[509]), .A(S), .Z(O[509]) );
  ANDN U59 ( .B(A[508]), .A(S), .Z(O[508]) );
  ANDN U60 ( .B(A[507]), .A(S), .Z(O[507]) );
  ANDN U61 ( .B(A[506]), .A(S), .Z(O[506]) );
  ANDN U62 ( .B(A[505]), .A(S), .Z(O[505]) );
  ANDN U63 ( .B(A[504]), .A(S), .Z(O[504]) );
  ANDN U64 ( .B(A[503]), .A(S), .Z(O[503]) );
  ANDN U65 ( .B(A[502]), .A(S), .Z(O[502]) );
  ANDN U66 ( .B(A[501]), .A(S), .Z(O[501]) );
  ANDN U67 ( .B(A[500]), .A(S), .Z(O[500]) );
  ANDN U68 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U69 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U70 ( .B(A[499]), .A(S), .Z(O[499]) );
  ANDN U71 ( .B(A[498]), .A(S), .Z(O[498]) );
  ANDN U72 ( .B(A[497]), .A(S), .Z(O[497]) );
  ANDN U73 ( .B(A[496]), .A(S), .Z(O[496]) );
  ANDN U74 ( .B(A[495]), .A(S), .Z(O[495]) );
  ANDN U75 ( .B(A[494]), .A(S), .Z(O[494]) );
  ANDN U76 ( .B(A[493]), .A(S), .Z(O[493]) );
  ANDN U77 ( .B(A[492]), .A(S), .Z(O[492]) );
  ANDN U78 ( .B(A[491]), .A(S), .Z(O[491]) );
  ANDN U79 ( .B(A[490]), .A(S), .Z(O[490]) );
  ANDN U80 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U81 ( .B(A[489]), .A(S), .Z(O[489]) );
  ANDN U82 ( .B(A[488]), .A(S), .Z(O[488]) );
  ANDN U83 ( .B(A[487]), .A(S), .Z(O[487]) );
  ANDN U84 ( .B(A[486]), .A(S), .Z(O[486]) );
  ANDN U85 ( .B(A[485]), .A(S), .Z(O[485]) );
  ANDN U86 ( .B(A[484]), .A(S), .Z(O[484]) );
  ANDN U87 ( .B(A[483]), .A(S), .Z(O[483]) );
  ANDN U88 ( .B(A[482]), .A(S), .Z(O[482]) );
  ANDN U89 ( .B(A[481]), .A(S), .Z(O[481]) );
  ANDN U90 ( .B(A[480]), .A(S), .Z(O[480]) );
  ANDN U91 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U92 ( .B(A[479]), .A(S), .Z(O[479]) );
  ANDN U93 ( .B(A[478]), .A(S), .Z(O[478]) );
  ANDN U94 ( .B(A[477]), .A(S), .Z(O[477]) );
  ANDN U95 ( .B(A[476]), .A(S), .Z(O[476]) );
  ANDN U96 ( .B(A[475]), .A(S), .Z(O[475]) );
  ANDN U97 ( .B(A[474]), .A(S), .Z(O[474]) );
  ANDN U98 ( .B(A[473]), .A(S), .Z(O[473]) );
  ANDN U99 ( .B(A[472]), .A(S), .Z(O[472]) );
  ANDN U100 ( .B(A[471]), .A(S), .Z(O[471]) );
  ANDN U101 ( .B(A[470]), .A(S), .Z(O[470]) );
  ANDN U102 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U103 ( .B(A[469]), .A(S), .Z(O[469]) );
  ANDN U104 ( .B(A[468]), .A(S), .Z(O[468]) );
  ANDN U105 ( .B(A[467]), .A(S), .Z(O[467]) );
  ANDN U106 ( .B(A[466]), .A(S), .Z(O[466]) );
  ANDN U107 ( .B(A[465]), .A(S), .Z(O[465]) );
  ANDN U108 ( .B(A[464]), .A(S), .Z(O[464]) );
  ANDN U109 ( .B(A[463]), .A(S), .Z(O[463]) );
  ANDN U110 ( .B(A[462]), .A(S), .Z(O[462]) );
  ANDN U111 ( .B(A[461]), .A(S), .Z(O[461]) );
  ANDN U112 ( .B(A[460]), .A(S), .Z(O[460]) );
  ANDN U113 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U114 ( .B(A[459]), .A(S), .Z(O[459]) );
  ANDN U115 ( .B(A[458]), .A(S), .Z(O[458]) );
  ANDN U116 ( .B(A[457]), .A(S), .Z(O[457]) );
  ANDN U117 ( .B(A[456]), .A(S), .Z(O[456]) );
  ANDN U118 ( .B(A[455]), .A(S), .Z(O[455]) );
  ANDN U119 ( .B(A[454]), .A(S), .Z(O[454]) );
  ANDN U120 ( .B(A[453]), .A(S), .Z(O[453]) );
  ANDN U121 ( .B(A[452]), .A(S), .Z(O[452]) );
  ANDN U122 ( .B(A[451]), .A(S), .Z(O[451]) );
  ANDN U123 ( .B(A[450]), .A(S), .Z(O[450]) );
  ANDN U124 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U125 ( .B(A[449]), .A(S), .Z(O[449]) );
  ANDN U126 ( .B(A[448]), .A(S), .Z(O[448]) );
  ANDN U127 ( .B(A[447]), .A(S), .Z(O[447]) );
  ANDN U128 ( .B(A[446]), .A(S), .Z(O[446]) );
  ANDN U129 ( .B(A[445]), .A(S), .Z(O[445]) );
  ANDN U130 ( .B(A[444]), .A(S), .Z(O[444]) );
  ANDN U131 ( .B(A[443]), .A(S), .Z(O[443]) );
  ANDN U132 ( .B(A[442]), .A(S), .Z(O[442]) );
  ANDN U133 ( .B(A[441]), .A(S), .Z(O[441]) );
  ANDN U134 ( .B(A[440]), .A(S), .Z(O[440]) );
  ANDN U135 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U136 ( .B(A[439]), .A(S), .Z(O[439]) );
  ANDN U137 ( .B(A[438]), .A(S), .Z(O[438]) );
  ANDN U138 ( .B(A[437]), .A(S), .Z(O[437]) );
  ANDN U139 ( .B(A[436]), .A(S), .Z(O[436]) );
  ANDN U140 ( .B(A[435]), .A(S), .Z(O[435]) );
  ANDN U141 ( .B(A[434]), .A(S), .Z(O[434]) );
  ANDN U142 ( .B(A[433]), .A(S), .Z(O[433]) );
  ANDN U143 ( .B(A[432]), .A(S), .Z(O[432]) );
  ANDN U144 ( .B(A[431]), .A(S), .Z(O[431]) );
  ANDN U145 ( .B(A[430]), .A(S), .Z(O[430]) );
  ANDN U146 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U147 ( .B(A[429]), .A(S), .Z(O[429]) );
  ANDN U148 ( .B(A[428]), .A(S), .Z(O[428]) );
  ANDN U149 ( .B(A[427]), .A(S), .Z(O[427]) );
  ANDN U150 ( .B(A[426]), .A(S), .Z(O[426]) );
  ANDN U151 ( .B(A[425]), .A(S), .Z(O[425]) );
  ANDN U152 ( .B(A[424]), .A(S), .Z(O[424]) );
  ANDN U153 ( .B(A[423]), .A(S), .Z(O[423]) );
  ANDN U154 ( .B(A[422]), .A(S), .Z(O[422]) );
  ANDN U155 ( .B(A[421]), .A(S), .Z(O[421]) );
  ANDN U156 ( .B(A[420]), .A(S), .Z(O[420]) );
  ANDN U157 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U158 ( .B(A[419]), .A(S), .Z(O[419]) );
  ANDN U159 ( .B(A[418]), .A(S), .Z(O[418]) );
  ANDN U160 ( .B(A[417]), .A(S), .Z(O[417]) );
  ANDN U161 ( .B(A[416]), .A(S), .Z(O[416]) );
  ANDN U162 ( .B(A[415]), .A(S), .Z(O[415]) );
  ANDN U163 ( .B(A[414]), .A(S), .Z(O[414]) );
  ANDN U164 ( .B(A[413]), .A(S), .Z(O[413]) );
  ANDN U165 ( .B(A[412]), .A(S), .Z(O[412]) );
  ANDN U166 ( .B(A[411]), .A(S), .Z(O[411]) );
  ANDN U167 ( .B(A[410]), .A(S), .Z(O[410]) );
  ANDN U168 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U169 ( .B(A[409]), .A(S), .Z(O[409]) );
  ANDN U170 ( .B(A[408]), .A(S), .Z(O[408]) );
  ANDN U171 ( .B(A[407]), .A(S), .Z(O[407]) );
  ANDN U172 ( .B(A[406]), .A(S), .Z(O[406]) );
  ANDN U173 ( .B(A[405]), .A(S), .Z(O[405]) );
  ANDN U174 ( .B(A[404]), .A(S), .Z(O[404]) );
  ANDN U175 ( .B(A[403]), .A(S), .Z(O[403]) );
  ANDN U176 ( .B(A[402]), .A(S), .Z(O[402]) );
  ANDN U177 ( .B(A[401]), .A(S), .Z(O[401]) );
  ANDN U178 ( .B(A[400]), .A(S), .Z(O[400]) );
  ANDN U179 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U180 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U181 ( .B(A[399]), .A(S), .Z(O[399]) );
  ANDN U182 ( .B(A[398]), .A(S), .Z(O[398]) );
  ANDN U183 ( .B(A[397]), .A(S), .Z(O[397]) );
  ANDN U184 ( .B(A[396]), .A(S), .Z(O[396]) );
  ANDN U185 ( .B(A[395]), .A(S), .Z(O[395]) );
  ANDN U186 ( .B(A[394]), .A(S), .Z(O[394]) );
  ANDN U187 ( .B(A[393]), .A(S), .Z(O[393]) );
  ANDN U188 ( .B(A[392]), .A(S), .Z(O[392]) );
  ANDN U189 ( .B(A[391]), .A(S), .Z(O[391]) );
  ANDN U190 ( .B(A[390]), .A(S), .Z(O[390]) );
  ANDN U191 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U192 ( .B(A[389]), .A(S), .Z(O[389]) );
  ANDN U193 ( .B(A[388]), .A(S), .Z(O[388]) );
  ANDN U194 ( .B(A[387]), .A(S), .Z(O[387]) );
  ANDN U195 ( .B(A[386]), .A(S), .Z(O[386]) );
  ANDN U196 ( .B(A[385]), .A(S), .Z(O[385]) );
  ANDN U197 ( .B(A[384]), .A(S), .Z(O[384]) );
  ANDN U198 ( .B(A[383]), .A(S), .Z(O[383]) );
  ANDN U199 ( .B(A[382]), .A(S), .Z(O[382]) );
  ANDN U200 ( .B(A[381]), .A(S), .Z(O[381]) );
  ANDN U201 ( .B(A[380]), .A(S), .Z(O[380]) );
  ANDN U202 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U203 ( .B(A[379]), .A(S), .Z(O[379]) );
  ANDN U204 ( .B(A[378]), .A(S), .Z(O[378]) );
  ANDN U205 ( .B(A[377]), .A(S), .Z(O[377]) );
  ANDN U206 ( .B(A[376]), .A(S), .Z(O[376]) );
  ANDN U207 ( .B(A[375]), .A(S), .Z(O[375]) );
  ANDN U208 ( .B(A[374]), .A(S), .Z(O[374]) );
  ANDN U209 ( .B(A[373]), .A(S), .Z(O[373]) );
  ANDN U210 ( .B(A[372]), .A(S), .Z(O[372]) );
  ANDN U211 ( .B(A[371]), .A(S), .Z(O[371]) );
  ANDN U212 ( .B(A[370]), .A(S), .Z(O[370]) );
  ANDN U213 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U214 ( .B(A[369]), .A(S), .Z(O[369]) );
  ANDN U215 ( .B(A[368]), .A(S), .Z(O[368]) );
  ANDN U216 ( .B(A[367]), .A(S), .Z(O[367]) );
  ANDN U217 ( .B(A[366]), .A(S), .Z(O[366]) );
  ANDN U218 ( .B(A[365]), .A(S), .Z(O[365]) );
  ANDN U219 ( .B(A[364]), .A(S), .Z(O[364]) );
  ANDN U220 ( .B(A[363]), .A(S), .Z(O[363]) );
  ANDN U221 ( .B(A[362]), .A(S), .Z(O[362]) );
  ANDN U222 ( .B(A[361]), .A(S), .Z(O[361]) );
  ANDN U223 ( .B(A[360]), .A(S), .Z(O[360]) );
  ANDN U224 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U225 ( .B(A[359]), .A(S), .Z(O[359]) );
  ANDN U226 ( .B(A[358]), .A(S), .Z(O[358]) );
  ANDN U227 ( .B(A[357]), .A(S), .Z(O[357]) );
  ANDN U228 ( .B(A[356]), .A(S), .Z(O[356]) );
  ANDN U229 ( .B(A[355]), .A(S), .Z(O[355]) );
  ANDN U230 ( .B(A[354]), .A(S), .Z(O[354]) );
  ANDN U231 ( .B(A[353]), .A(S), .Z(O[353]) );
  ANDN U232 ( .B(A[352]), .A(S), .Z(O[352]) );
  ANDN U233 ( .B(A[351]), .A(S), .Z(O[351]) );
  ANDN U234 ( .B(A[350]), .A(S), .Z(O[350]) );
  ANDN U235 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U236 ( .B(A[349]), .A(S), .Z(O[349]) );
  ANDN U237 ( .B(A[348]), .A(S), .Z(O[348]) );
  ANDN U238 ( .B(A[347]), .A(S), .Z(O[347]) );
  ANDN U239 ( .B(A[346]), .A(S), .Z(O[346]) );
  ANDN U240 ( .B(A[345]), .A(S), .Z(O[345]) );
  ANDN U241 ( .B(A[344]), .A(S), .Z(O[344]) );
  ANDN U242 ( .B(A[343]), .A(S), .Z(O[343]) );
  ANDN U243 ( .B(A[342]), .A(S), .Z(O[342]) );
  ANDN U244 ( .B(A[341]), .A(S), .Z(O[341]) );
  ANDN U245 ( .B(A[340]), .A(S), .Z(O[340]) );
  ANDN U246 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U247 ( .B(A[339]), .A(S), .Z(O[339]) );
  ANDN U248 ( .B(A[338]), .A(S), .Z(O[338]) );
  ANDN U249 ( .B(A[337]), .A(S), .Z(O[337]) );
  ANDN U250 ( .B(A[336]), .A(S), .Z(O[336]) );
  ANDN U251 ( .B(A[335]), .A(S), .Z(O[335]) );
  ANDN U252 ( .B(A[334]), .A(S), .Z(O[334]) );
  ANDN U253 ( .B(A[333]), .A(S), .Z(O[333]) );
  ANDN U254 ( .B(A[332]), .A(S), .Z(O[332]) );
  ANDN U255 ( .B(A[331]), .A(S), .Z(O[331]) );
  ANDN U256 ( .B(A[330]), .A(S), .Z(O[330]) );
  ANDN U257 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U258 ( .B(A[329]), .A(S), .Z(O[329]) );
  ANDN U259 ( .B(A[328]), .A(S), .Z(O[328]) );
  ANDN U260 ( .B(A[327]), .A(S), .Z(O[327]) );
  ANDN U261 ( .B(A[326]), .A(S), .Z(O[326]) );
  ANDN U262 ( .B(A[325]), .A(S), .Z(O[325]) );
  ANDN U263 ( .B(A[324]), .A(S), .Z(O[324]) );
  ANDN U264 ( .B(A[323]), .A(S), .Z(O[323]) );
  ANDN U265 ( .B(A[322]), .A(S), .Z(O[322]) );
  ANDN U266 ( .B(A[321]), .A(S), .Z(O[321]) );
  ANDN U267 ( .B(A[320]), .A(S), .Z(O[320]) );
  ANDN U268 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U269 ( .B(A[319]), .A(S), .Z(O[319]) );
  ANDN U270 ( .B(A[318]), .A(S), .Z(O[318]) );
  ANDN U271 ( .B(A[317]), .A(S), .Z(O[317]) );
  ANDN U272 ( .B(A[316]), .A(S), .Z(O[316]) );
  ANDN U273 ( .B(A[315]), .A(S), .Z(O[315]) );
  ANDN U274 ( .B(A[314]), .A(S), .Z(O[314]) );
  ANDN U275 ( .B(A[313]), .A(S), .Z(O[313]) );
  ANDN U276 ( .B(A[312]), .A(S), .Z(O[312]) );
  ANDN U277 ( .B(A[311]), .A(S), .Z(O[311]) );
  ANDN U278 ( .B(A[310]), .A(S), .Z(O[310]) );
  ANDN U279 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U280 ( .B(A[309]), .A(S), .Z(O[309]) );
  ANDN U281 ( .B(A[308]), .A(S), .Z(O[308]) );
  ANDN U282 ( .B(A[307]), .A(S), .Z(O[307]) );
  ANDN U283 ( .B(A[306]), .A(S), .Z(O[306]) );
  ANDN U284 ( .B(A[305]), .A(S), .Z(O[305]) );
  ANDN U285 ( .B(A[304]), .A(S), .Z(O[304]) );
  ANDN U286 ( .B(A[303]), .A(S), .Z(O[303]) );
  ANDN U287 ( .B(A[302]), .A(S), .Z(O[302]) );
  ANDN U288 ( .B(A[301]), .A(S), .Z(O[301]) );
  ANDN U289 ( .B(A[300]), .A(S), .Z(O[300]) );
  ANDN U290 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U291 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U292 ( .B(A[299]), .A(S), .Z(O[299]) );
  ANDN U293 ( .B(A[298]), .A(S), .Z(O[298]) );
  ANDN U294 ( .B(A[297]), .A(S), .Z(O[297]) );
  ANDN U295 ( .B(A[296]), .A(S), .Z(O[296]) );
  ANDN U296 ( .B(A[295]), .A(S), .Z(O[295]) );
  ANDN U297 ( .B(A[294]), .A(S), .Z(O[294]) );
  ANDN U298 ( .B(A[293]), .A(S), .Z(O[293]) );
  ANDN U299 ( .B(A[292]), .A(S), .Z(O[292]) );
  ANDN U300 ( .B(A[291]), .A(S), .Z(O[291]) );
  ANDN U301 ( .B(A[290]), .A(S), .Z(O[290]) );
  ANDN U302 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U303 ( .B(A[289]), .A(S), .Z(O[289]) );
  ANDN U304 ( .B(A[288]), .A(S), .Z(O[288]) );
  ANDN U305 ( .B(A[287]), .A(S), .Z(O[287]) );
  ANDN U306 ( .B(A[286]), .A(S), .Z(O[286]) );
  ANDN U307 ( .B(A[285]), .A(S), .Z(O[285]) );
  ANDN U308 ( .B(A[284]), .A(S), .Z(O[284]) );
  ANDN U309 ( .B(A[283]), .A(S), .Z(O[283]) );
  ANDN U310 ( .B(A[282]), .A(S), .Z(O[282]) );
  ANDN U311 ( .B(A[281]), .A(S), .Z(O[281]) );
  ANDN U312 ( .B(A[280]), .A(S), .Z(O[280]) );
  ANDN U313 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U314 ( .B(A[279]), .A(S), .Z(O[279]) );
  ANDN U315 ( .B(A[278]), .A(S), .Z(O[278]) );
  ANDN U316 ( .B(A[277]), .A(S), .Z(O[277]) );
  ANDN U317 ( .B(A[276]), .A(S), .Z(O[276]) );
  ANDN U318 ( .B(A[275]), .A(S), .Z(O[275]) );
  ANDN U319 ( .B(A[274]), .A(S), .Z(O[274]) );
  ANDN U320 ( .B(A[273]), .A(S), .Z(O[273]) );
  ANDN U321 ( .B(A[272]), .A(S), .Z(O[272]) );
  ANDN U322 ( .B(A[271]), .A(S), .Z(O[271]) );
  ANDN U323 ( .B(A[270]), .A(S), .Z(O[270]) );
  ANDN U324 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U325 ( .B(A[269]), .A(S), .Z(O[269]) );
  ANDN U326 ( .B(A[268]), .A(S), .Z(O[268]) );
  ANDN U327 ( .B(A[267]), .A(S), .Z(O[267]) );
  ANDN U328 ( .B(A[266]), .A(S), .Z(O[266]) );
  ANDN U329 ( .B(A[265]), .A(S), .Z(O[265]) );
  ANDN U330 ( .B(A[264]), .A(S), .Z(O[264]) );
  ANDN U331 ( .B(A[263]), .A(S), .Z(O[263]) );
  ANDN U332 ( .B(A[262]), .A(S), .Z(O[262]) );
  ANDN U333 ( .B(A[261]), .A(S), .Z(O[261]) );
  ANDN U334 ( .B(A[260]), .A(S), .Z(O[260]) );
  ANDN U335 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U336 ( .B(A[259]), .A(S), .Z(O[259]) );
  ANDN U337 ( .B(A[258]), .A(S), .Z(O[258]) );
  ANDN U338 ( .B(A[257]), .A(S), .Z(O[257]) );
  ANDN U339 ( .B(A[256]), .A(S), .Z(O[256]) );
  ANDN U340 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U341 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U342 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U343 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U344 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U345 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U346 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U347 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U348 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U349 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U350 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U351 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U352 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U353 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U354 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U355 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U356 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U357 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U358 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U359 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U360 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U361 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U362 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U363 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U364 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U365 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U366 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U367 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U368 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U369 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U370 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U371 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U372 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U373 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U374 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U375 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U376 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U377 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U378 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U379 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U380 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U381 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U382 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U383 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U384 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U385 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U386 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U387 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U388 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U389 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U390 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U391 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U392 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U393 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U394 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U395 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U396 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U397 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U398 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U399 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U400 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U401 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U402 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U403 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U404 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U405 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U406 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U407 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U408 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U409 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U410 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U411 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U412 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U413 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U414 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U415 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U416 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U417 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U418 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U419 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U420 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U421 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U422 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U423 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U424 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U425 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U426 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U427 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U428 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U429 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U430 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U431 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U432 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U433 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U434 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U435 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U436 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U437 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U438 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U439 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U440 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U441 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U442 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U443 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U444 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U445 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U446 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U447 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U448 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U449 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U450 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U451 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U452 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U453 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U454 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U455 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U456 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U457 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U458 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U459 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U460 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U461 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U462 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U463 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U464 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U465 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U466 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U467 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U468 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U469 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U470 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U471 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U472 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U473 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U474 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U475 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U476 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U477 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U478 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U479 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U480 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U481 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U482 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U483 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U484 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U485 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U486 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U487 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U488 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U489 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U490 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U491 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U492 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U493 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U494 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U495 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U496 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U497 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U498 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U499 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U500 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U501 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U502 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U503 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U504 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U505 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U506 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U507 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U508 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U509 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U510 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U511 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U512 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module FA_1290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_5924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_5925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  ANDN U1 ( .B(CI), .A(S), .Z(CO) );
  XOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_5926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N514 ( A, B, CI, S, CO );
  input [513:0] A;
  input [513:0] B;
  output [513:0] S;
  input CI;
  output CO;

  wire   [513:1] C;

  FA_1290 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(1'b0), .B(B[0]), .CI(1'b0), .S(
        S[0]) );
  FA_6436 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(
        S[1]), .CO(C[2]) );
  FA_6435 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(
        S[2]), .CO(C[3]) );
  FA_6434 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(
        S[3]), .CO(C[4]) );
  FA_6433 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(
        S[4]), .CO(C[5]) );
  FA_6432 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(
        S[5]), .CO(C[6]) );
  FA_6431 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(
        S[6]), .CO(C[7]) );
  FA_6430 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(
        S[7]), .CO(C[8]) );
  FA_6429 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(
        S[8]), .CO(C[9]) );
  FA_6428 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(
        S[9]), .CO(C[10]) );
  FA_6427 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_6426 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_6425 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_6424 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_6423 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_6422 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_6421 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_6420 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_6419 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_6418 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_6417 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_6416 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_6415 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_6414 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_6413 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_6412 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_6411 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_6410 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_6409 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_6408 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_6407 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_6406 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_6405 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(B[32]), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_6404 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(B[33]), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_6403 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(B[34]), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_6402 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(B[35]), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_6401 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(B[36]), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_6400 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(B[37]), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_6399 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(B[38]), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_6398 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(B[39]), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_6397 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(B[40]), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_6396 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(B[41]), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_6395 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(B[42]), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_6394 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(B[43]), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_6393 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(B[44]), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_6392 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(B[45]), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_6391 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(B[46]), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_6390 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(B[47]), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_6389 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(B[48]), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_6388 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(B[49]), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_6387 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(B[50]), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_6386 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(B[51]), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_6385 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(B[52]), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_6384 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(B[53]), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_6383 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(B[54]), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_6382 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(B[55]), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_6381 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(B[56]), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_6380 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(B[57]), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_6379 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(B[58]), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_6378 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(B[59]), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_6377 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(B[60]), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_6376 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(B[61]), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_6375 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(B[62]), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_6374 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(B[63]), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_6373 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(B[64]), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_6372 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(B[65]), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_6371 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(B[66]), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_6370 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(B[67]), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_6369 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(B[68]), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_6368 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(B[69]), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_6367 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(B[70]), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_6366 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(B[71]), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_6365 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(B[72]), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_6364 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(B[73]), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_6363 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(B[74]), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_6362 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(B[75]), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_6361 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(B[76]), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_6360 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(B[77]), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_6359 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(B[78]), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_6358 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(B[79]), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_6357 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(B[80]), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_6356 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(B[81]), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_6355 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(B[82]), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_6354 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(B[83]), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_6353 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(B[84]), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_6352 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(B[85]), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_6351 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(B[86]), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_6350 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(B[87]), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_6349 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(B[88]), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_6348 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(B[89]), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_6347 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(B[90]), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_6346 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(B[91]), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_6345 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(B[92]), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_6344 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(B[93]), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_6343 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(B[94]), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_6342 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(B[95]), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_6341 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(B[96]), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_6340 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(B[97]), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_6339 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(B[98]), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_6338 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(B[99]), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_6337 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(B[100]), .CI(
        C[100]), .S(S[100]), .CO(C[101]) );
  FA_6336 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(B[101]), .CI(
        C[101]), .S(S[101]), .CO(C[102]) );
  FA_6335 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(B[102]), .CI(
        C[102]), .S(S[102]), .CO(C[103]) );
  FA_6334 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(B[103]), .CI(
        C[103]), .S(S[103]), .CO(C[104]) );
  FA_6333 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(B[104]), .CI(
        C[104]), .S(S[104]), .CO(C[105]) );
  FA_6332 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(B[105]), .CI(
        C[105]), .S(S[105]), .CO(C[106]) );
  FA_6331 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(B[106]), .CI(
        C[106]), .S(S[106]), .CO(C[107]) );
  FA_6330 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(B[107]), .CI(
        C[107]), .S(S[107]), .CO(C[108]) );
  FA_6329 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(B[108]), .CI(
        C[108]), .S(S[108]), .CO(C[109]) );
  FA_6328 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(B[109]), .CI(
        C[109]), .S(S[109]), .CO(C[110]) );
  FA_6327 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(B[110]), .CI(
        C[110]), .S(S[110]), .CO(C[111]) );
  FA_6326 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(B[111]), .CI(
        C[111]), .S(S[111]), .CO(C[112]) );
  FA_6325 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(B[112]), .CI(
        C[112]), .S(S[112]), .CO(C[113]) );
  FA_6324 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(B[113]), .CI(
        C[113]), .S(S[113]), .CO(C[114]) );
  FA_6323 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(B[114]), .CI(
        C[114]), .S(S[114]), .CO(C[115]) );
  FA_6322 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(B[115]), .CI(
        C[115]), .S(S[115]), .CO(C[116]) );
  FA_6321 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(B[116]), .CI(
        C[116]), .S(S[116]), .CO(C[117]) );
  FA_6320 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(B[117]), .CI(
        C[117]), .S(S[117]), .CO(C[118]) );
  FA_6319 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(B[118]), .CI(
        C[118]), .S(S[118]), .CO(C[119]) );
  FA_6318 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(B[119]), .CI(
        C[119]), .S(S[119]), .CO(C[120]) );
  FA_6317 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(B[120]), .CI(
        C[120]), .S(S[120]), .CO(C[121]) );
  FA_6316 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(B[121]), .CI(
        C[121]), .S(S[121]), .CO(C[122]) );
  FA_6315 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(B[122]), .CI(
        C[122]), .S(S[122]), .CO(C[123]) );
  FA_6314 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(B[123]), .CI(
        C[123]), .S(S[123]), .CO(C[124]) );
  FA_6313 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(B[124]), .CI(
        C[124]), .S(S[124]), .CO(C[125]) );
  FA_6312 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(B[125]), .CI(
        C[125]), .S(S[125]), .CO(C[126]) );
  FA_6311 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(B[126]), .CI(
        C[126]), .S(S[126]), .CO(C[127]) );
  FA_6310 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(B[127]), .CI(
        C[127]), .S(S[127]), .CO(C[128]) );
  FA_6309 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(B[128]), .CI(
        C[128]), .S(S[128]), .CO(C[129]) );
  FA_6308 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(B[129]), .CI(
        C[129]), .S(S[129]), .CO(C[130]) );
  FA_6307 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(B[130]), .CI(
        C[130]), .S(S[130]), .CO(C[131]) );
  FA_6306 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(B[131]), .CI(
        C[131]), .S(S[131]), .CO(C[132]) );
  FA_6305 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(B[132]), .CI(
        C[132]), .S(S[132]), .CO(C[133]) );
  FA_6304 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(B[133]), .CI(
        C[133]), .S(S[133]), .CO(C[134]) );
  FA_6303 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(B[134]), .CI(
        C[134]), .S(S[134]), .CO(C[135]) );
  FA_6302 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(B[135]), .CI(
        C[135]), .S(S[135]), .CO(C[136]) );
  FA_6301 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(B[136]), .CI(
        C[136]), .S(S[136]), .CO(C[137]) );
  FA_6300 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(B[137]), .CI(
        C[137]), .S(S[137]), .CO(C[138]) );
  FA_6299 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(B[138]), .CI(
        C[138]), .S(S[138]), .CO(C[139]) );
  FA_6298 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(B[139]), .CI(
        C[139]), .S(S[139]), .CO(C[140]) );
  FA_6297 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(B[140]), .CI(
        C[140]), .S(S[140]), .CO(C[141]) );
  FA_6296 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(B[141]), .CI(
        C[141]), .S(S[141]), .CO(C[142]) );
  FA_6295 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(B[142]), .CI(
        C[142]), .S(S[142]), .CO(C[143]) );
  FA_6294 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(B[143]), .CI(
        C[143]), .S(S[143]), .CO(C[144]) );
  FA_6293 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(B[144]), .CI(
        C[144]), .S(S[144]), .CO(C[145]) );
  FA_6292 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(B[145]), .CI(
        C[145]), .S(S[145]), .CO(C[146]) );
  FA_6291 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(B[146]), .CI(
        C[146]), .S(S[146]), .CO(C[147]) );
  FA_6290 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(B[147]), .CI(
        C[147]), .S(S[147]), .CO(C[148]) );
  FA_6289 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(B[148]), .CI(
        C[148]), .S(S[148]), .CO(C[149]) );
  FA_6288 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(B[149]), .CI(
        C[149]), .S(S[149]), .CO(C[150]) );
  FA_6287 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(B[150]), .CI(
        C[150]), .S(S[150]), .CO(C[151]) );
  FA_6286 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(B[151]), .CI(
        C[151]), .S(S[151]), .CO(C[152]) );
  FA_6285 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(B[152]), .CI(
        C[152]), .S(S[152]), .CO(C[153]) );
  FA_6284 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(B[153]), .CI(
        C[153]), .S(S[153]), .CO(C[154]) );
  FA_6283 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(B[154]), .CI(
        C[154]), .S(S[154]), .CO(C[155]) );
  FA_6282 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(B[155]), .CI(
        C[155]), .S(S[155]), .CO(C[156]) );
  FA_6281 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(B[156]), .CI(
        C[156]), .S(S[156]), .CO(C[157]) );
  FA_6280 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(B[157]), .CI(
        C[157]), .S(S[157]), .CO(C[158]) );
  FA_6279 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(B[158]), .CI(
        C[158]), .S(S[158]), .CO(C[159]) );
  FA_6278 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(B[159]), .CI(
        C[159]), .S(S[159]), .CO(C[160]) );
  FA_6277 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(B[160]), .CI(
        C[160]), .S(S[160]), .CO(C[161]) );
  FA_6276 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(B[161]), .CI(
        C[161]), .S(S[161]), .CO(C[162]) );
  FA_6275 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(B[162]), .CI(
        C[162]), .S(S[162]), .CO(C[163]) );
  FA_6274 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(B[163]), .CI(
        C[163]), .S(S[163]), .CO(C[164]) );
  FA_6273 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(B[164]), .CI(
        C[164]), .S(S[164]), .CO(C[165]) );
  FA_6272 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(B[165]), .CI(
        C[165]), .S(S[165]), .CO(C[166]) );
  FA_6271 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(B[166]), .CI(
        C[166]), .S(S[166]), .CO(C[167]) );
  FA_6270 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(B[167]), .CI(
        C[167]), .S(S[167]), .CO(C[168]) );
  FA_6269 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(B[168]), .CI(
        C[168]), .S(S[168]), .CO(C[169]) );
  FA_6268 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(B[169]), .CI(
        C[169]), .S(S[169]), .CO(C[170]) );
  FA_6267 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(B[170]), .CI(
        C[170]), .S(S[170]), .CO(C[171]) );
  FA_6266 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(B[171]), .CI(
        C[171]), .S(S[171]), .CO(C[172]) );
  FA_6265 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(B[172]), .CI(
        C[172]), .S(S[172]), .CO(C[173]) );
  FA_6264 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(B[173]), .CI(
        C[173]), .S(S[173]), .CO(C[174]) );
  FA_6263 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(B[174]), .CI(
        C[174]), .S(S[174]), .CO(C[175]) );
  FA_6262 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(B[175]), .CI(
        C[175]), .S(S[175]), .CO(C[176]) );
  FA_6261 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(B[176]), .CI(
        C[176]), .S(S[176]), .CO(C[177]) );
  FA_6260 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(B[177]), .CI(
        C[177]), .S(S[177]), .CO(C[178]) );
  FA_6259 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(B[178]), .CI(
        C[178]), .S(S[178]), .CO(C[179]) );
  FA_6258 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(B[179]), .CI(
        C[179]), .S(S[179]), .CO(C[180]) );
  FA_6257 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(B[180]), .CI(
        C[180]), .S(S[180]), .CO(C[181]) );
  FA_6256 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(B[181]), .CI(
        C[181]), .S(S[181]), .CO(C[182]) );
  FA_6255 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(B[182]), .CI(
        C[182]), .S(S[182]), .CO(C[183]) );
  FA_6254 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(B[183]), .CI(
        C[183]), .S(S[183]), .CO(C[184]) );
  FA_6253 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(B[184]), .CI(
        C[184]), .S(S[184]), .CO(C[185]) );
  FA_6252 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(B[185]), .CI(
        C[185]), .S(S[185]), .CO(C[186]) );
  FA_6251 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(B[186]), .CI(
        C[186]), .S(S[186]), .CO(C[187]) );
  FA_6250 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(B[187]), .CI(
        C[187]), .S(S[187]), .CO(C[188]) );
  FA_6249 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(B[188]), .CI(
        C[188]), .S(S[188]), .CO(C[189]) );
  FA_6248 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(B[189]), .CI(
        C[189]), .S(S[189]), .CO(C[190]) );
  FA_6247 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(B[190]), .CI(
        C[190]), .S(S[190]), .CO(C[191]) );
  FA_6246 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(B[191]), .CI(
        C[191]), .S(S[191]), .CO(C[192]) );
  FA_6245 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(B[192]), .CI(
        C[192]), .S(S[192]), .CO(C[193]) );
  FA_6244 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(B[193]), .CI(
        C[193]), .S(S[193]), .CO(C[194]) );
  FA_6243 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(B[194]), .CI(
        C[194]), .S(S[194]), .CO(C[195]) );
  FA_6242 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(B[195]), .CI(
        C[195]), .S(S[195]), .CO(C[196]) );
  FA_6241 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(B[196]), .CI(
        C[196]), .S(S[196]), .CO(C[197]) );
  FA_6240 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(B[197]), .CI(
        C[197]), .S(S[197]), .CO(C[198]) );
  FA_6239 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(B[198]), .CI(
        C[198]), .S(S[198]), .CO(C[199]) );
  FA_6238 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(B[199]), .CI(
        C[199]), .S(S[199]), .CO(C[200]) );
  FA_6237 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(B[200]), .CI(
        C[200]), .S(S[200]), .CO(C[201]) );
  FA_6236 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(B[201]), .CI(
        C[201]), .S(S[201]), .CO(C[202]) );
  FA_6235 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(B[202]), .CI(
        C[202]), .S(S[202]), .CO(C[203]) );
  FA_6234 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(B[203]), .CI(
        C[203]), .S(S[203]), .CO(C[204]) );
  FA_6233 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(B[204]), .CI(
        C[204]), .S(S[204]), .CO(C[205]) );
  FA_6232 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(B[205]), .CI(
        C[205]), .S(S[205]), .CO(C[206]) );
  FA_6231 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(B[206]), .CI(
        C[206]), .S(S[206]), .CO(C[207]) );
  FA_6230 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(B[207]), .CI(
        C[207]), .S(S[207]), .CO(C[208]) );
  FA_6229 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(B[208]), .CI(
        C[208]), .S(S[208]), .CO(C[209]) );
  FA_6228 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(B[209]), .CI(
        C[209]), .S(S[209]), .CO(C[210]) );
  FA_6227 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(B[210]), .CI(
        C[210]), .S(S[210]), .CO(C[211]) );
  FA_6226 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(B[211]), .CI(
        C[211]), .S(S[211]), .CO(C[212]) );
  FA_6225 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(B[212]), .CI(
        C[212]), .S(S[212]), .CO(C[213]) );
  FA_6224 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(B[213]), .CI(
        C[213]), .S(S[213]), .CO(C[214]) );
  FA_6223 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(B[214]), .CI(
        C[214]), .S(S[214]), .CO(C[215]) );
  FA_6222 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(B[215]), .CI(
        C[215]), .S(S[215]), .CO(C[216]) );
  FA_6221 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(B[216]), .CI(
        C[216]), .S(S[216]), .CO(C[217]) );
  FA_6220 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(B[217]), .CI(
        C[217]), .S(S[217]), .CO(C[218]) );
  FA_6219 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(B[218]), .CI(
        C[218]), .S(S[218]), .CO(C[219]) );
  FA_6218 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(B[219]), .CI(
        C[219]), .S(S[219]), .CO(C[220]) );
  FA_6217 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(B[220]), .CI(
        C[220]), .S(S[220]), .CO(C[221]) );
  FA_6216 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(B[221]), .CI(
        C[221]), .S(S[221]), .CO(C[222]) );
  FA_6215 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(B[222]), .CI(
        C[222]), .S(S[222]), .CO(C[223]) );
  FA_6214 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(B[223]), .CI(
        C[223]), .S(S[223]), .CO(C[224]) );
  FA_6213 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(B[224]), .CI(
        C[224]), .S(S[224]), .CO(C[225]) );
  FA_6212 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(B[225]), .CI(
        C[225]), .S(S[225]), .CO(C[226]) );
  FA_6211 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(B[226]), .CI(
        C[226]), .S(S[226]), .CO(C[227]) );
  FA_6210 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(B[227]), .CI(
        C[227]), .S(S[227]), .CO(C[228]) );
  FA_6209 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(B[228]), .CI(
        C[228]), .S(S[228]), .CO(C[229]) );
  FA_6208 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(B[229]), .CI(
        C[229]), .S(S[229]), .CO(C[230]) );
  FA_6207 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(B[230]), .CI(
        C[230]), .S(S[230]), .CO(C[231]) );
  FA_6206 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(B[231]), .CI(
        C[231]), .S(S[231]), .CO(C[232]) );
  FA_6205 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(B[232]), .CI(
        C[232]), .S(S[232]), .CO(C[233]) );
  FA_6204 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(B[233]), .CI(
        C[233]), .S(S[233]), .CO(C[234]) );
  FA_6203 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(B[234]), .CI(
        C[234]), .S(S[234]), .CO(C[235]) );
  FA_6202 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(B[235]), .CI(
        C[235]), .S(S[235]), .CO(C[236]) );
  FA_6201 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(B[236]), .CI(
        C[236]), .S(S[236]), .CO(C[237]) );
  FA_6200 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(B[237]), .CI(
        C[237]), .S(S[237]), .CO(C[238]) );
  FA_6199 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(B[238]), .CI(
        C[238]), .S(S[238]), .CO(C[239]) );
  FA_6198 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(B[239]), .CI(
        C[239]), .S(S[239]), .CO(C[240]) );
  FA_6197 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(B[240]), .CI(
        C[240]), .S(S[240]), .CO(C[241]) );
  FA_6196 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(B[241]), .CI(
        C[241]), .S(S[241]), .CO(C[242]) );
  FA_6195 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(B[242]), .CI(
        C[242]), .S(S[242]), .CO(C[243]) );
  FA_6194 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(B[243]), .CI(
        C[243]), .S(S[243]), .CO(C[244]) );
  FA_6193 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(B[244]), .CI(
        C[244]), .S(S[244]), .CO(C[245]) );
  FA_6192 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(B[245]), .CI(
        C[245]), .S(S[245]), .CO(C[246]) );
  FA_6191 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(B[246]), .CI(
        C[246]), .S(S[246]), .CO(C[247]) );
  FA_6190 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(B[247]), .CI(
        C[247]), .S(S[247]), .CO(C[248]) );
  FA_6189 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(B[248]), .CI(
        C[248]), .S(S[248]), .CO(C[249]) );
  FA_6188 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(B[249]), .CI(
        C[249]), .S(S[249]), .CO(C[250]) );
  FA_6187 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(B[250]), .CI(
        C[250]), .S(S[250]), .CO(C[251]) );
  FA_6186 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(B[251]), .CI(
        C[251]), .S(S[251]), .CO(C[252]) );
  FA_6185 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(B[252]), .CI(
        C[252]), .S(S[252]), .CO(C[253]) );
  FA_6184 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(B[253]), .CI(
        C[253]), .S(S[253]), .CO(C[254]) );
  FA_6183 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(B[254]), .CI(
        C[254]), .S(S[254]), .CO(C[255]) );
  FA_6182 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(B[255]), .CI(
        C[255]), .S(S[255]), .CO(C[256]) );
  FA_6181 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(B[256]), .CI(
        C[256]), .S(S[256]), .CO(C[257]) );
  FA_6180 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(B[257]), .CI(
        C[257]), .S(S[257]), .CO(C[258]) );
  FA_6179 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(B[258]), .CI(
        C[258]), .S(S[258]), .CO(C[259]) );
  FA_6178 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(B[259]), .CI(
        C[259]), .S(S[259]), .CO(C[260]) );
  FA_6177 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(B[260]), .CI(
        C[260]), .S(S[260]), .CO(C[261]) );
  FA_6176 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(B[261]), .CI(
        C[261]), .S(S[261]), .CO(C[262]) );
  FA_6175 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(B[262]), .CI(
        C[262]), .S(S[262]), .CO(C[263]) );
  FA_6174 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(B[263]), .CI(
        C[263]), .S(S[263]), .CO(C[264]) );
  FA_6173 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(B[264]), .CI(
        C[264]), .S(S[264]), .CO(C[265]) );
  FA_6172 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(B[265]), .CI(
        C[265]), .S(S[265]), .CO(C[266]) );
  FA_6171 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(B[266]), .CI(
        C[266]), .S(S[266]), .CO(C[267]) );
  FA_6170 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(B[267]), .CI(
        C[267]), .S(S[267]), .CO(C[268]) );
  FA_6169 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(B[268]), .CI(
        C[268]), .S(S[268]), .CO(C[269]) );
  FA_6168 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(B[269]), .CI(
        C[269]), .S(S[269]), .CO(C[270]) );
  FA_6167 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(B[270]), .CI(
        C[270]), .S(S[270]), .CO(C[271]) );
  FA_6166 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(B[271]), .CI(
        C[271]), .S(S[271]), .CO(C[272]) );
  FA_6165 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(B[272]), .CI(
        C[272]), .S(S[272]), .CO(C[273]) );
  FA_6164 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(B[273]), .CI(
        C[273]), .S(S[273]), .CO(C[274]) );
  FA_6163 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(B[274]), .CI(
        C[274]), .S(S[274]), .CO(C[275]) );
  FA_6162 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(B[275]), .CI(
        C[275]), .S(S[275]), .CO(C[276]) );
  FA_6161 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(B[276]), .CI(
        C[276]), .S(S[276]), .CO(C[277]) );
  FA_6160 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(B[277]), .CI(
        C[277]), .S(S[277]), .CO(C[278]) );
  FA_6159 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(B[278]), .CI(
        C[278]), .S(S[278]), .CO(C[279]) );
  FA_6158 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(B[279]), .CI(
        C[279]), .S(S[279]), .CO(C[280]) );
  FA_6157 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(B[280]), .CI(
        C[280]), .S(S[280]), .CO(C[281]) );
  FA_6156 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(B[281]), .CI(
        C[281]), .S(S[281]), .CO(C[282]) );
  FA_6155 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(B[282]), .CI(
        C[282]), .S(S[282]), .CO(C[283]) );
  FA_6154 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(B[283]), .CI(
        C[283]), .S(S[283]), .CO(C[284]) );
  FA_6153 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(B[284]), .CI(
        C[284]), .S(S[284]), .CO(C[285]) );
  FA_6152 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(B[285]), .CI(
        C[285]), .S(S[285]), .CO(C[286]) );
  FA_6151 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(B[286]), .CI(
        C[286]), .S(S[286]), .CO(C[287]) );
  FA_6150 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(B[287]), .CI(
        C[287]), .S(S[287]), .CO(C[288]) );
  FA_6149 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(B[288]), .CI(
        C[288]), .S(S[288]), .CO(C[289]) );
  FA_6148 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(B[289]), .CI(
        C[289]), .S(S[289]), .CO(C[290]) );
  FA_6147 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(B[290]), .CI(
        C[290]), .S(S[290]), .CO(C[291]) );
  FA_6146 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(B[291]), .CI(
        C[291]), .S(S[291]), .CO(C[292]) );
  FA_6145 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(B[292]), .CI(
        C[292]), .S(S[292]), .CO(C[293]) );
  FA_6144 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(B[293]), .CI(
        C[293]), .S(S[293]), .CO(C[294]) );
  FA_6143 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(B[294]), .CI(
        C[294]), .S(S[294]), .CO(C[295]) );
  FA_6142 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(B[295]), .CI(
        C[295]), .S(S[295]), .CO(C[296]) );
  FA_6141 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(B[296]), .CI(
        C[296]), .S(S[296]), .CO(C[297]) );
  FA_6140 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(B[297]), .CI(
        C[297]), .S(S[297]), .CO(C[298]) );
  FA_6139 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(B[298]), .CI(
        C[298]), .S(S[298]), .CO(C[299]) );
  FA_6138 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(B[299]), .CI(
        C[299]), .S(S[299]), .CO(C[300]) );
  FA_6137 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(B[300]), .CI(
        C[300]), .S(S[300]), .CO(C[301]) );
  FA_6136 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(B[301]), .CI(
        C[301]), .S(S[301]), .CO(C[302]) );
  FA_6135 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(B[302]), .CI(
        C[302]), .S(S[302]), .CO(C[303]) );
  FA_6134 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(B[303]), .CI(
        C[303]), .S(S[303]), .CO(C[304]) );
  FA_6133 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(B[304]), .CI(
        C[304]), .S(S[304]), .CO(C[305]) );
  FA_6132 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(B[305]), .CI(
        C[305]), .S(S[305]), .CO(C[306]) );
  FA_6131 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(B[306]), .CI(
        C[306]), .S(S[306]), .CO(C[307]) );
  FA_6130 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(B[307]), .CI(
        C[307]), .S(S[307]), .CO(C[308]) );
  FA_6129 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(B[308]), .CI(
        C[308]), .S(S[308]), .CO(C[309]) );
  FA_6128 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(B[309]), .CI(
        C[309]), .S(S[309]), .CO(C[310]) );
  FA_6127 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(B[310]), .CI(
        C[310]), .S(S[310]), .CO(C[311]) );
  FA_6126 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(B[311]), .CI(
        C[311]), .S(S[311]), .CO(C[312]) );
  FA_6125 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(B[312]), .CI(
        C[312]), .S(S[312]), .CO(C[313]) );
  FA_6124 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(B[313]), .CI(
        C[313]), .S(S[313]), .CO(C[314]) );
  FA_6123 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(B[314]), .CI(
        C[314]), .S(S[314]), .CO(C[315]) );
  FA_6122 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(B[315]), .CI(
        C[315]), .S(S[315]), .CO(C[316]) );
  FA_6121 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(B[316]), .CI(
        C[316]), .S(S[316]), .CO(C[317]) );
  FA_6120 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(B[317]), .CI(
        C[317]), .S(S[317]), .CO(C[318]) );
  FA_6119 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(B[318]), .CI(
        C[318]), .S(S[318]), .CO(C[319]) );
  FA_6118 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(B[319]), .CI(
        C[319]), .S(S[319]), .CO(C[320]) );
  FA_6117 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(B[320]), .CI(
        C[320]), .S(S[320]), .CO(C[321]) );
  FA_6116 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(B[321]), .CI(
        C[321]), .S(S[321]), .CO(C[322]) );
  FA_6115 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(B[322]), .CI(
        C[322]), .S(S[322]), .CO(C[323]) );
  FA_6114 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(B[323]), .CI(
        C[323]), .S(S[323]), .CO(C[324]) );
  FA_6113 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(B[324]), .CI(
        C[324]), .S(S[324]), .CO(C[325]) );
  FA_6112 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(B[325]), .CI(
        C[325]), .S(S[325]), .CO(C[326]) );
  FA_6111 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(B[326]), .CI(
        C[326]), .S(S[326]), .CO(C[327]) );
  FA_6110 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(B[327]), .CI(
        C[327]), .S(S[327]), .CO(C[328]) );
  FA_6109 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(B[328]), .CI(
        C[328]), .S(S[328]), .CO(C[329]) );
  FA_6108 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(B[329]), .CI(
        C[329]), .S(S[329]), .CO(C[330]) );
  FA_6107 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(B[330]), .CI(
        C[330]), .S(S[330]), .CO(C[331]) );
  FA_6106 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(B[331]), .CI(
        C[331]), .S(S[331]), .CO(C[332]) );
  FA_6105 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(B[332]), .CI(
        C[332]), .S(S[332]), .CO(C[333]) );
  FA_6104 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(B[333]), .CI(
        C[333]), .S(S[333]), .CO(C[334]) );
  FA_6103 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(B[334]), .CI(
        C[334]), .S(S[334]), .CO(C[335]) );
  FA_6102 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(B[335]), .CI(
        C[335]), .S(S[335]), .CO(C[336]) );
  FA_6101 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(B[336]), .CI(
        C[336]), .S(S[336]), .CO(C[337]) );
  FA_6100 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(B[337]), .CI(
        C[337]), .S(S[337]), .CO(C[338]) );
  FA_6099 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(B[338]), .CI(
        C[338]), .S(S[338]), .CO(C[339]) );
  FA_6098 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(B[339]), .CI(
        C[339]), .S(S[339]), .CO(C[340]) );
  FA_6097 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(B[340]), .CI(
        C[340]), .S(S[340]), .CO(C[341]) );
  FA_6096 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(B[341]), .CI(
        C[341]), .S(S[341]), .CO(C[342]) );
  FA_6095 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(B[342]), .CI(
        C[342]), .S(S[342]), .CO(C[343]) );
  FA_6094 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(B[343]), .CI(
        C[343]), .S(S[343]), .CO(C[344]) );
  FA_6093 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(B[344]), .CI(
        C[344]), .S(S[344]), .CO(C[345]) );
  FA_6092 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(B[345]), .CI(
        C[345]), .S(S[345]), .CO(C[346]) );
  FA_6091 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(B[346]), .CI(
        C[346]), .S(S[346]), .CO(C[347]) );
  FA_6090 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(B[347]), .CI(
        C[347]), .S(S[347]), .CO(C[348]) );
  FA_6089 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(B[348]), .CI(
        C[348]), .S(S[348]), .CO(C[349]) );
  FA_6088 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(B[349]), .CI(
        C[349]), .S(S[349]), .CO(C[350]) );
  FA_6087 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(B[350]), .CI(
        C[350]), .S(S[350]), .CO(C[351]) );
  FA_6086 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(B[351]), .CI(
        C[351]), .S(S[351]), .CO(C[352]) );
  FA_6085 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(B[352]), .CI(
        C[352]), .S(S[352]), .CO(C[353]) );
  FA_6084 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(B[353]), .CI(
        C[353]), .S(S[353]), .CO(C[354]) );
  FA_6083 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(B[354]), .CI(
        C[354]), .S(S[354]), .CO(C[355]) );
  FA_6082 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(B[355]), .CI(
        C[355]), .S(S[355]), .CO(C[356]) );
  FA_6081 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(B[356]), .CI(
        C[356]), .S(S[356]), .CO(C[357]) );
  FA_6080 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(B[357]), .CI(
        C[357]), .S(S[357]), .CO(C[358]) );
  FA_6079 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(B[358]), .CI(
        C[358]), .S(S[358]), .CO(C[359]) );
  FA_6078 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(B[359]), .CI(
        C[359]), .S(S[359]), .CO(C[360]) );
  FA_6077 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(B[360]), .CI(
        C[360]), .S(S[360]), .CO(C[361]) );
  FA_6076 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(B[361]), .CI(
        C[361]), .S(S[361]), .CO(C[362]) );
  FA_6075 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(B[362]), .CI(
        C[362]), .S(S[362]), .CO(C[363]) );
  FA_6074 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(B[363]), .CI(
        C[363]), .S(S[363]), .CO(C[364]) );
  FA_6073 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(B[364]), .CI(
        C[364]), .S(S[364]), .CO(C[365]) );
  FA_6072 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(B[365]), .CI(
        C[365]), .S(S[365]), .CO(C[366]) );
  FA_6071 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(B[366]), .CI(
        C[366]), .S(S[366]), .CO(C[367]) );
  FA_6070 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(B[367]), .CI(
        C[367]), .S(S[367]), .CO(C[368]) );
  FA_6069 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(B[368]), .CI(
        C[368]), .S(S[368]), .CO(C[369]) );
  FA_6068 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(B[369]), .CI(
        C[369]), .S(S[369]), .CO(C[370]) );
  FA_6067 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(B[370]), .CI(
        C[370]), .S(S[370]), .CO(C[371]) );
  FA_6066 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(B[371]), .CI(
        C[371]), .S(S[371]), .CO(C[372]) );
  FA_6065 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(B[372]), .CI(
        C[372]), .S(S[372]), .CO(C[373]) );
  FA_6064 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(B[373]), .CI(
        C[373]), .S(S[373]), .CO(C[374]) );
  FA_6063 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(B[374]), .CI(
        C[374]), .S(S[374]), .CO(C[375]) );
  FA_6062 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(B[375]), .CI(
        C[375]), .S(S[375]), .CO(C[376]) );
  FA_6061 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(B[376]), .CI(
        C[376]), .S(S[376]), .CO(C[377]) );
  FA_6060 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(B[377]), .CI(
        C[377]), .S(S[377]), .CO(C[378]) );
  FA_6059 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(B[378]), .CI(
        C[378]), .S(S[378]), .CO(C[379]) );
  FA_6058 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(B[379]), .CI(
        C[379]), .S(S[379]), .CO(C[380]) );
  FA_6057 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(B[380]), .CI(
        C[380]), .S(S[380]), .CO(C[381]) );
  FA_6056 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(B[381]), .CI(
        C[381]), .S(S[381]), .CO(C[382]) );
  FA_6055 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(B[382]), .CI(
        C[382]), .S(S[382]), .CO(C[383]) );
  FA_6054 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(B[383]), .CI(
        C[383]), .S(S[383]), .CO(C[384]) );
  FA_6053 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(B[384]), .CI(
        C[384]), .S(S[384]), .CO(C[385]) );
  FA_6052 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(B[385]), .CI(
        C[385]), .S(S[385]), .CO(C[386]) );
  FA_6051 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(B[386]), .CI(
        C[386]), .S(S[386]), .CO(C[387]) );
  FA_6050 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(B[387]), .CI(
        C[387]), .S(S[387]), .CO(C[388]) );
  FA_6049 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(B[388]), .CI(
        C[388]), .S(S[388]), .CO(C[389]) );
  FA_6048 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(B[389]), .CI(
        C[389]), .S(S[389]), .CO(C[390]) );
  FA_6047 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(B[390]), .CI(
        C[390]), .S(S[390]), .CO(C[391]) );
  FA_6046 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(B[391]), .CI(
        C[391]), .S(S[391]), .CO(C[392]) );
  FA_6045 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(B[392]), .CI(
        C[392]), .S(S[392]), .CO(C[393]) );
  FA_6044 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(B[393]), .CI(
        C[393]), .S(S[393]), .CO(C[394]) );
  FA_6043 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(B[394]), .CI(
        C[394]), .S(S[394]), .CO(C[395]) );
  FA_6042 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(B[395]), .CI(
        C[395]), .S(S[395]), .CO(C[396]) );
  FA_6041 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(B[396]), .CI(
        C[396]), .S(S[396]), .CO(C[397]) );
  FA_6040 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(B[397]), .CI(
        C[397]), .S(S[397]), .CO(C[398]) );
  FA_6039 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(B[398]), .CI(
        C[398]), .S(S[398]), .CO(C[399]) );
  FA_6038 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(B[399]), .CI(
        C[399]), .S(S[399]), .CO(C[400]) );
  FA_6037 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(B[400]), .CI(
        C[400]), .S(S[400]), .CO(C[401]) );
  FA_6036 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(B[401]), .CI(
        C[401]), .S(S[401]), .CO(C[402]) );
  FA_6035 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(B[402]), .CI(
        C[402]), .S(S[402]), .CO(C[403]) );
  FA_6034 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(B[403]), .CI(
        C[403]), .S(S[403]), .CO(C[404]) );
  FA_6033 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(B[404]), .CI(
        C[404]), .S(S[404]), .CO(C[405]) );
  FA_6032 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(B[405]), .CI(
        C[405]), .S(S[405]), .CO(C[406]) );
  FA_6031 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(B[406]), .CI(
        C[406]), .S(S[406]), .CO(C[407]) );
  FA_6030 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(B[407]), .CI(
        C[407]), .S(S[407]), .CO(C[408]) );
  FA_6029 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(B[408]), .CI(
        C[408]), .S(S[408]), .CO(C[409]) );
  FA_6028 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(B[409]), .CI(
        C[409]), .S(S[409]), .CO(C[410]) );
  FA_6027 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(B[410]), .CI(
        C[410]), .S(S[410]), .CO(C[411]) );
  FA_6026 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(B[411]), .CI(
        C[411]), .S(S[411]), .CO(C[412]) );
  FA_6025 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(B[412]), .CI(
        C[412]), .S(S[412]), .CO(C[413]) );
  FA_6024 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(B[413]), .CI(
        C[413]), .S(S[413]), .CO(C[414]) );
  FA_6023 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(B[414]), .CI(
        C[414]), .S(S[414]), .CO(C[415]) );
  FA_6022 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(B[415]), .CI(
        C[415]), .S(S[415]), .CO(C[416]) );
  FA_6021 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(B[416]), .CI(
        C[416]), .S(S[416]), .CO(C[417]) );
  FA_6020 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(B[417]), .CI(
        C[417]), .S(S[417]), .CO(C[418]) );
  FA_6019 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(B[418]), .CI(
        C[418]), .S(S[418]), .CO(C[419]) );
  FA_6018 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(B[419]), .CI(
        C[419]), .S(S[419]), .CO(C[420]) );
  FA_6017 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(B[420]), .CI(
        C[420]), .S(S[420]), .CO(C[421]) );
  FA_6016 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(B[421]), .CI(
        C[421]), .S(S[421]), .CO(C[422]) );
  FA_6015 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(B[422]), .CI(
        C[422]), .S(S[422]), .CO(C[423]) );
  FA_6014 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(B[423]), .CI(
        C[423]), .S(S[423]), .CO(C[424]) );
  FA_6013 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(B[424]), .CI(
        C[424]), .S(S[424]), .CO(C[425]) );
  FA_6012 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(B[425]), .CI(
        C[425]), .S(S[425]), .CO(C[426]) );
  FA_6011 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(B[426]), .CI(
        C[426]), .S(S[426]), .CO(C[427]) );
  FA_6010 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(B[427]), .CI(
        C[427]), .S(S[427]), .CO(C[428]) );
  FA_6009 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(B[428]), .CI(
        C[428]), .S(S[428]), .CO(C[429]) );
  FA_6008 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(B[429]), .CI(
        C[429]), .S(S[429]), .CO(C[430]) );
  FA_6007 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(B[430]), .CI(
        C[430]), .S(S[430]), .CO(C[431]) );
  FA_6006 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(B[431]), .CI(
        C[431]), .S(S[431]), .CO(C[432]) );
  FA_6005 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(B[432]), .CI(
        C[432]), .S(S[432]), .CO(C[433]) );
  FA_6004 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(B[433]), .CI(
        C[433]), .S(S[433]), .CO(C[434]) );
  FA_6003 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(B[434]), .CI(
        C[434]), .S(S[434]), .CO(C[435]) );
  FA_6002 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(B[435]), .CI(
        C[435]), .S(S[435]), .CO(C[436]) );
  FA_6001 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(B[436]), .CI(
        C[436]), .S(S[436]), .CO(C[437]) );
  FA_6000 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(B[437]), .CI(
        C[437]), .S(S[437]), .CO(C[438]) );
  FA_5999 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(B[438]), .CI(
        C[438]), .S(S[438]), .CO(C[439]) );
  FA_5998 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(B[439]), .CI(
        C[439]), .S(S[439]), .CO(C[440]) );
  FA_5997 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(B[440]), .CI(
        C[440]), .S(S[440]), .CO(C[441]) );
  FA_5996 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(B[441]), .CI(
        C[441]), .S(S[441]), .CO(C[442]) );
  FA_5995 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(B[442]), .CI(
        C[442]), .S(S[442]), .CO(C[443]) );
  FA_5994 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(B[443]), .CI(
        C[443]), .S(S[443]), .CO(C[444]) );
  FA_5993 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(B[444]), .CI(
        C[444]), .S(S[444]), .CO(C[445]) );
  FA_5992 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(B[445]), .CI(
        C[445]), .S(S[445]), .CO(C[446]) );
  FA_5991 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(B[446]), .CI(
        C[446]), .S(S[446]), .CO(C[447]) );
  FA_5990 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(B[447]), .CI(
        C[447]), .S(S[447]), .CO(C[448]) );
  FA_5989 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(B[448]), .CI(
        C[448]), .S(S[448]), .CO(C[449]) );
  FA_5988 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(B[449]), .CI(
        C[449]), .S(S[449]), .CO(C[450]) );
  FA_5987 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(B[450]), .CI(
        C[450]), .S(S[450]), .CO(C[451]) );
  FA_5986 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(B[451]), .CI(
        C[451]), .S(S[451]), .CO(C[452]) );
  FA_5985 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(B[452]), .CI(
        C[452]), .S(S[452]), .CO(C[453]) );
  FA_5984 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(B[453]), .CI(
        C[453]), .S(S[453]), .CO(C[454]) );
  FA_5983 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(B[454]), .CI(
        C[454]), .S(S[454]), .CO(C[455]) );
  FA_5982 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(B[455]), .CI(
        C[455]), .S(S[455]), .CO(C[456]) );
  FA_5981 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(B[456]), .CI(
        C[456]), .S(S[456]), .CO(C[457]) );
  FA_5980 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(B[457]), .CI(
        C[457]), .S(S[457]), .CO(C[458]) );
  FA_5979 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(B[458]), .CI(
        C[458]), .S(S[458]), .CO(C[459]) );
  FA_5978 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(B[459]), .CI(
        C[459]), .S(S[459]), .CO(C[460]) );
  FA_5977 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(B[460]), .CI(
        C[460]), .S(S[460]), .CO(C[461]) );
  FA_5976 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(B[461]), .CI(
        C[461]), .S(S[461]), .CO(C[462]) );
  FA_5975 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(B[462]), .CI(
        C[462]), .S(S[462]), .CO(C[463]) );
  FA_5974 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(B[463]), .CI(
        C[463]), .S(S[463]), .CO(C[464]) );
  FA_5973 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(B[464]), .CI(
        C[464]), .S(S[464]), .CO(C[465]) );
  FA_5972 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(B[465]), .CI(
        C[465]), .S(S[465]), .CO(C[466]) );
  FA_5971 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(B[466]), .CI(
        C[466]), .S(S[466]), .CO(C[467]) );
  FA_5970 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(B[467]), .CI(
        C[467]), .S(S[467]), .CO(C[468]) );
  FA_5969 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(B[468]), .CI(
        C[468]), .S(S[468]), .CO(C[469]) );
  FA_5968 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(B[469]), .CI(
        C[469]), .S(S[469]), .CO(C[470]) );
  FA_5967 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(B[470]), .CI(
        C[470]), .S(S[470]), .CO(C[471]) );
  FA_5966 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(B[471]), .CI(
        C[471]), .S(S[471]), .CO(C[472]) );
  FA_5965 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(B[472]), .CI(
        C[472]), .S(S[472]), .CO(C[473]) );
  FA_5964 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(B[473]), .CI(
        C[473]), .S(S[473]), .CO(C[474]) );
  FA_5963 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(B[474]), .CI(
        C[474]), .S(S[474]), .CO(C[475]) );
  FA_5962 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(B[475]), .CI(
        C[475]), .S(S[475]), .CO(C[476]) );
  FA_5961 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(B[476]), .CI(
        C[476]), .S(S[476]), .CO(C[477]) );
  FA_5960 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(B[477]), .CI(
        C[477]), .S(S[477]), .CO(C[478]) );
  FA_5959 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(B[478]), .CI(
        C[478]), .S(S[478]), .CO(C[479]) );
  FA_5958 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(B[479]), .CI(
        C[479]), .S(S[479]), .CO(C[480]) );
  FA_5957 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(B[480]), .CI(
        C[480]), .S(S[480]), .CO(C[481]) );
  FA_5956 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(B[481]), .CI(
        C[481]), .S(S[481]), .CO(C[482]) );
  FA_5955 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(B[482]), .CI(
        C[482]), .S(S[482]), .CO(C[483]) );
  FA_5954 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(B[483]), .CI(
        C[483]), .S(S[483]), .CO(C[484]) );
  FA_5953 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(B[484]), .CI(
        C[484]), .S(S[484]), .CO(C[485]) );
  FA_5952 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(B[485]), .CI(
        C[485]), .S(S[485]), .CO(C[486]) );
  FA_5951 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(B[486]), .CI(
        C[486]), .S(S[486]), .CO(C[487]) );
  FA_5950 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(B[487]), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_5949 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(B[488]), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_5948 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(B[489]), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_5947 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(B[490]), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_5946 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(B[491]), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_5945 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(B[492]), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_5944 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(B[493]), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_5943 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(B[494]), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_5942 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(B[495]), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_5941 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(B[496]), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_5940 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(B[497]), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_5939 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(B[498]), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_5938 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(B[499]), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_5937 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(B[500]), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_5936 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(B[501]), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_5935 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(B[502]), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_5934 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(B[503]), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_5933 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(B[504]), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_5932 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(B[505]), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_5931 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(B[506]), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_5930 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(B[507]), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_5929 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(B[508]), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_5928 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(B[509]), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_5927 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(B[510]), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_5926 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(B[511]), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_5925 \FA_INST_1[512].FA_  ( .A(A[512]), .B(1'b0), .CI(C[512]), .S(S[512]), 
        .CO(C[513]) );
  FA_5924 \FA_INST_1[513].FA_  ( .A(A[513]), .B(1'b0), .CI(C[513]), .S(S[513])
         );
endmodule


module FA_5410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_5411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_5412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_5923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N514_0 ( A, B, O );
  input [513:0] A;
  input [513:0] B;
  output O;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514;
  wire   [513:1] C;

  FA_5923 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n514), .CI(1'b1), 
        .CO(C[1]) );
  FA_5922 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n513), .CI(C[1]), 
        .CO(C[2]) );
  FA_5921 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n512), .CI(C[2]), 
        .CO(C[3]) );
  FA_5920 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n511), .CI(C[3]), 
        .CO(C[4]) );
  FA_5919 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n510), .CI(C[4]), 
        .CO(C[5]) );
  FA_5918 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n509), .CI(C[5]), 
        .CO(C[6]) );
  FA_5917 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n508), .CI(C[6]), 
        .CO(C[7]) );
  FA_5916 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n507), .CI(C[7]), 
        .CO(C[8]) );
  FA_5915 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n506), .CI(C[8]), 
        .CO(C[9]) );
  FA_5914 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n505), .CI(C[9]), 
        .CO(C[10]) );
  FA_5913 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n504), .CI(C[10]), 
        .CO(C[11]) );
  FA_5912 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n503), .CI(C[11]), 
        .CO(C[12]) );
  FA_5911 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n502), .CI(C[12]), 
        .CO(C[13]) );
  FA_5910 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n501), .CI(C[13]), 
        .CO(C[14]) );
  FA_5909 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n500), .CI(C[14]), 
        .CO(C[15]) );
  FA_5908 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n499), .CI(C[15]), 
        .CO(C[16]) );
  FA_5907 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n498), .CI(C[16]), 
        .CO(C[17]) );
  FA_5906 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n497), .CI(C[17]), 
        .CO(C[18]) );
  FA_5905 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n496), .CI(C[18]), 
        .CO(C[19]) );
  FA_5904 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n495), .CI(C[19]), 
        .CO(C[20]) );
  FA_5903 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n494), .CI(C[20]), 
        .CO(C[21]) );
  FA_5902 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n493), .CI(C[21]), 
        .CO(C[22]) );
  FA_5901 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n492), .CI(C[22]), 
        .CO(C[23]) );
  FA_5900 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n491), .CI(C[23]), 
        .CO(C[24]) );
  FA_5899 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n490), .CI(C[24]), 
        .CO(C[25]) );
  FA_5898 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n489), .CI(C[25]), 
        .CO(C[26]) );
  FA_5897 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n488), .CI(C[26]), 
        .CO(C[27]) );
  FA_5896 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n487), .CI(C[27]), 
        .CO(C[28]) );
  FA_5895 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n486), .CI(C[28]), 
        .CO(C[29]) );
  FA_5894 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n485), .CI(C[29]), 
        .CO(C[30]) );
  FA_5893 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n484), .CI(C[30]), 
        .CO(C[31]) );
  FA_5892 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n483), .CI(C[31]), 
        .CO(C[32]) );
  FA_5891 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n482), .CI(C[32]), 
        .CO(C[33]) );
  FA_5890 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n481), .CI(C[33]), 
        .CO(C[34]) );
  FA_5889 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n480), .CI(C[34]), 
        .CO(C[35]) );
  FA_5888 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n479), .CI(C[35]), 
        .CO(C[36]) );
  FA_5887 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n478), .CI(C[36]), 
        .CO(C[37]) );
  FA_5886 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n477), .CI(C[37]), 
        .CO(C[38]) );
  FA_5885 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n476), .CI(C[38]), 
        .CO(C[39]) );
  FA_5884 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n475), .CI(C[39]), 
        .CO(C[40]) );
  FA_5883 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n474), .CI(C[40]), 
        .CO(C[41]) );
  FA_5882 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n473), .CI(C[41]), 
        .CO(C[42]) );
  FA_5881 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n472), .CI(C[42]), 
        .CO(C[43]) );
  FA_5880 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n471), .CI(C[43]), 
        .CO(C[44]) );
  FA_5879 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n470), .CI(C[44]), 
        .CO(C[45]) );
  FA_5878 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n469), .CI(C[45]), 
        .CO(C[46]) );
  FA_5877 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n468), .CI(C[46]), 
        .CO(C[47]) );
  FA_5876 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n467), .CI(C[47]), 
        .CO(C[48]) );
  FA_5875 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n466), .CI(C[48]), 
        .CO(C[49]) );
  FA_5874 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n465), .CI(C[49]), 
        .CO(C[50]) );
  FA_5873 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n464), .CI(C[50]), 
        .CO(C[51]) );
  FA_5872 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n463), .CI(C[51]), 
        .CO(C[52]) );
  FA_5871 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n462), .CI(C[52]), 
        .CO(C[53]) );
  FA_5870 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n461), .CI(C[53]), 
        .CO(C[54]) );
  FA_5869 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n460), .CI(C[54]), 
        .CO(C[55]) );
  FA_5868 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n459), .CI(C[55]), 
        .CO(C[56]) );
  FA_5867 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n458), .CI(C[56]), 
        .CO(C[57]) );
  FA_5866 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n457), .CI(C[57]), 
        .CO(C[58]) );
  FA_5865 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n456), .CI(C[58]), 
        .CO(C[59]) );
  FA_5864 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n455), .CI(C[59]), 
        .CO(C[60]) );
  FA_5863 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n454), .CI(C[60]), 
        .CO(C[61]) );
  FA_5862 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n453), .CI(C[61]), 
        .CO(C[62]) );
  FA_5861 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n452), .CI(C[62]), 
        .CO(C[63]) );
  FA_5860 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n451), .CI(C[63]), 
        .CO(C[64]) );
  FA_5859 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n450), .CI(C[64]), 
        .CO(C[65]) );
  FA_5858 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n449), .CI(C[65]), 
        .CO(C[66]) );
  FA_5857 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n448), .CI(C[66]), 
        .CO(C[67]) );
  FA_5856 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n447), .CI(C[67]), 
        .CO(C[68]) );
  FA_5855 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n446), .CI(C[68]), 
        .CO(C[69]) );
  FA_5854 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n445), .CI(C[69]), 
        .CO(C[70]) );
  FA_5853 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n444), .CI(C[70]), 
        .CO(C[71]) );
  FA_5852 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n443), .CI(C[71]), 
        .CO(C[72]) );
  FA_5851 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n442), .CI(C[72]), 
        .CO(C[73]) );
  FA_5850 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n441), .CI(C[73]), 
        .CO(C[74]) );
  FA_5849 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n440), .CI(C[74]), 
        .CO(C[75]) );
  FA_5848 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n439), .CI(C[75]), 
        .CO(C[76]) );
  FA_5847 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n438), .CI(C[76]), 
        .CO(C[77]) );
  FA_5846 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n437), .CI(C[77]), 
        .CO(C[78]) );
  FA_5845 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n436), .CI(C[78]), 
        .CO(C[79]) );
  FA_5844 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n435), .CI(C[79]), 
        .CO(C[80]) );
  FA_5843 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n434), .CI(C[80]), 
        .CO(C[81]) );
  FA_5842 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n433), .CI(C[81]), 
        .CO(C[82]) );
  FA_5841 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n432), .CI(C[82]), 
        .CO(C[83]) );
  FA_5840 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n431), .CI(C[83]), 
        .CO(C[84]) );
  FA_5839 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n430), .CI(C[84]), 
        .CO(C[85]) );
  FA_5838 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n429), .CI(C[85]), 
        .CO(C[86]) );
  FA_5837 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n428), .CI(C[86]), 
        .CO(C[87]) );
  FA_5836 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n427), .CI(C[87]), 
        .CO(C[88]) );
  FA_5835 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n426), .CI(C[88]), 
        .CO(C[89]) );
  FA_5834 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n425), .CI(C[89]), 
        .CO(C[90]) );
  FA_5833 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n424), .CI(C[90]), 
        .CO(C[91]) );
  FA_5832 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n423), .CI(C[91]), 
        .CO(C[92]) );
  FA_5831 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n422), .CI(C[92]), 
        .CO(C[93]) );
  FA_5830 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n421), .CI(C[93]), 
        .CO(C[94]) );
  FA_5829 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n420), .CI(C[94]), 
        .CO(C[95]) );
  FA_5828 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n419), .CI(C[95]), 
        .CO(C[96]) );
  FA_5827 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n418), .CI(C[96]), 
        .CO(C[97]) );
  FA_5826 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n417), .CI(C[97]), 
        .CO(C[98]) );
  FA_5825 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n416), .CI(C[98]), 
        .CO(C[99]) );
  FA_5824 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n415), .CI(C[99]), 
        .CO(C[100]) );
  FA_5823 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n414), .CI(C[100]), .CO(C[101]) );
  FA_5822 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n413), .CI(C[101]), .CO(C[102]) );
  FA_5821 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n412), .CI(C[102]), .CO(C[103]) );
  FA_5820 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n411), .CI(C[103]), .CO(C[104]) );
  FA_5819 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n410), .CI(C[104]), .CO(C[105]) );
  FA_5818 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n409), .CI(C[105]), .CO(C[106]) );
  FA_5817 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n408), .CI(C[106]), .CO(C[107]) );
  FA_5816 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n407), .CI(C[107]), .CO(C[108]) );
  FA_5815 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n406), .CI(C[108]), .CO(C[109]) );
  FA_5814 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n405), .CI(C[109]), .CO(C[110]) );
  FA_5813 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n404), .CI(C[110]), .CO(C[111]) );
  FA_5812 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n403), .CI(C[111]), .CO(C[112]) );
  FA_5811 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n402), .CI(C[112]), .CO(C[113]) );
  FA_5810 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n401), .CI(C[113]), .CO(C[114]) );
  FA_5809 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n400), .CI(C[114]), .CO(C[115]) );
  FA_5808 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n399), .CI(C[115]), .CO(C[116]) );
  FA_5807 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n398), .CI(C[116]), .CO(C[117]) );
  FA_5806 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n397), .CI(C[117]), .CO(C[118]) );
  FA_5805 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n396), .CI(C[118]), .CO(C[119]) );
  FA_5804 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n395), .CI(C[119]), .CO(C[120]) );
  FA_5803 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n394), .CI(C[120]), .CO(C[121]) );
  FA_5802 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n393), .CI(C[121]), .CO(C[122]) );
  FA_5801 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n392), .CI(C[122]), .CO(C[123]) );
  FA_5800 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n391), .CI(C[123]), .CO(C[124]) );
  FA_5799 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n390), .CI(C[124]), .CO(C[125]) );
  FA_5798 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n389), .CI(C[125]), .CO(C[126]) );
  FA_5797 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n388), .CI(C[126]), .CO(C[127]) );
  FA_5796 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n387), .CI(C[127]), .CO(C[128]) );
  FA_5795 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n386), .CI(C[128]), .CO(C[129]) );
  FA_5794 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n385), .CI(C[129]), .CO(C[130]) );
  FA_5793 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n384), .CI(C[130]), .CO(C[131]) );
  FA_5792 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n383), .CI(C[131]), .CO(C[132]) );
  FA_5791 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n382), .CI(C[132]), .CO(C[133]) );
  FA_5790 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n381), .CI(C[133]), .CO(C[134]) );
  FA_5789 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n380), .CI(C[134]), .CO(C[135]) );
  FA_5788 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n379), .CI(C[135]), .CO(C[136]) );
  FA_5787 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n378), .CI(C[136]), .CO(C[137]) );
  FA_5786 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n377), .CI(C[137]), .CO(C[138]) );
  FA_5785 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n376), .CI(C[138]), .CO(C[139]) );
  FA_5784 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n375), .CI(C[139]), .CO(C[140]) );
  FA_5783 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n374), .CI(C[140]), .CO(C[141]) );
  FA_5782 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n373), .CI(C[141]), .CO(C[142]) );
  FA_5781 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n372), .CI(C[142]), .CO(C[143]) );
  FA_5780 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n371), .CI(C[143]), .CO(C[144]) );
  FA_5779 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n370), .CI(C[144]), .CO(C[145]) );
  FA_5778 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n369), .CI(C[145]), .CO(C[146]) );
  FA_5777 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n368), .CI(C[146]), .CO(C[147]) );
  FA_5776 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n367), .CI(C[147]), .CO(C[148]) );
  FA_5775 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n366), .CI(C[148]), .CO(C[149]) );
  FA_5774 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n365), .CI(C[149]), .CO(C[150]) );
  FA_5773 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n364), .CI(C[150]), .CO(C[151]) );
  FA_5772 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n363), .CI(C[151]), .CO(C[152]) );
  FA_5771 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n362), .CI(C[152]), .CO(C[153]) );
  FA_5770 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n361), .CI(C[153]), .CO(C[154]) );
  FA_5769 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n360), .CI(C[154]), .CO(C[155]) );
  FA_5768 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n359), .CI(C[155]), .CO(C[156]) );
  FA_5767 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n358), .CI(C[156]), .CO(C[157]) );
  FA_5766 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n357), .CI(C[157]), .CO(C[158]) );
  FA_5765 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n356), .CI(C[158]), .CO(C[159]) );
  FA_5764 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n355), .CI(C[159]), .CO(C[160]) );
  FA_5763 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n354), .CI(C[160]), .CO(C[161]) );
  FA_5762 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n353), .CI(C[161]), .CO(C[162]) );
  FA_5761 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n352), .CI(C[162]), .CO(C[163]) );
  FA_5760 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n351), .CI(C[163]), .CO(C[164]) );
  FA_5759 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n350), .CI(C[164]), .CO(C[165]) );
  FA_5758 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n349), .CI(C[165]), .CO(C[166]) );
  FA_5757 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n348), .CI(C[166]), .CO(C[167]) );
  FA_5756 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n347), .CI(C[167]), .CO(C[168]) );
  FA_5755 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n346), .CI(C[168]), .CO(C[169]) );
  FA_5754 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n345), .CI(C[169]), .CO(C[170]) );
  FA_5753 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n344), .CI(C[170]), .CO(C[171]) );
  FA_5752 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n343), .CI(C[171]), .CO(C[172]) );
  FA_5751 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n342), .CI(C[172]), .CO(C[173]) );
  FA_5750 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n341), .CI(C[173]), .CO(C[174]) );
  FA_5749 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n340), .CI(C[174]), .CO(C[175]) );
  FA_5748 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n339), .CI(C[175]), .CO(C[176]) );
  FA_5747 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n338), .CI(C[176]), .CO(C[177]) );
  FA_5746 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n337), .CI(C[177]), .CO(C[178]) );
  FA_5745 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n336), .CI(C[178]), .CO(C[179]) );
  FA_5744 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n335), .CI(C[179]), .CO(C[180]) );
  FA_5743 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n334), .CI(C[180]), .CO(C[181]) );
  FA_5742 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n333), .CI(C[181]), .CO(C[182]) );
  FA_5741 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n332), .CI(C[182]), .CO(C[183]) );
  FA_5740 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n331), .CI(C[183]), .CO(C[184]) );
  FA_5739 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n330), .CI(C[184]), .CO(C[185]) );
  FA_5738 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n329), .CI(C[185]), .CO(C[186]) );
  FA_5737 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n328), .CI(C[186]), .CO(C[187]) );
  FA_5736 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n327), .CI(C[187]), .CO(C[188]) );
  FA_5735 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n326), .CI(C[188]), .CO(C[189]) );
  FA_5734 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n325), .CI(C[189]), .CO(C[190]) );
  FA_5733 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n324), .CI(C[190]), .CO(C[191]) );
  FA_5732 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n323), .CI(C[191]), .CO(C[192]) );
  FA_5731 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n322), .CI(C[192]), .CO(C[193]) );
  FA_5730 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n321), .CI(C[193]), .CO(C[194]) );
  FA_5729 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n320), .CI(C[194]), .CO(C[195]) );
  FA_5728 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n319), .CI(C[195]), .CO(C[196]) );
  FA_5727 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n318), .CI(C[196]), .CO(C[197]) );
  FA_5726 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n317), .CI(C[197]), .CO(C[198]) );
  FA_5725 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n316), .CI(C[198]), .CO(C[199]) );
  FA_5724 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n315), .CI(C[199]), .CO(C[200]) );
  FA_5723 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n314), .CI(C[200]), .CO(C[201]) );
  FA_5722 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n313), .CI(C[201]), .CO(C[202]) );
  FA_5721 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n312), .CI(C[202]), .CO(C[203]) );
  FA_5720 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n311), .CI(C[203]), .CO(C[204]) );
  FA_5719 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n310), .CI(C[204]), .CO(C[205]) );
  FA_5718 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n309), .CI(C[205]), .CO(C[206]) );
  FA_5717 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n308), .CI(C[206]), .CO(C[207]) );
  FA_5716 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n307), .CI(C[207]), .CO(C[208]) );
  FA_5715 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n306), .CI(C[208]), .CO(C[209]) );
  FA_5714 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n305), .CI(C[209]), .CO(C[210]) );
  FA_5713 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n304), .CI(C[210]), .CO(C[211]) );
  FA_5712 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n303), .CI(C[211]), .CO(C[212]) );
  FA_5711 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n302), .CI(C[212]), .CO(C[213]) );
  FA_5710 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n301), .CI(C[213]), .CO(C[214]) );
  FA_5709 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n300), .CI(C[214]), .CO(C[215]) );
  FA_5708 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n299), .CI(C[215]), .CO(C[216]) );
  FA_5707 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n298), .CI(C[216]), .CO(C[217]) );
  FA_5706 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n297), .CI(C[217]), .CO(C[218]) );
  FA_5705 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n296), .CI(C[218]), .CO(C[219]) );
  FA_5704 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n295), .CI(C[219]), .CO(C[220]) );
  FA_5703 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n294), .CI(C[220]), .CO(C[221]) );
  FA_5702 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n293), .CI(C[221]), .CO(C[222]) );
  FA_5701 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n292), .CI(C[222]), .CO(C[223]) );
  FA_5700 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n291), .CI(C[223]), .CO(C[224]) );
  FA_5699 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n290), .CI(C[224]), .CO(C[225]) );
  FA_5698 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n289), .CI(C[225]), .CO(C[226]) );
  FA_5697 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n288), .CI(C[226]), .CO(C[227]) );
  FA_5696 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n287), .CI(C[227]), .CO(C[228]) );
  FA_5695 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n286), .CI(C[228]), .CO(C[229]) );
  FA_5694 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n285), .CI(C[229]), .CO(C[230]) );
  FA_5693 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n284), .CI(C[230]), .CO(C[231]) );
  FA_5692 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n283), .CI(C[231]), .CO(C[232]) );
  FA_5691 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n282), .CI(C[232]), .CO(C[233]) );
  FA_5690 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n281), .CI(C[233]), .CO(C[234]) );
  FA_5689 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n280), .CI(C[234]), .CO(C[235]) );
  FA_5688 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n279), .CI(C[235]), .CO(C[236]) );
  FA_5687 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n278), .CI(C[236]), .CO(C[237]) );
  FA_5686 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n277), .CI(C[237]), .CO(C[238]) );
  FA_5685 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n276), .CI(C[238]), .CO(C[239]) );
  FA_5684 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n275), .CI(C[239]), .CO(C[240]) );
  FA_5683 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n274), .CI(C[240]), .CO(C[241]) );
  FA_5682 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n273), .CI(C[241]), .CO(C[242]) );
  FA_5681 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n272), .CI(C[242]), .CO(C[243]) );
  FA_5680 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n271), .CI(C[243]), .CO(C[244]) );
  FA_5679 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n270), .CI(C[244]), .CO(C[245]) );
  FA_5678 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n269), .CI(C[245]), .CO(C[246]) );
  FA_5677 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n268), .CI(C[246]), .CO(C[247]) );
  FA_5676 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n267), .CI(C[247]), .CO(C[248]) );
  FA_5675 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n266), .CI(C[248]), .CO(C[249]) );
  FA_5674 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n265), .CI(C[249]), .CO(C[250]) );
  FA_5673 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n264), .CI(C[250]), .CO(C[251]) );
  FA_5672 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n263), .CI(C[251]), .CO(C[252]) );
  FA_5671 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n262), .CI(C[252]), .CO(C[253]) );
  FA_5670 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n261), .CI(C[253]), .CO(C[254]) );
  FA_5669 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n260), .CI(C[254]), .CO(C[255]) );
  FA_5668 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n259), .CI(C[255]), .CO(C[256]) );
  FA_5667 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n258), .CI(C[256]), .CO(C[257]) );
  FA_5666 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n257), .CI(C[257]), .CO(C[258]) );
  FA_5665 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n256), .CI(C[258]), .CO(C[259]) );
  FA_5664 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n255), .CI(C[259]), .CO(C[260]) );
  FA_5663 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n254), .CI(C[260]), .CO(C[261]) );
  FA_5662 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n253), .CI(C[261]), .CO(C[262]) );
  FA_5661 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n252), .CI(C[262]), .CO(C[263]) );
  FA_5660 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n251), .CI(C[263]), .CO(C[264]) );
  FA_5659 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n250), .CI(C[264]), .CO(C[265]) );
  FA_5658 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n249), .CI(C[265]), .CO(C[266]) );
  FA_5657 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n248), .CI(C[266]), .CO(C[267]) );
  FA_5656 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n247), .CI(C[267]), .CO(C[268]) );
  FA_5655 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n246), .CI(C[268]), .CO(C[269]) );
  FA_5654 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n245), .CI(C[269]), .CO(C[270]) );
  FA_5653 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n244), .CI(C[270]), .CO(C[271]) );
  FA_5652 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n243), .CI(C[271]), .CO(C[272]) );
  FA_5651 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n242), .CI(C[272]), .CO(C[273]) );
  FA_5650 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n241), .CI(C[273]), .CO(C[274]) );
  FA_5649 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n240), .CI(C[274]), .CO(C[275]) );
  FA_5648 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n239), .CI(C[275]), .CO(C[276]) );
  FA_5647 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n238), .CI(C[276]), .CO(C[277]) );
  FA_5646 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n237), .CI(C[277]), .CO(C[278]) );
  FA_5645 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n236), .CI(C[278]), .CO(C[279]) );
  FA_5644 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n235), .CI(C[279]), .CO(C[280]) );
  FA_5643 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n234), .CI(C[280]), .CO(C[281]) );
  FA_5642 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n233), .CI(C[281]), .CO(C[282]) );
  FA_5641 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n232), .CI(C[282]), .CO(C[283]) );
  FA_5640 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n231), .CI(C[283]), .CO(C[284]) );
  FA_5639 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n230), .CI(C[284]), .CO(C[285]) );
  FA_5638 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n229), .CI(C[285]), .CO(C[286]) );
  FA_5637 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n228), .CI(C[286]), .CO(C[287]) );
  FA_5636 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n227), .CI(C[287]), .CO(C[288]) );
  FA_5635 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n226), .CI(C[288]), .CO(C[289]) );
  FA_5634 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n225), .CI(C[289]), .CO(C[290]) );
  FA_5633 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n224), .CI(C[290]), .CO(C[291]) );
  FA_5632 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n223), .CI(C[291]), .CO(C[292]) );
  FA_5631 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n222), .CI(C[292]), .CO(C[293]) );
  FA_5630 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n221), .CI(C[293]), .CO(C[294]) );
  FA_5629 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n220), .CI(C[294]), .CO(C[295]) );
  FA_5628 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n219), .CI(C[295]), .CO(C[296]) );
  FA_5627 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n218), .CI(C[296]), .CO(C[297]) );
  FA_5626 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n217), .CI(C[297]), .CO(C[298]) );
  FA_5625 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n216), .CI(C[298]), .CO(C[299]) );
  FA_5624 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n215), .CI(C[299]), .CO(C[300]) );
  FA_5623 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n214), .CI(C[300]), .CO(C[301]) );
  FA_5622 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n213), .CI(C[301]), .CO(C[302]) );
  FA_5621 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n212), .CI(C[302]), .CO(C[303]) );
  FA_5620 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n211), .CI(C[303]), .CO(C[304]) );
  FA_5619 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n210), .CI(C[304]), .CO(C[305]) );
  FA_5618 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n209), .CI(C[305]), .CO(C[306]) );
  FA_5617 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n208), .CI(C[306]), .CO(C[307]) );
  FA_5616 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n207), .CI(C[307]), .CO(C[308]) );
  FA_5615 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n206), .CI(C[308]), .CO(C[309]) );
  FA_5614 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n205), .CI(C[309]), .CO(C[310]) );
  FA_5613 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n204), .CI(C[310]), .CO(C[311]) );
  FA_5612 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n203), .CI(C[311]), .CO(C[312]) );
  FA_5611 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n202), .CI(C[312]), .CO(C[313]) );
  FA_5610 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n201), .CI(C[313]), .CO(C[314]) );
  FA_5609 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n200), .CI(C[314]), .CO(C[315]) );
  FA_5608 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n199), .CI(C[315]), .CO(C[316]) );
  FA_5607 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n198), .CI(C[316]), .CO(C[317]) );
  FA_5606 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n197), .CI(C[317]), .CO(C[318]) );
  FA_5605 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n196), .CI(C[318]), .CO(C[319]) );
  FA_5604 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n195), .CI(C[319]), .CO(C[320]) );
  FA_5603 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n194), .CI(C[320]), .CO(C[321]) );
  FA_5602 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n193), .CI(C[321]), .CO(C[322]) );
  FA_5601 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n192), .CI(C[322]), .CO(C[323]) );
  FA_5600 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n191), .CI(C[323]), .CO(C[324]) );
  FA_5599 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n190), .CI(C[324]), .CO(C[325]) );
  FA_5598 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n189), .CI(C[325]), .CO(C[326]) );
  FA_5597 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n188), .CI(C[326]), .CO(C[327]) );
  FA_5596 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n187), .CI(C[327]), .CO(C[328]) );
  FA_5595 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n186), .CI(C[328]), .CO(C[329]) );
  FA_5594 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n185), .CI(C[329]), .CO(C[330]) );
  FA_5593 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n184), .CI(C[330]), .CO(C[331]) );
  FA_5592 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n183), .CI(C[331]), .CO(C[332]) );
  FA_5591 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n182), .CI(C[332]), .CO(C[333]) );
  FA_5590 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n181), .CI(C[333]), .CO(C[334]) );
  FA_5589 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n180), .CI(C[334]), .CO(C[335]) );
  FA_5588 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n179), .CI(C[335]), .CO(C[336]) );
  FA_5587 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n178), .CI(C[336]), .CO(C[337]) );
  FA_5586 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n177), .CI(C[337]), .CO(C[338]) );
  FA_5585 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n176), .CI(C[338]), .CO(C[339]) );
  FA_5584 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n175), .CI(C[339]), .CO(C[340]) );
  FA_5583 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n174), .CI(C[340]), .CO(C[341]) );
  FA_5582 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n173), .CI(C[341]), .CO(C[342]) );
  FA_5581 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n172), .CI(C[342]), .CO(C[343]) );
  FA_5580 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n171), .CI(C[343]), .CO(C[344]) );
  FA_5579 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n170), .CI(C[344]), .CO(C[345]) );
  FA_5578 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n169), .CI(C[345]), .CO(C[346]) );
  FA_5577 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n168), .CI(C[346]), .CO(C[347]) );
  FA_5576 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n167), .CI(C[347]), .CO(C[348]) );
  FA_5575 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n166), .CI(C[348]), .CO(C[349]) );
  FA_5574 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n165), .CI(C[349]), .CO(C[350]) );
  FA_5573 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n164), .CI(C[350]), .CO(C[351]) );
  FA_5572 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n163), .CI(C[351]), .CO(C[352]) );
  FA_5571 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n162), .CI(C[352]), .CO(C[353]) );
  FA_5570 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n161), .CI(C[353]), .CO(C[354]) );
  FA_5569 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n160), .CI(C[354]), .CO(C[355]) );
  FA_5568 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n159), .CI(C[355]), .CO(C[356]) );
  FA_5567 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n158), .CI(C[356]), .CO(C[357]) );
  FA_5566 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n157), .CI(C[357]), .CO(C[358]) );
  FA_5565 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n156), .CI(C[358]), .CO(C[359]) );
  FA_5564 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n155), .CI(C[359]), .CO(C[360]) );
  FA_5563 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n154), .CI(C[360]), .CO(C[361]) );
  FA_5562 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n153), .CI(C[361]), .CO(C[362]) );
  FA_5561 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n152), .CI(C[362]), .CO(C[363]) );
  FA_5560 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n151), .CI(C[363]), .CO(C[364]) );
  FA_5559 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n150), .CI(C[364]), .CO(C[365]) );
  FA_5558 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n149), .CI(C[365]), .CO(C[366]) );
  FA_5557 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n148), .CI(C[366]), .CO(C[367]) );
  FA_5556 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n147), .CI(C[367]), .CO(C[368]) );
  FA_5555 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n146), .CI(C[368]), .CO(C[369]) );
  FA_5554 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n145), .CI(C[369]), .CO(C[370]) );
  FA_5553 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n144), .CI(C[370]), .CO(C[371]) );
  FA_5552 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n143), .CI(C[371]), .CO(C[372]) );
  FA_5551 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n142), .CI(C[372]), .CO(C[373]) );
  FA_5550 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n141), .CI(C[373]), .CO(C[374]) );
  FA_5549 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n140), .CI(C[374]), .CO(C[375]) );
  FA_5548 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n139), .CI(C[375]), .CO(C[376]) );
  FA_5547 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n138), .CI(C[376]), .CO(C[377]) );
  FA_5546 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n137), .CI(C[377]), .CO(C[378]) );
  FA_5545 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n136), .CI(C[378]), .CO(C[379]) );
  FA_5544 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n135), .CI(C[379]), .CO(C[380]) );
  FA_5543 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n134), .CI(C[380]), .CO(C[381]) );
  FA_5542 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n133), .CI(C[381]), .CO(C[382]) );
  FA_5541 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n132), .CI(C[382]), .CO(C[383]) );
  FA_5540 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n131), .CI(C[383]), .CO(C[384]) );
  FA_5539 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n130), .CI(C[384]), .CO(C[385]) );
  FA_5538 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n129), .CI(C[385]), .CO(C[386]) );
  FA_5537 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n128), .CI(C[386]), .CO(C[387]) );
  FA_5536 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n127), .CI(C[387]), .CO(C[388]) );
  FA_5535 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n126), .CI(C[388]), .CO(C[389]) );
  FA_5534 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n125), .CI(C[389]), .CO(C[390]) );
  FA_5533 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n124), .CI(C[390]), .CO(C[391]) );
  FA_5532 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n123), .CI(C[391]), .CO(C[392]) );
  FA_5531 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n122), .CI(C[392]), .CO(C[393]) );
  FA_5530 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n121), .CI(C[393]), .CO(C[394]) );
  FA_5529 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n120), .CI(C[394]), .CO(C[395]) );
  FA_5528 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n119), .CI(C[395]), .CO(C[396]) );
  FA_5527 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n118), .CI(C[396]), .CO(C[397]) );
  FA_5526 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n117), .CI(C[397]), .CO(C[398]) );
  FA_5525 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n116), .CI(C[398]), .CO(C[399]) );
  FA_5524 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n115), .CI(C[399]), .CO(C[400]) );
  FA_5523 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n114), .CI(C[400]), .CO(C[401]) );
  FA_5522 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n113), .CI(C[401]), .CO(C[402]) );
  FA_5521 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n112), .CI(C[402]), .CO(C[403]) );
  FA_5520 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n111), .CI(C[403]), .CO(C[404]) );
  FA_5519 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n110), .CI(C[404]), .CO(C[405]) );
  FA_5518 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n109), .CI(C[405]), .CO(C[406]) );
  FA_5517 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n108), .CI(C[406]), .CO(C[407]) );
  FA_5516 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n107), .CI(C[407]), .CO(C[408]) );
  FA_5515 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n106), .CI(C[408]), .CO(C[409]) );
  FA_5514 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n105), .CI(C[409]), .CO(C[410]) );
  FA_5513 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n104), .CI(C[410]), .CO(C[411]) );
  FA_5512 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n103), .CI(C[411]), .CO(C[412]) );
  FA_5511 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n102), .CI(C[412]), .CO(C[413]) );
  FA_5510 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n101), .CI(C[413]), .CO(C[414]) );
  FA_5509 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n100), .CI(C[414]), .CO(C[415]) );
  FA_5508 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n99), .CI(C[415]), 
        .CO(C[416]) );
  FA_5507 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n98), .CI(C[416]), 
        .CO(C[417]) );
  FA_5506 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n97), .CI(C[417]), 
        .CO(C[418]) );
  FA_5505 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n96), .CI(C[418]), 
        .CO(C[419]) );
  FA_5504 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n95), .CI(C[419]), 
        .CO(C[420]) );
  FA_5503 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n94), .CI(C[420]), 
        .CO(C[421]) );
  FA_5502 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n93), .CI(C[421]), 
        .CO(C[422]) );
  FA_5501 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n92), .CI(C[422]), 
        .CO(C[423]) );
  FA_5500 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n91), .CI(C[423]), 
        .CO(C[424]) );
  FA_5499 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n90), .CI(C[424]), 
        .CO(C[425]) );
  FA_5498 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n89), .CI(C[425]), 
        .CO(C[426]) );
  FA_5497 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n88), .CI(C[426]), 
        .CO(C[427]) );
  FA_5496 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n87), .CI(C[427]), 
        .CO(C[428]) );
  FA_5495 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n86), .CI(C[428]), 
        .CO(C[429]) );
  FA_5494 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n85), .CI(C[429]), 
        .CO(C[430]) );
  FA_5493 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n84), .CI(C[430]), 
        .CO(C[431]) );
  FA_5492 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n83), .CI(C[431]), 
        .CO(C[432]) );
  FA_5491 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n82), .CI(C[432]), 
        .CO(C[433]) );
  FA_5490 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n81), .CI(C[433]), 
        .CO(C[434]) );
  FA_5489 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n80), .CI(C[434]), 
        .CO(C[435]) );
  FA_5488 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n79), .CI(C[435]), 
        .CO(C[436]) );
  FA_5487 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n78), .CI(C[436]), 
        .CO(C[437]) );
  FA_5486 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n77), .CI(C[437]), 
        .CO(C[438]) );
  FA_5485 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n76), .CI(C[438]), 
        .CO(C[439]) );
  FA_5484 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n75), .CI(C[439]), 
        .CO(C[440]) );
  FA_5483 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n74), .CI(C[440]), 
        .CO(C[441]) );
  FA_5482 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n73), .CI(C[441]), 
        .CO(C[442]) );
  FA_5481 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n72), .CI(C[442]), 
        .CO(C[443]) );
  FA_5480 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n71), .CI(C[443]), 
        .CO(C[444]) );
  FA_5479 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n70), .CI(C[444]), 
        .CO(C[445]) );
  FA_5478 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n69), .CI(C[445]), 
        .CO(C[446]) );
  FA_5477 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n68), .CI(C[446]), 
        .CO(C[447]) );
  FA_5476 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n67), .CI(C[447]), 
        .CO(C[448]) );
  FA_5475 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n66), .CI(C[448]), 
        .CO(C[449]) );
  FA_5474 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n65), .CI(C[449]), 
        .CO(C[450]) );
  FA_5473 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n64), .CI(C[450]), 
        .CO(C[451]) );
  FA_5472 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n63), .CI(C[451]), 
        .CO(C[452]) );
  FA_5471 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n62), .CI(C[452]), 
        .CO(C[453]) );
  FA_5470 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n61), .CI(C[453]), 
        .CO(C[454]) );
  FA_5469 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n60), .CI(C[454]), 
        .CO(C[455]) );
  FA_5468 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n59), .CI(C[455]), 
        .CO(C[456]) );
  FA_5467 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n58), .CI(C[456]), 
        .CO(C[457]) );
  FA_5466 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n57), .CI(C[457]), 
        .CO(C[458]) );
  FA_5465 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n56), .CI(C[458]), 
        .CO(C[459]) );
  FA_5464 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n55), .CI(C[459]), 
        .CO(C[460]) );
  FA_5463 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n54), .CI(C[460]), 
        .CO(C[461]) );
  FA_5462 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n53), .CI(C[461]), 
        .CO(C[462]) );
  FA_5461 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n52), .CI(C[462]), 
        .CO(C[463]) );
  FA_5460 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n51), .CI(C[463]), 
        .CO(C[464]) );
  FA_5459 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n50), .CI(C[464]), 
        .CO(C[465]) );
  FA_5458 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n49), .CI(C[465]), 
        .CO(C[466]) );
  FA_5457 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n48), .CI(C[466]), 
        .CO(C[467]) );
  FA_5456 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n47), .CI(C[467]), 
        .CO(C[468]) );
  FA_5455 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n46), .CI(C[468]), 
        .CO(C[469]) );
  FA_5454 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n45), .CI(C[469]), 
        .CO(C[470]) );
  FA_5453 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n44), .CI(C[470]), 
        .CO(C[471]) );
  FA_5452 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n43), .CI(C[471]), 
        .CO(C[472]) );
  FA_5451 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n42), .CI(C[472]), 
        .CO(C[473]) );
  FA_5450 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n41), .CI(C[473]), 
        .CO(C[474]) );
  FA_5449 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n40), .CI(C[474]), 
        .CO(C[475]) );
  FA_5448 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n39), .CI(C[475]), 
        .CO(C[476]) );
  FA_5447 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n38), .CI(C[476]), 
        .CO(C[477]) );
  FA_5446 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n37), .CI(C[477]), 
        .CO(C[478]) );
  FA_5445 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n36), .CI(C[478]), 
        .CO(C[479]) );
  FA_5444 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n35), .CI(C[479]), 
        .CO(C[480]) );
  FA_5443 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n34), .CI(C[480]), 
        .CO(C[481]) );
  FA_5442 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n33), .CI(C[481]), 
        .CO(C[482]) );
  FA_5441 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n32), .CI(C[482]), 
        .CO(C[483]) );
  FA_5440 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n31), .CI(C[483]), 
        .CO(C[484]) );
  FA_5439 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n30), .CI(C[484]), 
        .CO(C[485]) );
  FA_5438 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n29), .CI(C[485]), 
        .CO(C[486]) );
  FA_5437 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n28), .CI(C[486]), 
        .CO(C[487]) );
  FA_5436 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n27), .CI(C[487]), 
        .CO(C[488]) );
  FA_5435 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n26), .CI(C[488]), 
        .CO(C[489]) );
  FA_5434 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n25), .CI(C[489]), 
        .CO(C[490]) );
  FA_5433 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n24), .CI(C[490]), 
        .CO(C[491]) );
  FA_5432 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n23), .CI(C[491]), 
        .CO(C[492]) );
  FA_5431 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n22), .CI(C[492]), 
        .CO(C[493]) );
  FA_5430 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n21), .CI(C[493]), 
        .CO(C[494]) );
  FA_5429 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n20), .CI(C[494]), 
        .CO(C[495]) );
  FA_5428 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n19), .CI(C[495]), 
        .CO(C[496]) );
  FA_5427 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n18), .CI(C[496]), 
        .CO(C[497]) );
  FA_5426 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n17), .CI(C[497]), 
        .CO(C[498]) );
  FA_5425 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n16), .CI(C[498]), 
        .CO(C[499]) );
  FA_5424 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n15), .CI(C[499]), 
        .CO(C[500]) );
  FA_5423 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n14), .CI(C[500]), 
        .CO(C[501]) );
  FA_5422 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n13), .CI(C[501]), 
        .CO(C[502]) );
  FA_5421 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n12), .CI(C[502]), 
        .CO(C[503]) );
  FA_5420 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n11), .CI(C[503]), 
        .CO(C[504]) );
  FA_5419 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n10), .CI(C[504]), 
        .CO(C[505]) );
  FA_5418 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n9), .CI(C[505]), 
        .CO(C[506]) );
  FA_5417 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n8), .CI(C[506]), 
        .CO(C[507]) );
  FA_5416 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n7), .CI(C[507]), 
        .CO(C[508]) );
  FA_5415 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n6), .CI(C[508]), 
        .CO(C[509]) );
  FA_5414 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n5), .CI(C[509]), 
        .CO(C[510]) );
  FA_5413 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n4), .CI(C[510]), 
        .CO(C[511]) );
  FA_5412 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n3), .CI(C[511]), 
        .CO(C[512]) );
  FA_5411 \FA_INST_1[512].FA_  ( .A(A[512]), .B(1'b1), .CI(C[512]), .CO(C[513]) );
  FA_5410 \FA_INST_1[513].FA_  ( .A(A[513]), .B(1'b1), .CI(C[513]), .CO(O) );
  IV U2 ( .A(B[415]), .Z(n99) );
  IV U3 ( .A(B[416]), .Z(n98) );
  IV U4 ( .A(B[417]), .Z(n97) );
  IV U5 ( .A(B[418]), .Z(n96) );
  IV U6 ( .A(B[419]), .Z(n95) );
  IV U7 ( .A(B[420]), .Z(n94) );
  IV U8 ( .A(B[421]), .Z(n93) );
  IV U9 ( .A(B[422]), .Z(n92) );
  IV U10 ( .A(B[423]), .Z(n91) );
  IV U11 ( .A(B[424]), .Z(n90) );
  IV U12 ( .A(B[505]), .Z(n9) );
  IV U13 ( .A(B[425]), .Z(n89) );
  IV U14 ( .A(B[426]), .Z(n88) );
  IV U15 ( .A(B[427]), .Z(n87) );
  IV U16 ( .A(B[428]), .Z(n86) );
  IV U17 ( .A(B[429]), .Z(n85) );
  IV U18 ( .A(B[430]), .Z(n84) );
  IV U19 ( .A(B[431]), .Z(n83) );
  IV U20 ( .A(B[432]), .Z(n82) );
  IV U21 ( .A(B[433]), .Z(n81) );
  IV U22 ( .A(B[434]), .Z(n80) );
  IV U23 ( .A(B[506]), .Z(n8) );
  IV U24 ( .A(B[435]), .Z(n79) );
  IV U25 ( .A(B[436]), .Z(n78) );
  IV U26 ( .A(B[437]), .Z(n77) );
  IV U27 ( .A(B[438]), .Z(n76) );
  IV U28 ( .A(B[439]), .Z(n75) );
  IV U29 ( .A(B[440]), .Z(n74) );
  IV U30 ( .A(B[441]), .Z(n73) );
  IV U31 ( .A(B[442]), .Z(n72) );
  IV U32 ( .A(B[443]), .Z(n71) );
  IV U33 ( .A(B[444]), .Z(n70) );
  IV U34 ( .A(B[507]), .Z(n7) );
  IV U35 ( .A(B[445]), .Z(n69) );
  IV U36 ( .A(B[446]), .Z(n68) );
  IV U37 ( .A(B[447]), .Z(n67) );
  IV U38 ( .A(B[448]), .Z(n66) );
  IV U39 ( .A(B[449]), .Z(n65) );
  IV U40 ( .A(B[450]), .Z(n64) );
  IV U41 ( .A(B[451]), .Z(n63) );
  IV U42 ( .A(B[452]), .Z(n62) );
  IV U43 ( .A(B[453]), .Z(n61) );
  IV U44 ( .A(B[454]), .Z(n60) );
  IV U45 ( .A(B[508]), .Z(n6) );
  IV U46 ( .A(B[455]), .Z(n59) );
  IV U47 ( .A(B[456]), .Z(n58) );
  IV U48 ( .A(B[457]), .Z(n57) );
  IV U49 ( .A(B[458]), .Z(n56) );
  IV U50 ( .A(B[459]), .Z(n55) );
  IV U51 ( .A(B[460]), .Z(n54) );
  IV U52 ( .A(B[461]), .Z(n53) );
  IV U53 ( .A(B[462]), .Z(n52) );
  IV U54 ( .A(B[0]), .Z(n514) );
  IV U55 ( .A(B[1]), .Z(n513) );
  IV U56 ( .A(B[2]), .Z(n512) );
  IV U57 ( .A(B[3]), .Z(n511) );
  IV U58 ( .A(B[4]), .Z(n510) );
  IV U59 ( .A(B[463]), .Z(n51) );
  IV U60 ( .A(B[5]), .Z(n509) );
  IV U61 ( .A(B[6]), .Z(n508) );
  IV U62 ( .A(B[7]), .Z(n507) );
  IV U63 ( .A(B[8]), .Z(n506) );
  IV U64 ( .A(B[9]), .Z(n505) );
  IV U65 ( .A(B[10]), .Z(n504) );
  IV U66 ( .A(B[11]), .Z(n503) );
  IV U67 ( .A(B[12]), .Z(n502) );
  IV U68 ( .A(B[13]), .Z(n501) );
  IV U69 ( .A(B[14]), .Z(n500) );
  IV U70 ( .A(B[464]), .Z(n50) );
  IV U71 ( .A(B[509]), .Z(n5) );
  IV U72 ( .A(B[15]), .Z(n499) );
  IV U73 ( .A(B[16]), .Z(n498) );
  IV U74 ( .A(B[17]), .Z(n497) );
  IV U75 ( .A(B[18]), .Z(n496) );
  IV U76 ( .A(B[19]), .Z(n495) );
  IV U77 ( .A(B[20]), .Z(n494) );
  IV U78 ( .A(B[21]), .Z(n493) );
  IV U79 ( .A(B[22]), .Z(n492) );
  IV U80 ( .A(B[23]), .Z(n491) );
  IV U81 ( .A(B[24]), .Z(n490) );
  IV U82 ( .A(B[465]), .Z(n49) );
  IV U83 ( .A(B[25]), .Z(n489) );
  IV U84 ( .A(B[26]), .Z(n488) );
  IV U85 ( .A(B[27]), .Z(n487) );
  IV U86 ( .A(B[28]), .Z(n486) );
  IV U87 ( .A(B[29]), .Z(n485) );
  IV U88 ( .A(B[30]), .Z(n484) );
  IV U89 ( .A(B[31]), .Z(n483) );
  IV U90 ( .A(B[32]), .Z(n482) );
  IV U91 ( .A(B[33]), .Z(n481) );
  IV U92 ( .A(B[34]), .Z(n480) );
  IV U93 ( .A(B[466]), .Z(n48) );
  IV U94 ( .A(B[35]), .Z(n479) );
  IV U95 ( .A(B[36]), .Z(n478) );
  IV U96 ( .A(B[37]), .Z(n477) );
  IV U97 ( .A(B[38]), .Z(n476) );
  IV U98 ( .A(B[39]), .Z(n475) );
  IV U99 ( .A(B[40]), .Z(n474) );
  IV U100 ( .A(B[41]), .Z(n473) );
  IV U101 ( .A(B[42]), .Z(n472) );
  IV U102 ( .A(B[43]), .Z(n471) );
  IV U103 ( .A(B[44]), .Z(n470) );
  IV U104 ( .A(B[467]), .Z(n47) );
  IV U105 ( .A(B[45]), .Z(n469) );
  IV U106 ( .A(B[46]), .Z(n468) );
  IV U107 ( .A(B[47]), .Z(n467) );
  IV U108 ( .A(B[48]), .Z(n466) );
  IV U109 ( .A(B[49]), .Z(n465) );
  IV U110 ( .A(B[50]), .Z(n464) );
  IV U111 ( .A(B[51]), .Z(n463) );
  IV U112 ( .A(B[52]), .Z(n462) );
  IV U113 ( .A(B[53]), .Z(n461) );
  IV U114 ( .A(B[54]), .Z(n460) );
  IV U115 ( .A(B[468]), .Z(n46) );
  IV U116 ( .A(B[55]), .Z(n459) );
  IV U117 ( .A(B[56]), .Z(n458) );
  IV U118 ( .A(B[57]), .Z(n457) );
  IV U119 ( .A(B[58]), .Z(n456) );
  IV U120 ( .A(B[59]), .Z(n455) );
  IV U121 ( .A(B[60]), .Z(n454) );
  IV U122 ( .A(B[61]), .Z(n453) );
  IV U123 ( .A(B[62]), .Z(n452) );
  IV U124 ( .A(B[63]), .Z(n451) );
  IV U125 ( .A(B[64]), .Z(n450) );
  IV U126 ( .A(B[469]), .Z(n45) );
  IV U127 ( .A(B[65]), .Z(n449) );
  IV U128 ( .A(B[66]), .Z(n448) );
  IV U129 ( .A(B[67]), .Z(n447) );
  IV U130 ( .A(B[68]), .Z(n446) );
  IV U131 ( .A(B[69]), .Z(n445) );
  IV U132 ( .A(B[70]), .Z(n444) );
  IV U133 ( .A(B[71]), .Z(n443) );
  IV U134 ( .A(B[72]), .Z(n442) );
  IV U135 ( .A(B[73]), .Z(n441) );
  IV U136 ( .A(B[74]), .Z(n440) );
  IV U137 ( .A(B[470]), .Z(n44) );
  IV U138 ( .A(B[75]), .Z(n439) );
  IV U139 ( .A(B[76]), .Z(n438) );
  IV U140 ( .A(B[77]), .Z(n437) );
  IV U141 ( .A(B[78]), .Z(n436) );
  IV U142 ( .A(B[79]), .Z(n435) );
  IV U143 ( .A(B[80]), .Z(n434) );
  IV U144 ( .A(B[81]), .Z(n433) );
  IV U145 ( .A(B[82]), .Z(n432) );
  IV U146 ( .A(B[83]), .Z(n431) );
  IV U147 ( .A(B[84]), .Z(n430) );
  IV U148 ( .A(B[471]), .Z(n43) );
  IV U149 ( .A(B[85]), .Z(n429) );
  IV U150 ( .A(B[86]), .Z(n428) );
  IV U151 ( .A(B[87]), .Z(n427) );
  IV U152 ( .A(B[88]), .Z(n426) );
  IV U153 ( .A(B[89]), .Z(n425) );
  IV U154 ( .A(B[90]), .Z(n424) );
  IV U155 ( .A(B[91]), .Z(n423) );
  IV U156 ( .A(B[92]), .Z(n422) );
  IV U157 ( .A(B[93]), .Z(n421) );
  IV U158 ( .A(B[94]), .Z(n420) );
  IV U159 ( .A(B[472]), .Z(n42) );
  IV U160 ( .A(B[95]), .Z(n419) );
  IV U161 ( .A(B[96]), .Z(n418) );
  IV U162 ( .A(B[97]), .Z(n417) );
  IV U163 ( .A(B[98]), .Z(n416) );
  IV U164 ( .A(B[99]), .Z(n415) );
  IV U165 ( .A(B[100]), .Z(n414) );
  IV U166 ( .A(B[101]), .Z(n413) );
  IV U167 ( .A(B[102]), .Z(n412) );
  IV U168 ( .A(B[103]), .Z(n411) );
  IV U169 ( .A(B[104]), .Z(n410) );
  IV U170 ( .A(B[473]), .Z(n41) );
  IV U171 ( .A(B[105]), .Z(n409) );
  IV U172 ( .A(B[106]), .Z(n408) );
  IV U173 ( .A(B[107]), .Z(n407) );
  IV U174 ( .A(B[108]), .Z(n406) );
  IV U175 ( .A(B[109]), .Z(n405) );
  IV U176 ( .A(B[110]), .Z(n404) );
  IV U177 ( .A(B[111]), .Z(n403) );
  IV U178 ( .A(B[112]), .Z(n402) );
  IV U179 ( .A(B[113]), .Z(n401) );
  IV U180 ( .A(B[114]), .Z(n400) );
  IV U181 ( .A(B[474]), .Z(n40) );
  IV U182 ( .A(B[510]), .Z(n4) );
  IV U183 ( .A(B[115]), .Z(n399) );
  IV U184 ( .A(B[116]), .Z(n398) );
  IV U185 ( .A(B[117]), .Z(n397) );
  IV U186 ( .A(B[118]), .Z(n396) );
  IV U187 ( .A(B[119]), .Z(n395) );
  IV U188 ( .A(B[120]), .Z(n394) );
  IV U189 ( .A(B[121]), .Z(n393) );
  IV U190 ( .A(B[122]), .Z(n392) );
  IV U191 ( .A(B[123]), .Z(n391) );
  IV U192 ( .A(B[124]), .Z(n390) );
  IV U193 ( .A(B[475]), .Z(n39) );
  IV U194 ( .A(B[125]), .Z(n389) );
  IV U195 ( .A(B[126]), .Z(n388) );
  IV U196 ( .A(B[127]), .Z(n387) );
  IV U197 ( .A(B[128]), .Z(n386) );
  IV U198 ( .A(B[129]), .Z(n385) );
  IV U199 ( .A(B[130]), .Z(n384) );
  IV U200 ( .A(B[131]), .Z(n383) );
  IV U201 ( .A(B[132]), .Z(n382) );
  IV U202 ( .A(B[133]), .Z(n381) );
  IV U203 ( .A(B[134]), .Z(n380) );
  IV U204 ( .A(B[476]), .Z(n38) );
  IV U205 ( .A(B[135]), .Z(n379) );
  IV U206 ( .A(B[136]), .Z(n378) );
  IV U207 ( .A(B[137]), .Z(n377) );
  IV U208 ( .A(B[138]), .Z(n376) );
  IV U209 ( .A(B[139]), .Z(n375) );
  IV U210 ( .A(B[140]), .Z(n374) );
  IV U211 ( .A(B[141]), .Z(n373) );
  IV U212 ( .A(B[142]), .Z(n372) );
  IV U213 ( .A(B[143]), .Z(n371) );
  IV U214 ( .A(B[144]), .Z(n370) );
  IV U215 ( .A(B[477]), .Z(n37) );
  IV U216 ( .A(B[145]), .Z(n369) );
  IV U217 ( .A(B[146]), .Z(n368) );
  IV U218 ( .A(B[147]), .Z(n367) );
  IV U219 ( .A(B[148]), .Z(n366) );
  IV U220 ( .A(B[149]), .Z(n365) );
  IV U221 ( .A(B[150]), .Z(n364) );
  IV U222 ( .A(B[151]), .Z(n363) );
  IV U223 ( .A(B[152]), .Z(n362) );
  IV U224 ( .A(B[153]), .Z(n361) );
  IV U225 ( .A(B[154]), .Z(n360) );
  IV U226 ( .A(B[478]), .Z(n36) );
  IV U227 ( .A(B[155]), .Z(n359) );
  IV U228 ( .A(B[156]), .Z(n358) );
  IV U229 ( .A(B[157]), .Z(n357) );
  IV U230 ( .A(B[158]), .Z(n356) );
  IV U231 ( .A(B[159]), .Z(n355) );
  IV U232 ( .A(B[160]), .Z(n354) );
  IV U233 ( .A(B[161]), .Z(n353) );
  IV U234 ( .A(B[162]), .Z(n352) );
  IV U235 ( .A(B[163]), .Z(n351) );
  IV U236 ( .A(B[164]), .Z(n350) );
  IV U237 ( .A(B[479]), .Z(n35) );
  IV U238 ( .A(B[165]), .Z(n349) );
  IV U239 ( .A(B[166]), .Z(n348) );
  IV U240 ( .A(B[167]), .Z(n347) );
  IV U241 ( .A(B[168]), .Z(n346) );
  IV U242 ( .A(B[169]), .Z(n345) );
  IV U243 ( .A(B[170]), .Z(n344) );
  IV U244 ( .A(B[171]), .Z(n343) );
  IV U245 ( .A(B[172]), .Z(n342) );
  IV U246 ( .A(B[173]), .Z(n341) );
  IV U247 ( .A(B[174]), .Z(n340) );
  IV U248 ( .A(B[480]), .Z(n34) );
  IV U249 ( .A(B[175]), .Z(n339) );
  IV U250 ( .A(B[176]), .Z(n338) );
  IV U251 ( .A(B[177]), .Z(n337) );
  IV U252 ( .A(B[178]), .Z(n336) );
  IV U253 ( .A(B[179]), .Z(n335) );
  IV U254 ( .A(B[180]), .Z(n334) );
  IV U255 ( .A(B[181]), .Z(n333) );
  IV U256 ( .A(B[182]), .Z(n332) );
  IV U257 ( .A(B[183]), .Z(n331) );
  IV U258 ( .A(B[184]), .Z(n330) );
  IV U259 ( .A(B[481]), .Z(n33) );
  IV U260 ( .A(B[185]), .Z(n329) );
  IV U261 ( .A(B[186]), .Z(n328) );
  IV U262 ( .A(B[187]), .Z(n327) );
  IV U263 ( .A(B[188]), .Z(n326) );
  IV U264 ( .A(B[189]), .Z(n325) );
  IV U265 ( .A(B[190]), .Z(n324) );
  IV U266 ( .A(B[191]), .Z(n323) );
  IV U267 ( .A(B[192]), .Z(n322) );
  IV U268 ( .A(B[193]), .Z(n321) );
  IV U269 ( .A(B[194]), .Z(n320) );
  IV U270 ( .A(B[482]), .Z(n32) );
  IV U271 ( .A(B[195]), .Z(n319) );
  IV U272 ( .A(B[196]), .Z(n318) );
  IV U273 ( .A(B[197]), .Z(n317) );
  IV U274 ( .A(B[198]), .Z(n316) );
  IV U275 ( .A(B[199]), .Z(n315) );
  IV U276 ( .A(B[200]), .Z(n314) );
  IV U277 ( .A(B[201]), .Z(n313) );
  IV U278 ( .A(B[202]), .Z(n312) );
  IV U279 ( .A(B[203]), .Z(n311) );
  IV U280 ( .A(B[204]), .Z(n310) );
  IV U281 ( .A(B[483]), .Z(n31) );
  IV U282 ( .A(B[205]), .Z(n309) );
  IV U283 ( .A(B[206]), .Z(n308) );
  IV U284 ( .A(B[207]), .Z(n307) );
  IV U285 ( .A(B[208]), .Z(n306) );
  IV U286 ( .A(B[209]), .Z(n305) );
  IV U287 ( .A(B[210]), .Z(n304) );
  IV U288 ( .A(B[211]), .Z(n303) );
  IV U289 ( .A(B[212]), .Z(n302) );
  IV U290 ( .A(B[213]), .Z(n301) );
  IV U291 ( .A(B[214]), .Z(n300) );
  IV U292 ( .A(B[484]), .Z(n30) );
  IV U293 ( .A(B[511]), .Z(n3) );
  IV U294 ( .A(B[215]), .Z(n299) );
  IV U295 ( .A(B[216]), .Z(n298) );
  IV U296 ( .A(B[217]), .Z(n297) );
  IV U297 ( .A(B[218]), .Z(n296) );
  IV U298 ( .A(B[219]), .Z(n295) );
  IV U299 ( .A(B[220]), .Z(n294) );
  IV U300 ( .A(B[221]), .Z(n293) );
  IV U301 ( .A(B[222]), .Z(n292) );
  IV U302 ( .A(B[223]), .Z(n291) );
  IV U303 ( .A(B[224]), .Z(n290) );
  IV U304 ( .A(B[485]), .Z(n29) );
  IV U305 ( .A(B[225]), .Z(n289) );
  IV U306 ( .A(B[226]), .Z(n288) );
  IV U307 ( .A(B[227]), .Z(n287) );
  IV U308 ( .A(B[228]), .Z(n286) );
  IV U309 ( .A(B[229]), .Z(n285) );
  IV U310 ( .A(B[230]), .Z(n284) );
  IV U311 ( .A(B[231]), .Z(n283) );
  IV U312 ( .A(B[232]), .Z(n282) );
  IV U313 ( .A(B[233]), .Z(n281) );
  IV U314 ( .A(B[234]), .Z(n280) );
  IV U315 ( .A(B[486]), .Z(n28) );
  IV U316 ( .A(B[235]), .Z(n279) );
  IV U317 ( .A(B[236]), .Z(n278) );
  IV U318 ( .A(B[237]), .Z(n277) );
  IV U319 ( .A(B[238]), .Z(n276) );
  IV U320 ( .A(B[239]), .Z(n275) );
  IV U321 ( .A(B[240]), .Z(n274) );
  IV U322 ( .A(B[241]), .Z(n273) );
  IV U323 ( .A(B[242]), .Z(n272) );
  IV U324 ( .A(B[243]), .Z(n271) );
  IV U325 ( .A(B[244]), .Z(n270) );
  IV U326 ( .A(B[487]), .Z(n27) );
  IV U327 ( .A(B[245]), .Z(n269) );
  IV U328 ( .A(B[246]), .Z(n268) );
  IV U329 ( .A(B[247]), .Z(n267) );
  IV U330 ( .A(B[248]), .Z(n266) );
  IV U331 ( .A(B[249]), .Z(n265) );
  IV U332 ( .A(B[250]), .Z(n264) );
  IV U333 ( .A(B[251]), .Z(n263) );
  IV U334 ( .A(B[252]), .Z(n262) );
  IV U335 ( .A(B[253]), .Z(n261) );
  IV U336 ( .A(B[254]), .Z(n260) );
  IV U337 ( .A(B[488]), .Z(n26) );
  IV U338 ( .A(B[255]), .Z(n259) );
  IV U339 ( .A(B[256]), .Z(n258) );
  IV U340 ( .A(B[257]), .Z(n257) );
  IV U341 ( .A(B[258]), .Z(n256) );
  IV U342 ( .A(B[259]), .Z(n255) );
  IV U343 ( .A(B[260]), .Z(n254) );
  IV U344 ( .A(B[261]), .Z(n253) );
  IV U345 ( .A(B[262]), .Z(n252) );
  IV U346 ( .A(B[263]), .Z(n251) );
  IV U347 ( .A(B[264]), .Z(n250) );
  IV U348 ( .A(B[489]), .Z(n25) );
  IV U349 ( .A(B[265]), .Z(n249) );
  IV U350 ( .A(B[266]), .Z(n248) );
  IV U351 ( .A(B[267]), .Z(n247) );
  IV U352 ( .A(B[268]), .Z(n246) );
  IV U353 ( .A(B[269]), .Z(n245) );
  IV U354 ( .A(B[270]), .Z(n244) );
  IV U355 ( .A(B[271]), .Z(n243) );
  IV U356 ( .A(B[272]), .Z(n242) );
  IV U357 ( .A(B[273]), .Z(n241) );
  IV U358 ( .A(B[274]), .Z(n240) );
  IV U359 ( .A(B[490]), .Z(n24) );
  IV U360 ( .A(B[275]), .Z(n239) );
  IV U361 ( .A(B[276]), .Z(n238) );
  IV U362 ( .A(B[277]), .Z(n237) );
  IV U363 ( .A(B[278]), .Z(n236) );
  IV U364 ( .A(B[279]), .Z(n235) );
  IV U365 ( .A(B[280]), .Z(n234) );
  IV U366 ( .A(B[281]), .Z(n233) );
  IV U367 ( .A(B[282]), .Z(n232) );
  IV U368 ( .A(B[283]), .Z(n231) );
  IV U369 ( .A(B[284]), .Z(n230) );
  IV U370 ( .A(B[491]), .Z(n23) );
  IV U371 ( .A(B[285]), .Z(n229) );
  IV U372 ( .A(B[286]), .Z(n228) );
  IV U373 ( .A(B[287]), .Z(n227) );
  IV U374 ( .A(B[288]), .Z(n226) );
  IV U375 ( .A(B[289]), .Z(n225) );
  IV U376 ( .A(B[290]), .Z(n224) );
  IV U377 ( .A(B[291]), .Z(n223) );
  IV U378 ( .A(B[292]), .Z(n222) );
  IV U379 ( .A(B[293]), .Z(n221) );
  IV U380 ( .A(B[294]), .Z(n220) );
  IV U381 ( .A(B[492]), .Z(n22) );
  IV U382 ( .A(B[295]), .Z(n219) );
  IV U383 ( .A(B[296]), .Z(n218) );
  IV U384 ( .A(B[297]), .Z(n217) );
  IV U385 ( .A(B[298]), .Z(n216) );
  IV U386 ( .A(B[299]), .Z(n215) );
  IV U387 ( .A(B[300]), .Z(n214) );
  IV U388 ( .A(B[301]), .Z(n213) );
  IV U389 ( .A(B[302]), .Z(n212) );
  IV U390 ( .A(B[303]), .Z(n211) );
  IV U391 ( .A(B[304]), .Z(n210) );
  IV U392 ( .A(B[493]), .Z(n21) );
  IV U393 ( .A(B[305]), .Z(n209) );
  IV U394 ( .A(B[306]), .Z(n208) );
  IV U395 ( .A(B[307]), .Z(n207) );
  IV U396 ( .A(B[308]), .Z(n206) );
  IV U397 ( .A(B[309]), .Z(n205) );
  IV U398 ( .A(B[310]), .Z(n204) );
  IV U399 ( .A(B[311]), .Z(n203) );
  IV U400 ( .A(B[312]), .Z(n202) );
  IV U401 ( .A(B[313]), .Z(n201) );
  IV U402 ( .A(B[314]), .Z(n200) );
  IV U403 ( .A(B[494]), .Z(n20) );
  IV U404 ( .A(B[315]), .Z(n199) );
  IV U405 ( .A(B[316]), .Z(n198) );
  IV U406 ( .A(B[317]), .Z(n197) );
  IV U407 ( .A(B[318]), .Z(n196) );
  IV U408 ( .A(B[319]), .Z(n195) );
  IV U409 ( .A(B[320]), .Z(n194) );
  IV U410 ( .A(B[321]), .Z(n193) );
  IV U411 ( .A(B[322]), .Z(n192) );
  IV U412 ( .A(B[323]), .Z(n191) );
  IV U413 ( .A(B[324]), .Z(n190) );
  IV U414 ( .A(B[495]), .Z(n19) );
  IV U415 ( .A(B[325]), .Z(n189) );
  IV U416 ( .A(B[326]), .Z(n188) );
  IV U417 ( .A(B[327]), .Z(n187) );
  IV U418 ( .A(B[328]), .Z(n186) );
  IV U419 ( .A(B[329]), .Z(n185) );
  IV U420 ( .A(B[330]), .Z(n184) );
  IV U421 ( .A(B[331]), .Z(n183) );
  IV U422 ( .A(B[332]), .Z(n182) );
  IV U423 ( .A(B[333]), .Z(n181) );
  IV U424 ( .A(B[334]), .Z(n180) );
  IV U425 ( .A(B[496]), .Z(n18) );
  IV U426 ( .A(B[335]), .Z(n179) );
  IV U427 ( .A(B[336]), .Z(n178) );
  IV U428 ( .A(B[337]), .Z(n177) );
  IV U429 ( .A(B[338]), .Z(n176) );
  IV U430 ( .A(B[339]), .Z(n175) );
  IV U431 ( .A(B[340]), .Z(n174) );
  IV U432 ( .A(B[341]), .Z(n173) );
  IV U433 ( .A(B[342]), .Z(n172) );
  IV U434 ( .A(B[343]), .Z(n171) );
  IV U435 ( .A(B[344]), .Z(n170) );
  IV U436 ( .A(B[497]), .Z(n17) );
  IV U437 ( .A(B[345]), .Z(n169) );
  IV U438 ( .A(B[346]), .Z(n168) );
  IV U439 ( .A(B[347]), .Z(n167) );
  IV U440 ( .A(B[348]), .Z(n166) );
  IV U441 ( .A(B[349]), .Z(n165) );
  IV U442 ( .A(B[350]), .Z(n164) );
  IV U443 ( .A(B[351]), .Z(n163) );
  IV U444 ( .A(B[352]), .Z(n162) );
  IV U445 ( .A(B[353]), .Z(n161) );
  IV U446 ( .A(B[354]), .Z(n160) );
  IV U447 ( .A(B[498]), .Z(n16) );
  IV U448 ( .A(B[355]), .Z(n159) );
  IV U449 ( .A(B[356]), .Z(n158) );
  IV U450 ( .A(B[357]), .Z(n157) );
  IV U451 ( .A(B[358]), .Z(n156) );
  IV U452 ( .A(B[359]), .Z(n155) );
  IV U453 ( .A(B[360]), .Z(n154) );
  IV U454 ( .A(B[361]), .Z(n153) );
  IV U455 ( .A(B[362]), .Z(n152) );
  IV U456 ( .A(B[363]), .Z(n151) );
  IV U457 ( .A(B[364]), .Z(n150) );
  IV U458 ( .A(B[499]), .Z(n15) );
  IV U459 ( .A(B[365]), .Z(n149) );
  IV U460 ( .A(B[366]), .Z(n148) );
  IV U461 ( .A(B[367]), .Z(n147) );
  IV U462 ( .A(B[368]), .Z(n146) );
  IV U463 ( .A(B[369]), .Z(n145) );
  IV U464 ( .A(B[370]), .Z(n144) );
  IV U465 ( .A(B[371]), .Z(n143) );
  IV U466 ( .A(B[372]), .Z(n142) );
  IV U467 ( .A(B[373]), .Z(n141) );
  IV U468 ( .A(B[374]), .Z(n140) );
  IV U469 ( .A(B[500]), .Z(n14) );
  IV U470 ( .A(B[375]), .Z(n139) );
  IV U471 ( .A(B[376]), .Z(n138) );
  IV U472 ( .A(B[377]), .Z(n137) );
  IV U473 ( .A(B[378]), .Z(n136) );
  IV U474 ( .A(B[379]), .Z(n135) );
  IV U475 ( .A(B[380]), .Z(n134) );
  IV U476 ( .A(B[381]), .Z(n133) );
  IV U477 ( .A(B[382]), .Z(n132) );
  IV U478 ( .A(B[383]), .Z(n131) );
  IV U479 ( .A(B[384]), .Z(n130) );
  IV U480 ( .A(B[501]), .Z(n13) );
  IV U481 ( .A(B[385]), .Z(n129) );
  IV U482 ( .A(B[386]), .Z(n128) );
  IV U483 ( .A(B[387]), .Z(n127) );
  IV U484 ( .A(B[388]), .Z(n126) );
  IV U485 ( .A(B[389]), .Z(n125) );
  IV U486 ( .A(B[390]), .Z(n124) );
  IV U487 ( .A(B[391]), .Z(n123) );
  IV U488 ( .A(B[392]), .Z(n122) );
  IV U489 ( .A(B[393]), .Z(n121) );
  IV U490 ( .A(B[394]), .Z(n120) );
  IV U491 ( .A(B[502]), .Z(n12) );
  IV U492 ( .A(B[395]), .Z(n119) );
  IV U493 ( .A(B[396]), .Z(n118) );
  IV U494 ( .A(B[397]), .Z(n117) );
  IV U495 ( .A(B[398]), .Z(n116) );
  IV U496 ( .A(B[399]), .Z(n115) );
  IV U497 ( .A(B[400]), .Z(n114) );
  IV U498 ( .A(B[401]), .Z(n113) );
  IV U499 ( .A(B[402]), .Z(n112) );
  IV U500 ( .A(B[403]), .Z(n111) );
  IV U501 ( .A(B[404]), .Z(n110) );
  IV U502 ( .A(B[503]), .Z(n11) );
  IV U503 ( .A(B[405]), .Z(n109) );
  IV U504 ( .A(B[406]), .Z(n108) );
  IV U505 ( .A(B[407]), .Z(n107) );
  IV U506 ( .A(B[408]), .Z(n106) );
  IV U507 ( .A(B[409]), .Z(n105) );
  IV U508 ( .A(B[410]), .Z(n104) );
  IV U509 ( .A(B[411]), .Z(n103) );
  IV U510 ( .A(B[412]), .Z(n102) );
  IV U511 ( .A(B[413]), .Z(n101) );
  IV U512 ( .A(B[414]), .Z(n100) );
  IV U513 ( .A(B[504]), .Z(n10) );
endmodule


module FA_4896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_4897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  NANDN U1 ( .A(CI), .B(S), .Z(CO) );
  XNOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_4898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N514_0 ( A, B, S, CO );
  input [513:0] A;
  input [513:0] B;
  output [513:0] S;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514;
  wire   [513:1] C;

  FA_5409 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n514), .CI(1'b1), .S(
        S[0]), .CO(C[1]) );
  FA_5408 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n513), .CI(C[1]), .S(
        S[1]), .CO(C[2]) );
  FA_5407 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n512), .CI(C[2]), .S(
        S[2]), .CO(C[3]) );
  FA_5406 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n511), .CI(C[3]), .S(
        S[3]), .CO(C[4]) );
  FA_5405 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n510), .CI(C[4]), .S(
        S[4]), .CO(C[5]) );
  FA_5404 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n509), .CI(C[5]), .S(
        S[5]), .CO(C[6]) );
  FA_5403 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n508), .CI(C[6]), .S(
        S[6]), .CO(C[7]) );
  FA_5402 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n507), .CI(C[7]), .S(
        S[7]), .CO(C[8]) );
  FA_5401 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n506), .CI(C[8]), .S(
        S[8]), .CO(C[9]) );
  FA_5400 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n505), .CI(C[9]), .S(
        S[9]), .CO(C[10]) );
  FA_5399 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n504), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_5398 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n503), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_5397 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n502), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_5396 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n501), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_5395 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n500), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_5394 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n499), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_5393 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n498), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_5392 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n497), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_5391 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n496), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_5390 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n495), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_5389 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n494), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_5388 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n493), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_5387 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n492), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_5386 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n491), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_5385 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n490), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_5384 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n489), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_5383 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n488), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_5382 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n487), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_5381 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n486), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_5380 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n485), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_5379 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n484), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_5378 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n483), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_5377 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n482), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_5376 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n481), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_5375 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n480), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_5374 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n479), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_5373 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n478), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_5372 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n477), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_5371 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n476), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_5370 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n475), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_5369 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n474), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_5368 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n473), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_5367 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n472), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_5366 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n471), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_5365 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n470), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_5364 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n469), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_5363 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n468), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_5362 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n467), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_5361 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n466), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_5360 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n465), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_5359 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n464), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_5358 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n463), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_5357 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n462), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_5356 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n461), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_5355 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n460), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_5354 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n459), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_5353 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n458), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_5352 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n457), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_5351 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n456), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_5350 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n455), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_5349 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n454), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_5348 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n453), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_5347 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n452), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_5346 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n451), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_5345 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n450), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_5344 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n449), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_5343 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n448), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_5342 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n447), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_5341 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n446), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_5340 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n445), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_5339 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n444), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_5338 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n443), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_5337 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n442), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_5336 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n441), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_5335 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n440), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_5334 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n439), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_5333 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n438), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_5332 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n437), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_5331 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n436), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_5330 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n435), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_5329 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n434), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_5328 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n433), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_5327 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n432), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_5326 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n431), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_5325 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n430), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_5324 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n429), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_5323 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n428), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_5322 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n427), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_5321 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n426), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_5320 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n425), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_5319 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n424), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_5318 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n423), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_5317 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n422), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_5316 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n421), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_5315 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n420), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_5314 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n419), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_5313 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n418), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_5312 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n417), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_5311 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n416), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_5310 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n415), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_5309 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n414), .CI(C[100]), .S(S[100]), .CO(C[101]) );
  FA_5308 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n413), .CI(C[101]), .S(S[101]), .CO(C[102]) );
  FA_5307 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n412), .CI(C[102]), .S(S[102]), .CO(C[103]) );
  FA_5306 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n411), .CI(C[103]), .S(S[103]), .CO(C[104]) );
  FA_5305 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n410), .CI(C[104]), .S(S[104]), .CO(C[105]) );
  FA_5304 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n409), .CI(C[105]), .S(S[105]), .CO(C[106]) );
  FA_5303 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n408), .CI(C[106]), .S(S[106]), .CO(C[107]) );
  FA_5302 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n407), .CI(C[107]), .S(S[107]), .CO(C[108]) );
  FA_5301 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n406), .CI(C[108]), .S(S[108]), .CO(C[109]) );
  FA_5300 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n405), .CI(C[109]), .S(S[109]), .CO(C[110]) );
  FA_5299 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n404), .CI(C[110]), .S(S[110]), .CO(C[111]) );
  FA_5298 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n403), .CI(C[111]), .S(S[111]), .CO(C[112]) );
  FA_5297 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n402), .CI(C[112]), .S(S[112]), .CO(C[113]) );
  FA_5296 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n401), .CI(C[113]), .S(S[113]), .CO(C[114]) );
  FA_5295 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n400), .CI(C[114]), .S(S[114]), .CO(C[115]) );
  FA_5294 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n399), .CI(C[115]), .S(S[115]), .CO(C[116]) );
  FA_5293 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n398), .CI(C[116]), .S(S[116]), .CO(C[117]) );
  FA_5292 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n397), .CI(C[117]), .S(S[117]), .CO(C[118]) );
  FA_5291 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n396), .CI(C[118]), .S(S[118]), .CO(C[119]) );
  FA_5290 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n395), .CI(C[119]), .S(S[119]), .CO(C[120]) );
  FA_5289 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n394), .CI(C[120]), .S(S[120]), .CO(C[121]) );
  FA_5288 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n393), .CI(C[121]), .S(S[121]), .CO(C[122]) );
  FA_5287 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n392), .CI(C[122]), .S(S[122]), .CO(C[123]) );
  FA_5286 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n391), .CI(C[123]), .S(S[123]), .CO(C[124]) );
  FA_5285 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n390), .CI(C[124]), .S(S[124]), .CO(C[125]) );
  FA_5284 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n389), .CI(C[125]), .S(S[125]), .CO(C[126]) );
  FA_5283 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n388), .CI(C[126]), .S(S[126]), .CO(C[127]) );
  FA_5282 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n387), .CI(C[127]), .S(S[127]), .CO(C[128]) );
  FA_5281 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n386), .CI(C[128]), .S(S[128]), .CO(C[129]) );
  FA_5280 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n385), .CI(C[129]), .S(S[129]), .CO(C[130]) );
  FA_5279 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n384), .CI(C[130]), .S(S[130]), .CO(C[131]) );
  FA_5278 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n383), .CI(C[131]), .S(S[131]), .CO(C[132]) );
  FA_5277 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n382), .CI(C[132]), .S(S[132]), .CO(C[133]) );
  FA_5276 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n381), .CI(C[133]), .S(S[133]), .CO(C[134]) );
  FA_5275 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n380), .CI(C[134]), .S(S[134]), .CO(C[135]) );
  FA_5274 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n379), .CI(C[135]), .S(S[135]), .CO(C[136]) );
  FA_5273 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n378), .CI(C[136]), .S(S[136]), .CO(C[137]) );
  FA_5272 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n377), .CI(C[137]), .S(S[137]), .CO(C[138]) );
  FA_5271 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n376), .CI(C[138]), .S(S[138]), .CO(C[139]) );
  FA_5270 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n375), .CI(C[139]), .S(S[139]), .CO(C[140]) );
  FA_5269 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n374), .CI(C[140]), .S(S[140]), .CO(C[141]) );
  FA_5268 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n373), .CI(C[141]), .S(S[141]), .CO(C[142]) );
  FA_5267 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n372), .CI(C[142]), .S(S[142]), .CO(C[143]) );
  FA_5266 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n371), .CI(C[143]), .S(S[143]), .CO(C[144]) );
  FA_5265 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n370), .CI(C[144]), .S(S[144]), .CO(C[145]) );
  FA_5264 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n369), .CI(C[145]), .S(S[145]), .CO(C[146]) );
  FA_5263 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n368), .CI(C[146]), .S(S[146]), .CO(C[147]) );
  FA_5262 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n367), .CI(C[147]), .S(S[147]), .CO(C[148]) );
  FA_5261 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n366), .CI(C[148]), .S(S[148]), .CO(C[149]) );
  FA_5260 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n365), .CI(C[149]), .S(S[149]), .CO(C[150]) );
  FA_5259 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n364), .CI(C[150]), .S(S[150]), .CO(C[151]) );
  FA_5258 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n363), .CI(C[151]), .S(S[151]), .CO(C[152]) );
  FA_5257 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n362), .CI(C[152]), .S(S[152]), .CO(C[153]) );
  FA_5256 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n361), .CI(C[153]), .S(S[153]), .CO(C[154]) );
  FA_5255 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n360), .CI(C[154]), .S(S[154]), .CO(C[155]) );
  FA_5254 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n359), .CI(C[155]), .S(S[155]), .CO(C[156]) );
  FA_5253 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n358), .CI(C[156]), .S(S[156]), .CO(C[157]) );
  FA_5252 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n357), .CI(C[157]), .S(S[157]), .CO(C[158]) );
  FA_5251 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n356), .CI(C[158]), .S(S[158]), .CO(C[159]) );
  FA_5250 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n355), .CI(C[159]), .S(S[159]), .CO(C[160]) );
  FA_5249 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n354), .CI(C[160]), .S(S[160]), .CO(C[161]) );
  FA_5248 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n353), .CI(C[161]), .S(S[161]), .CO(C[162]) );
  FA_5247 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n352), .CI(C[162]), .S(S[162]), .CO(C[163]) );
  FA_5246 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n351), .CI(C[163]), .S(S[163]), .CO(C[164]) );
  FA_5245 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n350), .CI(C[164]), .S(S[164]), .CO(C[165]) );
  FA_5244 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n349), .CI(C[165]), .S(S[165]), .CO(C[166]) );
  FA_5243 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n348), .CI(C[166]), .S(S[166]), .CO(C[167]) );
  FA_5242 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n347), .CI(C[167]), .S(S[167]), .CO(C[168]) );
  FA_5241 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n346), .CI(C[168]), .S(S[168]), .CO(C[169]) );
  FA_5240 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n345), .CI(C[169]), .S(S[169]), .CO(C[170]) );
  FA_5239 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n344), .CI(C[170]), .S(S[170]), .CO(C[171]) );
  FA_5238 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n343), .CI(C[171]), .S(S[171]), .CO(C[172]) );
  FA_5237 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n342), .CI(C[172]), .S(S[172]), .CO(C[173]) );
  FA_5236 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n341), .CI(C[173]), .S(S[173]), .CO(C[174]) );
  FA_5235 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n340), .CI(C[174]), .S(S[174]), .CO(C[175]) );
  FA_5234 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n339), .CI(C[175]), .S(S[175]), .CO(C[176]) );
  FA_5233 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n338), .CI(C[176]), .S(S[176]), .CO(C[177]) );
  FA_5232 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n337), .CI(C[177]), .S(S[177]), .CO(C[178]) );
  FA_5231 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n336), .CI(C[178]), .S(S[178]), .CO(C[179]) );
  FA_5230 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n335), .CI(C[179]), .S(S[179]), .CO(C[180]) );
  FA_5229 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n334), .CI(C[180]), .S(S[180]), .CO(C[181]) );
  FA_5228 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n333), .CI(C[181]), .S(S[181]), .CO(C[182]) );
  FA_5227 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n332), .CI(C[182]), .S(S[182]), .CO(C[183]) );
  FA_5226 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n331), .CI(C[183]), .S(S[183]), .CO(C[184]) );
  FA_5225 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n330), .CI(C[184]), .S(S[184]), .CO(C[185]) );
  FA_5224 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n329), .CI(C[185]), .S(S[185]), .CO(C[186]) );
  FA_5223 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n328), .CI(C[186]), .S(S[186]), .CO(C[187]) );
  FA_5222 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n327), .CI(C[187]), .S(S[187]), .CO(C[188]) );
  FA_5221 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n326), .CI(C[188]), .S(S[188]), .CO(C[189]) );
  FA_5220 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n325), .CI(C[189]), .S(S[189]), .CO(C[190]) );
  FA_5219 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n324), .CI(C[190]), .S(S[190]), .CO(C[191]) );
  FA_5218 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n323), .CI(C[191]), .S(S[191]), .CO(C[192]) );
  FA_5217 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n322), .CI(C[192]), .S(S[192]), .CO(C[193]) );
  FA_5216 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n321), .CI(C[193]), .S(S[193]), .CO(C[194]) );
  FA_5215 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n320), .CI(C[194]), .S(S[194]), .CO(C[195]) );
  FA_5214 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n319), .CI(C[195]), .S(S[195]), .CO(C[196]) );
  FA_5213 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n318), .CI(C[196]), .S(S[196]), .CO(C[197]) );
  FA_5212 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n317), .CI(C[197]), .S(S[197]), .CO(C[198]) );
  FA_5211 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n316), .CI(C[198]), .S(S[198]), .CO(C[199]) );
  FA_5210 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n315), .CI(C[199]), .S(S[199]), .CO(C[200]) );
  FA_5209 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n314), .CI(C[200]), .S(S[200]), .CO(C[201]) );
  FA_5208 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n313), .CI(C[201]), .S(S[201]), .CO(C[202]) );
  FA_5207 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n312), .CI(C[202]), .S(S[202]), .CO(C[203]) );
  FA_5206 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n311), .CI(C[203]), .S(S[203]), .CO(C[204]) );
  FA_5205 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n310), .CI(C[204]), .S(S[204]), .CO(C[205]) );
  FA_5204 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n309), .CI(C[205]), .S(S[205]), .CO(C[206]) );
  FA_5203 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n308), .CI(C[206]), .S(S[206]), .CO(C[207]) );
  FA_5202 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n307), .CI(C[207]), .S(S[207]), .CO(C[208]) );
  FA_5201 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n306), .CI(C[208]), .S(S[208]), .CO(C[209]) );
  FA_5200 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n305), .CI(C[209]), .S(S[209]), .CO(C[210]) );
  FA_5199 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n304), .CI(C[210]), .S(S[210]), .CO(C[211]) );
  FA_5198 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n303), .CI(C[211]), .S(S[211]), .CO(C[212]) );
  FA_5197 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n302), .CI(C[212]), .S(S[212]), .CO(C[213]) );
  FA_5196 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n301), .CI(C[213]), .S(S[213]), .CO(C[214]) );
  FA_5195 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n300), .CI(C[214]), .S(S[214]), .CO(C[215]) );
  FA_5194 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n299), .CI(C[215]), .S(S[215]), .CO(C[216]) );
  FA_5193 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n298), .CI(C[216]), .S(S[216]), .CO(C[217]) );
  FA_5192 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n297), .CI(C[217]), .S(S[217]), .CO(C[218]) );
  FA_5191 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n296), .CI(C[218]), .S(S[218]), .CO(C[219]) );
  FA_5190 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n295), .CI(C[219]), .S(S[219]), .CO(C[220]) );
  FA_5189 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n294), .CI(C[220]), .S(S[220]), .CO(C[221]) );
  FA_5188 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n293), .CI(C[221]), .S(S[221]), .CO(C[222]) );
  FA_5187 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n292), .CI(C[222]), .S(S[222]), .CO(C[223]) );
  FA_5186 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n291), .CI(C[223]), .S(S[223]), .CO(C[224]) );
  FA_5185 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n290), .CI(C[224]), .S(S[224]), .CO(C[225]) );
  FA_5184 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n289), .CI(C[225]), .S(S[225]), .CO(C[226]) );
  FA_5183 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n288), .CI(C[226]), .S(S[226]), .CO(C[227]) );
  FA_5182 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n287), .CI(C[227]), .S(S[227]), .CO(C[228]) );
  FA_5181 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n286), .CI(C[228]), .S(S[228]), .CO(C[229]) );
  FA_5180 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n285), .CI(C[229]), .S(S[229]), .CO(C[230]) );
  FA_5179 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n284), .CI(C[230]), .S(S[230]), .CO(C[231]) );
  FA_5178 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n283), .CI(C[231]), .S(S[231]), .CO(C[232]) );
  FA_5177 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n282), .CI(C[232]), .S(S[232]), .CO(C[233]) );
  FA_5176 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n281), .CI(C[233]), .S(S[233]), .CO(C[234]) );
  FA_5175 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n280), .CI(C[234]), .S(S[234]), .CO(C[235]) );
  FA_5174 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n279), .CI(C[235]), .S(S[235]), .CO(C[236]) );
  FA_5173 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n278), .CI(C[236]), .S(S[236]), .CO(C[237]) );
  FA_5172 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n277), .CI(C[237]), .S(S[237]), .CO(C[238]) );
  FA_5171 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n276), .CI(C[238]), .S(S[238]), .CO(C[239]) );
  FA_5170 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n275), .CI(C[239]), .S(S[239]), .CO(C[240]) );
  FA_5169 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n274), .CI(C[240]), .S(S[240]), .CO(C[241]) );
  FA_5168 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n273), .CI(C[241]), .S(S[241]), .CO(C[242]) );
  FA_5167 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n272), .CI(C[242]), .S(S[242]), .CO(C[243]) );
  FA_5166 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n271), .CI(C[243]), .S(S[243]), .CO(C[244]) );
  FA_5165 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n270), .CI(C[244]), .S(S[244]), .CO(C[245]) );
  FA_5164 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n269), .CI(C[245]), .S(S[245]), .CO(C[246]) );
  FA_5163 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n268), .CI(C[246]), .S(S[246]), .CO(C[247]) );
  FA_5162 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n267), .CI(C[247]), .S(S[247]), .CO(C[248]) );
  FA_5161 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n266), .CI(C[248]), .S(S[248]), .CO(C[249]) );
  FA_5160 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n265), .CI(C[249]), .S(S[249]), .CO(C[250]) );
  FA_5159 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n264), .CI(C[250]), .S(S[250]), .CO(C[251]) );
  FA_5158 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n263), .CI(C[251]), .S(S[251]), .CO(C[252]) );
  FA_5157 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n262), .CI(C[252]), .S(S[252]), .CO(C[253]) );
  FA_5156 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n261), .CI(C[253]), .S(S[253]), .CO(C[254]) );
  FA_5155 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n260), .CI(C[254]), .S(S[254]), .CO(C[255]) );
  FA_5154 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n259), .CI(C[255]), .S(S[255]), .CO(C[256]) );
  FA_5153 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n258), .CI(C[256]), .S(S[256]), .CO(C[257]) );
  FA_5152 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n257), .CI(C[257]), .S(S[257]), .CO(C[258]) );
  FA_5151 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n256), .CI(C[258]), .S(S[258]), .CO(C[259]) );
  FA_5150 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n255), .CI(C[259]), .S(S[259]), .CO(C[260]) );
  FA_5149 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n254), .CI(C[260]), .S(S[260]), .CO(C[261]) );
  FA_5148 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n253), .CI(C[261]), .S(S[261]), .CO(C[262]) );
  FA_5147 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n252), .CI(C[262]), .S(S[262]), .CO(C[263]) );
  FA_5146 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n251), .CI(C[263]), .S(S[263]), .CO(C[264]) );
  FA_5145 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n250), .CI(C[264]), .S(S[264]), .CO(C[265]) );
  FA_5144 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n249), .CI(C[265]), .S(S[265]), .CO(C[266]) );
  FA_5143 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n248), .CI(C[266]), .S(S[266]), .CO(C[267]) );
  FA_5142 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n247), .CI(C[267]), .S(S[267]), .CO(C[268]) );
  FA_5141 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n246), .CI(C[268]), .S(S[268]), .CO(C[269]) );
  FA_5140 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n245), .CI(C[269]), .S(S[269]), .CO(C[270]) );
  FA_5139 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n244), .CI(C[270]), .S(S[270]), .CO(C[271]) );
  FA_5138 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n243), .CI(C[271]), .S(S[271]), .CO(C[272]) );
  FA_5137 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n242), .CI(C[272]), .S(S[272]), .CO(C[273]) );
  FA_5136 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n241), .CI(C[273]), .S(S[273]), .CO(C[274]) );
  FA_5135 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n240), .CI(C[274]), .S(S[274]), .CO(C[275]) );
  FA_5134 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n239), .CI(C[275]), .S(S[275]), .CO(C[276]) );
  FA_5133 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n238), .CI(C[276]), .S(S[276]), .CO(C[277]) );
  FA_5132 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n237), .CI(C[277]), .S(S[277]), .CO(C[278]) );
  FA_5131 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n236), .CI(C[278]), .S(S[278]), .CO(C[279]) );
  FA_5130 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n235), .CI(C[279]), .S(S[279]), .CO(C[280]) );
  FA_5129 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n234), .CI(C[280]), .S(S[280]), .CO(C[281]) );
  FA_5128 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n233), .CI(C[281]), .S(S[281]), .CO(C[282]) );
  FA_5127 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n232), .CI(C[282]), .S(S[282]), .CO(C[283]) );
  FA_5126 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n231), .CI(C[283]), .S(S[283]), .CO(C[284]) );
  FA_5125 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n230), .CI(C[284]), .S(S[284]), .CO(C[285]) );
  FA_5124 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n229), .CI(C[285]), .S(S[285]), .CO(C[286]) );
  FA_5123 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n228), .CI(C[286]), .S(S[286]), .CO(C[287]) );
  FA_5122 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n227), .CI(C[287]), .S(S[287]), .CO(C[288]) );
  FA_5121 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n226), .CI(C[288]), .S(S[288]), .CO(C[289]) );
  FA_5120 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n225), .CI(C[289]), .S(S[289]), .CO(C[290]) );
  FA_5119 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n224), .CI(C[290]), .S(S[290]), .CO(C[291]) );
  FA_5118 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n223), .CI(C[291]), .S(S[291]), .CO(C[292]) );
  FA_5117 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n222), .CI(C[292]), .S(S[292]), .CO(C[293]) );
  FA_5116 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n221), .CI(C[293]), .S(S[293]), .CO(C[294]) );
  FA_5115 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n220), .CI(C[294]), .S(S[294]), .CO(C[295]) );
  FA_5114 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n219), .CI(C[295]), .S(S[295]), .CO(C[296]) );
  FA_5113 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n218), .CI(C[296]), .S(S[296]), .CO(C[297]) );
  FA_5112 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n217), .CI(C[297]), .S(S[297]), .CO(C[298]) );
  FA_5111 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n216), .CI(C[298]), .S(S[298]), .CO(C[299]) );
  FA_5110 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n215), .CI(C[299]), .S(S[299]), .CO(C[300]) );
  FA_5109 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n214), .CI(C[300]), .S(S[300]), .CO(C[301]) );
  FA_5108 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n213), .CI(C[301]), .S(S[301]), .CO(C[302]) );
  FA_5107 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n212), .CI(C[302]), .S(S[302]), .CO(C[303]) );
  FA_5106 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n211), .CI(C[303]), .S(S[303]), .CO(C[304]) );
  FA_5105 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n210), .CI(C[304]), .S(S[304]), .CO(C[305]) );
  FA_5104 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n209), .CI(C[305]), .S(S[305]), .CO(C[306]) );
  FA_5103 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n208), .CI(C[306]), .S(S[306]), .CO(C[307]) );
  FA_5102 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n207), .CI(C[307]), .S(S[307]), .CO(C[308]) );
  FA_5101 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n206), .CI(C[308]), .S(S[308]), .CO(C[309]) );
  FA_5100 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n205), .CI(C[309]), .S(S[309]), .CO(C[310]) );
  FA_5099 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n204), .CI(C[310]), .S(S[310]), .CO(C[311]) );
  FA_5098 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n203), .CI(C[311]), .S(S[311]), .CO(C[312]) );
  FA_5097 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n202), .CI(C[312]), .S(S[312]), .CO(C[313]) );
  FA_5096 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n201), .CI(C[313]), .S(S[313]), .CO(C[314]) );
  FA_5095 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n200), .CI(C[314]), .S(S[314]), .CO(C[315]) );
  FA_5094 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n199), .CI(C[315]), .S(S[315]), .CO(C[316]) );
  FA_5093 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n198), .CI(C[316]), .S(S[316]), .CO(C[317]) );
  FA_5092 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n197), .CI(C[317]), .S(S[317]), .CO(C[318]) );
  FA_5091 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n196), .CI(C[318]), .S(S[318]), .CO(C[319]) );
  FA_5090 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n195), .CI(C[319]), .S(S[319]), .CO(C[320]) );
  FA_5089 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n194), .CI(C[320]), .S(S[320]), .CO(C[321]) );
  FA_5088 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n193), .CI(C[321]), .S(S[321]), .CO(C[322]) );
  FA_5087 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n192), .CI(C[322]), .S(S[322]), .CO(C[323]) );
  FA_5086 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n191), .CI(C[323]), .S(S[323]), .CO(C[324]) );
  FA_5085 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n190), .CI(C[324]), .S(S[324]), .CO(C[325]) );
  FA_5084 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n189), .CI(C[325]), .S(S[325]), .CO(C[326]) );
  FA_5083 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n188), .CI(C[326]), .S(S[326]), .CO(C[327]) );
  FA_5082 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n187), .CI(C[327]), .S(S[327]), .CO(C[328]) );
  FA_5081 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n186), .CI(C[328]), .S(S[328]), .CO(C[329]) );
  FA_5080 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n185), .CI(C[329]), .S(S[329]), .CO(C[330]) );
  FA_5079 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n184), .CI(C[330]), .S(S[330]), .CO(C[331]) );
  FA_5078 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n183), .CI(C[331]), .S(S[331]), .CO(C[332]) );
  FA_5077 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n182), .CI(C[332]), .S(S[332]), .CO(C[333]) );
  FA_5076 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n181), .CI(C[333]), .S(S[333]), .CO(C[334]) );
  FA_5075 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n180), .CI(C[334]), .S(S[334]), .CO(C[335]) );
  FA_5074 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n179), .CI(C[335]), .S(S[335]), .CO(C[336]) );
  FA_5073 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n178), .CI(C[336]), .S(S[336]), .CO(C[337]) );
  FA_5072 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n177), .CI(C[337]), .S(S[337]), .CO(C[338]) );
  FA_5071 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n176), .CI(C[338]), .S(S[338]), .CO(C[339]) );
  FA_5070 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n175), .CI(C[339]), .S(S[339]), .CO(C[340]) );
  FA_5069 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n174), .CI(C[340]), .S(S[340]), .CO(C[341]) );
  FA_5068 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n173), .CI(C[341]), .S(S[341]), .CO(C[342]) );
  FA_5067 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n172), .CI(C[342]), .S(S[342]), .CO(C[343]) );
  FA_5066 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n171), .CI(C[343]), .S(S[343]), .CO(C[344]) );
  FA_5065 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n170), .CI(C[344]), .S(S[344]), .CO(C[345]) );
  FA_5064 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n169), .CI(C[345]), .S(S[345]), .CO(C[346]) );
  FA_5063 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n168), .CI(C[346]), .S(S[346]), .CO(C[347]) );
  FA_5062 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n167), .CI(C[347]), .S(S[347]), .CO(C[348]) );
  FA_5061 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n166), .CI(C[348]), .S(S[348]), .CO(C[349]) );
  FA_5060 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n165), .CI(C[349]), .S(S[349]), .CO(C[350]) );
  FA_5059 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n164), .CI(C[350]), .S(S[350]), .CO(C[351]) );
  FA_5058 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n163), .CI(C[351]), .S(S[351]), .CO(C[352]) );
  FA_5057 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n162), .CI(C[352]), .S(S[352]), .CO(C[353]) );
  FA_5056 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n161), .CI(C[353]), .S(S[353]), .CO(C[354]) );
  FA_5055 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n160), .CI(C[354]), .S(S[354]), .CO(C[355]) );
  FA_5054 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n159), .CI(C[355]), .S(S[355]), .CO(C[356]) );
  FA_5053 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n158), .CI(C[356]), .S(S[356]), .CO(C[357]) );
  FA_5052 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n157), .CI(C[357]), .S(S[357]), .CO(C[358]) );
  FA_5051 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n156), .CI(C[358]), .S(S[358]), .CO(C[359]) );
  FA_5050 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n155), .CI(C[359]), .S(S[359]), .CO(C[360]) );
  FA_5049 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n154), .CI(C[360]), .S(S[360]), .CO(C[361]) );
  FA_5048 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n153), .CI(C[361]), .S(S[361]), .CO(C[362]) );
  FA_5047 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n152), .CI(C[362]), .S(S[362]), .CO(C[363]) );
  FA_5046 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n151), .CI(C[363]), .S(S[363]), .CO(C[364]) );
  FA_5045 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n150), .CI(C[364]), .S(S[364]), .CO(C[365]) );
  FA_5044 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n149), .CI(C[365]), .S(S[365]), .CO(C[366]) );
  FA_5043 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n148), .CI(C[366]), .S(S[366]), .CO(C[367]) );
  FA_5042 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n147), .CI(C[367]), .S(S[367]), .CO(C[368]) );
  FA_5041 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n146), .CI(C[368]), .S(S[368]), .CO(C[369]) );
  FA_5040 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n145), .CI(C[369]), .S(S[369]), .CO(C[370]) );
  FA_5039 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n144), .CI(C[370]), .S(S[370]), .CO(C[371]) );
  FA_5038 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n143), .CI(C[371]), .S(S[371]), .CO(C[372]) );
  FA_5037 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n142), .CI(C[372]), .S(S[372]), .CO(C[373]) );
  FA_5036 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n141), .CI(C[373]), .S(S[373]), .CO(C[374]) );
  FA_5035 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n140), .CI(C[374]), .S(S[374]), .CO(C[375]) );
  FA_5034 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n139), .CI(C[375]), .S(S[375]), .CO(C[376]) );
  FA_5033 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n138), .CI(C[376]), .S(S[376]), .CO(C[377]) );
  FA_5032 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n137), .CI(C[377]), .S(S[377]), .CO(C[378]) );
  FA_5031 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n136), .CI(C[378]), .S(S[378]), .CO(C[379]) );
  FA_5030 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n135), .CI(C[379]), .S(S[379]), .CO(C[380]) );
  FA_5029 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n134), .CI(C[380]), .S(S[380]), .CO(C[381]) );
  FA_5028 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n133), .CI(C[381]), .S(S[381]), .CO(C[382]) );
  FA_5027 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n132), .CI(C[382]), .S(S[382]), .CO(C[383]) );
  FA_5026 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n131), .CI(C[383]), .S(S[383]), .CO(C[384]) );
  FA_5025 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n130), .CI(C[384]), .S(S[384]), .CO(C[385]) );
  FA_5024 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n129), .CI(C[385]), .S(S[385]), .CO(C[386]) );
  FA_5023 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n128), .CI(C[386]), .S(S[386]), .CO(C[387]) );
  FA_5022 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n127), .CI(C[387]), .S(S[387]), .CO(C[388]) );
  FA_5021 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n126), .CI(C[388]), .S(S[388]), .CO(C[389]) );
  FA_5020 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n125), .CI(C[389]), .S(S[389]), .CO(C[390]) );
  FA_5019 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n124), .CI(C[390]), .S(S[390]), .CO(C[391]) );
  FA_5018 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n123), .CI(C[391]), .S(S[391]), .CO(C[392]) );
  FA_5017 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n122), .CI(C[392]), .S(S[392]), .CO(C[393]) );
  FA_5016 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n121), .CI(C[393]), .S(S[393]), .CO(C[394]) );
  FA_5015 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n120), .CI(C[394]), .S(S[394]), .CO(C[395]) );
  FA_5014 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n119), .CI(C[395]), .S(S[395]), .CO(C[396]) );
  FA_5013 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n118), .CI(C[396]), .S(S[396]), .CO(C[397]) );
  FA_5012 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n117), .CI(C[397]), .S(S[397]), .CO(C[398]) );
  FA_5011 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n116), .CI(C[398]), .S(S[398]), .CO(C[399]) );
  FA_5010 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n115), .CI(C[399]), .S(S[399]), .CO(C[400]) );
  FA_5009 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n114), .CI(C[400]), .S(S[400]), .CO(C[401]) );
  FA_5008 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n113), .CI(C[401]), .S(S[401]), .CO(C[402]) );
  FA_5007 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n112), .CI(C[402]), .S(S[402]), .CO(C[403]) );
  FA_5006 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n111), .CI(C[403]), .S(S[403]), .CO(C[404]) );
  FA_5005 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n110), .CI(C[404]), .S(S[404]), .CO(C[405]) );
  FA_5004 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n109), .CI(C[405]), .S(S[405]), .CO(C[406]) );
  FA_5003 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n108), .CI(C[406]), .S(S[406]), .CO(C[407]) );
  FA_5002 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n107), .CI(C[407]), .S(S[407]), .CO(C[408]) );
  FA_5001 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n106), .CI(C[408]), .S(S[408]), .CO(C[409]) );
  FA_5000 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n105), .CI(C[409]), .S(S[409]), .CO(C[410]) );
  FA_4999 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n104), .CI(C[410]), .S(S[410]), .CO(C[411]) );
  FA_4998 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n103), .CI(C[411]), .S(S[411]), .CO(C[412]) );
  FA_4997 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n102), .CI(C[412]), .S(S[412]), .CO(C[413]) );
  FA_4996 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n101), .CI(C[413]), .S(S[413]), .CO(C[414]) );
  FA_4995 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n100), .CI(C[414]), .S(S[414]), .CO(C[415]) );
  FA_4994 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n99), .CI(C[415]), 
        .S(S[415]), .CO(C[416]) );
  FA_4993 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n98), .CI(C[416]), 
        .S(S[416]), .CO(C[417]) );
  FA_4992 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n97), .CI(C[417]), 
        .S(S[417]), .CO(C[418]) );
  FA_4991 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n96), .CI(C[418]), 
        .S(S[418]), .CO(C[419]) );
  FA_4990 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n95), .CI(C[419]), 
        .S(S[419]), .CO(C[420]) );
  FA_4989 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n94), .CI(C[420]), 
        .S(S[420]), .CO(C[421]) );
  FA_4988 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n93), .CI(C[421]), 
        .S(S[421]), .CO(C[422]) );
  FA_4987 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n92), .CI(C[422]), 
        .S(S[422]), .CO(C[423]) );
  FA_4986 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n91), .CI(C[423]), 
        .S(S[423]), .CO(C[424]) );
  FA_4985 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n90), .CI(C[424]), 
        .S(S[424]), .CO(C[425]) );
  FA_4984 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n89), .CI(C[425]), 
        .S(S[425]), .CO(C[426]) );
  FA_4983 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n88), .CI(C[426]), 
        .S(S[426]), .CO(C[427]) );
  FA_4982 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n87), .CI(C[427]), 
        .S(S[427]), .CO(C[428]) );
  FA_4981 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n86), .CI(C[428]), 
        .S(S[428]), .CO(C[429]) );
  FA_4980 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n85), .CI(C[429]), 
        .S(S[429]), .CO(C[430]) );
  FA_4979 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n84), .CI(C[430]), 
        .S(S[430]), .CO(C[431]) );
  FA_4978 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n83), .CI(C[431]), 
        .S(S[431]), .CO(C[432]) );
  FA_4977 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n82), .CI(C[432]), 
        .S(S[432]), .CO(C[433]) );
  FA_4976 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n81), .CI(C[433]), 
        .S(S[433]), .CO(C[434]) );
  FA_4975 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n80), .CI(C[434]), 
        .S(S[434]), .CO(C[435]) );
  FA_4974 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n79), .CI(C[435]), 
        .S(S[435]), .CO(C[436]) );
  FA_4973 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n78), .CI(C[436]), 
        .S(S[436]), .CO(C[437]) );
  FA_4972 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n77), .CI(C[437]), 
        .S(S[437]), .CO(C[438]) );
  FA_4971 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n76), .CI(C[438]), 
        .S(S[438]), .CO(C[439]) );
  FA_4970 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n75), .CI(C[439]), 
        .S(S[439]), .CO(C[440]) );
  FA_4969 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n74), .CI(C[440]), 
        .S(S[440]), .CO(C[441]) );
  FA_4968 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n73), .CI(C[441]), 
        .S(S[441]), .CO(C[442]) );
  FA_4967 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n72), .CI(C[442]), 
        .S(S[442]), .CO(C[443]) );
  FA_4966 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n71), .CI(C[443]), 
        .S(S[443]), .CO(C[444]) );
  FA_4965 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n70), .CI(C[444]), 
        .S(S[444]), .CO(C[445]) );
  FA_4964 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n69), .CI(C[445]), 
        .S(S[445]), .CO(C[446]) );
  FA_4963 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n68), .CI(C[446]), 
        .S(S[446]), .CO(C[447]) );
  FA_4962 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n67), .CI(C[447]), 
        .S(S[447]), .CO(C[448]) );
  FA_4961 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n66), .CI(C[448]), 
        .S(S[448]), .CO(C[449]) );
  FA_4960 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n65), .CI(C[449]), 
        .S(S[449]), .CO(C[450]) );
  FA_4959 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n64), .CI(C[450]), 
        .S(S[450]), .CO(C[451]) );
  FA_4958 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n63), .CI(C[451]), 
        .S(S[451]), .CO(C[452]) );
  FA_4957 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n62), .CI(C[452]), 
        .S(S[452]), .CO(C[453]) );
  FA_4956 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n61), .CI(C[453]), 
        .S(S[453]), .CO(C[454]) );
  FA_4955 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n60), .CI(C[454]), 
        .S(S[454]), .CO(C[455]) );
  FA_4954 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n59), .CI(C[455]), 
        .S(S[455]), .CO(C[456]) );
  FA_4953 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n58), .CI(C[456]), 
        .S(S[456]), .CO(C[457]) );
  FA_4952 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n57), .CI(C[457]), 
        .S(S[457]), .CO(C[458]) );
  FA_4951 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n56), .CI(C[458]), 
        .S(S[458]), .CO(C[459]) );
  FA_4950 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n55), .CI(C[459]), 
        .S(S[459]), .CO(C[460]) );
  FA_4949 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n54), .CI(C[460]), 
        .S(S[460]), .CO(C[461]) );
  FA_4948 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n53), .CI(C[461]), 
        .S(S[461]), .CO(C[462]) );
  FA_4947 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n52), .CI(C[462]), 
        .S(S[462]), .CO(C[463]) );
  FA_4946 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n51), .CI(C[463]), 
        .S(S[463]), .CO(C[464]) );
  FA_4945 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n50), .CI(C[464]), 
        .S(S[464]), .CO(C[465]) );
  FA_4944 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n49), .CI(C[465]), 
        .S(S[465]), .CO(C[466]) );
  FA_4943 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n48), .CI(C[466]), 
        .S(S[466]), .CO(C[467]) );
  FA_4942 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n47), .CI(C[467]), 
        .S(S[467]), .CO(C[468]) );
  FA_4941 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n46), .CI(C[468]), 
        .S(S[468]), .CO(C[469]) );
  FA_4940 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n45), .CI(C[469]), 
        .S(S[469]), .CO(C[470]) );
  FA_4939 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n44), .CI(C[470]), 
        .S(S[470]), .CO(C[471]) );
  FA_4938 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n43), .CI(C[471]), 
        .S(S[471]), .CO(C[472]) );
  FA_4937 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n42), .CI(C[472]), 
        .S(S[472]), .CO(C[473]) );
  FA_4936 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n41), .CI(C[473]), 
        .S(S[473]), .CO(C[474]) );
  FA_4935 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n40), .CI(C[474]), 
        .S(S[474]), .CO(C[475]) );
  FA_4934 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n39), .CI(C[475]), 
        .S(S[475]), .CO(C[476]) );
  FA_4933 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n38), .CI(C[476]), 
        .S(S[476]), .CO(C[477]) );
  FA_4932 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n37), .CI(C[477]), 
        .S(S[477]), .CO(C[478]) );
  FA_4931 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n36), .CI(C[478]), 
        .S(S[478]), .CO(C[479]) );
  FA_4930 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n35), .CI(C[479]), 
        .S(S[479]), .CO(C[480]) );
  FA_4929 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n34), .CI(C[480]), 
        .S(S[480]), .CO(C[481]) );
  FA_4928 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n33), .CI(C[481]), 
        .S(S[481]), .CO(C[482]) );
  FA_4927 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n32), .CI(C[482]), 
        .S(S[482]), .CO(C[483]) );
  FA_4926 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n31), .CI(C[483]), 
        .S(S[483]), .CO(C[484]) );
  FA_4925 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n30), .CI(C[484]), 
        .S(S[484]), .CO(C[485]) );
  FA_4924 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n29), .CI(C[485]), 
        .S(S[485]), .CO(C[486]) );
  FA_4923 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n28), .CI(C[486]), 
        .S(S[486]), .CO(C[487]) );
  FA_4922 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n27), .CI(C[487]), 
        .S(S[487]), .CO(C[488]) );
  FA_4921 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n26), .CI(C[488]), 
        .S(S[488]), .CO(C[489]) );
  FA_4920 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n25), .CI(C[489]), 
        .S(S[489]), .CO(C[490]) );
  FA_4919 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n24), .CI(C[490]), 
        .S(S[490]), .CO(C[491]) );
  FA_4918 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n23), .CI(C[491]), 
        .S(S[491]), .CO(C[492]) );
  FA_4917 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n22), .CI(C[492]), 
        .S(S[492]), .CO(C[493]) );
  FA_4916 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n21), .CI(C[493]), 
        .S(S[493]), .CO(C[494]) );
  FA_4915 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n20), .CI(C[494]), 
        .S(S[494]), .CO(C[495]) );
  FA_4914 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n19), .CI(C[495]), 
        .S(S[495]), .CO(C[496]) );
  FA_4913 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n18), .CI(C[496]), 
        .S(S[496]), .CO(C[497]) );
  FA_4912 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n17), .CI(C[497]), 
        .S(S[497]), .CO(C[498]) );
  FA_4911 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n16), .CI(C[498]), 
        .S(S[498]), .CO(C[499]) );
  FA_4910 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n15), .CI(C[499]), 
        .S(S[499]), .CO(C[500]) );
  FA_4909 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n14), .CI(C[500]), 
        .S(S[500]), .CO(C[501]) );
  FA_4908 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n13), .CI(C[501]), 
        .S(S[501]), .CO(C[502]) );
  FA_4907 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n12), .CI(C[502]), 
        .S(S[502]), .CO(C[503]) );
  FA_4906 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n11), .CI(C[503]), 
        .S(S[503]), .CO(C[504]) );
  FA_4905 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n10), .CI(C[504]), 
        .S(S[504]), .CO(C[505]) );
  FA_4904 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n9), .CI(C[505]), 
        .S(S[505]), .CO(C[506]) );
  FA_4903 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n8), .CI(C[506]), 
        .S(S[506]), .CO(C[507]) );
  FA_4902 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n7), .CI(C[507]), 
        .S(S[507]), .CO(C[508]) );
  FA_4901 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n6), .CI(C[508]), 
        .S(S[508]), .CO(C[509]) );
  FA_4900 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n5), .CI(C[509]), 
        .S(S[509]), .CO(C[510]) );
  FA_4899 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n4), .CI(C[510]), 
        .S(S[510]), .CO(C[511]) );
  FA_4898 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n3), .CI(C[511]), 
        .S(S[511]), .CO(C[512]) );
  FA_4897 \FA_INST_1[512].FA_  ( .A(A[512]), .B(1'b1), .CI(C[512]), .S(S[512]), 
        .CO(C[513]) );
  FA_4896 \FA_INST_1[513].FA_  ( .A(A[513]), .B(1'b1), .CI(C[513]), .S(S[513])
         );
  IV U2 ( .A(B[415]), .Z(n99) );
  IV U3 ( .A(B[416]), .Z(n98) );
  IV U4 ( .A(B[417]), .Z(n97) );
  IV U5 ( .A(B[418]), .Z(n96) );
  IV U6 ( .A(B[419]), .Z(n95) );
  IV U7 ( .A(B[420]), .Z(n94) );
  IV U8 ( .A(B[421]), .Z(n93) );
  IV U9 ( .A(B[422]), .Z(n92) );
  IV U10 ( .A(B[423]), .Z(n91) );
  IV U11 ( .A(B[424]), .Z(n90) );
  IV U12 ( .A(B[505]), .Z(n9) );
  IV U13 ( .A(B[425]), .Z(n89) );
  IV U14 ( .A(B[426]), .Z(n88) );
  IV U15 ( .A(B[427]), .Z(n87) );
  IV U16 ( .A(B[428]), .Z(n86) );
  IV U17 ( .A(B[429]), .Z(n85) );
  IV U18 ( .A(B[430]), .Z(n84) );
  IV U19 ( .A(B[431]), .Z(n83) );
  IV U20 ( .A(B[432]), .Z(n82) );
  IV U21 ( .A(B[433]), .Z(n81) );
  IV U22 ( .A(B[434]), .Z(n80) );
  IV U23 ( .A(B[506]), .Z(n8) );
  IV U24 ( .A(B[435]), .Z(n79) );
  IV U25 ( .A(B[436]), .Z(n78) );
  IV U26 ( .A(B[437]), .Z(n77) );
  IV U27 ( .A(B[438]), .Z(n76) );
  IV U28 ( .A(B[439]), .Z(n75) );
  IV U29 ( .A(B[440]), .Z(n74) );
  IV U30 ( .A(B[441]), .Z(n73) );
  IV U31 ( .A(B[442]), .Z(n72) );
  IV U32 ( .A(B[443]), .Z(n71) );
  IV U33 ( .A(B[444]), .Z(n70) );
  IV U34 ( .A(B[507]), .Z(n7) );
  IV U35 ( .A(B[445]), .Z(n69) );
  IV U36 ( .A(B[446]), .Z(n68) );
  IV U37 ( .A(B[447]), .Z(n67) );
  IV U38 ( .A(B[448]), .Z(n66) );
  IV U39 ( .A(B[449]), .Z(n65) );
  IV U40 ( .A(B[450]), .Z(n64) );
  IV U41 ( .A(B[451]), .Z(n63) );
  IV U42 ( .A(B[452]), .Z(n62) );
  IV U43 ( .A(B[453]), .Z(n61) );
  IV U44 ( .A(B[454]), .Z(n60) );
  IV U45 ( .A(B[508]), .Z(n6) );
  IV U46 ( .A(B[455]), .Z(n59) );
  IV U47 ( .A(B[456]), .Z(n58) );
  IV U48 ( .A(B[457]), .Z(n57) );
  IV U49 ( .A(B[458]), .Z(n56) );
  IV U50 ( .A(B[459]), .Z(n55) );
  IV U51 ( .A(B[460]), .Z(n54) );
  IV U52 ( .A(B[461]), .Z(n53) );
  IV U53 ( .A(B[462]), .Z(n52) );
  IV U54 ( .A(B[0]), .Z(n514) );
  IV U55 ( .A(B[1]), .Z(n513) );
  IV U56 ( .A(B[2]), .Z(n512) );
  IV U57 ( .A(B[3]), .Z(n511) );
  IV U58 ( .A(B[4]), .Z(n510) );
  IV U59 ( .A(B[463]), .Z(n51) );
  IV U60 ( .A(B[5]), .Z(n509) );
  IV U61 ( .A(B[6]), .Z(n508) );
  IV U62 ( .A(B[7]), .Z(n507) );
  IV U63 ( .A(B[8]), .Z(n506) );
  IV U64 ( .A(B[9]), .Z(n505) );
  IV U65 ( .A(B[10]), .Z(n504) );
  IV U66 ( .A(B[11]), .Z(n503) );
  IV U67 ( .A(B[12]), .Z(n502) );
  IV U68 ( .A(B[13]), .Z(n501) );
  IV U69 ( .A(B[14]), .Z(n500) );
  IV U70 ( .A(B[464]), .Z(n50) );
  IV U71 ( .A(B[509]), .Z(n5) );
  IV U72 ( .A(B[15]), .Z(n499) );
  IV U73 ( .A(B[16]), .Z(n498) );
  IV U74 ( .A(B[17]), .Z(n497) );
  IV U75 ( .A(B[18]), .Z(n496) );
  IV U76 ( .A(B[19]), .Z(n495) );
  IV U77 ( .A(B[20]), .Z(n494) );
  IV U78 ( .A(B[21]), .Z(n493) );
  IV U79 ( .A(B[22]), .Z(n492) );
  IV U80 ( .A(B[23]), .Z(n491) );
  IV U81 ( .A(B[24]), .Z(n490) );
  IV U82 ( .A(B[465]), .Z(n49) );
  IV U83 ( .A(B[25]), .Z(n489) );
  IV U84 ( .A(B[26]), .Z(n488) );
  IV U85 ( .A(B[27]), .Z(n487) );
  IV U86 ( .A(B[28]), .Z(n486) );
  IV U87 ( .A(B[29]), .Z(n485) );
  IV U88 ( .A(B[30]), .Z(n484) );
  IV U89 ( .A(B[31]), .Z(n483) );
  IV U90 ( .A(B[32]), .Z(n482) );
  IV U91 ( .A(B[33]), .Z(n481) );
  IV U92 ( .A(B[34]), .Z(n480) );
  IV U93 ( .A(B[466]), .Z(n48) );
  IV U94 ( .A(B[35]), .Z(n479) );
  IV U95 ( .A(B[36]), .Z(n478) );
  IV U96 ( .A(B[37]), .Z(n477) );
  IV U97 ( .A(B[38]), .Z(n476) );
  IV U98 ( .A(B[39]), .Z(n475) );
  IV U99 ( .A(B[40]), .Z(n474) );
  IV U100 ( .A(B[41]), .Z(n473) );
  IV U101 ( .A(B[42]), .Z(n472) );
  IV U102 ( .A(B[43]), .Z(n471) );
  IV U103 ( .A(B[44]), .Z(n470) );
  IV U104 ( .A(B[467]), .Z(n47) );
  IV U105 ( .A(B[45]), .Z(n469) );
  IV U106 ( .A(B[46]), .Z(n468) );
  IV U107 ( .A(B[47]), .Z(n467) );
  IV U108 ( .A(B[48]), .Z(n466) );
  IV U109 ( .A(B[49]), .Z(n465) );
  IV U110 ( .A(B[50]), .Z(n464) );
  IV U111 ( .A(B[51]), .Z(n463) );
  IV U112 ( .A(B[52]), .Z(n462) );
  IV U113 ( .A(B[53]), .Z(n461) );
  IV U114 ( .A(B[54]), .Z(n460) );
  IV U115 ( .A(B[468]), .Z(n46) );
  IV U116 ( .A(B[55]), .Z(n459) );
  IV U117 ( .A(B[56]), .Z(n458) );
  IV U118 ( .A(B[57]), .Z(n457) );
  IV U119 ( .A(B[58]), .Z(n456) );
  IV U120 ( .A(B[59]), .Z(n455) );
  IV U121 ( .A(B[60]), .Z(n454) );
  IV U122 ( .A(B[61]), .Z(n453) );
  IV U123 ( .A(B[62]), .Z(n452) );
  IV U124 ( .A(B[63]), .Z(n451) );
  IV U125 ( .A(B[64]), .Z(n450) );
  IV U126 ( .A(B[469]), .Z(n45) );
  IV U127 ( .A(B[65]), .Z(n449) );
  IV U128 ( .A(B[66]), .Z(n448) );
  IV U129 ( .A(B[67]), .Z(n447) );
  IV U130 ( .A(B[68]), .Z(n446) );
  IV U131 ( .A(B[69]), .Z(n445) );
  IV U132 ( .A(B[70]), .Z(n444) );
  IV U133 ( .A(B[71]), .Z(n443) );
  IV U134 ( .A(B[72]), .Z(n442) );
  IV U135 ( .A(B[73]), .Z(n441) );
  IV U136 ( .A(B[74]), .Z(n440) );
  IV U137 ( .A(B[470]), .Z(n44) );
  IV U138 ( .A(B[75]), .Z(n439) );
  IV U139 ( .A(B[76]), .Z(n438) );
  IV U140 ( .A(B[77]), .Z(n437) );
  IV U141 ( .A(B[78]), .Z(n436) );
  IV U142 ( .A(B[79]), .Z(n435) );
  IV U143 ( .A(B[80]), .Z(n434) );
  IV U144 ( .A(B[81]), .Z(n433) );
  IV U145 ( .A(B[82]), .Z(n432) );
  IV U146 ( .A(B[83]), .Z(n431) );
  IV U147 ( .A(B[84]), .Z(n430) );
  IV U148 ( .A(B[471]), .Z(n43) );
  IV U149 ( .A(B[85]), .Z(n429) );
  IV U150 ( .A(B[86]), .Z(n428) );
  IV U151 ( .A(B[87]), .Z(n427) );
  IV U152 ( .A(B[88]), .Z(n426) );
  IV U153 ( .A(B[89]), .Z(n425) );
  IV U154 ( .A(B[90]), .Z(n424) );
  IV U155 ( .A(B[91]), .Z(n423) );
  IV U156 ( .A(B[92]), .Z(n422) );
  IV U157 ( .A(B[93]), .Z(n421) );
  IV U158 ( .A(B[94]), .Z(n420) );
  IV U159 ( .A(B[472]), .Z(n42) );
  IV U160 ( .A(B[95]), .Z(n419) );
  IV U161 ( .A(B[96]), .Z(n418) );
  IV U162 ( .A(B[97]), .Z(n417) );
  IV U163 ( .A(B[98]), .Z(n416) );
  IV U164 ( .A(B[99]), .Z(n415) );
  IV U165 ( .A(B[100]), .Z(n414) );
  IV U166 ( .A(B[101]), .Z(n413) );
  IV U167 ( .A(B[102]), .Z(n412) );
  IV U168 ( .A(B[103]), .Z(n411) );
  IV U169 ( .A(B[104]), .Z(n410) );
  IV U170 ( .A(B[473]), .Z(n41) );
  IV U171 ( .A(B[105]), .Z(n409) );
  IV U172 ( .A(B[106]), .Z(n408) );
  IV U173 ( .A(B[107]), .Z(n407) );
  IV U174 ( .A(B[108]), .Z(n406) );
  IV U175 ( .A(B[109]), .Z(n405) );
  IV U176 ( .A(B[110]), .Z(n404) );
  IV U177 ( .A(B[111]), .Z(n403) );
  IV U178 ( .A(B[112]), .Z(n402) );
  IV U179 ( .A(B[113]), .Z(n401) );
  IV U180 ( .A(B[114]), .Z(n400) );
  IV U181 ( .A(B[474]), .Z(n40) );
  IV U182 ( .A(B[510]), .Z(n4) );
  IV U183 ( .A(B[115]), .Z(n399) );
  IV U184 ( .A(B[116]), .Z(n398) );
  IV U185 ( .A(B[117]), .Z(n397) );
  IV U186 ( .A(B[118]), .Z(n396) );
  IV U187 ( .A(B[119]), .Z(n395) );
  IV U188 ( .A(B[120]), .Z(n394) );
  IV U189 ( .A(B[121]), .Z(n393) );
  IV U190 ( .A(B[122]), .Z(n392) );
  IV U191 ( .A(B[123]), .Z(n391) );
  IV U192 ( .A(B[124]), .Z(n390) );
  IV U193 ( .A(B[475]), .Z(n39) );
  IV U194 ( .A(B[125]), .Z(n389) );
  IV U195 ( .A(B[126]), .Z(n388) );
  IV U196 ( .A(B[127]), .Z(n387) );
  IV U197 ( .A(B[128]), .Z(n386) );
  IV U198 ( .A(B[129]), .Z(n385) );
  IV U199 ( .A(B[130]), .Z(n384) );
  IV U200 ( .A(B[131]), .Z(n383) );
  IV U201 ( .A(B[132]), .Z(n382) );
  IV U202 ( .A(B[133]), .Z(n381) );
  IV U203 ( .A(B[134]), .Z(n380) );
  IV U204 ( .A(B[476]), .Z(n38) );
  IV U205 ( .A(B[135]), .Z(n379) );
  IV U206 ( .A(B[136]), .Z(n378) );
  IV U207 ( .A(B[137]), .Z(n377) );
  IV U208 ( .A(B[138]), .Z(n376) );
  IV U209 ( .A(B[139]), .Z(n375) );
  IV U210 ( .A(B[140]), .Z(n374) );
  IV U211 ( .A(B[141]), .Z(n373) );
  IV U212 ( .A(B[142]), .Z(n372) );
  IV U213 ( .A(B[143]), .Z(n371) );
  IV U214 ( .A(B[144]), .Z(n370) );
  IV U215 ( .A(B[477]), .Z(n37) );
  IV U216 ( .A(B[145]), .Z(n369) );
  IV U217 ( .A(B[146]), .Z(n368) );
  IV U218 ( .A(B[147]), .Z(n367) );
  IV U219 ( .A(B[148]), .Z(n366) );
  IV U220 ( .A(B[149]), .Z(n365) );
  IV U221 ( .A(B[150]), .Z(n364) );
  IV U222 ( .A(B[151]), .Z(n363) );
  IV U223 ( .A(B[152]), .Z(n362) );
  IV U224 ( .A(B[153]), .Z(n361) );
  IV U225 ( .A(B[154]), .Z(n360) );
  IV U226 ( .A(B[478]), .Z(n36) );
  IV U227 ( .A(B[155]), .Z(n359) );
  IV U228 ( .A(B[156]), .Z(n358) );
  IV U229 ( .A(B[157]), .Z(n357) );
  IV U230 ( .A(B[158]), .Z(n356) );
  IV U231 ( .A(B[159]), .Z(n355) );
  IV U232 ( .A(B[160]), .Z(n354) );
  IV U233 ( .A(B[161]), .Z(n353) );
  IV U234 ( .A(B[162]), .Z(n352) );
  IV U235 ( .A(B[163]), .Z(n351) );
  IV U236 ( .A(B[164]), .Z(n350) );
  IV U237 ( .A(B[479]), .Z(n35) );
  IV U238 ( .A(B[165]), .Z(n349) );
  IV U239 ( .A(B[166]), .Z(n348) );
  IV U240 ( .A(B[167]), .Z(n347) );
  IV U241 ( .A(B[168]), .Z(n346) );
  IV U242 ( .A(B[169]), .Z(n345) );
  IV U243 ( .A(B[170]), .Z(n344) );
  IV U244 ( .A(B[171]), .Z(n343) );
  IV U245 ( .A(B[172]), .Z(n342) );
  IV U246 ( .A(B[173]), .Z(n341) );
  IV U247 ( .A(B[174]), .Z(n340) );
  IV U248 ( .A(B[480]), .Z(n34) );
  IV U249 ( .A(B[175]), .Z(n339) );
  IV U250 ( .A(B[176]), .Z(n338) );
  IV U251 ( .A(B[177]), .Z(n337) );
  IV U252 ( .A(B[178]), .Z(n336) );
  IV U253 ( .A(B[179]), .Z(n335) );
  IV U254 ( .A(B[180]), .Z(n334) );
  IV U255 ( .A(B[181]), .Z(n333) );
  IV U256 ( .A(B[182]), .Z(n332) );
  IV U257 ( .A(B[183]), .Z(n331) );
  IV U258 ( .A(B[184]), .Z(n330) );
  IV U259 ( .A(B[481]), .Z(n33) );
  IV U260 ( .A(B[185]), .Z(n329) );
  IV U261 ( .A(B[186]), .Z(n328) );
  IV U262 ( .A(B[187]), .Z(n327) );
  IV U263 ( .A(B[188]), .Z(n326) );
  IV U264 ( .A(B[189]), .Z(n325) );
  IV U265 ( .A(B[190]), .Z(n324) );
  IV U266 ( .A(B[191]), .Z(n323) );
  IV U267 ( .A(B[192]), .Z(n322) );
  IV U268 ( .A(B[193]), .Z(n321) );
  IV U269 ( .A(B[194]), .Z(n320) );
  IV U270 ( .A(B[482]), .Z(n32) );
  IV U271 ( .A(B[195]), .Z(n319) );
  IV U272 ( .A(B[196]), .Z(n318) );
  IV U273 ( .A(B[197]), .Z(n317) );
  IV U274 ( .A(B[198]), .Z(n316) );
  IV U275 ( .A(B[199]), .Z(n315) );
  IV U276 ( .A(B[200]), .Z(n314) );
  IV U277 ( .A(B[201]), .Z(n313) );
  IV U278 ( .A(B[202]), .Z(n312) );
  IV U279 ( .A(B[203]), .Z(n311) );
  IV U280 ( .A(B[204]), .Z(n310) );
  IV U281 ( .A(B[483]), .Z(n31) );
  IV U282 ( .A(B[205]), .Z(n309) );
  IV U283 ( .A(B[206]), .Z(n308) );
  IV U284 ( .A(B[207]), .Z(n307) );
  IV U285 ( .A(B[208]), .Z(n306) );
  IV U286 ( .A(B[209]), .Z(n305) );
  IV U287 ( .A(B[210]), .Z(n304) );
  IV U288 ( .A(B[211]), .Z(n303) );
  IV U289 ( .A(B[212]), .Z(n302) );
  IV U290 ( .A(B[213]), .Z(n301) );
  IV U291 ( .A(B[214]), .Z(n300) );
  IV U292 ( .A(B[484]), .Z(n30) );
  IV U293 ( .A(B[511]), .Z(n3) );
  IV U294 ( .A(B[215]), .Z(n299) );
  IV U295 ( .A(B[216]), .Z(n298) );
  IV U296 ( .A(B[217]), .Z(n297) );
  IV U297 ( .A(B[218]), .Z(n296) );
  IV U298 ( .A(B[219]), .Z(n295) );
  IV U299 ( .A(B[220]), .Z(n294) );
  IV U300 ( .A(B[221]), .Z(n293) );
  IV U301 ( .A(B[222]), .Z(n292) );
  IV U302 ( .A(B[223]), .Z(n291) );
  IV U303 ( .A(B[224]), .Z(n290) );
  IV U304 ( .A(B[485]), .Z(n29) );
  IV U305 ( .A(B[225]), .Z(n289) );
  IV U306 ( .A(B[226]), .Z(n288) );
  IV U307 ( .A(B[227]), .Z(n287) );
  IV U308 ( .A(B[228]), .Z(n286) );
  IV U309 ( .A(B[229]), .Z(n285) );
  IV U310 ( .A(B[230]), .Z(n284) );
  IV U311 ( .A(B[231]), .Z(n283) );
  IV U312 ( .A(B[232]), .Z(n282) );
  IV U313 ( .A(B[233]), .Z(n281) );
  IV U314 ( .A(B[234]), .Z(n280) );
  IV U315 ( .A(B[486]), .Z(n28) );
  IV U316 ( .A(B[235]), .Z(n279) );
  IV U317 ( .A(B[236]), .Z(n278) );
  IV U318 ( .A(B[237]), .Z(n277) );
  IV U319 ( .A(B[238]), .Z(n276) );
  IV U320 ( .A(B[239]), .Z(n275) );
  IV U321 ( .A(B[240]), .Z(n274) );
  IV U322 ( .A(B[241]), .Z(n273) );
  IV U323 ( .A(B[242]), .Z(n272) );
  IV U324 ( .A(B[243]), .Z(n271) );
  IV U325 ( .A(B[244]), .Z(n270) );
  IV U326 ( .A(B[487]), .Z(n27) );
  IV U327 ( .A(B[245]), .Z(n269) );
  IV U328 ( .A(B[246]), .Z(n268) );
  IV U329 ( .A(B[247]), .Z(n267) );
  IV U330 ( .A(B[248]), .Z(n266) );
  IV U331 ( .A(B[249]), .Z(n265) );
  IV U332 ( .A(B[250]), .Z(n264) );
  IV U333 ( .A(B[251]), .Z(n263) );
  IV U334 ( .A(B[252]), .Z(n262) );
  IV U335 ( .A(B[253]), .Z(n261) );
  IV U336 ( .A(B[254]), .Z(n260) );
  IV U337 ( .A(B[488]), .Z(n26) );
  IV U338 ( .A(B[255]), .Z(n259) );
  IV U339 ( .A(B[256]), .Z(n258) );
  IV U340 ( .A(B[257]), .Z(n257) );
  IV U341 ( .A(B[258]), .Z(n256) );
  IV U342 ( .A(B[259]), .Z(n255) );
  IV U343 ( .A(B[260]), .Z(n254) );
  IV U344 ( .A(B[261]), .Z(n253) );
  IV U345 ( .A(B[262]), .Z(n252) );
  IV U346 ( .A(B[263]), .Z(n251) );
  IV U347 ( .A(B[264]), .Z(n250) );
  IV U348 ( .A(B[489]), .Z(n25) );
  IV U349 ( .A(B[265]), .Z(n249) );
  IV U350 ( .A(B[266]), .Z(n248) );
  IV U351 ( .A(B[267]), .Z(n247) );
  IV U352 ( .A(B[268]), .Z(n246) );
  IV U353 ( .A(B[269]), .Z(n245) );
  IV U354 ( .A(B[270]), .Z(n244) );
  IV U355 ( .A(B[271]), .Z(n243) );
  IV U356 ( .A(B[272]), .Z(n242) );
  IV U357 ( .A(B[273]), .Z(n241) );
  IV U358 ( .A(B[274]), .Z(n240) );
  IV U359 ( .A(B[490]), .Z(n24) );
  IV U360 ( .A(B[275]), .Z(n239) );
  IV U361 ( .A(B[276]), .Z(n238) );
  IV U362 ( .A(B[277]), .Z(n237) );
  IV U363 ( .A(B[278]), .Z(n236) );
  IV U364 ( .A(B[279]), .Z(n235) );
  IV U365 ( .A(B[280]), .Z(n234) );
  IV U366 ( .A(B[281]), .Z(n233) );
  IV U367 ( .A(B[282]), .Z(n232) );
  IV U368 ( .A(B[283]), .Z(n231) );
  IV U369 ( .A(B[284]), .Z(n230) );
  IV U370 ( .A(B[491]), .Z(n23) );
  IV U371 ( .A(B[285]), .Z(n229) );
  IV U372 ( .A(B[286]), .Z(n228) );
  IV U373 ( .A(B[287]), .Z(n227) );
  IV U374 ( .A(B[288]), .Z(n226) );
  IV U375 ( .A(B[289]), .Z(n225) );
  IV U376 ( .A(B[290]), .Z(n224) );
  IV U377 ( .A(B[291]), .Z(n223) );
  IV U378 ( .A(B[292]), .Z(n222) );
  IV U379 ( .A(B[293]), .Z(n221) );
  IV U380 ( .A(B[294]), .Z(n220) );
  IV U381 ( .A(B[492]), .Z(n22) );
  IV U382 ( .A(B[295]), .Z(n219) );
  IV U383 ( .A(B[296]), .Z(n218) );
  IV U384 ( .A(B[297]), .Z(n217) );
  IV U385 ( .A(B[298]), .Z(n216) );
  IV U386 ( .A(B[299]), .Z(n215) );
  IV U387 ( .A(B[300]), .Z(n214) );
  IV U388 ( .A(B[301]), .Z(n213) );
  IV U389 ( .A(B[302]), .Z(n212) );
  IV U390 ( .A(B[303]), .Z(n211) );
  IV U391 ( .A(B[304]), .Z(n210) );
  IV U392 ( .A(B[493]), .Z(n21) );
  IV U393 ( .A(B[305]), .Z(n209) );
  IV U394 ( .A(B[306]), .Z(n208) );
  IV U395 ( .A(B[307]), .Z(n207) );
  IV U396 ( .A(B[308]), .Z(n206) );
  IV U397 ( .A(B[309]), .Z(n205) );
  IV U398 ( .A(B[310]), .Z(n204) );
  IV U399 ( .A(B[311]), .Z(n203) );
  IV U400 ( .A(B[312]), .Z(n202) );
  IV U401 ( .A(B[313]), .Z(n201) );
  IV U402 ( .A(B[314]), .Z(n200) );
  IV U403 ( .A(B[494]), .Z(n20) );
  IV U404 ( .A(B[315]), .Z(n199) );
  IV U405 ( .A(B[316]), .Z(n198) );
  IV U406 ( .A(B[317]), .Z(n197) );
  IV U407 ( .A(B[318]), .Z(n196) );
  IV U408 ( .A(B[319]), .Z(n195) );
  IV U409 ( .A(B[320]), .Z(n194) );
  IV U410 ( .A(B[321]), .Z(n193) );
  IV U411 ( .A(B[322]), .Z(n192) );
  IV U412 ( .A(B[323]), .Z(n191) );
  IV U413 ( .A(B[324]), .Z(n190) );
  IV U414 ( .A(B[495]), .Z(n19) );
  IV U415 ( .A(B[325]), .Z(n189) );
  IV U416 ( .A(B[326]), .Z(n188) );
  IV U417 ( .A(B[327]), .Z(n187) );
  IV U418 ( .A(B[328]), .Z(n186) );
  IV U419 ( .A(B[329]), .Z(n185) );
  IV U420 ( .A(B[330]), .Z(n184) );
  IV U421 ( .A(B[331]), .Z(n183) );
  IV U422 ( .A(B[332]), .Z(n182) );
  IV U423 ( .A(B[333]), .Z(n181) );
  IV U424 ( .A(B[334]), .Z(n180) );
  IV U425 ( .A(B[496]), .Z(n18) );
  IV U426 ( .A(B[335]), .Z(n179) );
  IV U427 ( .A(B[336]), .Z(n178) );
  IV U428 ( .A(B[337]), .Z(n177) );
  IV U429 ( .A(B[338]), .Z(n176) );
  IV U430 ( .A(B[339]), .Z(n175) );
  IV U431 ( .A(B[340]), .Z(n174) );
  IV U432 ( .A(B[341]), .Z(n173) );
  IV U433 ( .A(B[342]), .Z(n172) );
  IV U434 ( .A(B[343]), .Z(n171) );
  IV U435 ( .A(B[344]), .Z(n170) );
  IV U436 ( .A(B[497]), .Z(n17) );
  IV U437 ( .A(B[345]), .Z(n169) );
  IV U438 ( .A(B[346]), .Z(n168) );
  IV U439 ( .A(B[347]), .Z(n167) );
  IV U440 ( .A(B[348]), .Z(n166) );
  IV U441 ( .A(B[349]), .Z(n165) );
  IV U442 ( .A(B[350]), .Z(n164) );
  IV U443 ( .A(B[351]), .Z(n163) );
  IV U444 ( .A(B[352]), .Z(n162) );
  IV U445 ( .A(B[353]), .Z(n161) );
  IV U446 ( .A(B[354]), .Z(n160) );
  IV U447 ( .A(B[498]), .Z(n16) );
  IV U448 ( .A(B[355]), .Z(n159) );
  IV U449 ( .A(B[356]), .Z(n158) );
  IV U450 ( .A(B[357]), .Z(n157) );
  IV U451 ( .A(B[358]), .Z(n156) );
  IV U452 ( .A(B[359]), .Z(n155) );
  IV U453 ( .A(B[360]), .Z(n154) );
  IV U454 ( .A(B[361]), .Z(n153) );
  IV U455 ( .A(B[362]), .Z(n152) );
  IV U456 ( .A(B[363]), .Z(n151) );
  IV U457 ( .A(B[364]), .Z(n150) );
  IV U458 ( .A(B[499]), .Z(n15) );
  IV U459 ( .A(B[365]), .Z(n149) );
  IV U460 ( .A(B[366]), .Z(n148) );
  IV U461 ( .A(B[367]), .Z(n147) );
  IV U462 ( .A(B[368]), .Z(n146) );
  IV U463 ( .A(B[369]), .Z(n145) );
  IV U464 ( .A(B[370]), .Z(n144) );
  IV U465 ( .A(B[371]), .Z(n143) );
  IV U466 ( .A(B[372]), .Z(n142) );
  IV U467 ( .A(B[373]), .Z(n141) );
  IV U468 ( .A(B[374]), .Z(n140) );
  IV U469 ( .A(B[500]), .Z(n14) );
  IV U470 ( .A(B[375]), .Z(n139) );
  IV U471 ( .A(B[376]), .Z(n138) );
  IV U472 ( .A(B[377]), .Z(n137) );
  IV U473 ( .A(B[378]), .Z(n136) );
  IV U474 ( .A(B[379]), .Z(n135) );
  IV U475 ( .A(B[380]), .Z(n134) );
  IV U476 ( .A(B[381]), .Z(n133) );
  IV U477 ( .A(B[382]), .Z(n132) );
  IV U478 ( .A(B[383]), .Z(n131) );
  IV U479 ( .A(B[384]), .Z(n130) );
  IV U480 ( .A(B[501]), .Z(n13) );
  IV U481 ( .A(B[385]), .Z(n129) );
  IV U482 ( .A(B[386]), .Z(n128) );
  IV U483 ( .A(B[387]), .Z(n127) );
  IV U484 ( .A(B[388]), .Z(n126) );
  IV U485 ( .A(B[389]), .Z(n125) );
  IV U486 ( .A(B[390]), .Z(n124) );
  IV U487 ( .A(B[391]), .Z(n123) );
  IV U488 ( .A(B[392]), .Z(n122) );
  IV U489 ( .A(B[393]), .Z(n121) );
  IV U490 ( .A(B[394]), .Z(n120) );
  IV U491 ( .A(B[502]), .Z(n12) );
  IV U492 ( .A(B[395]), .Z(n119) );
  IV U493 ( .A(B[396]), .Z(n118) );
  IV U494 ( .A(B[397]), .Z(n117) );
  IV U495 ( .A(B[398]), .Z(n116) );
  IV U496 ( .A(B[399]), .Z(n115) );
  IV U497 ( .A(B[400]), .Z(n114) );
  IV U498 ( .A(B[401]), .Z(n113) );
  IV U499 ( .A(B[402]), .Z(n112) );
  IV U500 ( .A(B[403]), .Z(n111) );
  IV U501 ( .A(B[404]), .Z(n110) );
  IV U502 ( .A(B[503]), .Z(n11) );
  IV U503 ( .A(B[405]), .Z(n109) );
  IV U504 ( .A(B[406]), .Z(n108) );
  IV U505 ( .A(B[407]), .Z(n107) );
  IV U506 ( .A(B[408]), .Z(n106) );
  IV U507 ( .A(B[409]), .Z(n105) );
  IV U508 ( .A(B[410]), .Z(n104) );
  IV U509 ( .A(B[411]), .Z(n103) );
  IV U510 ( .A(B[412]), .Z(n102) );
  IV U511 ( .A(B[413]), .Z(n101) );
  IV U512 ( .A(B[414]), .Z(n100) );
  IV U513 ( .A(B[504]), .Z(n10) );
endmodule


module MUX_N514_1 ( A, B, S, O );
  input [513:0] A;
  input [513:0] B;
  output [513:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[511]), .A(S), .Z(O[511]) );
  ANDN U56 ( .B(A[510]), .A(S), .Z(O[510]) );
  ANDN U57 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U58 ( .B(A[509]), .A(S), .Z(O[509]) );
  ANDN U59 ( .B(A[508]), .A(S), .Z(O[508]) );
  ANDN U60 ( .B(A[507]), .A(S), .Z(O[507]) );
  ANDN U61 ( .B(A[506]), .A(S), .Z(O[506]) );
  ANDN U62 ( .B(A[505]), .A(S), .Z(O[505]) );
  ANDN U63 ( .B(A[504]), .A(S), .Z(O[504]) );
  ANDN U64 ( .B(A[503]), .A(S), .Z(O[503]) );
  ANDN U65 ( .B(A[502]), .A(S), .Z(O[502]) );
  ANDN U66 ( .B(A[501]), .A(S), .Z(O[501]) );
  ANDN U67 ( .B(A[500]), .A(S), .Z(O[500]) );
  ANDN U68 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U69 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U70 ( .B(A[499]), .A(S), .Z(O[499]) );
  ANDN U71 ( .B(A[498]), .A(S), .Z(O[498]) );
  ANDN U72 ( .B(A[497]), .A(S), .Z(O[497]) );
  ANDN U73 ( .B(A[496]), .A(S), .Z(O[496]) );
  ANDN U74 ( .B(A[495]), .A(S), .Z(O[495]) );
  ANDN U75 ( .B(A[494]), .A(S), .Z(O[494]) );
  ANDN U76 ( .B(A[493]), .A(S), .Z(O[493]) );
  ANDN U77 ( .B(A[492]), .A(S), .Z(O[492]) );
  ANDN U78 ( .B(A[491]), .A(S), .Z(O[491]) );
  ANDN U79 ( .B(A[490]), .A(S), .Z(O[490]) );
  ANDN U80 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U81 ( .B(A[489]), .A(S), .Z(O[489]) );
  ANDN U82 ( .B(A[488]), .A(S), .Z(O[488]) );
  ANDN U83 ( .B(A[487]), .A(S), .Z(O[487]) );
  ANDN U84 ( .B(A[486]), .A(S), .Z(O[486]) );
  ANDN U85 ( .B(A[485]), .A(S), .Z(O[485]) );
  ANDN U86 ( .B(A[484]), .A(S), .Z(O[484]) );
  ANDN U87 ( .B(A[483]), .A(S), .Z(O[483]) );
  ANDN U88 ( .B(A[482]), .A(S), .Z(O[482]) );
  ANDN U89 ( .B(A[481]), .A(S), .Z(O[481]) );
  ANDN U90 ( .B(A[480]), .A(S), .Z(O[480]) );
  ANDN U91 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U92 ( .B(A[479]), .A(S), .Z(O[479]) );
  ANDN U93 ( .B(A[478]), .A(S), .Z(O[478]) );
  ANDN U94 ( .B(A[477]), .A(S), .Z(O[477]) );
  ANDN U95 ( .B(A[476]), .A(S), .Z(O[476]) );
  ANDN U96 ( .B(A[475]), .A(S), .Z(O[475]) );
  ANDN U97 ( .B(A[474]), .A(S), .Z(O[474]) );
  ANDN U98 ( .B(A[473]), .A(S), .Z(O[473]) );
  ANDN U99 ( .B(A[472]), .A(S), .Z(O[472]) );
  ANDN U100 ( .B(A[471]), .A(S), .Z(O[471]) );
  ANDN U101 ( .B(A[470]), .A(S), .Z(O[470]) );
  ANDN U102 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U103 ( .B(A[469]), .A(S), .Z(O[469]) );
  ANDN U104 ( .B(A[468]), .A(S), .Z(O[468]) );
  ANDN U105 ( .B(A[467]), .A(S), .Z(O[467]) );
  ANDN U106 ( .B(A[466]), .A(S), .Z(O[466]) );
  ANDN U107 ( .B(A[465]), .A(S), .Z(O[465]) );
  ANDN U108 ( .B(A[464]), .A(S), .Z(O[464]) );
  ANDN U109 ( .B(A[463]), .A(S), .Z(O[463]) );
  ANDN U110 ( .B(A[462]), .A(S), .Z(O[462]) );
  ANDN U111 ( .B(A[461]), .A(S), .Z(O[461]) );
  ANDN U112 ( .B(A[460]), .A(S), .Z(O[460]) );
  ANDN U113 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U114 ( .B(A[459]), .A(S), .Z(O[459]) );
  ANDN U115 ( .B(A[458]), .A(S), .Z(O[458]) );
  ANDN U116 ( .B(A[457]), .A(S), .Z(O[457]) );
  ANDN U117 ( .B(A[456]), .A(S), .Z(O[456]) );
  ANDN U118 ( .B(A[455]), .A(S), .Z(O[455]) );
  ANDN U119 ( .B(A[454]), .A(S), .Z(O[454]) );
  ANDN U120 ( .B(A[453]), .A(S), .Z(O[453]) );
  ANDN U121 ( .B(A[452]), .A(S), .Z(O[452]) );
  ANDN U122 ( .B(A[451]), .A(S), .Z(O[451]) );
  ANDN U123 ( .B(A[450]), .A(S), .Z(O[450]) );
  ANDN U124 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U125 ( .B(A[449]), .A(S), .Z(O[449]) );
  ANDN U126 ( .B(A[448]), .A(S), .Z(O[448]) );
  ANDN U127 ( .B(A[447]), .A(S), .Z(O[447]) );
  ANDN U128 ( .B(A[446]), .A(S), .Z(O[446]) );
  ANDN U129 ( .B(A[445]), .A(S), .Z(O[445]) );
  ANDN U130 ( .B(A[444]), .A(S), .Z(O[444]) );
  ANDN U131 ( .B(A[443]), .A(S), .Z(O[443]) );
  ANDN U132 ( .B(A[442]), .A(S), .Z(O[442]) );
  ANDN U133 ( .B(A[441]), .A(S), .Z(O[441]) );
  ANDN U134 ( .B(A[440]), .A(S), .Z(O[440]) );
  ANDN U135 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U136 ( .B(A[439]), .A(S), .Z(O[439]) );
  ANDN U137 ( .B(A[438]), .A(S), .Z(O[438]) );
  ANDN U138 ( .B(A[437]), .A(S), .Z(O[437]) );
  ANDN U139 ( .B(A[436]), .A(S), .Z(O[436]) );
  ANDN U140 ( .B(A[435]), .A(S), .Z(O[435]) );
  ANDN U141 ( .B(A[434]), .A(S), .Z(O[434]) );
  ANDN U142 ( .B(A[433]), .A(S), .Z(O[433]) );
  ANDN U143 ( .B(A[432]), .A(S), .Z(O[432]) );
  ANDN U144 ( .B(A[431]), .A(S), .Z(O[431]) );
  ANDN U145 ( .B(A[430]), .A(S), .Z(O[430]) );
  ANDN U146 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U147 ( .B(A[429]), .A(S), .Z(O[429]) );
  ANDN U148 ( .B(A[428]), .A(S), .Z(O[428]) );
  ANDN U149 ( .B(A[427]), .A(S), .Z(O[427]) );
  ANDN U150 ( .B(A[426]), .A(S), .Z(O[426]) );
  ANDN U151 ( .B(A[425]), .A(S), .Z(O[425]) );
  ANDN U152 ( .B(A[424]), .A(S), .Z(O[424]) );
  ANDN U153 ( .B(A[423]), .A(S), .Z(O[423]) );
  ANDN U154 ( .B(A[422]), .A(S), .Z(O[422]) );
  ANDN U155 ( .B(A[421]), .A(S), .Z(O[421]) );
  ANDN U156 ( .B(A[420]), .A(S), .Z(O[420]) );
  ANDN U157 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U158 ( .B(A[419]), .A(S), .Z(O[419]) );
  ANDN U159 ( .B(A[418]), .A(S), .Z(O[418]) );
  ANDN U160 ( .B(A[417]), .A(S), .Z(O[417]) );
  ANDN U161 ( .B(A[416]), .A(S), .Z(O[416]) );
  ANDN U162 ( .B(A[415]), .A(S), .Z(O[415]) );
  ANDN U163 ( .B(A[414]), .A(S), .Z(O[414]) );
  ANDN U164 ( .B(A[413]), .A(S), .Z(O[413]) );
  ANDN U165 ( .B(A[412]), .A(S), .Z(O[412]) );
  ANDN U166 ( .B(A[411]), .A(S), .Z(O[411]) );
  ANDN U167 ( .B(A[410]), .A(S), .Z(O[410]) );
  ANDN U168 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U169 ( .B(A[409]), .A(S), .Z(O[409]) );
  ANDN U170 ( .B(A[408]), .A(S), .Z(O[408]) );
  ANDN U171 ( .B(A[407]), .A(S), .Z(O[407]) );
  ANDN U172 ( .B(A[406]), .A(S), .Z(O[406]) );
  ANDN U173 ( .B(A[405]), .A(S), .Z(O[405]) );
  ANDN U174 ( .B(A[404]), .A(S), .Z(O[404]) );
  ANDN U175 ( .B(A[403]), .A(S), .Z(O[403]) );
  ANDN U176 ( .B(A[402]), .A(S), .Z(O[402]) );
  ANDN U177 ( .B(A[401]), .A(S), .Z(O[401]) );
  ANDN U178 ( .B(A[400]), .A(S), .Z(O[400]) );
  ANDN U179 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U180 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U181 ( .B(A[399]), .A(S), .Z(O[399]) );
  ANDN U182 ( .B(A[398]), .A(S), .Z(O[398]) );
  ANDN U183 ( .B(A[397]), .A(S), .Z(O[397]) );
  ANDN U184 ( .B(A[396]), .A(S), .Z(O[396]) );
  ANDN U185 ( .B(A[395]), .A(S), .Z(O[395]) );
  ANDN U186 ( .B(A[394]), .A(S), .Z(O[394]) );
  ANDN U187 ( .B(A[393]), .A(S), .Z(O[393]) );
  ANDN U188 ( .B(A[392]), .A(S), .Z(O[392]) );
  ANDN U189 ( .B(A[391]), .A(S), .Z(O[391]) );
  ANDN U190 ( .B(A[390]), .A(S), .Z(O[390]) );
  ANDN U191 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U192 ( .B(A[389]), .A(S), .Z(O[389]) );
  ANDN U193 ( .B(A[388]), .A(S), .Z(O[388]) );
  ANDN U194 ( .B(A[387]), .A(S), .Z(O[387]) );
  ANDN U195 ( .B(A[386]), .A(S), .Z(O[386]) );
  ANDN U196 ( .B(A[385]), .A(S), .Z(O[385]) );
  ANDN U197 ( .B(A[384]), .A(S), .Z(O[384]) );
  ANDN U198 ( .B(A[383]), .A(S), .Z(O[383]) );
  ANDN U199 ( .B(A[382]), .A(S), .Z(O[382]) );
  ANDN U200 ( .B(A[381]), .A(S), .Z(O[381]) );
  ANDN U201 ( .B(A[380]), .A(S), .Z(O[380]) );
  ANDN U202 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U203 ( .B(A[379]), .A(S), .Z(O[379]) );
  ANDN U204 ( .B(A[378]), .A(S), .Z(O[378]) );
  ANDN U205 ( .B(A[377]), .A(S), .Z(O[377]) );
  ANDN U206 ( .B(A[376]), .A(S), .Z(O[376]) );
  ANDN U207 ( .B(A[375]), .A(S), .Z(O[375]) );
  ANDN U208 ( .B(A[374]), .A(S), .Z(O[374]) );
  ANDN U209 ( .B(A[373]), .A(S), .Z(O[373]) );
  ANDN U210 ( .B(A[372]), .A(S), .Z(O[372]) );
  ANDN U211 ( .B(A[371]), .A(S), .Z(O[371]) );
  ANDN U212 ( .B(A[370]), .A(S), .Z(O[370]) );
  ANDN U213 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U214 ( .B(A[369]), .A(S), .Z(O[369]) );
  ANDN U215 ( .B(A[368]), .A(S), .Z(O[368]) );
  ANDN U216 ( .B(A[367]), .A(S), .Z(O[367]) );
  ANDN U217 ( .B(A[366]), .A(S), .Z(O[366]) );
  ANDN U218 ( .B(A[365]), .A(S), .Z(O[365]) );
  ANDN U219 ( .B(A[364]), .A(S), .Z(O[364]) );
  ANDN U220 ( .B(A[363]), .A(S), .Z(O[363]) );
  ANDN U221 ( .B(A[362]), .A(S), .Z(O[362]) );
  ANDN U222 ( .B(A[361]), .A(S), .Z(O[361]) );
  ANDN U223 ( .B(A[360]), .A(S), .Z(O[360]) );
  ANDN U224 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U225 ( .B(A[359]), .A(S), .Z(O[359]) );
  ANDN U226 ( .B(A[358]), .A(S), .Z(O[358]) );
  ANDN U227 ( .B(A[357]), .A(S), .Z(O[357]) );
  ANDN U228 ( .B(A[356]), .A(S), .Z(O[356]) );
  ANDN U229 ( .B(A[355]), .A(S), .Z(O[355]) );
  ANDN U230 ( .B(A[354]), .A(S), .Z(O[354]) );
  ANDN U231 ( .B(A[353]), .A(S), .Z(O[353]) );
  ANDN U232 ( .B(A[352]), .A(S), .Z(O[352]) );
  ANDN U233 ( .B(A[351]), .A(S), .Z(O[351]) );
  ANDN U234 ( .B(A[350]), .A(S), .Z(O[350]) );
  ANDN U235 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U236 ( .B(A[349]), .A(S), .Z(O[349]) );
  ANDN U237 ( .B(A[348]), .A(S), .Z(O[348]) );
  ANDN U238 ( .B(A[347]), .A(S), .Z(O[347]) );
  ANDN U239 ( .B(A[346]), .A(S), .Z(O[346]) );
  ANDN U240 ( .B(A[345]), .A(S), .Z(O[345]) );
  ANDN U241 ( .B(A[344]), .A(S), .Z(O[344]) );
  ANDN U242 ( .B(A[343]), .A(S), .Z(O[343]) );
  ANDN U243 ( .B(A[342]), .A(S), .Z(O[342]) );
  ANDN U244 ( .B(A[341]), .A(S), .Z(O[341]) );
  ANDN U245 ( .B(A[340]), .A(S), .Z(O[340]) );
  ANDN U246 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U247 ( .B(A[339]), .A(S), .Z(O[339]) );
  ANDN U248 ( .B(A[338]), .A(S), .Z(O[338]) );
  ANDN U249 ( .B(A[337]), .A(S), .Z(O[337]) );
  ANDN U250 ( .B(A[336]), .A(S), .Z(O[336]) );
  ANDN U251 ( .B(A[335]), .A(S), .Z(O[335]) );
  ANDN U252 ( .B(A[334]), .A(S), .Z(O[334]) );
  ANDN U253 ( .B(A[333]), .A(S), .Z(O[333]) );
  ANDN U254 ( .B(A[332]), .A(S), .Z(O[332]) );
  ANDN U255 ( .B(A[331]), .A(S), .Z(O[331]) );
  ANDN U256 ( .B(A[330]), .A(S), .Z(O[330]) );
  ANDN U257 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U258 ( .B(A[329]), .A(S), .Z(O[329]) );
  ANDN U259 ( .B(A[328]), .A(S), .Z(O[328]) );
  ANDN U260 ( .B(A[327]), .A(S), .Z(O[327]) );
  ANDN U261 ( .B(A[326]), .A(S), .Z(O[326]) );
  ANDN U262 ( .B(A[325]), .A(S), .Z(O[325]) );
  ANDN U263 ( .B(A[324]), .A(S), .Z(O[324]) );
  ANDN U264 ( .B(A[323]), .A(S), .Z(O[323]) );
  ANDN U265 ( .B(A[322]), .A(S), .Z(O[322]) );
  ANDN U266 ( .B(A[321]), .A(S), .Z(O[321]) );
  ANDN U267 ( .B(A[320]), .A(S), .Z(O[320]) );
  ANDN U268 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U269 ( .B(A[319]), .A(S), .Z(O[319]) );
  ANDN U270 ( .B(A[318]), .A(S), .Z(O[318]) );
  ANDN U271 ( .B(A[317]), .A(S), .Z(O[317]) );
  ANDN U272 ( .B(A[316]), .A(S), .Z(O[316]) );
  ANDN U273 ( .B(A[315]), .A(S), .Z(O[315]) );
  ANDN U274 ( .B(A[314]), .A(S), .Z(O[314]) );
  ANDN U275 ( .B(A[313]), .A(S), .Z(O[313]) );
  ANDN U276 ( .B(A[312]), .A(S), .Z(O[312]) );
  ANDN U277 ( .B(A[311]), .A(S), .Z(O[311]) );
  ANDN U278 ( .B(A[310]), .A(S), .Z(O[310]) );
  ANDN U279 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U280 ( .B(A[309]), .A(S), .Z(O[309]) );
  ANDN U281 ( .B(A[308]), .A(S), .Z(O[308]) );
  ANDN U282 ( .B(A[307]), .A(S), .Z(O[307]) );
  ANDN U283 ( .B(A[306]), .A(S), .Z(O[306]) );
  ANDN U284 ( .B(A[305]), .A(S), .Z(O[305]) );
  ANDN U285 ( .B(A[304]), .A(S), .Z(O[304]) );
  ANDN U286 ( .B(A[303]), .A(S), .Z(O[303]) );
  ANDN U287 ( .B(A[302]), .A(S), .Z(O[302]) );
  ANDN U288 ( .B(A[301]), .A(S), .Z(O[301]) );
  ANDN U289 ( .B(A[300]), .A(S), .Z(O[300]) );
  ANDN U290 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U291 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U292 ( .B(A[299]), .A(S), .Z(O[299]) );
  ANDN U293 ( .B(A[298]), .A(S), .Z(O[298]) );
  ANDN U294 ( .B(A[297]), .A(S), .Z(O[297]) );
  ANDN U295 ( .B(A[296]), .A(S), .Z(O[296]) );
  ANDN U296 ( .B(A[295]), .A(S), .Z(O[295]) );
  ANDN U297 ( .B(A[294]), .A(S), .Z(O[294]) );
  ANDN U298 ( .B(A[293]), .A(S), .Z(O[293]) );
  ANDN U299 ( .B(A[292]), .A(S), .Z(O[292]) );
  ANDN U300 ( .B(A[291]), .A(S), .Z(O[291]) );
  ANDN U301 ( .B(A[290]), .A(S), .Z(O[290]) );
  ANDN U302 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U303 ( .B(A[289]), .A(S), .Z(O[289]) );
  ANDN U304 ( .B(A[288]), .A(S), .Z(O[288]) );
  ANDN U305 ( .B(A[287]), .A(S), .Z(O[287]) );
  ANDN U306 ( .B(A[286]), .A(S), .Z(O[286]) );
  ANDN U307 ( .B(A[285]), .A(S), .Z(O[285]) );
  ANDN U308 ( .B(A[284]), .A(S), .Z(O[284]) );
  ANDN U309 ( .B(A[283]), .A(S), .Z(O[283]) );
  ANDN U310 ( .B(A[282]), .A(S), .Z(O[282]) );
  ANDN U311 ( .B(A[281]), .A(S), .Z(O[281]) );
  ANDN U312 ( .B(A[280]), .A(S), .Z(O[280]) );
  ANDN U313 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U314 ( .B(A[279]), .A(S), .Z(O[279]) );
  ANDN U315 ( .B(A[278]), .A(S), .Z(O[278]) );
  ANDN U316 ( .B(A[277]), .A(S), .Z(O[277]) );
  ANDN U317 ( .B(A[276]), .A(S), .Z(O[276]) );
  ANDN U318 ( .B(A[275]), .A(S), .Z(O[275]) );
  ANDN U319 ( .B(A[274]), .A(S), .Z(O[274]) );
  ANDN U320 ( .B(A[273]), .A(S), .Z(O[273]) );
  ANDN U321 ( .B(A[272]), .A(S), .Z(O[272]) );
  ANDN U322 ( .B(A[271]), .A(S), .Z(O[271]) );
  ANDN U323 ( .B(A[270]), .A(S), .Z(O[270]) );
  ANDN U324 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U325 ( .B(A[269]), .A(S), .Z(O[269]) );
  ANDN U326 ( .B(A[268]), .A(S), .Z(O[268]) );
  ANDN U327 ( .B(A[267]), .A(S), .Z(O[267]) );
  ANDN U328 ( .B(A[266]), .A(S), .Z(O[266]) );
  ANDN U329 ( .B(A[265]), .A(S), .Z(O[265]) );
  ANDN U330 ( .B(A[264]), .A(S), .Z(O[264]) );
  ANDN U331 ( .B(A[263]), .A(S), .Z(O[263]) );
  ANDN U332 ( .B(A[262]), .A(S), .Z(O[262]) );
  ANDN U333 ( .B(A[261]), .A(S), .Z(O[261]) );
  ANDN U334 ( .B(A[260]), .A(S), .Z(O[260]) );
  ANDN U335 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U336 ( .B(A[259]), .A(S), .Z(O[259]) );
  ANDN U337 ( .B(A[258]), .A(S), .Z(O[258]) );
  ANDN U338 ( .B(A[257]), .A(S), .Z(O[257]) );
  ANDN U339 ( .B(A[256]), .A(S), .Z(O[256]) );
  ANDN U340 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U341 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U342 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U343 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U344 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U345 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U346 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U347 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U348 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U349 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U350 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U351 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U352 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U353 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U354 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U355 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U356 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U357 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U358 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U359 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U360 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U361 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U362 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U363 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U364 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U365 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U366 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U367 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U368 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U369 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U370 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U371 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U372 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U373 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U374 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U375 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U376 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U377 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U378 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U379 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U380 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U381 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U382 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U383 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U384 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U385 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U386 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U387 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U388 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U389 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U390 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U391 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U392 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U393 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U394 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U395 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U396 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U397 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U398 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U399 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U400 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U401 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U402 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U403 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U404 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U405 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U406 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U407 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U408 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U409 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U410 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U411 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U412 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U413 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U414 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U415 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U416 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U417 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U418 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U419 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U420 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U421 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U422 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U423 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U424 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U425 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U426 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U427 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U428 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U429 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U430 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U431 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U432 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U433 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U434 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U435 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U436 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U437 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U438 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U439 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U440 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U441 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U442 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U443 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U444 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U445 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U446 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U447 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U448 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U449 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U450 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U451 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U452 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U453 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U454 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U455 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U456 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U457 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U458 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U459 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U460 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U461 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U462 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U463 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U464 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U465 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U466 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U467 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U468 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U469 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U470 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U471 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U472 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U473 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U474 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U475 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U476 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U477 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U478 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U479 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U480 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U481 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U482 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U483 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U484 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U485 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U486 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U487 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U488 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U489 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U490 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U491 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U492 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U493 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U494 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U495 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U496 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U497 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U498 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U499 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U500 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U501 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U502 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U503 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U504 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U505 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U506 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U507 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U508 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U509 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U510 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U511 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U512 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module MUX_N514_2 ( A, B, S, O );
  input [513:0] A;
  input [513:0] B;
  output [513:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[511]), .A(S), .Z(O[511]) );
  ANDN U56 ( .B(A[510]), .A(S), .Z(O[510]) );
  ANDN U57 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U58 ( .B(A[509]), .A(S), .Z(O[509]) );
  ANDN U59 ( .B(A[508]), .A(S), .Z(O[508]) );
  ANDN U60 ( .B(A[507]), .A(S), .Z(O[507]) );
  ANDN U61 ( .B(A[506]), .A(S), .Z(O[506]) );
  ANDN U62 ( .B(A[505]), .A(S), .Z(O[505]) );
  ANDN U63 ( .B(A[504]), .A(S), .Z(O[504]) );
  ANDN U64 ( .B(A[503]), .A(S), .Z(O[503]) );
  ANDN U65 ( .B(A[502]), .A(S), .Z(O[502]) );
  ANDN U66 ( .B(A[501]), .A(S), .Z(O[501]) );
  ANDN U67 ( .B(A[500]), .A(S), .Z(O[500]) );
  ANDN U68 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U69 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U70 ( .B(A[499]), .A(S), .Z(O[499]) );
  ANDN U71 ( .B(A[498]), .A(S), .Z(O[498]) );
  ANDN U72 ( .B(A[497]), .A(S), .Z(O[497]) );
  ANDN U73 ( .B(A[496]), .A(S), .Z(O[496]) );
  ANDN U74 ( .B(A[495]), .A(S), .Z(O[495]) );
  ANDN U75 ( .B(A[494]), .A(S), .Z(O[494]) );
  ANDN U76 ( .B(A[493]), .A(S), .Z(O[493]) );
  ANDN U77 ( .B(A[492]), .A(S), .Z(O[492]) );
  ANDN U78 ( .B(A[491]), .A(S), .Z(O[491]) );
  ANDN U79 ( .B(A[490]), .A(S), .Z(O[490]) );
  ANDN U80 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U81 ( .B(A[489]), .A(S), .Z(O[489]) );
  ANDN U82 ( .B(A[488]), .A(S), .Z(O[488]) );
  ANDN U83 ( .B(A[487]), .A(S), .Z(O[487]) );
  ANDN U84 ( .B(A[486]), .A(S), .Z(O[486]) );
  ANDN U85 ( .B(A[485]), .A(S), .Z(O[485]) );
  ANDN U86 ( .B(A[484]), .A(S), .Z(O[484]) );
  ANDN U87 ( .B(A[483]), .A(S), .Z(O[483]) );
  ANDN U88 ( .B(A[482]), .A(S), .Z(O[482]) );
  ANDN U89 ( .B(A[481]), .A(S), .Z(O[481]) );
  ANDN U90 ( .B(A[480]), .A(S), .Z(O[480]) );
  ANDN U91 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U92 ( .B(A[479]), .A(S), .Z(O[479]) );
  ANDN U93 ( .B(A[478]), .A(S), .Z(O[478]) );
  ANDN U94 ( .B(A[477]), .A(S), .Z(O[477]) );
  ANDN U95 ( .B(A[476]), .A(S), .Z(O[476]) );
  ANDN U96 ( .B(A[475]), .A(S), .Z(O[475]) );
  ANDN U97 ( .B(A[474]), .A(S), .Z(O[474]) );
  ANDN U98 ( .B(A[473]), .A(S), .Z(O[473]) );
  ANDN U99 ( .B(A[472]), .A(S), .Z(O[472]) );
  ANDN U100 ( .B(A[471]), .A(S), .Z(O[471]) );
  ANDN U101 ( .B(A[470]), .A(S), .Z(O[470]) );
  ANDN U102 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U103 ( .B(A[469]), .A(S), .Z(O[469]) );
  ANDN U104 ( .B(A[468]), .A(S), .Z(O[468]) );
  ANDN U105 ( .B(A[467]), .A(S), .Z(O[467]) );
  ANDN U106 ( .B(A[466]), .A(S), .Z(O[466]) );
  ANDN U107 ( .B(A[465]), .A(S), .Z(O[465]) );
  ANDN U108 ( .B(A[464]), .A(S), .Z(O[464]) );
  ANDN U109 ( .B(A[463]), .A(S), .Z(O[463]) );
  ANDN U110 ( .B(A[462]), .A(S), .Z(O[462]) );
  ANDN U111 ( .B(A[461]), .A(S), .Z(O[461]) );
  ANDN U112 ( .B(A[460]), .A(S), .Z(O[460]) );
  ANDN U113 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U114 ( .B(A[459]), .A(S), .Z(O[459]) );
  ANDN U115 ( .B(A[458]), .A(S), .Z(O[458]) );
  ANDN U116 ( .B(A[457]), .A(S), .Z(O[457]) );
  ANDN U117 ( .B(A[456]), .A(S), .Z(O[456]) );
  ANDN U118 ( .B(A[455]), .A(S), .Z(O[455]) );
  ANDN U119 ( .B(A[454]), .A(S), .Z(O[454]) );
  ANDN U120 ( .B(A[453]), .A(S), .Z(O[453]) );
  ANDN U121 ( .B(A[452]), .A(S), .Z(O[452]) );
  ANDN U122 ( .B(A[451]), .A(S), .Z(O[451]) );
  ANDN U123 ( .B(A[450]), .A(S), .Z(O[450]) );
  ANDN U124 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U125 ( .B(A[449]), .A(S), .Z(O[449]) );
  ANDN U126 ( .B(A[448]), .A(S), .Z(O[448]) );
  ANDN U127 ( .B(A[447]), .A(S), .Z(O[447]) );
  ANDN U128 ( .B(A[446]), .A(S), .Z(O[446]) );
  ANDN U129 ( .B(A[445]), .A(S), .Z(O[445]) );
  ANDN U130 ( .B(A[444]), .A(S), .Z(O[444]) );
  ANDN U131 ( .B(A[443]), .A(S), .Z(O[443]) );
  ANDN U132 ( .B(A[442]), .A(S), .Z(O[442]) );
  ANDN U133 ( .B(A[441]), .A(S), .Z(O[441]) );
  ANDN U134 ( .B(A[440]), .A(S), .Z(O[440]) );
  ANDN U135 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U136 ( .B(A[439]), .A(S), .Z(O[439]) );
  ANDN U137 ( .B(A[438]), .A(S), .Z(O[438]) );
  ANDN U138 ( .B(A[437]), .A(S), .Z(O[437]) );
  ANDN U139 ( .B(A[436]), .A(S), .Z(O[436]) );
  ANDN U140 ( .B(A[435]), .A(S), .Z(O[435]) );
  ANDN U141 ( .B(A[434]), .A(S), .Z(O[434]) );
  ANDN U142 ( .B(A[433]), .A(S), .Z(O[433]) );
  ANDN U143 ( .B(A[432]), .A(S), .Z(O[432]) );
  ANDN U144 ( .B(A[431]), .A(S), .Z(O[431]) );
  ANDN U145 ( .B(A[430]), .A(S), .Z(O[430]) );
  ANDN U146 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U147 ( .B(A[429]), .A(S), .Z(O[429]) );
  ANDN U148 ( .B(A[428]), .A(S), .Z(O[428]) );
  ANDN U149 ( .B(A[427]), .A(S), .Z(O[427]) );
  ANDN U150 ( .B(A[426]), .A(S), .Z(O[426]) );
  ANDN U151 ( .B(A[425]), .A(S), .Z(O[425]) );
  ANDN U152 ( .B(A[424]), .A(S), .Z(O[424]) );
  ANDN U153 ( .B(A[423]), .A(S), .Z(O[423]) );
  ANDN U154 ( .B(A[422]), .A(S), .Z(O[422]) );
  ANDN U155 ( .B(A[421]), .A(S), .Z(O[421]) );
  ANDN U156 ( .B(A[420]), .A(S), .Z(O[420]) );
  ANDN U157 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U158 ( .B(A[419]), .A(S), .Z(O[419]) );
  ANDN U159 ( .B(A[418]), .A(S), .Z(O[418]) );
  ANDN U160 ( .B(A[417]), .A(S), .Z(O[417]) );
  ANDN U161 ( .B(A[416]), .A(S), .Z(O[416]) );
  ANDN U162 ( .B(A[415]), .A(S), .Z(O[415]) );
  ANDN U163 ( .B(A[414]), .A(S), .Z(O[414]) );
  ANDN U164 ( .B(A[413]), .A(S), .Z(O[413]) );
  ANDN U165 ( .B(A[412]), .A(S), .Z(O[412]) );
  ANDN U166 ( .B(A[411]), .A(S), .Z(O[411]) );
  ANDN U167 ( .B(A[410]), .A(S), .Z(O[410]) );
  ANDN U168 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U169 ( .B(A[409]), .A(S), .Z(O[409]) );
  ANDN U170 ( .B(A[408]), .A(S), .Z(O[408]) );
  ANDN U171 ( .B(A[407]), .A(S), .Z(O[407]) );
  ANDN U172 ( .B(A[406]), .A(S), .Z(O[406]) );
  ANDN U173 ( .B(A[405]), .A(S), .Z(O[405]) );
  ANDN U174 ( .B(A[404]), .A(S), .Z(O[404]) );
  ANDN U175 ( .B(A[403]), .A(S), .Z(O[403]) );
  ANDN U176 ( .B(A[402]), .A(S), .Z(O[402]) );
  ANDN U177 ( .B(A[401]), .A(S), .Z(O[401]) );
  ANDN U178 ( .B(A[400]), .A(S), .Z(O[400]) );
  ANDN U179 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U180 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U181 ( .B(A[399]), .A(S), .Z(O[399]) );
  ANDN U182 ( .B(A[398]), .A(S), .Z(O[398]) );
  ANDN U183 ( .B(A[397]), .A(S), .Z(O[397]) );
  ANDN U184 ( .B(A[396]), .A(S), .Z(O[396]) );
  ANDN U185 ( .B(A[395]), .A(S), .Z(O[395]) );
  ANDN U186 ( .B(A[394]), .A(S), .Z(O[394]) );
  ANDN U187 ( .B(A[393]), .A(S), .Z(O[393]) );
  ANDN U188 ( .B(A[392]), .A(S), .Z(O[392]) );
  ANDN U189 ( .B(A[391]), .A(S), .Z(O[391]) );
  ANDN U190 ( .B(A[390]), .A(S), .Z(O[390]) );
  ANDN U191 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U192 ( .B(A[389]), .A(S), .Z(O[389]) );
  ANDN U193 ( .B(A[388]), .A(S), .Z(O[388]) );
  ANDN U194 ( .B(A[387]), .A(S), .Z(O[387]) );
  ANDN U195 ( .B(A[386]), .A(S), .Z(O[386]) );
  ANDN U196 ( .B(A[385]), .A(S), .Z(O[385]) );
  ANDN U197 ( .B(A[384]), .A(S), .Z(O[384]) );
  ANDN U198 ( .B(A[383]), .A(S), .Z(O[383]) );
  ANDN U199 ( .B(A[382]), .A(S), .Z(O[382]) );
  ANDN U200 ( .B(A[381]), .A(S), .Z(O[381]) );
  ANDN U201 ( .B(A[380]), .A(S), .Z(O[380]) );
  ANDN U202 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U203 ( .B(A[379]), .A(S), .Z(O[379]) );
  ANDN U204 ( .B(A[378]), .A(S), .Z(O[378]) );
  ANDN U205 ( .B(A[377]), .A(S), .Z(O[377]) );
  ANDN U206 ( .B(A[376]), .A(S), .Z(O[376]) );
  ANDN U207 ( .B(A[375]), .A(S), .Z(O[375]) );
  ANDN U208 ( .B(A[374]), .A(S), .Z(O[374]) );
  ANDN U209 ( .B(A[373]), .A(S), .Z(O[373]) );
  ANDN U210 ( .B(A[372]), .A(S), .Z(O[372]) );
  ANDN U211 ( .B(A[371]), .A(S), .Z(O[371]) );
  ANDN U212 ( .B(A[370]), .A(S), .Z(O[370]) );
  ANDN U213 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U214 ( .B(A[369]), .A(S), .Z(O[369]) );
  ANDN U215 ( .B(A[368]), .A(S), .Z(O[368]) );
  ANDN U216 ( .B(A[367]), .A(S), .Z(O[367]) );
  ANDN U217 ( .B(A[366]), .A(S), .Z(O[366]) );
  ANDN U218 ( .B(A[365]), .A(S), .Z(O[365]) );
  ANDN U219 ( .B(A[364]), .A(S), .Z(O[364]) );
  ANDN U220 ( .B(A[363]), .A(S), .Z(O[363]) );
  ANDN U221 ( .B(A[362]), .A(S), .Z(O[362]) );
  ANDN U222 ( .B(A[361]), .A(S), .Z(O[361]) );
  ANDN U223 ( .B(A[360]), .A(S), .Z(O[360]) );
  ANDN U224 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U225 ( .B(A[359]), .A(S), .Z(O[359]) );
  ANDN U226 ( .B(A[358]), .A(S), .Z(O[358]) );
  ANDN U227 ( .B(A[357]), .A(S), .Z(O[357]) );
  ANDN U228 ( .B(A[356]), .A(S), .Z(O[356]) );
  ANDN U229 ( .B(A[355]), .A(S), .Z(O[355]) );
  ANDN U230 ( .B(A[354]), .A(S), .Z(O[354]) );
  ANDN U231 ( .B(A[353]), .A(S), .Z(O[353]) );
  ANDN U232 ( .B(A[352]), .A(S), .Z(O[352]) );
  ANDN U233 ( .B(A[351]), .A(S), .Z(O[351]) );
  ANDN U234 ( .B(A[350]), .A(S), .Z(O[350]) );
  ANDN U235 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U236 ( .B(A[349]), .A(S), .Z(O[349]) );
  ANDN U237 ( .B(A[348]), .A(S), .Z(O[348]) );
  ANDN U238 ( .B(A[347]), .A(S), .Z(O[347]) );
  ANDN U239 ( .B(A[346]), .A(S), .Z(O[346]) );
  ANDN U240 ( .B(A[345]), .A(S), .Z(O[345]) );
  ANDN U241 ( .B(A[344]), .A(S), .Z(O[344]) );
  ANDN U242 ( .B(A[343]), .A(S), .Z(O[343]) );
  ANDN U243 ( .B(A[342]), .A(S), .Z(O[342]) );
  ANDN U244 ( .B(A[341]), .A(S), .Z(O[341]) );
  ANDN U245 ( .B(A[340]), .A(S), .Z(O[340]) );
  ANDN U246 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U247 ( .B(A[339]), .A(S), .Z(O[339]) );
  ANDN U248 ( .B(A[338]), .A(S), .Z(O[338]) );
  ANDN U249 ( .B(A[337]), .A(S), .Z(O[337]) );
  ANDN U250 ( .B(A[336]), .A(S), .Z(O[336]) );
  ANDN U251 ( .B(A[335]), .A(S), .Z(O[335]) );
  ANDN U252 ( .B(A[334]), .A(S), .Z(O[334]) );
  ANDN U253 ( .B(A[333]), .A(S), .Z(O[333]) );
  ANDN U254 ( .B(A[332]), .A(S), .Z(O[332]) );
  ANDN U255 ( .B(A[331]), .A(S), .Z(O[331]) );
  ANDN U256 ( .B(A[330]), .A(S), .Z(O[330]) );
  ANDN U257 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U258 ( .B(A[329]), .A(S), .Z(O[329]) );
  ANDN U259 ( .B(A[328]), .A(S), .Z(O[328]) );
  ANDN U260 ( .B(A[327]), .A(S), .Z(O[327]) );
  ANDN U261 ( .B(A[326]), .A(S), .Z(O[326]) );
  ANDN U262 ( .B(A[325]), .A(S), .Z(O[325]) );
  ANDN U263 ( .B(A[324]), .A(S), .Z(O[324]) );
  ANDN U264 ( .B(A[323]), .A(S), .Z(O[323]) );
  ANDN U265 ( .B(A[322]), .A(S), .Z(O[322]) );
  ANDN U266 ( .B(A[321]), .A(S), .Z(O[321]) );
  ANDN U267 ( .B(A[320]), .A(S), .Z(O[320]) );
  ANDN U268 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U269 ( .B(A[319]), .A(S), .Z(O[319]) );
  ANDN U270 ( .B(A[318]), .A(S), .Z(O[318]) );
  ANDN U271 ( .B(A[317]), .A(S), .Z(O[317]) );
  ANDN U272 ( .B(A[316]), .A(S), .Z(O[316]) );
  ANDN U273 ( .B(A[315]), .A(S), .Z(O[315]) );
  ANDN U274 ( .B(A[314]), .A(S), .Z(O[314]) );
  ANDN U275 ( .B(A[313]), .A(S), .Z(O[313]) );
  ANDN U276 ( .B(A[312]), .A(S), .Z(O[312]) );
  ANDN U277 ( .B(A[311]), .A(S), .Z(O[311]) );
  ANDN U278 ( .B(A[310]), .A(S), .Z(O[310]) );
  ANDN U279 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U280 ( .B(A[309]), .A(S), .Z(O[309]) );
  ANDN U281 ( .B(A[308]), .A(S), .Z(O[308]) );
  ANDN U282 ( .B(A[307]), .A(S), .Z(O[307]) );
  ANDN U283 ( .B(A[306]), .A(S), .Z(O[306]) );
  ANDN U284 ( .B(A[305]), .A(S), .Z(O[305]) );
  ANDN U285 ( .B(A[304]), .A(S), .Z(O[304]) );
  ANDN U286 ( .B(A[303]), .A(S), .Z(O[303]) );
  ANDN U287 ( .B(A[302]), .A(S), .Z(O[302]) );
  ANDN U288 ( .B(A[301]), .A(S), .Z(O[301]) );
  ANDN U289 ( .B(A[300]), .A(S), .Z(O[300]) );
  ANDN U290 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U291 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U292 ( .B(A[299]), .A(S), .Z(O[299]) );
  ANDN U293 ( .B(A[298]), .A(S), .Z(O[298]) );
  ANDN U294 ( .B(A[297]), .A(S), .Z(O[297]) );
  ANDN U295 ( .B(A[296]), .A(S), .Z(O[296]) );
  ANDN U296 ( .B(A[295]), .A(S), .Z(O[295]) );
  ANDN U297 ( .B(A[294]), .A(S), .Z(O[294]) );
  ANDN U298 ( .B(A[293]), .A(S), .Z(O[293]) );
  ANDN U299 ( .B(A[292]), .A(S), .Z(O[292]) );
  ANDN U300 ( .B(A[291]), .A(S), .Z(O[291]) );
  ANDN U301 ( .B(A[290]), .A(S), .Z(O[290]) );
  ANDN U302 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U303 ( .B(A[289]), .A(S), .Z(O[289]) );
  ANDN U304 ( .B(A[288]), .A(S), .Z(O[288]) );
  ANDN U305 ( .B(A[287]), .A(S), .Z(O[287]) );
  ANDN U306 ( .B(A[286]), .A(S), .Z(O[286]) );
  ANDN U307 ( .B(A[285]), .A(S), .Z(O[285]) );
  ANDN U308 ( .B(A[284]), .A(S), .Z(O[284]) );
  ANDN U309 ( .B(A[283]), .A(S), .Z(O[283]) );
  ANDN U310 ( .B(A[282]), .A(S), .Z(O[282]) );
  ANDN U311 ( .B(A[281]), .A(S), .Z(O[281]) );
  ANDN U312 ( .B(A[280]), .A(S), .Z(O[280]) );
  ANDN U313 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U314 ( .B(A[279]), .A(S), .Z(O[279]) );
  ANDN U315 ( .B(A[278]), .A(S), .Z(O[278]) );
  ANDN U316 ( .B(A[277]), .A(S), .Z(O[277]) );
  ANDN U317 ( .B(A[276]), .A(S), .Z(O[276]) );
  ANDN U318 ( .B(A[275]), .A(S), .Z(O[275]) );
  ANDN U319 ( .B(A[274]), .A(S), .Z(O[274]) );
  ANDN U320 ( .B(A[273]), .A(S), .Z(O[273]) );
  ANDN U321 ( .B(A[272]), .A(S), .Z(O[272]) );
  ANDN U322 ( .B(A[271]), .A(S), .Z(O[271]) );
  ANDN U323 ( .B(A[270]), .A(S), .Z(O[270]) );
  ANDN U324 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U325 ( .B(A[269]), .A(S), .Z(O[269]) );
  ANDN U326 ( .B(A[268]), .A(S), .Z(O[268]) );
  ANDN U327 ( .B(A[267]), .A(S), .Z(O[267]) );
  ANDN U328 ( .B(A[266]), .A(S), .Z(O[266]) );
  ANDN U329 ( .B(A[265]), .A(S), .Z(O[265]) );
  ANDN U330 ( .B(A[264]), .A(S), .Z(O[264]) );
  ANDN U331 ( .B(A[263]), .A(S), .Z(O[263]) );
  ANDN U332 ( .B(A[262]), .A(S), .Z(O[262]) );
  ANDN U333 ( .B(A[261]), .A(S), .Z(O[261]) );
  ANDN U334 ( .B(A[260]), .A(S), .Z(O[260]) );
  ANDN U335 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U336 ( .B(A[259]), .A(S), .Z(O[259]) );
  ANDN U337 ( .B(A[258]), .A(S), .Z(O[258]) );
  ANDN U338 ( .B(A[257]), .A(S), .Z(O[257]) );
  ANDN U339 ( .B(A[256]), .A(S), .Z(O[256]) );
  ANDN U340 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U341 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U342 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U343 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U344 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U345 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U346 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U347 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U348 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U349 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U350 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U351 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U352 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U353 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U354 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U355 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U356 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U357 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U358 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U359 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U360 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U361 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U362 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U363 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U364 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U365 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U366 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U367 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U368 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U369 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U370 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U371 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U372 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U373 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U374 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U375 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U376 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U377 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U378 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U379 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U380 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U381 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U382 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U383 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U384 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U385 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U386 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U387 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U388 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U389 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U390 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U391 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U392 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U393 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U394 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U395 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U396 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U397 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U398 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U399 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U400 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U401 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U402 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U403 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U404 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U405 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U406 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U407 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U408 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U409 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U410 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U411 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U412 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U413 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U414 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U415 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U416 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U417 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U418 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U419 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U420 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U421 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U422 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U423 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U424 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U425 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U426 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U427 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U428 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U429 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U430 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U431 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U432 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U433 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U434 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U435 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U436 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U437 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U438 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U439 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U440 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U441 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U442 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U443 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U444 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U445 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U446 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U447 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U448 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U449 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U450 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U451 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U452 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U453 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U454 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U455 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U456 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U457 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U458 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U459 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U460 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U461 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U462 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U463 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U464 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U465 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U466 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U467 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U468 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U469 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U470 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U471 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U472 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U473 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U474 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U475 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U476 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U477 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U478 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U479 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U480 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U481 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U482 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U483 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U484 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U485 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U486 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U487 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U488 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U489 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U490 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U491 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U492 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U493 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U494 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U495 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U496 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U497 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U498 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U499 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U500 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U501 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U502 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U503 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U504 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U505 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U506 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U507 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U508 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U509 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U510 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U511 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U512 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module FA_4382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_4383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_4384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_4895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N514_1 ( A, B, O );
  input [513:0] A;
  input [513:0] B;
  output O;
  wire   n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  wire   [513:1] C;

  FA_4895 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n516), .CI(1'b1), 
        .CO(C[1]) );
  FA_4894 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n517), .CI(C[1]), 
        .CO(C[2]) );
  FA_4893 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n518), .CI(C[2]), 
        .CO(C[3]) );
  FA_4892 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n519), .CI(C[3]), 
        .CO(C[4]) );
  FA_4891 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n520), .CI(C[4]), 
        .CO(C[5]) );
  FA_4890 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n521), .CI(C[5]), 
        .CO(C[6]) );
  FA_4889 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n522), .CI(C[6]), 
        .CO(C[7]) );
  FA_4888 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n523), .CI(C[7]), 
        .CO(C[8]) );
  FA_4887 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n524), .CI(C[8]), 
        .CO(C[9]) );
  FA_4886 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n525), .CI(C[9]), 
        .CO(C[10]) );
  FA_4885 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n526), .CI(C[10]), 
        .CO(C[11]) );
  FA_4884 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n527), .CI(C[11]), 
        .CO(C[12]) );
  FA_4883 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n528), .CI(C[12]), 
        .CO(C[13]) );
  FA_4882 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n529), .CI(C[13]), 
        .CO(C[14]) );
  FA_4881 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n530), .CI(C[14]), 
        .CO(C[15]) );
  FA_4880 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n531), .CI(C[15]), 
        .CO(C[16]) );
  FA_4879 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n532), .CI(C[16]), 
        .CO(C[17]) );
  FA_4878 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n533), .CI(C[17]), 
        .CO(C[18]) );
  FA_4877 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n534), .CI(C[18]), 
        .CO(C[19]) );
  FA_4876 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n535), .CI(C[19]), 
        .CO(C[20]) );
  FA_4875 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n536), .CI(C[20]), 
        .CO(C[21]) );
  FA_4874 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n537), .CI(C[21]), 
        .CO(C[22]) );
  FA_4873 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n538), .CI(C[22]), 
        .CO(C[23]) );
  FA_4872 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n539), .CI(C[23]), 
        .CO(C[24]) );
  FA_4871 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n540), .CI(C[24]), 
        .CO(C[25]) );
  FA_4870 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n541), .CI(C[25]), 
        .CO(C[26]) );
  FA_4869 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n542), .CI(C[26]), 
        .CO(C[27]) );
  FA_4868 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n543), .CI(C[27]), 
        .CO(C[28]) );
  FA_4867 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n544), .CI(C[28]), 
        .CO(C[29]) );
  FA_4866 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n545), .CI(C[29]), 
        .CO(C[30]) );
  FA_4865 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n546), .CI(C[30]), 
        .CO(C[31]) );
  FA_4864 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n547), .CI(C[31]), 
        .CO(C[32]) );
  FA_4863 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n548), .CI(C[32]), 
        .CO(C[33]) );
  FA_4862 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n549), .CI(C[33]), 
        .CO(C[34]) );
  FA_4861 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n550), .CI(C[34]), 
        .CO(C[35]) );
  FA_4860 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n551), .CI(C[35]), 
        .CO(C[36]) );
  FA_4859 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n552), .CI(C[36]), 
        .CO(C[37]) );
  FA_4858 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n553), .CI(C[37]), 
        .CO(C[38]) );
  FA_4857 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n554), .CI(C[38]), 
        .CO(C[39]) );
  FA_4856 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n555), .CI(C[39]), 
        .CO(C[40]) );
  FA_4855 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n556), .CI(C[40]), 
        .CO(C[41]) );
  FA_4854 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n557), .CI(C[41]), 
        .CO(C[42]) );
  FA_4853 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n558), .CI(C[42]), 
        .CO(C[43]) );
  FA_4852 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n559), .CI(C[43]), 
        .CO(C[44]) );
  FA_4851 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n560), .CI(C[44]), 
        .CO(C[45]) );
  FA_4850 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n561), .CI(C[45]), 
        .CO(C[46]) );
  FA_4849 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n562), .CI(C[46]), 
        .CO(C[47]) );
  FA_4848 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n563), .CI(C[47]), 
        .CO(C[48]) );
  FA_4847 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n564), .CI(C[48]), 
        .CO(C[49]) );
  FA_4846 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n565), .CI(C[49]), 
        .CO(C[50]) );
  FA_4845 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n566), .CI(C[50]), 
        .CO(C[51]) );
  FA_4844 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n567), .CI(C[51]), 
        .CO(C[52]) );
  FA_4843 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n568), .CI(C[52]), 
        .CO(C[53]) );
  FA_4842 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n569), .CI(C[53]), 
        .CO(C[54]) );
  FA_4841 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n570), .CI(C[54]), 
        .CO(C[55]) );
  FA_4840 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n571), .CI(C[55]), 
        .CO(C[56]) );
  FA_4839 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n572), .CI(C[56]), 
        .CO(C[57]) );
  FA_4838 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n573), .CI(C[57]), 
        .CO(C[58]) );
  FA_4837 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n574), .CI(C[58]), 
        .CO(C[59]) );
  FA_4836 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n575), .CI(C[59]), 
        .CO(C[60]) );
  FA_4835 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n576), .CI(C[60]), 
        .CO(C[61]) );
  FA_4834 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n577), .CI(C[61]), 
        .CO(C[62]) );
  FA_4833 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n578), .CI(C[62]), 
        .CO(C[63]) );
  FA_4832 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n579), .CI(C[63]), 
        .CO(C[64]) );
  FA_4831 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n580), .CI(C[64]), 
        .CO(C[65]) );
  FA_4830 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n581), .CI(C[65]), 
        .CO(C[66]) );
  FA_4829 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n582), .CI(C[66]), 
        .CO(C[67]) );
  FA_4828 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n583), .CI(C[67]), 
        .CO(C[68]) );
  FA_4827 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n584), .CI(C[68]), 
        .CO(C[69]) );
  FA_4826 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n585), .CI(C[69]), 
        .CO(C[70]) );
  FA_4825 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n586), .CI(C[70]), 
        .CO(C[71]) );
  FA_4824 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n587), .CI(C[71]), 
        .CO(C[72]) );
  FA_4823 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n588), .CI(C[72]), 
        .CO(C[73]) );
  FA_4822 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n589), .CI(C[73]), 
        .CO(C[74]) );
  FA_4821 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n590), .CI(C[74]), 
        .CO(C[75]) );
  FA_4820 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n591), .CI(C[75]), 
        .CO(C[76]) );
  FA_4819 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n592), .CI(C[76]), 
        .CO(C[77]) );
  FA_4818 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n593), .CI(C[77]), 
        .CO(C[78]) );
  FA_4817 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n594), .CI(C[78]), 
        .CO(C[79]) );
  FA_4816 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n595), .CI(C[79]), 
        .CO(C[80]) );
  FA_4815 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n596), .CI(C[80]), 
        .CO(C[81]) );
  FA_4814 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n597), .CI(C[81]), 
        .CO(C[82]) );
  FA_4813 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n598), .CI(C[82]), 
        .CO(C[83]) );
  FA_4812 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n599), .CI(C[83]), 
        .CO(C[84]) );
  FA_4811 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n600), .CI(C[84]), 
        .CO(C[85]) );
  FA_4810 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n601), .CI(C[85]), 
        .CO(C[86]) );
  FA_4809 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n602), .CI(C[86]), 
        .CO(C[87]) );
  FA_4808 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n603), .CI(C[87]), 
        .CO(C[88]) );
  FA_4807 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n604), .CI(C[88]), 
        .CO(C[89]) );
  FA_4806 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n605), .CI(C[89]), 
        .CO(C[90]) );
  FA_4805 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n606), .CI(C[90]), 
        .CO(C[91]) );
  FA_4804 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n607), .CI(C[91]), 
        .CO(C[92]) );
  FA_4803 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n608), .CI(C[92]), 
        .CO(C[93]) );
  FA_4802 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n609), .CI(C[93]), 
        .CO(C[94]) );
  FA_4801 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n610), .CI(C[94]), 
        .CO(C[95]) );
  FA_4800 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n611), .CI(C[95]), 
        .CO(C[96]) );
  FA_4799 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n612), .CI(C[96]), 
        .CO(C[97]) );
  FA_4798 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n613), .CI(C[97]), 
        .CO(C[98]) );
  FA_4797 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n614), .CI(C[98]), 
        .CO(C[99]) );
  FA_4796 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n615), .CI(C[99]), 
        .CO(C[100]) );
  FA_4795 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n616), .CI(C[100]), .CO(C[101]) );
  FA_4794 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n617), .CI(C[101]), .CO(C[102]) );
  FA_4793 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n618), .CI(C[102]), .CO(C[103]) );
  FA_4792 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n619), .CI(C[103]), .CO(C[104]) );
  FA_4791 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n620), .CI(C[104]), .CO(C[105]) );
  FA_4790 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n621), .CI(C[105]), .CO(C[106]) );
  FA_4789 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n622), .CI(C[106]), .CO(C[107]) );
  FA_4788 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n623), .CI(C[107]), .CO(C[108]) );
  FA_4787 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n624), .CI(C[108]), .CO(C[109]) );
  FA_4786 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n625), .CI(C[109]), .CO(C[110]) );
  FA_4785 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n626), .CI(C[110]), .CO(C[111]) );
  FA_4784 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n627), .CI(C[111]), .CO(C[112]) );
  FA_4783 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n628), .CI(C[112]), .CO(C[113]) );
  FA_4782 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n629), .CI(C[113]), .CO(C[114]) );
  FA_4781 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n630), .CI(C[114]), .CO(C[115]) );
  FA_4780 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n631), .CI(C[115]), .CO(C[116]) );
  FA_4779 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n632), .CI(C[116]), .CO(C[117]) );
  FA_4778 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n633), .CI(C[117]), .CO(C[118]) );
  FA_4777 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n634), .CI(C[118]), .CO(C[119]) );
  FA_4776 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n635), .CI(C[119]), .CO(C[120]) );
  FA_4775 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n636), .CI(C[120]), .CO(C[121]) );
  FA_4774 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n637), .CI(C[121]), .CO(C[122]) );
  FA_4773 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n638), .CI(C[122]), .CO(C[123]) );
  FA_4772 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n639), .CI(C[123]), .CO(C[124]) );
  FA_4771 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n640), .CI(C[124]), .CO(C[125]) );
  FA_4770 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n641), .CI(C[125]), .CO(C[126]) );
  FA_4769 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n642), .CI(C[126]), .CO(C[127]) );
  FA_4768 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n643), .CI(C[127]), .CO(C[128]) );
  FA_4767 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n644), .CI(C[128]), .CO(C[129]) );
  FA_4766 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n645), .CI(C[129]), .CO(C[130]) );
  FA_4765 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n646), .CI(C[130]), .CO(C[131]) );
  FA_4764 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n647), .CI(C[131]), .CO(C[132]) );
  FA_4763 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n648), .CI(C[132]), .CO(C[133]) );
  FA_4762 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n649), .CI(C[133]), .CO(C[134]) );
  FA_4761 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n650), .CI(C[134]), .CO(C[135]) );
  FA_4760 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n651), .CI(C[135]), .CO(C[136]) );
  FA_4759 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n652), .CI(C[136]), .CO(C[137]) );
  FA_4758 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n653), .CI(C[137]), .CO(C[138]) );
  FA_4757 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n654), .CI(C[138]), .CO(C[139]) );
  FA_4756 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n655), .CI(C[139]), .CO(C[140]) );
  FA_4755 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n656), .CI(C[140]), .CO(C[141]) );
  FA_4754 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n657), .CI(C[141]), .CO(C[142]) );
  FA_4753 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n658), .CI(C[142]), .CO(C[143]) );
  FA_4752 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n659), .CI(C[143]), .CO(C[144]) );
  FA_4751 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n660), .CI(C[144]), .CO(C[145]) );
  FA_4750 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n661), .CI(C[145]), .CO(C[146]) );
  FA_4749 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n662), .CI(C[146]), .CO(C[147]) );
  FA_4748 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n663), .CI(C[147]), .CO(C[148]) );
  FA_4747 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n664), .CI(C[148]), .CO(C[149]) );
  FA_4746 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n665), .CI(C[149]), .CO(C[150]) );
  FA_4745 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n666), .CI(C[150]), .CO(C[151]) );
  FA_4744 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n667), .CI(C[151]), .CO(C[152]) );
  FA_4743 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n668), .CI(C[152]), .CO(C[153]) );
  FA_4742 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n669), .CI(C[153]), .CO(C[154]) );
  FA_4741 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n670), .CI(C[154]), .CO(C[155]) );
  FA_4740 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n671), .CI(C[155]), .CO(C[156]) );
  FA_4739 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n672), .CI(C[156]), .CO(C[157]) );
  FA_4738 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n673), .CI(C[157]), .CO(C[158]) );
  FA_4737 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n674), .CI(C[158]), .CO(C[159]) );
  FA_4736 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n675), .CI(C[159]), .CO(C[160]) );
  FA_4735 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n676), .CI(C[160]), .CO(C[161]) );
  FA_4734 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n677), .CI(C[161]), .CO(C[162]) );
  FA_4733 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n678), .CI(C[162]), .CO(C[163]) );
  FA_4732 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n679), .CI(C[163]), .CO(C[164]) );
  FA_4731 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n680), .CI(C[164]), .CO(C[165]) );
  FA_4730 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n681), .CI(C[165]), .CO(C[166]) );
  FA_4729 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n682), .CI(C[166]), .CO(C[167]) );
  FA_4728 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n683), .CI(C[167]), .CO(C[168]) );
  FA_4727 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n684), .CI(C[168]), .CO(C[169]) );
  FA_4726 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n685), .CI(C[169]), .CO(C[170]) );
  FA_4725 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n686), .CI(C[170]), .CO(C[171]) );
  FA_4724 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n687), .CI(C[171]), .CO(C[172]) );
  FA_4723 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n688), .CI(C[172]), .CO(C[173]) );
  FA_4722 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n689), .CI(C[173]), .CO(C[174]) );
  FA_4721 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n690), .CI(C[174]), .CO(C[175]) );
  FA_4720 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n691), .CI(C[175]), .CO(C[176]) );
  FA_4719 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n692), .CI(C[176]), .CO(C[177]) );
  FA_4718 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n693), .CI(C[177]), .CO(C[178]) );
  FA_4717 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n694), .CI(C[178]), .CO(C[179]) );
  FA_4716 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n695), .CI(C[179]), .CO(C[180]) );
  FA_4715 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n696), .CI(C[180]), .CO(C[181]) );
  FA_4714 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n697), .CI(C[181]), .CO(C[182]) );
  FA_4713 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n698), .CI(C[182]), .CO(C[183]) );
  FA_4712 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n699), .CI(C[183]), .CO(C[184]) );
  FA_4711 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n700), .CI(C[184]), .CO(C[185]) );
  FA_4710 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n701), .CI(C[185]), .CO(C[186]) );
  FA_4709 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n702), .CI(C[186]), .CO(C[187]) );
  FA_4708 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n703), .CI(C[187]), .CO(C[188]) );
  FA_4707 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n704), .CI(C[188]), .CO(C[189]) );
  FA_4706 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n705), .CI(C[189]), .CO(C[190]) );
  FA_4705 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n706), .CI(C[190]), .CO(C[191]) );
  FA_4704 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n707), .CI(C[191]), .CO(C[192]) );
  FA_4703 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n708), .CI(C[192]), .CO(C[193]) );
  FA_4702 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n709), .CI(C[193]), .CO(C[194]) );
  FA_4701 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n710), .CI(C[194]), .CO(C[195]) );
  FA_4700 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n711), .CI(C[195]), .CO(C[196]) );
  FA_4699 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n712), .CI(C[196]), .CO(C[197]) );
  FA_4698 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n713), .CI(C[197]), .CO(C[198]) );
  FA_4697 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n714), .CI(C[198]), .CO(C[199]) );
  FA_4696 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n715), .CI(C[199]), .CO(C[200]) );
  FA_4695 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n716), .CI(C[200]), .CO(C[201]) );
  FA_4694 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n717), .CI(C[201]), .CO(C[202]) );
  FA_4693 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n718), .CI(C[202]), .CO(C[203]) );
  FA_4692 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n719), .CI(C[203]), .CO(C[204]) );
  FA_4691 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n720), .CI(C[204]), .CO(C[205]) );
  FA_4690 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n721), .CI(C[205]), .CO(C[206]) );
  FA_4689 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n722), .CI(C[206]), .CO(C[207]) );
  FA_4688 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n723), .CI(C[207]), .CO(C[208]) );
  FA_4687 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n724), .CI(C[208]), .CO(C[209]) );
  FA_4686 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n725), .CI(C[209]), .CO(C[210]) );
  FA_4685 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n726), .CI(C[210]), .CO(C[211]) );
  FA_4684 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n727), .CI(C[211]), .CO(C[212]) );
  FA_4683 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n728), .CI(C[212]), .CO(C[213]) );
  FA_4682 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n729), .CI(C[213]), .CO(C[214]) );
  FA_4681 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n730), .CI(C[214]), .CO(C[215]) );
  FA_4680 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n731), .CI(C[215]), .CO(C[216]) );
  FA_4679 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n732), .CI(C[216]), .CO(C[217]) );
  FA_4678 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n733), .CI(C[217]), .CO(C[218]) );
  FA_4677 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n734), .CI(C[218]), .CO(C[219]) );
  FA_4676 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n735), .CI(C[219]), .CO(C[220]) );
  FA_4675 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n736), .CI(C[220]), .CO(C[221]) );
  FA_4674 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n737), .CI(C[221]), .CO(C[222]) );
  FA_4673 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n738), .CI(C[222]), .CO(C[223]) );
  FA_4672 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n739), .CI(C[223]), .CO(C[224]) );
  FA_4671 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n740), .CI(C[224]), .CO(C[225]) );
  FA_4670 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n741), .CI(C[225]), .CO(C[226]) );
  FA_4669 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n742), .CI(C[226]), .CO(C[227]) );
  FA_4668 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n743), .CI(C[227]), .CO(C[228]) );
  FA_4667 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n744), .CI(C[228]), .CO(C[229]) );
  FA_4666 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n745), .CI(C[229]), .CO(C[230]) );
  FA_4665 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n746), .CI(C[230]), .CO(C[231]) );
  FA_4664 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n747), .CI(C[231]), .CO(C[232]) );
  FA_4663 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n748), .CI(C[232]), .CO(C[233]) );
  FA_4662 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n749), .CI(C[233]), .CO(C[234]) );
  FA_4661 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n750), .CI(C[234]), .CO(C[235]) );
  FA_4660 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n751), .CI(C[235]), .CO(C[236]) );
  FA_4659 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n752), .CI(C[236]), .CO(C[237]) );
  FA_4658 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n753), .CI(C[237]), .CO(C[238]) );
  FA_4657 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n754), .CI(C[238]), .CO(C[239]) );
  FA_4656 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n755), .CI(C[239]), .CO(C[240]) );
  FA_4655 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n756), .CI(C[240]), .CO(C[241]) );
  FA_4654 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n757), .CI(C[241]), .CO(C[242]) );
  FA_4653 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n758), .CI(C[242]), .CO(C[243]) );
  FA_4652 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n759), .CI(C[243]), .CO(C[244]) );
  FA_4651 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n760), .CI(C[244]), .CO(C[245]) );
  FA_4650 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n761), .CI(C[245]), .CO(C[246]) );
  FA_4649 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n762), .CI(C[246]), .CO(C[247]) );
  FA_4648 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n763), .CI(C[247]), .CO(C[248]) );
  FA_4647 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n764), .CI(C[248]), .CO(C[249]) );
  FA_4646 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n765), .CI(C[249]), .CO(C[250]) );
  FA_4645 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n766), .CI(C[250]), .CO(C[251]) );
  FA_4644 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n767), .CI(C[251]), .CO(C[252]) );
  FA_4643 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n768), .CI(C[252]), .CO(C[253]) );
  FA_4642 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n769), .CI(C[253]), .CO(C[254]) );
  FA_4641 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n770), .CI(C[254]), .CO(C[255]) );
  FA_4640 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n771), .CI(C[255]), .CO(C[256]) );
  FA_4639 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n772), .CI(C[256]), .CO(C[257]) );
  FA_4638 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n773), .CI(C[257]), .CO(C[258]) );
  FA_4637 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n774), .CI(C[258]), .CO(C[259]) );
  FA_4636 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n775), .CI(C[259]), .CO(C[260]) );
  FA_4635 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n776), .CI(C[260]), .CO(C[261]) );
  FA_4634 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n777), .CI(C[261]), .CO(C[262]) );
  FA_4633 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n778), .CI(C[262]), .CO(C[263]) );
  FA_4632 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n779), .CI(C[263]), .CO(C[264]) );
  FA_4631 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n780), .CI(C[264]), .CO(C[265]) );
  FA_4630 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n781), .CI(C[265]), .CO(C[266]) );
  FA_4629 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n782), .CI(C[266]), .CO(C[267]) );
  FA_4628 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n783), .CI(C[267]), .CO(C[268]) );
  FA_4627 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n784), .CI(C[268]), .CO(C[269]) );
  FA_4626 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n785), .CI(C[269]), .CO(C[270]) );
  FA_4625 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n786), .CI(C[270]), .CO(C[271]) );
  FA_4624 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n787), .CI(C[271]), .CO(C[272]) );
  FA_4623 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n788), .CI(C[272]), .CO(C[273]) );
  FA_4622 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n789), .CI(C[273]), .CO(C[274]) );
  FA_4621 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n790), .CI(C[274]), .CO(C[275]) );
  FA_4620 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n791), .CI(C[275]), .CO(C[276]) );
  FA_4619 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n792), .CI(C[276]), .CO(C[277]) );
  FA_4618 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n793), .CI(C[277]), .CO(C[278]) );
  FA_4617 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n794), .CI(C[278]), .CO(C[279]) );
  FA_4616 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n795), .CI(C[279]), .CO(C[280]) );
  FA_4615 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n796), .CI(C[280]), .CO(C[281]) );
  FA_4614 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n797), .CI(C[281]), .CO(C[282]) );
  FA_4613 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n798), .CI(C[282]), .CO(C[283]) );
  FA_4612 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n799), .CI(C[283]), .CO(C[284]) );
  FA_4611 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n800), .CI(C[284]), .CO(C[285]) );
  FA_4610 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n801), .CI(C[285]), .CO(C[286]) );
  FA_4609 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n802), .CI(C[286]), .CO(C[287]) );
  FA_4608 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n803), .CI(C[287]), .CO(C[288]) );
  FA_4607 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n804), .CI(C[288]), .CO(C[289]) );
  FA_4606 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n805), .CI(C[289]), .CO(C[290]) );
  FA_4605 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n806), .CI(C[290]), .CO(C[291]) );
  FA_4604 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n807), .CI(C[291]), .CO(C[292]) );
  FA_4603 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n808), .CI(C[292]), .CO(C[293]) );
  FA_4602 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n809), .CI(C[293]), .CO(C[294]) );
  FA_4601 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n810), .CI(C[294]), .CO(C[295]) );
  FA_4600 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n811), .CI(C[295]), .CO(C[296]) );
  FA_4599 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n812), .CI(C[296]), .CO(C[297]) );
  FA_4598 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n813), .CI(C[297]), .CO(C[298]) );
  FA_4597 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n814), .CI(C[298]), .CO(C[299]) );
  FA_4596 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n815), .CI(C[299]), .CO(C[300]) );
  FA_4595 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n816), .CI(C[300]), .CO(C[301]) );
  FA_4594 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n817), .CI(C[301]), .CO(C[302]) );
  FA_4593 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n818), .CI(C[302]), .CO(C[303]) );
  FA_4592 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n819), .CI(C[303]), .CO(C[304]) );
  FA_4591 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n820), .CI(C[304]), .CO(C[305]) );
  FA_4590 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n821), .CI(C[305]), .CO(C[306]) );
  FA_4589 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n822), .CI(C[306]), .CO(C[307]) );
  FA_4588 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n823), .CI(C[307]), .CO(C[308]) );
  FA_4587 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n824), .CI(C[308]), .CO(C[309]) );
  FA_4586 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n825), .CI(C[309]), .CO(C[310]) );
  FA_4585 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n826), .CI(C[310]), .CO(C[311]) );
  FA_4584 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n827), .CI(C[311]), .CO(C[312]) );
  FA_4583 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n828), .CI(C[312]), .CO(C[313]) );
  FA_4582 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n829), .CI(C[313]), .CO(C[314]) );
  FA_4581 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n830), .CI(C[314]), .CO(C[315]) );
  FA_4580 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n831), .CI(C[315]), .CO(C[316]) );
  FA_4579 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n832), .CI(C[316]), .CO(C[317]) );
  FA_4578 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n833), .CI(C[317]), .CO(C[318]) );
  FA_4577 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n834), .CI(C[318]), .CO(C[319]) );
  FA_4576 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n835), .CI(C[319]), .CO(C[320]) );
  FA_4575 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n836), .CI(C[320]), .CO(C[321]) );
  FA_4574 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n837), .CI(C[321]), .CO(C[322]) );
  FA_4573 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n838), .CI(C[322]), .CO(C[323]) );
  FA_4572 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n839), .CI(C[323]), .CO(C[324]) );
  FA_4571 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n840), .CI(C[324]), .CO(C[325]) );
  FA_4570 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n841), .CI(C[325]), .CO(C[326]) );
  FA_4569 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n842), .CI(C[326]), .CO(C[327]) );
  FA_4568 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n843), .CI(C[327]), .CO(C[328]) );
  FA_4567 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n844), .CI(C[328]), .CO(C[329]) );
  FA_4566 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n845), .CI(C[329]), .CO(C[330]) );
  FA_4565 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n846), .CI(C[330]), .CO(C[331]) );
  FA_4564 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n847), .CI(C[331]), .CO(C[332]) );
  FA_4563 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n848), .CI(C[332]), .CO(C[333]) );
  FA_4562 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n849), .CI(C[333]), .CO(C[334]) );
  FA_4561 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n850), .CI(C[334]), .CO(C[335]) );
  FA_4560 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n851), .CI(C[335]), .CO(C[336]) );
  FA_4559 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n852), .CI(C[336]), .CO(C[337]) );
  FA_4558 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n853), .CI(C[337]), .CO(C[338]) );
  FA_4557 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n854), .CI(C[338]), .CO(C[339]) );
  FA_4556 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n855), .CI(C[339]), .CO(C[340]) );
  FA_4555 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n856), .CI(C[340]), .CO(C[341]) );
  FA_4554 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n857), .CI(C[341]), .CO(C[342]) );
  FA_4553 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n858), .CI(C[342]), .CO(C[343]) );
  FA_4552 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n859), .CI(C[343]), .CO(C[344]) );
  FA_4551 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n860), .CI(C[344]), .CO(C[345]) );
  FA_4550 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n861), .CI(C[345]), .CO(C[346]) );
  FA_4549 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n862), .CI(C[346]), .CO(C[347]) );
  FA_4548 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n863), .CI(C[347]), .CO(C[348]) );
  FA_4547 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n864), .CI(C[348]), .CO(C[349]) );
  FA_4546 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n865), .CI(C[349]), .CO(C[350]) );
  FA_4545 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n866), .CI(C[350]), .CO(C[351]) );
  FA_4544 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n867), .CI(C[351]), .CO(C[352]) );
  FA_4543 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n868), .CI(C[352]), .CO(C[353]) );
  FA_4542 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n869), .CI(C[353]), .CO(C[354]) );
  FA_4541 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n870), .CI(C[354]), .CO(C[355]) );
  FA_4540 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n871), .CI(C[355]), .CO(C[356]) );
  FA_4539 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n872), .CI(C[356]), .CO(C[357]) );
  FA_4538 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n873), .CI(C[357]), .CO(C[358]) );
  FA_4537 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n874), .CI(C[358]), .CO(C[359]) );
  FA_4536 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n875), .CI(C[359]), .CO(C[360]) );
  FA_4535 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n876), .CI(C[360]), .CO(C[361]) );
  FA_4534 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n877), .CI(C[361]), .CO(C[362]) );
  FA_4533 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n878), .CI(C[362]), .CO(C[363]) );
  FA_4532 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n879), .CI(C[363]), .CO(C[364]) );
  FA_4531 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n880), .CI(C[364]), .CO(C[365]) );
  FA_4530 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n881), .CI(C[365]), .CO(C[366]) );
  FA_4529 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n882), .CI(C[366]), .CO(C[367]) );
  FA_4528 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n883), .CI(C[367]), .CO(C[368]) );
  FA_4527 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n884), .CI(C[368]), .CO(C[369]) );
  FA_4526 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n885), .CI(C[369]), .CO(C[370]) );
  FA_4525 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n886), .CI(C[370]), .CO(C[371]) );
  FA_4524 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n887), .CI(C[371]), .CO(C[372]) );
  FA_4523 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n888), .CI(C[372]), .CO(C[373]) );
  FA_4522 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n889), .CI(C[373]), .CO(C[374]) );
  FA_4521 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n890), .CI(C[374]), .CO(C[375]) );
  FA_4520 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n891), .CI(C[375]), .CO(C[376]) );
  FA_4519 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n892), .CI(C[376]), .CO(C[377]) );
  FA_4518 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n893), .CI(C[377]), .CO(C[378]) );
  FA_4517 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n894), .CI(C[378]), .CO(C[379]) );
  FA_4516 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n895), .CI(C[379]), .CO(C[380]) );
  FA_4515 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n896), .CI(C[380]), .CO(C[381]) );
  FA_4514 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n897), .CI(C[381]), .CO(C[382]) );
  FA_4513 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n898), .CI(C[382]), .CO(C[383]) );
  FA_4512 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n899), .CI(C[383]), .CO(C[384]) );
  FA_4511 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n900), .CI(C[384]), .CO(C[385]) );
  FA_4510 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n901), .CI(C[385]), .CO(C[386]) );
  FA_4509 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n902), .CI(C[386]), .CO(C[387]) );
  FA_4508 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n903), .CI(C[387]), .CO(C[388]) );
  FA_4507 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n904), .CI(C[388]), .CO(C[389]) );
  FA_4506 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n905), .CI(C[389]), .CO(C[390]) );
  FA_4505 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n906), .CI(C[390]), .CO(C[391]) );
  FA_4504 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n907), .CI(C[391]), .CO(C[392]) );
  FA_4503 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n908), .CI(C[392]), .CO(C[393]) );
  FA_4502 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n909), .CI(C[393]), .CO(C[394]) );
  FA_4501 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n910), .CI(C[394]), .CO(C[395]) );
  FA_4500 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n911), .CI(C[395]), .CO(C[396]) );
  FA_4499 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n912), .CI(C[396]), .CO(C[397]) );
  FA_4498 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n913), .CI(C[397]), .CO(C[398]) );
  FA_4497 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n914), .CI(C[398]), .CO(C[399]) );
  FA_4496 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n915), .CI(C[399]), .CO(C[400]) );
  FA_4495 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n916), .CI(C[400]), .CO(C[401]) );
  FA_4494 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n917), .CI(C[401]), .CO(C[402]) );
  FA_4493 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n918), .CI(C[402]), .CO(C[403]) );
  FA_4492 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n919), .CI(C[403]), .CO(C[404]) );
  FA_4491 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n920), .CI(C[404]), .CO(C[405]) );
  FA_4490 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n921), .CI(C[405]), .CO(C[406]) );
  FA_4489 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n922), .CI(C[406]), .CO(C[407]) );
  FA_4488 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n923), .CI(C[407]), .CO(C[408]) );
  FA_4487 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n924), .CI(C[408]), .CO(C[409]) );
  FA_4486 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n925), .CI(C[409]), .CO(C[410]) );
  FA_4485 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n926), .CI(C[410]), .CO(C[411]) );
  FA_4484 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n927), .CI(C[411]), .CO(C[412]) );
  FA_4483 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n928), .CI(C[412]), .CO(C[413]) );
  FA_4482 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n929), .CI(C[413]), .CO(C[414]) );
  FA_4481 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n930), .CI(C[414]), .CO(C[415]) );
  FA_4480 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n931), .CI(C[415]), .CO(C[416]) );
  FA_4479 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n932), .CI(C[416]), .CO(C[417]) );
  FA_4478 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n933), .CI(C[417]), .CO(C[418]) );
  FA_4477 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n934), .CI(C[418]), .CO(C[419]) );
  FA_4476 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n935), .CI(C[419]), .CO(C[420]) );
  FA_4475 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n936), .CI(C[420]), .CO(C[421]) );
  FA_4474 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n937), .CI(C[421]), .CO(C[422]) );
  FA_4473 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n938), .CI(C[422]), .CO(C[423]) );
  FA_4472 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n939), .CI(C[423]), .CO(C[424]) );
  FA_4471 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n940), .CI(C[424]), .CO(C[425]) );
  FA_4470 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n941), .CI(C[425]), .CO(C[426]) );
  FA_4469 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n942), .CI(C[426]), .CO(C[427]) );
  FA_4468 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n943), .CI(C[427]), .CO(C[428]) );
  FA_4467 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n944), .CI(C[428]), .CO(C[429]) );
  FA_4466 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n945), .CI(C[429]), .CO(C[430]) );
  FA_4465 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n946), .CI(C[430]), .CO(C[431]) );
  FA_4464 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n947), .CI(C[431]), .CO(C[432]) );
  FA_4463 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n948), .CI(C[432]), .CO(C[433]) );
  FA_4462 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n949), .CI(C[433]), .CO(C[434]) );
  FA_4461 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n950), .CI(C[434]), .CO(C[435]) );
  FA_4460 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n951), .CI(C[435]), .CO(C[436]) );
  FA_4459 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n952), .CI(C[436]), .CO(C[437]) );
  FA_4458 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n953), .CI(C[437]), .CO(C[438]) );
  FA_4457 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n954), .CI(C[438]), .CO(C[439]) );
  FA_4456 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n955), .CI(C[439]), .CO(C[440]) );
  FA_4455 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n956), .CI(C[440]), .CO(C[441]) );
  FA_4454 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n957), .CI(C[441]), .CO(C[442]) );
  FA_4453 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n958), .CI(C[442]), .CO(C[443]) );
  FA_4452 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n959), .CI(C[443]), .CO(C[444]) );
  FA_4451 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n960), .CI(C[444]), .CO(C[445]) );
  FA_4450 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n961), .CI(C[445]), .CO(C[446]) );
  FA_4449 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n962), .CI(C[446]), .CO(C[447]) );
  FA_4448 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n963), .CI(C[447]), .CO(C[448]) );
  FA_4447 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n964), .CI(C[448]), .CO(C[449]) );
  FA_4446 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n965), .CI(C[449]), .CO(C[450]) );
  FA_4445 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n966), .CI(C[450]), .CO(C[451]) );
  FA_4444 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n967), .CI(C[451]), .CO(C[452]) );
  FA_4443 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n968), .CI(C[452]), .CO(C[453]) );
  FA_4442 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n969), .CI(C[453]), .CO(C[454]) );
  FA_4441 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n970), .CI(C[454]), .CO(C[455]) );
  FA_4440 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n971), .CI(C[455]), .CO(C[456]) );
  FA_4439 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n972), .CI(C[456]), .CO(C[457]) );
  FA_4438 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n973), .CI(C[457]), .CO(C[458]) );
  FA_4437 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n974), .CI(C[458]), .CO(C[459]) );
  FA_4436 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n975), .CI(C[459]), .CO(C[460]) );
  FA_4435 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n976), .CI(C[460]), .CO(C[461]) );
  FA_4434 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n977), .CI(C[461]), .CO(C[462]) );
  FA_4433 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n978), .CI(C[462]), .CO(C[463]) );
  FA_4432 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n979), .CI(C[463]), .CO(C[464]) );
  FA_4431 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n980), .CI(C[464]), .CO(C[465]) );
  FA_4430 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n981), .CI(C[465]), .CO(C[466]) );
  FA_4429 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n982), .CI(C[466]), .CO(C[467]) );
  FA_4428 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n983), .CI(C[467]), .CO(C[468]) );
  FA_4427 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n984), .CI(C[468]), .CO(C[469]) );
  FA_4426 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n985), .CI(C[469]), .CO(C[470]) );
  FA_4425 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n986), .CI(C[470]), .CO(C[471]) );
  FA_4424 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n987), .CI(C[471]), .CO(C[472]) );
  FA_4423 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n988), .CI(C[472]), .CO(C[473]) );
  FA_4422 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n989), .CI(C[473]), .CO(C[474]) );
  FA_4421 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n990), .CI(C[474]), .CO(C[475]) );
  FA_4420 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n991), .CI(C[475]), .CO(C[476]) );
  FA_4419 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n992), .CI(C[476]), .CO(C[477]) );
  FA_4418 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n993), .CI(C[477]), .CO(C[478]) );
  FA_4417 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n994), .CI(C[478]), .CO(C[479]) );
  FA_4416 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n995), .CI(C[479]), .CO(C[480]) );
  FA_4415 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n996), .CI(C[480]), .CO(C[481]) );
  FA_4414 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n997), .CI(C[481]), .CO(C[482]) );
  FA_4413 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n998), .CI(C[482]), .CO(C[483]) );
  FA_4412 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n999), .CI(C[483]), .CO(C[484]) );
  FA_4411 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n1000), .CI(
        C[484]), .CO(C[485]) );
  FA_4410 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n1001), .CI(
        C[485]), .CO(C[486]) );
  FA_4409 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n1002), .CI(
        C[486]), .CO(C[487]) );
  FA_4408 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n1003), .CI(
        C[487]), .CO(C[488]) );
  FA_4407 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n1004), .CI(
        C[488]), .CO(C[489]) );
  FA_4406 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n1005), .CI(
        C[489]), .CO(C[490]) );
  FA_4405 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n1006), .CI(
        C[490]), .CO(C[491]) );
  FA_4404 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n1007), .CI(
        C[491]), .CO(C[492]) );
  FA_4403 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n1008), .CI(
        C[492]), .CO(C[493]) );
  FA_4402 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n1009), .CI(
        C[493]), .CO(C[494]) );
  FA_4401 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n1010), .CI(
        C[494]), .CO(C[495]) );
  FA_4400 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n1011), .CI(
        C[495]), .CO(C[496]) );
  FA_4399 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n1012), .CI(
        C[496]), .CO(C[497]) );
  FA_4398 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n1013), .CI(
        C[497]), .CO(C[498]) );
  FA_4397 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n1014), .CI(
        C[498]), .CO(C[499]) );
  FA_4396 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n1015), .CI(
        C[499]), .CO(C[500]) );
  FA_4395 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n1016), .CI(
        C[500]), .CO(C[501]) );
  FA_4394 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n1017), .CI(
        C[501]), .CO(C[502]) );
  FA_4393 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n1018), .CI(
        C[502]), .CO(C[503]) );
  FA_4392 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n1019), .CI(
        C[503]), .CO(C[504]) );
  FA_4391 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n1020), .CI(
        C[504]), .CO(C[505]) );
  FA_4390 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n1021), .CI(
        C[505]), .CO(C[506]) );
  FA_4389 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n1022), .CI(
        C[506]), .CO(C[507]) );
  FA_4388 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n1023), .CI(
        C[507]), .CO(C[508]) );
  FA_4387 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n1024), .CI(
        C[508]), .CO(C[509]) );
  FA_4386 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n1025), .CI(
        C[509]), .CO(C[510]) );
  FA_4385 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n1026), .CI(
        C[510]), .CO(C[511]) );
  FA_4384 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n1027), .CI(
        C[511]), .CO(C[512]) );
  FA_4383 \FA_INST_1[512].FA_  ( .A(1'b0), .B(n1028), .CI(C[512]), .CO(C[513])
         );
  FA_4382 \FA_INST_1[513].FA_  ( .A(1'b0), .B(n1029), .CI(C[513]), .CO(O) );
  IV U2 ( .A(B[415]), .Z(n931) );
  IV U3 ( .A(B[416]), .Z(n932) );
  IV U4 ( .A(B[417]), .Z(n933) );
  IV U5 ( .A(B[418]), .Z(n934) );
  IV U6 ( .A(B[419]), .Z(n935) );
  IV U7 ( .A(B[420]), .Z(n936) );
  IV U8 ( .A(B[421]), .Z(n937) );
  IV U9 ( .A(B[422]), .Z(n938) );
  IV U10 ( .A(B[423]), .Z(n939) );
  IV U11 ( .A(B[424]), .Z(n940) );
  IV U12 ( .A(B[505]), .Z(n1021) );
  IV U13 ( .A(B[425]), .Z(n941) );
  IV U14 ( .A(B[426]), .Z(n942) );
  IV U15 ( .A(B[427]), .Z(n943) );
  IV U16 ( .A(B[428]), .Z(n944) );
  IV U17 ( .A(B[429]), .Z(n945) );
  IV U18 ( .A(B[430]), .Z(n946) );
  IV U19 ( .A(B[431]), .Z(n947) );
  IV U20 ( .A(B[432]), .Z(n948) );
  IV U21 ( .A(B[433]), .Z(n949) );
  IV U22 ( .A(B[434]), .Z(n950) );
  IV U23 ( .A(B[506]), .Z(n1022) );
  IV U24 ( .A(B[435]), .Z(n951) );
  IV U25 ( .A(B[436]), .Z(n952) );
  IV U26 ( .A(B[437]), .Z(n953) );
  IV U27 ( .A(B[438]), .Z(n954) );
  IV U28 ( .A(B[439]), .Z(n955) );
  IV U29 ( .A(B[440]), .Z(n956) );
  IV U30 ( .A(B[441]), .Z(n957) );
  IV U31 ( .A(B[442]), .Z(n958) );
  IV U32 ( .A(B[443]), .Z(n959) );
  IV U33 ( .A(B[444]), .Z(n960) );
  IV U34 ( .A(B[507]), .Z(n1023) );
  IV U35 ( .A(B[445]), .Z(n961) );
  IV U36 ( .A(B[446]), .Z(n962) );
  IV U37 ( .A(B[447]), .Z(n963) );
  IV U38 ( .A(B[448]), .Z(n964) );
  IV U39 ( .A(B[449]), .Z(n965) );
  IV U40 ( .A(B[450]), .Z(n966) );
  IV U41 ( .A(B[451]), .Z(n967) );
  IV U42 ( .A(B[452]), .Z(n968) );
  IV U43 ( .A(B[453]), .Z(n969) );
  IV U44 ( .A(B[454]), .Z(n970) );
  IV U45 ( .A(B[508]), .Z(n1024) );
  IV U46 ( .A(B[455]), .Z(n971) );
  IV U47 ( .A(B[456]), .Z(n972) );
  IV U48 ( .A(B[457]), .Z(n973) );
  IV U49 ( .A(B[458]), .Z(n974) );
  IV U50 ( .A(B[459]), .Z(n975) );
  IV U51 ( .A(B[460]), .Z(n976) );
  IV U52 ( .A(B[461]), .Z(n977) );
  IV U53 ( .A(B[462]), .Z(n978) );
  IV U54 ( .A(B[0]), .Z(n516) );
  IV U55 ( .A(B[1]), .Z(n517) );
  IV U56 ( .A(B[2]), .Z(n518) );
  IV U57 ( .A(B[3]), .Z(n519) );
  IV U58 ( .A(B[4]), .Z(n520) );
  IV U59 ( .A(B[463]), .Z(n979) );
  IV U60 ( .A(B[5]), .Z(n521) );
  IV U61 ( .A(B[6]), .Z(n522) );
  IV U62 ( .A(B[7]), .Z(n523) );
  IV U63 ( .A(B[8]), .Z(n524) );
  IV U64 ( .A(B[9]), .Z(n525) );
  IV U65 ( .A(B[10]), .Z(n526) );
  IV U66 ( .A(B[11]), .Z(n527) );
  IV U67 ( .A(B[12]), .Z(n528) );
  IV U68 ( .A(B[13]), .Z(n529) );
  IV U69 ( .A(B[14]), .Z(n530) );
  IV U70 ( .A(B[464]), .Z(n980) );
  IV U71 ( .A(B[509]), .Z(n1025) );
  IV U72 ( .A(B[15]), .Z(n531) );
  IV U73 ( .A(B[16]), .Z(n532) );
  IV U74 ( .A(B[17]), .Z(n533) );
  IV U75 ( .A(B[18]), .Z(n534) );
  IV U76 ( .A(B[19]), .Z(n535) );
  IV U77 ( .A(B[20]), .Z(n536) );
  IV U78 ( .A(B[21]), .Z(n537) );
  IV U79 ( .A(B[22]), .Z(n538) );
  IV U80 ( .A(B[23]), .Z(n539) );
  IV U81 ( .A(B[24]), .Z(n540) );
  IV U82 ( .A(B[465]), .Z(n981) );
  IV U83 ( .A(B[25]), .Z(n541) );
  IV U84 ( .A(B[26]), .Z(n542) );
  IV U85 ( .A(B[27]), .Z(n543) );
  IV U86 ( .A(B[28]), .Z(n544) );
  IV U87 ( .A(B[29]), .Z(n545) );
  IV U88 ( .A(B[30]), .Z(n546) );
  IV U89 ( .A(B[31]), .Z(n547) );
  IV U90 ( .A(B[32]), .Z(n548) );
  IV U91 ( .A(B[33]), .Z(n549) );
  IV U92 ( .A(B[34]), .Z(n550) );
  IV U93 ( .A(B[466]), .Z(n982) );
  IV U94 ( .A(B[35]), .Z(n551) );
  IV U95 ( .A(B[36]), .Z(n552) );
  IV U96 ( .A(B[37]), .Z(n553) );
  IV U97 ( .A(B[38]), .Z(n554) );
  IV U98 ( .A(B[39]), .Z(n555) );
  IV U99 ( .A(B[40]), .Z(n556) );
  IV U100 ( .A(B[41]), .Z(n557) );
  IV U101 ( .A(B[42]), .Z(n558) );
  IV U102 ( .A(B[43]), .Z(n559) );
  IV U103 ( .A(B[44]), .Z(n560) );
  IV U104 ( .A(B[467]), .Z(n983) );
  IV U105 ( .A(B[45]), .Z(n561) );
  IV U106 ( .A(B[46]), .Z(n562) );
  IV U107 ( .A(B[47]), .Z(n563) );
  IV U108 ( .A(B[48]), .Z(n564) );
  IV U109 ( .A(B[49]), .Z(n565) );
  IV U110 ( .A(B[50]), .Z(n566) );
  IV U111 ( .A(B[51]), .Z(n567) );
  IV U112 ( .A(B[52]), .Z(n568) );
  IV U113 ( .A(B[53]), .Z(n569) );
  IV U114 ( .A(B[54]), .Z(n570) );
  IV U115 ( .A(B[468]), .Z(n984) );
  IV U116 ( .A(B[55]), .Z(n571) );
  IV U117 ( .A(B[56]), .Z(n572) );
  IV U118 ( .A(B[57]), .Z(n573) );
  IV U119 ( .A(B[58]), .Z(n574) );
  IV U120 ( .A(B[59]), .Z(n575) );
  IV U121 ( .A(B[60]), .Z(n576) );
  IV U122 ( .A(B[61]), .Z(n577) );
  IV U123 ( .A(B[62]), .Z(n578) );
  IV U124 ( .A(B[63]), .Z(n579) );
  IV U125 ( .A(B[64]), .Z(n580) );
  IV U126 ( .A(B[469]), .Z(n985) );
  IV U127 ( .A(B[65]), .Z(n581) );
  IV U128 ( .A(B[66]), .Z(n582) );
  IV U129 ( .A(B[67]), .Z(n583) );
  IV U130 ( .A(B[68]), .Z(n584) );
  IV U131 ( .A(B[69]), .Z(n585) );
  IV U132 ( .A(B[70]), .Z(n586) );
  IV U133 ( .A(B[71]), .Z(n587) );
  IV U134 ( .A(B[72]), .Z(n588) );
  IV U135 ( .A(B[73]), .Z(n589) );
  IV U136 ( .A(B[74]), .Z(n590) );
  IV U137 ( .A(B[470]), .Z(n986) );
  IV U138 ( .A(B[75]), .Z(n591) );
  IV U139 ( .A(B[76]), .Z(n592) );
  IV U140 ( .A(B[77]), .Z(n593) );
  IV U141 ( .A(B[78]), .Z(n594) );
  IV U142 ( .A(B[79]), .Z(n595) );
  IV U143 ( .A(B[80]), .Z(n596) );
  IV U144 ( .A(B[81]), .Z(n597) );
  IV U145 ( .A(B[82]), .Z(n598) );
  IV U146 ( .A(B[83]), .Z(n599) );
  IV U147 ( .A(B[84]), .Z(n600) );
  IV U148 ( .A(B[471]), .Z(n987) );
  IV U149 ( .A(B[85]), .Z(n601) );
  IV U150 ( .A(B[86]), .Z(n602) );
  IV U151 ( .A(B[87]), .Z(n603) );
  IV U152 ( .A(B[88]), .Z(n604) );
  IV U153 ( .A(B[89]), .Z(n605) );
  IV U154 ( .A(B[90]), .Z(n606) );
  IV U155 ( .A(B[91]), .Z(n607) );
  IV U156 ( .A(B[92]), .Z(n608) );
  IV U157 ( .A(B[93]), .Z(n609) );
  IV U158 ( .A(B[94]), .Z(n610) );
  IV U159 ( .A(B[472]), .Z(n988) );
  IV U160 ( .A(B[95]), .Z(n611) );
  IV U161 ( .A(B[96]), .Z(n612) );
  IV U162 ( .A(B[97]), .Z(n613) );
  IV U163 ( .A(B[98]), .Z(n614) );
  IV U164 ( .A(B[99]), .Z(n615) );
  IV U165 ( .A(B[100]), .Z(n616) );
  IV U166 ( .A(B[101]), .Z(n617) );
  IV U167 ( .A(B[102]), .Z(n618) );
  IV U168 ( .A(B[103]), .Z(n619) );
  IV U169 ( .A(B[104]), .Z(n620) );
  IV U170 ( .A(B[473]), .Z(n989) );
  IV U171 ( .A(B[105]), .Z(n621) );
  IV U172 ( .A(B[106]), .Z(n622) );
  IV U173 ( .A(B[107]), .Z(n623) );
  IV U174 ( .A(B[108]), .Z(n624) );
  IV U175 ( .A(B[109]), .Z(n625) );
  IV U176 ( .A(B[110]), .Z(n626) );
  IV U177 ( .A(B[111]), .Z(n627) );
  IV U178 ( .A(B[112]), .Z(n628) );
  IV U179 ( .A(B[113]), .Z(n629) );
  IV U180 ( .A(B[114]), .Z(n630) );
  IV U181 ( .A(B[474]), .Z(n990) );
  IV U182 ( .A(B[510]), .Z(n1026) );
  IV U183 ( .A(B[115]), .Z(n631) );
  IV U184 ( .A(B[116]), .Z(n632) );
  IV U185 ( .A(B[117]), .Z(n633) );
  IV U186 ( .A(B[118]), .Z(n634) );
  IV U187 ( .A(B[119]), .Z(n635) );
  IV U188 ( .A(B[120]), .Z(n636) );
  IV U189 ( .A(B[121]), .Z(n637) );
  IV U190 ( .A(B[122]), .Z(n638) );
  IV U191 ( .A(B[123]), .Z(n639) );
  IV U192 ( .A(B[124]), .Z(n640) );
  IV U193 ( .A(B[475]), .Z(n991) );
  IV U194 ( .A(B[125]), .Z(n641) );
  IV U195 ( .A(B[126]), .Z(n642) );
  IV U196 ( .A(B[127]), .Z(n643) );
  IV U197 ( .A(B[128]), .Z(n644) );
  IV U198 ( .A(B[129]), .Z(n645) );
  IV U199 ( .A(B[130]), .Z(n646) );
  IV U200 ( .A(B[131]), .Z(n647) );
  IV U201 ( .A(B[132]), .Z(n648) );
  IV U202 ( .A(B[133]), .Z(n649) );
  IV U203 ( .A(B[134]), .Z(n650) );
  IV U204 ( .A(B[476]), .Z(n992) );
  IV U205 ( .A(B[135]), .Z(n651) );
  IV U206 ( .A(B[136]), .Z(n652) );
  IV U207 ( .A(B[137]), .Z(n653) );
  IV U208 ( .A(B[138]), .Z(n654) );
  IV U209 ( .A(B[139]), .Z(n655) );
  IV U210 ( .A(B[140]), .Z(n656) );
  IV U211 ( .A(B[141]), .Z(n657) );
  IV U212 ( .A(B[142]), .Z(n658) );
  IV U213 ( .A(B[143]), .Z(n659) );
  IV U214 ( .A(B[144]), .Z(n660) );
  IV U215 ( .A(B[477]), .Z(n993) );
  IV U216 ( .A(B[145]), .Z(n661) );
  IV U217 ( .A(B[146]), .Z(n662) );
  IV U218 ( .A(B[147]), .Z(n663) );
  IV U219 ( .A(B[148]), .Z(n664) );
  IV U220 ( .A(B[149]), .Z(n665) );
  IV U221 ( .A(B[150]), .Z(n666) );
  IV U222 ( .A(B[151]), .Z(n667) );
  IV U223 ( .A(B[152]), .Z(n668) );
  IV U224 ( .A(B[153]), .Z(n669) );
  IV U225 ( .A(B[154]), .Z(n670) );
  IV U226 ( .A(B[478]), .Z(n994) );
  IV U227 ( .A(B[155]), .Z(n671) );
  IV U228 ( .A(B[156]), .Z(n672) );
  IV U229 ( .A(B[157]), .Z(n673) );
  IV U230 ( .A(B[158]), .Z(n674) );
  IV U231 ( .A(B[159]), .Z(n675) );
  IV U232 ( .A(B[160]), .Z(n676) );
  IV U233 ( .A(B[161]), .Z(n677) );
  IV U234 ( .A(B[162]), .Z(n678) );
  IV U235 ( .A(B[163]), .Z(n679) );
  IV U236 ( .A(B[164]), .Z(n680) );
  IV U237 ( .A(B[479]), .Z(n995) );
  IV U238 ( .A(B[165]), .Z(n681) );
  IV U239 ( .A(B[166]), .Z(n682) );
  IV U240 ( .A(B[167]), .Z(n683) );
  IV U241 ( .A(B[168]), .Z(n684) );
  IV U242 ( .A(B[169]), .Z(n685) );
  IV U243 ( .A(B[170]), .Z(n686) );
  IV U244 ( .A(B[171]), .Z(n687) );
  IV U245 ( .A(B[172]), .Z(n688) );
  IV U246 ( .A(B[173]), .Z(n689) );
  IV U247 ( .A(B[174]), .Z(n690) );
  IV U248 ( .A(B[480]), .Z(n996) );
  IV U249 ( .A(B[175]), .Z(n691) );
  IV U250 ( .A(B[176]), .Z(n692) );
  IV U251 ( .A(B[177]), .Z(n693) );
  IV U252 ( .A(B[178]), .Z(n694) );
  IV U253 ( .A(B[179]), .Z(n695) );
  IV U254 ( .A(B[180]), .Z(n696) );
  IV U255 ( .A(B[181]), .Z(n697) );
  IV U256 ( .A(B[182]), .Z(n698) );
  IV U257 ( .A(B[183]), .Z(n699) );
  IV U258 ( .A(B[184]), .Z(n700) );
  IV U259 ( .A(B[481]), .Z(n997) );
  IV U260 ( .A(B[185]), .Z(n701) );
  IV U261 ( .A(B[186]), .Z(n702) );
  IV U262 ( .A(B[187]), .Z(n703) );
  IV U263 ( .A(B[188]), .Z(n704) );
  IV U264 ( .A(B[189]), .Z(n705) );
  IV U265 ( .A(B[190]), .Z(n706) );
  IV U266 ( .A(B[191]), .Z(n707) );
  IV U267 ( .A(B[192]), .Z(n708) );
  IV U268 ( .A(B[193]), .Z(n709) );
  IV U269 ( .A(B[194]), .Z(n710) );
  IV U270 ( .A(B[482]), .Z(n998) );
  IV U271 ( .A(B[195]), .Z(n711) );
  IV U272 ( .A(B[196]), .Z(n712) );
  IV U273 ( .A(B[197]), .Z(n713) );
  IV U274 ( .A(B[198]), .Z(n714) );
  IV U275 ( .A(B[199]), .Z(n715) );
  IV U276 ( .A(B[200]), .Z(n716) );
  IV U277 ( .A(B[201]), .Z(n717) );
  IV U278 ( .A(B[202]), .Z(n718) );
  IV U279 ( .A(B[203]), .Z(n719) );
  IV U280 ( .A(B[204]), .Z(n720) );
  IV U281 ( .A(B[483]), .Z(n999) );
  IV U282 ( .A(B[205]), .Z(n721) );
  IV U283 ( .A(B[206]), .Z(n722) );
  IV U284 ( .A(B[207]), .Z(n723) );
  IV U285 ( .A(B[208]), .Z(n724) );
  IV U286 ( .A(B[209]), .Z(n725) );
  IV U287 ( .A(B[210]), .Z(n726) );
  IV U288 ( .A(B[211]), .Z(n727) );
  IV U289 ( .A(B[212]), .Z(n728) );
  IV U290 ( .A(B[213]), .Z(n729) );
  IV U291 ( .A(B[214]), .Z(n730) );
  IV U292 ( .A(B[484]), .Z(n1000) );
  IV U293 ( .A(B[511]), .Z(n1027) );
  IV U294 ( .A(B[215]), .Z(n731) );
  IV U295 ( .A(B[216]), .Z(n732) );
  IV U296 ( .A(B[217]), .Z(n733) );
  IV U297 ( .A(B[218]), .Z(n734) );
  IV U298 ( .A(B[219]), .Z(n735) );
  IV U299 ( .A(B[220]), .Z(n736) );
  IV U300 ( .A(B[221]), .Z(n737) );
  IV U301 ( .A(B[222]), .Z(n738) );
  IV U302 ( .A(B[223]), .Z(n739) );
  IV U303 ( .A(B[224]), .Z(n740) );
  IV U304 ( .A(B[485]), .Z(n1001) );
  IV U305 ( .A(B[225]), .Z(n741) );
  IV U306 ( .A(B[226]), .Z(n742) );
  IV U307 ( .A(B[227]), .Z(n743) );
  IV U308 ( .A(B[228]), .Z(n744) );
  IV U309 ( .A(B[229]), .Z(n745) );
  IV U310 ( .A(B[230]), .Z(n746) );
  IV U311 ( .A(B[231]), .Z(n747) );
  IV U312 ( .A(B[232]), .Z(n748) );
  IV U313 ( .A(B[233]), .Z(n749) );
  IV U314 ( .A(B[234]), .Z(n750) );
  IV U315 ( .A(B[486]), .Z(n1002) );
  IV U316 ( .A(B[235]), .Z(n751) );
  IV U317 ( .A(B[236]), .Z(n752) );
  IV U318 ( .A(B[237]), .Z(n753) );
  IV U319 ( .A(B[238]), .Z(n754) );
  IV U320 ( .A(B[239]), .Z(n755) );
  IV U321 ( .A(B[240]), .Z(n756) );
  IV U322 ( .A(B[241]), .Z(n757) );
  IV U323 ( .A(B[242]), .Z(n758) );
  IV U324 ( .A(B[243]), .Z(n759) );
  IV U325 ( .A(B[244]), .Z(n760) );
  IV U326 ( .A(B[487]), .Z(n1003) );
  IV U327 ( .A(B[245]), .Z(n761) );
  IV U328 ( .A(B[246]), .Z(n762) );
  IV U329 ( .A(B[247]), .Z(n763) );
  IV U330 ( .A(B[248]), .Z(n764) );
  IV U331 ( .A(B[249]), .Z(n765) );
  IV U332 ( .A(B[250]), .Z(n766) );
  IV U333 ( .A(B[251]), .Z(n767) );
  IV U334 ( .A(B[252]), .Z(n768) );
  IV U335 ( .A(B[253]), .Z(n769) );
  IV U336 ( .A(B[254]), .Z(n770) );
  IV U337 ( .A(B[488]), .Z(n1004) );
  IV U338 ( .A(B[255]), .Z(n771) );
  IV U339 ( .A(B[256]), .Z(n772) );
  IV U340 ( .A(B[257]), .Z(n773) );
  IV U341 ( .A(B[258]), .Z(n774) );
  IV U342 ( .A(B[259]), .Z(n775) );
  IV U343 ( .A(B[260]), .Z(n776) );
  IV U344 ( .A(B[261]), .Z(n777) );
  IV U345 ( .A(B[262]), .Z(n778) );
  IV U346 ( .A(B[263]), .Z(n779) );
  IV U347 ( .A(B[264]), .Z(n780) );
  IV U348 ( .A(B[489]), .Z(n1005) );
  IV U349 ( .A(B[265]), .Z(n781) );
  IV U350 ( .A(B[266]), .Z(n782) );
  IV U351 ( .A(B[267]), .Z(n783) );
  IV U352 ( .A(B[268]), .Z(n784) );
  IV U353 ( .A(B[269]), .Z(n785) );
  IV U354 ( .A(B[270]), .Z(n786) );
  IV U355 ( .A(B[271]), .Z(n787) );
  IV U356 ( .A(B[272]), .Z(n788) );
  IV U357 ( .A(B[273]), .Z(n789) );
  IV U358 ( .A(B[274]), .Z(n790) );
  IV U359 ( .A(B[490]), .Z(n1006) );
  IV U360 ( .A(B[275]), .Z(n791) );
  IV U361 ( .A(B[276]), .Z(n792) );
  IV U362 ( .A(B[277]), .Z(n793) );
  IV U363 ( .A(B[278]), .Z(n794) );
  IV U364 ( .A(B[279]), .Z(n795) );
  IV U365 ( .A(B[280]), .Z(n796) );
  IV U366 ( .A(B[281]), .Z(n797) );
  IV U367 ( .A(B[282]), .Z(n798) );
  IV U368 ( .A(B[283]), .Z(n799) );
  IV U369 ( .A(B[284]), .Z(n800) );
  IV U370 ( .A(B[491]), .Z(n1007) );
  IV U371 ( .A(B[285]), .Z(n801) );
  IV U372 ( .A(B[286]), .Z(n802) );
  IV U373 ( .A(B[287]), .Z(n803) );
  IV U374 ( .A(B[288]), .Z(n804) );
  IV U375 ( .A(B[289]), .Z(n805) );
  IV U376 ( .A(B[290]), .Z(n806) );
  IV U377 ( .A(B[291]), .Z(n807) );
  IV U378 ( .A(B[292]), .Z(n808) );
  IV U379 ( .A(B[293]), .Z(n809) );
  IV U380 ( .A(B[294]), .Z(n810) );
  IV U381 ( .A(B[492]), .Z(n1008) );
  IV U382 ( .A(B[295]), .Z(n811) );
  IV U383 ( .A(B[296]), .Z(n812) );
  IV U384 ( .A(B[297]), .Z(n813) );
  IV U385 ( .A(B[298]), .Z(n814) );
  IV U386 ( .A(B[299]), .Z(n815) );
  IV U387 ( .A(B[300]), .Z(n816) );
  IV U388 ( .A(B[301]), .Z(n817) );
  IV U389 ( .A(B[302]), .Z(n818) );
  IV U390 ( .A(B[303]), .Z(n819) );
  IV U391 ( .A(B[304]), .Z(n820) );
  IV U392 ( .A(B[493]), .Z(n1009) );
  IV U393 ( .A(B[305]), .Z(n821) );
  IV U394 ( .A(B[306]), .Z(n822) );
  IV U395 ( .A(B[307]), .Z(n823) );
  IV U396 ( .A(B[308]), .Z(n824) );
  IV U397 ( .A(B[309]), .Z(n825) );
  IV U398 ( .A(B[310]), .Z(n826) );
  IV U399 ( .A(B[311]), .Z(n827) );
  IV U400 ( .A(B[312]), .Z(n828) );
  IV U401 ( .A(B[313]), .Z(n829) );
  IV U402 ( .A(B[314]), .Z(n830) );
  IV U403 ( .A(B[494]), .Z(n1010) );
  IV U404 ( .A(B[512]), .Z(n1028) );
  IV U405 ( .A(B[315]), .Z(n831) );
  IV U406 ( .A(B[316]), .Z(n832) );
  IV U407 ( .A(B[317]), .Z(n833) );
  IV U408 ( .A(B[318]), .Z(n834) );
  IV U409 ( .A(B[319]), .Z(n835) );
  IV U410 ( .A(B[320]), .Z(n836) );
  IV U411 ( .A(B[321]), .Z(n837) );
  IV U412 ( .A(B[322]), .Z(n838) );
  IV U413 ( .A(B[323]), .Z(n839) );
  IV U414 ( .A(B[324]), .Z(n840) );
  IV U415 ( .A(B[495]), .Z(n1011) );
  IV U416 ( .A(B[325]), .Z(n841) );
  IV U417 ( .A(B[326]), .Z(n842) );
  IV U418 ( .A(B[327]), .Z(n843) );
  IV U419 ( .A(B[328]), .Z(n844) );
  IV U420 ( .A(B[329]), .Z(n845) );
  IV U421 ( .A(B[330]), .Z(n846) );
  IV U422 ( .A(B[331]), .Z(n847) );
  IV U423 ( .A(B[332]), .Z(n848) );
  IV U424 ( .A(B[333]), .Z(n849) );
  IV U425 ( .A(B[334]), .Z(n850) );
  IV U426 ( .A(B[496]), .Z(n1012) );
  IV U427 ( .A(B[335]), .Z(n851) );
  IV U428 ( .A(B[336]), .Z(n852) );
  IV U429 ( .A(B[337]), .Z(n853) );
  IV U430 ( .A(B[338]), .Z(n854) );
  IV U431 ( .A(B[339]), .Z(n855) );
  IV U432 ( .A(B[340]), .Z(n856) );
  IV U433 ( .A(B[341]), .Z(n857) );
  IV U434 ( .A(B[342]), .Z(n858) );
  IV U435 ( .A(B[343]), .Z(n859) );
  IV U436 ( .A(B[344]), .Z(n860) );
  IV U437 ( .A(B[497]), .Z(n1013) );
  IV U438 ( .A(B[345]), .Z(n861) );
  IV U439 ( .A(B[346]), .Z(n862) );
  IV U440 ( .A(B[347]), .Z(n863) );
  IV U441 ( .A(B[348]), .Z(n864) );
  IV U442 ( .A(B[349]), .Z(n865) );
  IV U443 ( .A(B[350]), .Z(n866) );
  IV U444 ( .A(B[351]), .Z(n867) );
  IV U445 ( .A(B[352]), .Z(n868) );
  IV U446 ( .A(B[353]), .Z(n869) );
  IV U447 ( .A(B[354]), .Z(n870) );
  IV U448 ( .A(B[498]), .Z(n1014) );
  IV U449 ( .A(B[355]), .Z(n871) );
  IV U450 ( .A(B[356]), .Z(n872) );
  IV U451 ( .A(B[357]), .Z(n873) );
  IV U452 ( .A(B[358]), .Z(n874) );
  IV U453 ( .A(B[359]), .Z(n875) );
  IV U454 ( .A(B[360]), .Z(n876) );
  IV U455 ( .A(B[361]), .Z(n877) );
  IV U456 ( .A(B[362]), .Z(n878) );
  IV U457 ( .A(B[363]), .Z(n879) );
  IV U458 ( .A(B[364]), .Z(n880) );
  IV U459 ( .A(B[499]), .Z(n1015) );
  IV U460 ( .A(B[365]), .Z(n881) );
  IV U461 ( .A(B[366]), .Z(n882) );
  IV U462 ( .A(B[367]), .Z(n883) );
  IV U463 ( .A(B[368]), .Z(n884) );
  IV U464 ( .A(B[369]), .Z(n885) );
  IV U465 ( .A(B[370]), .Z(n886) );
  IV U466 ( .A(B[371]), .Z(n887) );
  IV U467 ( .A(B[372]), .Z(n888) );
  IV U468 ( .A(B[373]), .Z(n889) );
  IV U469 ( .A(B[374]), .Z(n890) );
  IV U470 ( .A(B[500]), .Z(n1016) );
  IV U471 ( .A(B[375]), .Z(n891) );
  IV U472 ( .A(B[376]), .Z(n892) );
  IV U473 ( .A(B[377]), .Z(n893) );
  IV U474 ( .A(B[378]), .Z(n894) );
  IV U475 ( .A(B[379]), .Z(n895) );
  IV U476 ( .A(B[380]), .Z(n896) );
  IV U477 ( .A(B[381]), .Z(n897) );
  IV U478 ( .A(B[382]), .Z(n898) );
  IV U479 ( .A(B[383]), .Z(n899) );
  IV U480 ( .A(B[384]), .Z(n900) );
  IV U481 ( .A(B[501]), .Z(n1017) );
  IV U482 ( .A(B[385]), .Z(n901) );
  IV U483 ( .A(B[386]), .Z(n902) );
  IV U484 ( .A(B[387]), .Z(n903) );
  IV U485 ( .A(B[388]), .Z(n904) );
  IV U486 ( .A(B[389]), .Z(n905) );
  IV U487 ( .A(B[390]), .Z(n906) );
  IV U488 ( .A(B[391]), .Z(n907) );
  IV U489 ( .A(B[392]), .Z(n908) );
  IV U490 ( .A(B[393]), .Z(n909) );
  IV U491 ( .A(B[394]), .Z(n910) );
  IV U492 ( .A(B[502]), .Z(n1018) );
  IV U493 ( .A(B[395]), .Z(n911) );
  IV U494 ( .A(B[396]), .Z(n912) );
  IV U495 ( .A(B[397]), .Z(n913) );
  IV U496 ( .A(B[398]), .Z(n914) );
  IV U497 ( .A(B[399]), .Z(n915) );
  IV U498 ( .A(B[400]), .Z(n916) );
  IV U499 ( .A(B[401]), .Z(n917) );
  IV U500 ( .A(B[402]), .Z(n918) );
  IV U501 ( .A(B[403]), .Z(n919) );
  IV U502 ( .A(B[404]), .Z(n920) );
  IV U503 ( .A(B[503]), .Z(n1019) );
  IV U504 ( .A(B[405]), .Z(n921) );
  IV U505 ( .A(B[406]), .Z(n922) );
  IV U506 ( .A(B[407]), .Z(n923) );
  IV U507 ( .A(B[408]), .Z(n924) );
  IV U508 ( .A(B[409]), .Z(n925) );
  IV U509 ( .A(B[410]), .Z(n926) );
  IV U510 ( .A(B[411]), .Z(n927) );
  IV U511 ( .A(B[412]), .Z(n928) );
  IV U512 ( .A(B[413]), .Z(n929) );
  IV U513 ( .A(B[414]), .Z(n930) );
  IV U514 ( .A(B[504]), .Z(n1020) );
  IV U515 ( .A(B[513]), .Z(n1029) );
endmodule


module FA_3869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_3870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N514_1 ( A, B, S, CO );
  input [513:0] A;
  input [513:0] B;
  output [513:0] S;
  output CO;
  wire   n2, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  wire   [513:1] C;

  FA_4381 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n2), .CI(1'b1), .S(
        S[0]), .CO(C[1]) );
  FA_4380 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n514), .CI(C[1]), .S(
        S[1]), .CO(C[2]) );
  FA_4379 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n515), .CI(C[2]), .S(
        S[2]), .CO(C[3]) );
  FA_4378 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n516), .CI(C[3]), .S(
        S[3]), .CO(C[4]) );
  FA_4377 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n517), .CI(C[4]), .S(
        S[4]), .CO(C[5]) );
  FA_4376 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n518), .CI(C[5]), .S(
        S[5]), .CO(C[6]) );
  FA_4375 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n519), .CI(C[6]), .S(
        S[6]), .CO(C[7]) );
  FA_4374 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n520), .CI(C[7]), .S(
        S[7]), .CO(C[8]) );
  FA_4373 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n521), .CI(C[8]), .S(
        S[8]), .CO(C[9]) );
  FA_4372 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n522), .CI(C[9]), .S(
        S[9]), .CO(C[10]) );
  FA_4371 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n523), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_4370 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n524), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_4369 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n525), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_4368 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n526), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_4367 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n527), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_4366 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n528), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_4365 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n529), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_4364 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n530), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_4363 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n531), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_4362 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n532), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_4361 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n533), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_4360 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n534), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_4359 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n535), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_4358 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n536), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_4357 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n537), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_4356 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n538), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_4355 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n539), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_4354 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n540), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_4353 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n541), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_4352 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n542), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_4351 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n543), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_4350 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n544), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_4349 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n545), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_4348 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n546), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_4347 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n547), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_4346 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n548), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_4345 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n549), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_4344 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n550), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_4343 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n551), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_4342 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n552), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_4341 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n553), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_4340 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n554), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_4339 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n555), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_4338 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n556), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_4337 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n557), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_4336 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n558), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_4335 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n559), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_4334 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n560), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_4333 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n561), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_4332 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n562), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_4331 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n563), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_4330 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n564), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_4329 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n565), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_4328 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n566), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_4327 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n567), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_4326 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n568), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_4325 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n569), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_4324 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n570), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_4323 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n571), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_4322 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n572), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_4321 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n573), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_4320 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n574), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_4319 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n575), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_4318 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n576), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_4317 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n577), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_4316 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n578), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_4315 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n579), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_4314 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n580), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_4313 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n581), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_4312 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n582), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_4311 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n583), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_4310 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n584), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_4309 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n585), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_4308 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n586), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_4307 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n587), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_4306 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n588), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_4305 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n589), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_4304 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n590), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_4303 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n591), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_4302 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n592), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_4301 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n593), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_4300 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n594), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_4299 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n595), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_4298 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n596), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_4297 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n597), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_4296 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n598), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_4295 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n599), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_4294 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n600), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_4293 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n601), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_4292 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n602), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_4291 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n603), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_4290 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n604), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_4289 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n605), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_4288 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n606), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_4287 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n607), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_4286 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n608), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_4285 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n609), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_4284 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n610), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_4283 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n611), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_4282 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n612), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_4281 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n613), .CI(C[100]), .S(S[100]), .CO(C[101]) );
  FA_4280 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n614), .CI(C[101]), .S(S[101]), .CO(C[102]) );
  FA_4279 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n615), .CI(C[102]), .S(S[102]), .CO(C[103]) );
  FA_4278 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n616), .CI(C[103]), .S(S[103]), .CO(C[104]) );
  FA_4277 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n617), .CI(C[104]), .S(S[104]), .CO(C[105]) );
  FA_4276 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n618), .CI(C[105]), .S(S[105]), .CO(C[106]) );
  FA_4275 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n619), .CI(C[106]), .S(S[106]), .CO(C[107]) );
  FA_4274 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n620), .CI(C[107]), .S(S[107]), .CO(C[108]) );
  FA_4273 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n621), .CI(C[108]), .S(S[108]), .CO(C[109]) );
  FA_4272 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n622), .CI(C[109]), .S(S[109]), .CO(C[110]) );
  FA_4271 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n623), .CI(C[110]), .S(S[110]), .CO(C[111]) );
  FA_4270 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n624), .CI(C[111]), .S(S[111]), .CO(C[112]) );
  FA_4269 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n625), .CI(C[112]), .S(S[112]), .CO(C[113]) );
  FA_4268 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n626), .CI(C[113]), .S(S[113]), .CO(C[114]) );
  FA_4267 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n627), .CI(C[114]), .S(S[114]), .CO(C[115]) );
  FA_4266 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n628), .CI(C[115]), .S(S[115]), .CO(C[116]) );
  FA_4265 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n629), .CI(C[116]), .S(S[116]), .CO(C[117]) );
  FA_4264 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n630), .CI(C[117]), .S(S[117]), .CO(C[118]) );
  FA_4263 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n631), .CI(C[118]), .S(S[118]), .CO(C[119]) );
  FA_4262 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n632), .CI(C[119]), .S(S[119]), .CO(C[120]) );
  FA_4261 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n633), .CI(C[120]), .S(S[120]), .CO(C[121]) );
  FA_4260 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n634), .CI(C[121]), .S(S[121]), .CO(C[122]) );
  FA_4259 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n635), .CI(C[122]), .S(S[122]), .CO(C[123]) );
  FA_4258 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n636), .CI(C[123]), .S(S[123]), .CO(C[124]) );
  FA_4257 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n637), .CI(C[124]), .S(S[124]), .CO(C[125]) );
  FA_4256 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n638), .CI(C[125]), .S(S[125]), .CO(C[126]) );
  FA_4255 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n639), .CI(C[126]), .S(S[126]), .CO(C[127]) );
  FA_4254 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n640), .CI(C[127]), .S(S[127]), .CO(C[128]) );
  FA_4253 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n641), .CI(C[128]), .S(S[128]), .CO(C[129]) );
  FA_4252 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n642), .CI(C[129]), .S(S[129]), .CO(C[130]) );
  FA_4251 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n643), .CI(C[130]), .S(S[130]), .CO(C[131]) );
  FA_4250 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n644), .CI(C[131]), .S(S[131]), .CO(C[132]) );
  FA_4249 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n645), .CI(C[132]), .S(S[132]), .CO(C[133]) );
  FA_4248 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n646), .CI(C[133]), .S(S[133]), .CO(C[134]) );
  FA_4247 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n647), .CI(C[134]), .S(S[134]), .CO(C[135]) );
  FA_4246 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n648), .CI(C[135]), .S(S[135]), .CO(C[136]) );
  FA_4245 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n649), .CI(C[136]), .S(S[136]), .CO(C[137]) );
  FA_4244 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n650), .CI(C[137]), .S(S[137]), .CO(C[138]) );
  FA_4243 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n651), .CI(C[138]), .S(S[138]), .CO(C[139]) );
  FA_4242 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n652), .CI(C[139]), .S(S[139]), .CO(C[140]) );
  FA_4241 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n653), .CI(C[140]), .S(S[140]), .CO(C[141]) );
  FA_4240 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n654), .CI(C[141]), .S(S[141]), .CO(C[142]) );
  FA_4239 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n655), .CI(C[142]), .S(S[142]), .CO(C[143]) );
  FA_4238 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n656), .CI(C[143]), .S(S[143]), .CO(C[144]) );
  FA_4237 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n657), .CI(C[144]), .S(S[144]), .CO(C[145]) );
  FA_4236 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n658), .CI(C[145]), .S(S[145]), .CO(C[146]) );
  FA_4235 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n659), .CI(C[146]), .S(S[146]), .CO(C[147]) );
  FA_4234 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n660), .CI(C[147]), .S(S[147]), .CO(C[148]) );
  FA_4233 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n661), .CI(C[148]), .S(S[148]), .CO(C[149]) );
  FA_4232 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n662), .CI(C[149]), .S(S[149]), .CO(C[150]) );
  FA_4231 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n663), .CI(C[150]), .S(S[150]), .CO(C[151]) );
  FA_4230 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n664), .CI(C[151]), .S(S[151]), .CO(C[152]) );
  FA_4229 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n665), .CI(C[152]), .S(S[152]), .CO(C[153]) );
  FA_4228 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n666), .CI(C[153]), .S(S[153]), .CO(C[154]) );
  FA_4227 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n667), .CI(C[154]), .S(S[154]), .CO(C[155]) );
  FA_4226 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n668), .CI(C[155]), .S(S[155]), .CO(C[156]) );
  FA_4225 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n669), .CI(C[156]), .S(S[156]), .CO(C[157]) );
  FA_4224 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n670), .CI(C[157]), .S(S[157]), .CO(C[158]) );
  FA_4223 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n671), .CI(C[158]), .S(S[158]), .CO(C[159]) );
  FA_4222 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n672), .CI(C[159]), .S(S[159]), .CO(C[160]) );
  FA_4221 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n673), .CI(C[160]), .S(S[160]), .CO(C[161]) );
  FA_4220 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n674), .CI(C[161]), .S(S[161]), .CO(C[162]) );
  FA_4219 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n675), .CI(C[162]), .S(S[162]), .CO(C[163]) );
  FA_4218 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n676), .CI(C[163]), .S(S[163]), .CO(C[164]) );
  FA_4217 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n677), .CI(C[164]), .S(S[164]), .CO(C[165]) );
  FA_4216 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n678), .CI(C[165]), .S(S[165]), .CO(C[166]) );
  FA_4215 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n679), .CI(C[166]), .S(S[166]), .CO(C[167]) );
  FA_4214 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n680), .CI(C[167]), .S(S[167]), .CO(C[168]) );
  FA_4213 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n681), .CI(C[168]), .S(S[168]), .CO(C[169]) );
  FA_4212 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n682), .CI(C[169]), .S(S[169]), .CO(C[170]) );
  FA_4211 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n683), .CI(C[170]), .S(S[170]), .CO(C[171]) );
  FA_4210 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n684), .CI(C[171]), .S(S[171]), .CO(C[172]) );
  FA_4209 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n685), .CI(C[172]), .S(S[172]), .CO(C[173]) );
  FA_4208 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n686), .CI(C[173]), .S(S[173]), .CO(C[174]) );
  FA_4207 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n687), .CI(C[174]), .S(S[174]), .CO(C[175]) );
  FA_4206 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n688), .CI(C[175]), .S(S[175]), .CO(C[176]) );
  FA_4205 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n689), .CI(C[176]), .S(S[176]), .CO(C[177]) );
  FA_4204 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n690), .CI(C[177]), .S(S[177]), .CO(C[178]) );
  FA_4203 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n691), .CI(C[178]), .S(S[178]), .CO(C[179]) );
  FA_4202 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n692), .CI(C[179]), .S(S[179]), .CO(C[180]) );
  FA_4201 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n693), .CI(C[180]), .S(S[180]), .CO(C[181]) );
  FA_4200 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n694), .CI(C[181]), .S(S[181]), .CO(C[182]) );
  FA_4199 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n695), .CI(C[182]), .S(S[182]), .CO(C[183]) );
  FA_4198 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n696), .CI(C[183]), .S(S[183]), .CO(C[184]) );
  FA_4197 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n697), .CI(C[184]), .S(S[184]), .CO(C[185]) );
  FA_4196 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n698), .CI(C[185]), .S(S[185]), .CO(C[186]) );
  FA_4195 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n699), .CI(C[186]), .S(S[186]), .CO(C[187]) );
  FA_4194 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n700), .CI(C[187]), .S(S[187]), .CO(C[188]) );
  FA_4193 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n701), .CI(C[188]), .S(S[188]), .CO(C[189]) );
  FA_4192 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n702), .CI(C[189]), .S(S[189]), .CO(C[190]) );
  FA_4191 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n703), .CI(C[190]), .S(S[190]), .CO(C[191]) );
  FA_4190 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n704), .CI(C[191]), .S(S[191]), .CO(C[192]) );
  FA_4189 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n705), .CI(C[192]), .S(S[192]), .CO(C[193]) );
  FA_4188 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n706), .CI(C[193]), .S(S[193]), .CO(C[194]) );
  FA_4187 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n707), .CI(C[194]), .S(S[194]), .CO(C[195]) );
  FA_4186 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n708), .CI(C[195]), .S(S[195]), .CO(C[196]) );
  FA_4185 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n709), .CI(C[196]), .S(S[196]), .CO(C[197]) );
  FA_4184 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n710), .CI(C[197]), .S(S[197]), .CO(C[198]) );
  FA_4183 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n711), .CI(C[198]), .S(S[198]), .CO(C[199]) );
  FA_4182 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n712), .CI(C[199]), .S(S[199]), .CO(C[200]) );
  FA_4181 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n713), .CI(C[200]), .S(S[200]), .CO(C[201]) );
  FA_4180 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n714), .CI(C[201]), .S(S[201]), .CO(C[202]) );
  FA_4179 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n715), .CI(C[202]), .S(S[202]), .CO(C[203]) );
  FA_4178 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n716), .CI(C[203]), .S(S[203]), .CO(C[204]) );
  FA_4177 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n717), .CI(C[204]), .S(S[204]), .CO(C[205]) );
  FA_4176 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n718), .CI(C[205]), .S(S[205]), .CO(C[206]) );
  FA_4175 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n719), .CI(C[206]), .S(S[206]), .CO(C[207]) );
  FA_4174 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n720), .CI(C[207]), .S(S[207]), .CO(C[208]) );
  FA_4173 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n721), .CI(C[208]), .S(S[208]), .CO(C[209]) );
  FA_4172 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n722), .CI(C[209]), .S(S[209]), .CO(C[210]) );
  FA_4171 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n723), .CI(C[210]), .S(S[210]), .CO(C[211]) );
  FA_4170 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n724), .CI(C[211]), .S(S[211]), .CO(C[212]) );
  FA_4169 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n725), .CI(C[212]), .S(S[212]), .CO(C[213]) );
  FA_4168 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n726), .CI(C[213]), .S(S[213]), .CO(C[214]) );
  FA_4167 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n727), .CI(C[214]), .S(S[214]), .CO(C[215]) );
  FA_4166 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n728), .CI(C[215]), .S(S[215]), .CO(C[216]) );
  FA_4165 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n729), .CI(C[216]), .S(S[216]), .CO(C[217]) );
  FA_4164 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n730), .CI(C[217]), .S(S[217]), .CO(C[218]) );
  FA_4163 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n731), .CI(C[218]), .S(S[218]), .CO(C[219]) );
  FA_4162 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n732), .CI(C[219]), .S(S[219]), .CO(C[220]) );
  FA_4161 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n733), .CI(C[220]), .S(S[220]), .CO(C[221]) );
  FA_4160 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n734), .CI(C[221]), .S(S[221]), .CO(C[222]) );
  FA_4159 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n735), .CI(C[222]), .S(S[222]), .CO(C[223]) );
  FA_4158 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n736), .CI(C[223]), .S(S[223]), .CO(C[224]) );
  FA_4157 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n737), .CI(C[224]), .S(S[224]), .CO(C[225]) );
  FA_4156 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n738), .CI(C[225]), .S(S[225]), .CO(C[226]) );
  FA_4155 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n739), .CI(C[226]), .S(S[226]), .CO(C[227]) );
  FA_4154 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n740), .CI(C[227]), .S(S[227]), .CO(C[228]) );
  FA_4153 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n741), .CI(C[228]), .S(S[228]), .CO(C[229]) );
  FA_4152 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n742), .CI(C[229]), .S(S[229]), .CO(C[230]) );
  FA_4151 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n743), .CI(C[230]), .S(S[230]), .CO(C[231]) );
  FA_4150 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n744), .CI(C[231]), .S(S[231]), .CO(C[232]) );
  FA_4149 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n745), .CI(C[232]), .S(S[232]), .CO(C[233]) );
  FA_4148 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n746), .CI(C[233]), .S(S[233]), .CO(C[234]) );
  FA_4147 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n747), .CI(C[234]), .S(S[234]), .CO(C[235]) );
  FA_4146 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n748), .CI(C[235]), .S(S[235]), .CO(C[236]) );
  FA_4145 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n749), .CI(C[236]), .S(S[236]), .CO(C[237]) );
  FA_4144 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n750), .CI(C[237]), .S(S[237]), .CO(C[238]) );
  FA_4143 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n751), .CI(C[238]), .S(S[238]), .CO(C[239]) );
  FA_4142 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n752), .CI(C[239]), .S(S[239]), .CO(C[240]) );
  FA_4141 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n753), .CI(C[240]), .S(S[240]), .CO(C[241]) );
  FA_4140 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n754), .CI(C[241]), .S(S[241]), .CO(C[242]) );
  FA_4139 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n755), .CI(C[242]), .S(S[242]), .CO(C[243]) );
  FA_4138 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n756), .CI(C[243]), .S(S[243]), .CO(C[244]) );
  FA_4137 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n757), .CI(C[244]), .S(S[244]), .CO(C[245]) );
  FA_4136 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n758), .CI(C[245]), .S(S[245]), .CO(C[246]) );
  FA_4135 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n759), .CI(C[246]), .S(S[246]), .CO(C[247]) );
  FA_4134 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n760), .CI(C[247]), .S(S[247]), .CO(C[248]) );
  FA_4133 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n761), .CI(C[248]), .S(S[248]), .CO(C[249]) );
  FA_4132 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n762), .CI(C[249]), .S(S[249]), .CO(C[250]) );
  FA_4131 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n763), .CI(C[250]), .S(S[250]), .CO(C[251]) );
  FA_4130 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n764), .CI(C[251]), .S(S[251]), .CO(C[252]) );
  FA_4129 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n765), .CI(C[252]), .S(S[252]), .CO(C[253]) );
  FA_4128 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n766), .CI(C[253]), .S(S[253]), .CO(C[254]) );
  FA_4127 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n767), .CI(C[254]), .S(S[254]), .CO(C[255]) );
  FA_4126 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n768), .CI(C[255]), .S(S[255]), .CO(C[256]) );
  FA_4125 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n769), .CI(C[256]), .S(S[256]), .CO(C[257]) );
  FA_4124 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n770), .CI(C[257]), .S(S[257]), .CO(C[258]) );
  FA_4123 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n771), .CI(C[258]), .S(S[258]), .CO(C[259]) );
  FA_4122 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n772), .CI(C[259]), .S(S[259]), .CO(C[260]) );
  FA_4121 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n773), .CI(C[260]), .S(S[260]), .CO(C[261]) );
  FA_4120 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n774), .CI(C[261]), .S(S[261]), .CO(C[262]) );
  FA_4119 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n775), .CI(C[262]), .S(S[262]), .CO(C[263]) );
  FA_4118 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n776), .CI(C[263]), .S(S[263]), .CO(C[264]) );
  FA_4117 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n777), .CI(C[264]), .S(S[264]), .CO(C[265]) );
  FA_4116 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n778), .CI(C[265]), .S(S[265]), .CO(C[266]) );
  FA_4115 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n779), .CI(C[266]), .S(S[266]), .CO(C[267]) );
  FA_4114 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n780), .CI(C[267]), .S(S[267]), .CO(C[268]) );
  FA_4113 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n781), .CI(C[268]), .S(S[268]), .CO(C[269]) );
  FA_4112 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n782), .CI(C[269]), .S(S[269]), .CO(C[270]) );
  FA_4111 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n783), .CI(C[270]), .S(S[270]), .CO(C[271]) );
  FA_4110 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n784), .CI(C[271]), .S(S[271]), .CO(C[272]) );
  FA_4109 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n785), .CI(C[272]), .S(S[272]), .CO(C[273]) );
  FA_4108 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n786), .CI(C[273]), .S(S[273]), .CO(C[274]) );
  FA_4107 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n787), .CI(C[274]), .S(S[274]), .CO(C[275]) );
  FA_4106 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n788), .CI(C[275]), .S(S[275]), .CO(C[276]) );
  FA_4105 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n789), .CI(C[276]), .S(S[276]), .CO(C[277]) );
  FA_4104 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n790), .CI(C[277]), .S(S[277]), .CO(C[278]) );
  FA_4103 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n791), .CI(C[278]), .S(S[278]), .CO(C[279]) );
  FA_4102 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n792), .CI(C[279]), .S(S[279]), .CO(C[280]) );
  FA_4101 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n793), .CI(C[280]), .S(S[280]), .CO(C[281]) );
  FA_4100 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n794), .CI(C[281]), .S(S[281]), .CO(C[282]) );
  FA_4099 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n795), .CI(C[282]), .S(S[282]), .CO(C[283]) );
  FA_4098 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n796), .CI(C[283]), .S(S[283]), .CO(C[284]) );
  FA_4097 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n797), .CI(C[284]), .S(S[284]), .CO(C[285]) );
  FA_4096 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n798), .CI(C[285]), .S(S[285]), .CO(C[286]) );
  FA_4095 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n799), .CI(C[286]), .S(S[286]), .CO(C[287]) );
  FA_4094 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n800), .CI(C[287]), .S(S[287]), .CO(C[288]) );
  FA_4093 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n801), .CI(C[288]), .S(S[288]), .CO(C[289]) );
  FA_4092 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n802), .CI(C[289]), .S(S[289]), .CO(C[290]) );
  FA_4091 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n803), .CI(C[290]), .S(S[290]), .CO(C[291]) );
  FA_4090 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n804), .CI(C[291]), .S(S[291]), .CO(C[292]) );
  FA_4089 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n805), .CI(C[292]), .S(S[292]), .CO(C[293]) );
  FA_4088 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n806), .CI(C[293]), .S(S[293]), .CO(C[294]) );
  FA_4087 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n807), .CI(C[294]), .S(S[294]), .CO(C[295]) );
  FA_4086 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n808), .CI(C[295]), .S(S[295]), .CO(C[296]) );
  FA_4085 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n809), .CI(C[296]), .S(S[296]), .CO(C[297]) );
  FA_4084 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n810), .CI(C[297]), .S(S[297]), .CO(C[298]) );
  FA_4083 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n811), .CI(C[298]), .S(S[298]), .CO(C[299]) );
  FA_4082 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n812), .CI(C[299]), .S(S[299]), .CO(C[300]) );
  FA_4081 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n813), .CI(C[300]), .S(S[300]), .CO(C[301]) );
  FA_4080 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n814), .CI(C[301]), .S(S[301]), .CO(C[302]) );
  FA_4079 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n815), .CI(C[302]), .S(S[302]), .CO(C[303]) );
  FA_4078 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n816), .CI(C[303]), .S(S[303]), .CO(C[304]) );
  FA_4077 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n817), .CI(C[304]), .S(S[304]), .CO(C[305]) );
  FA_4076 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n818), .CI(C[305]), .S(S[305]), .CO(C[306]) );
  FA_4075 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n819), .CI(C[306]), .S(S[306]), .CO(C[307]) );
  FA_4074 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n820), .CI(C[307]), .S(S[307]), .CO(C[308]) );
  FA_4073 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n821), .CI(C[308]), .S(S[308]), .CO(C[309]) );
  FA_4072 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n822), .CI(C[309]), .S(S[309]), .CO(C[310]) );
  FA_4071 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n823), .CI(C[310]), .S(S[310]), .CO(C[311]) );
  FA_4070 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n824), .CI(C[311]), .S(S[311]), .CO(C[312]) );
  FA_4069 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n825), .CI(C[312]), .S(S[312]), .CO(C[313]) );
  FA_4068 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n826), .CI(C[313]), .S(S[313]), .CO(C[314]) );
  FA_4067 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n827), .CI(C[314]), .S(S[314]), .CO(C[315]) );
  FA_4066 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n828), .CI(C[315]), .S(S[315]), .CO(C[316]) );
  FA_4065 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n829), .CI(C[316]), .S(S[316]), .CO(C[317]) );
  FA_4064 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n830), .CI(C[317]), .S(S[317]), .CO(C[318]) );
  FA_4063 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n831), .CI(C[318]), .S(S[318]), .CO(C[319]) );
  FA_4062 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n832), .CI(C[319]), .S(S[319]), .CO(C[320]) );
  FA_4061 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n833), .CI(C[320]), .S(S[320]), .CO(C[321]) );
  FA_4060 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n834), .CI(C[321]), .S(S[321]), .CO(C[322]) );
  FA_4059 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n835), .CI(C[322]), .S(S[322]), .CO(C[323]) );
  FA_4058 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n836), .CI(C[323]), .S(S[323]), .CO(C[324]) );
  FA_4057 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n837), .CI(C[324]), .S(S[324]), .CO(C[325]) );
  FA_4056 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n838), .CI(C[325]), .S(S[325]), .CO(C[326]) );
  FA_4055 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n839), .CI(C[326]), .S(S[326]), .CO(C[327]) );
  FA_4054 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n840), .CI(C[327]), .S(S[327]), .CO(C[328]) );
  FA_4053 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n841), .CI(C[328]), .S(S[328]), .CO(C[329]) );
  FA_4052 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n842), .CI(C[329]), .S(S[329]), .CO(C[330]) );
  FA_4051 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n843), .CI(C[330]), .S(S[330]), .CO(C[331]) );
  FA_4050 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n844), .CI(C[331]), .S(S[331]), .CO(C[332]) );
  FA_4049 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n845), .CI(C[332]), .S(S[332]), .CO(C[333]) );
  FA_4048 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n846), .CI(C[333]), .S(S[333]), .CO(C[334]) );
  FA_4047 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n847), .CI(C[334]), .S(S[334]), .CO(C[335]) );
  FA_4046 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n848), .CI(C[335]), .S(S[335]), .CO(C[336]) );
  FA_4045 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n849), .CI(C[336]), .S(S[336]), .CO(C[337]) );
  FA_4044 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n850), .CI(C[337]), .S(S[337]), .CO(C[338]) );
  FA_4043 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n851), .CI(C[338]), .S(S[338]), .CO(C[339]) );
  FA_4042 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n852), .CI(C[339]), .S(S[339]), .CO(C[340]) );
  FA_4041 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n853), .CI(C[340]), .S(S[340]), .CO(C[341]) );
  FA_4040 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n854), .CI(C[341]), .S(S[341]), .CO(C[342]) );
  FA_4039 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n855), .CI(C[342]), .S(S[342]), .CO(C[343]) );
  FA_4038 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n856), .CI(C[343]), .S(S[343]), .CO(C[344]) );
  FA_4037 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n857), .CI(C[344]), .S(S[344]), .CO(C[345]) );
  FA_4036 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n858), .CI(C[345]), .S(S[345]), .CO(C[346]) );
  FA_4035 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n859), .CI(C[346]), .S(S[346]), .CO(C[347]) );
  FA_4034 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n860), .CI(C[347]), .S(S[347]), .CO(C[348]) );
  FA_4033 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n861), .CI(C[348]), .S(S[348]), .CO(C[349]) );
  FA_4032 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n862), .CI(C[349]), .S(S[349]), .CO(C[350]) );
  FA_4031 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n863), .CI(C[350]), .S(S[350]), .CO(C[351]) );
  FA_4030 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n864), .CI(C[351]), .S(S[351]), .CO(C[352]) );
  FA_4029 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n865), .CI(C[352]), .S(S[352]), .CO(C[353]) );
  FA_4028 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n866), .CI(C[353]), .S(S[353]), .CO(C[354]) );
  FA_4027 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n867), .CI(C[354]), .S(S[354]), .CO(C[355]) );
  FA_4026 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n868), .CI(C[355]), .S(S[355]), .CO(C[356]) );
  FA_4025 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n869), .CI(C[356]), .S(S[356]), .CO(C[357]) );
  FA_4024 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n870), .CI(C[357]), .S(S[357]), .CO(C[358]) );
  FA_4023 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n871), .CI(C[358]), .S(S[358]), .CO(C[359]) );
  FA_4022 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n872), .CI(C[359]), .S(S[359]), .CO(C[360]) );
  FA_4021 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n873), .CI(C[360]), .S(S[360]), .CO(C[361]) );
  FA_4020 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n874), .CI(C[361]), .S(S[361]), .CO(C[362]) );
  FA_4019 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n875), .CI(C[362]), .S(S[362]), .CO(C[363]) );
  FA_4018 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n876), .CI(C[363]), .S(S[363]), .CO(C[364]) );
  FA_4017 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n877), .CI(C[364]), .S(S[364]), .CO(C[365]) );
  FA_4016 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n878), .CI(C[365]), .S(S[365]), .CO(C[366]) );
  FA_4015 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n879), .CI(C[366]), .S(S[366]), .CO(C[367]) );
  FA_4014 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n880), .CI(C[367]), .S(S[367]), .CO(C[368]) );
  FA_4013 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n881), .CI(C[368]), .S(S[368]), .CO(C[369]) );
  FA_4012 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n882), .CI(C[369]), .S(S[369]), .CO(C[370]) );
  FA_4011 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n883), .CI(C[370]), .S(S[370]), .CO(C[371]) );
  FA_4010 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n884), .CI(C[371]), .S(S[371]), .CO(C[372]) );
  FA_4009 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n885), .CI(C[372]), .S(S[372]), .CO(C[373]) );
  FA_4008 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n886), .CI(C[373]), .S(S[373]), .CO(C[374]) );
  FA_4007 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n887), .CI(C[374]), .S(S[374]), .CO(C[375]) );
  FA_4006 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n888), .CI(C[375]), .S(S[375]), .CO(C[376]) );
  FA_4005 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n889), .CI(C[376]), .S(S[376]), .CO(C[377]) );
  FA_4004 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n890), .CI(C[377]), .S(S[377]), .CO(C[378]) );
  FA_4003 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n891), .CI(C[378]), .S(S[378]), .CO(C[379]) );
  FA_4002 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n892), .CI(C[379]), .S(S[379]), .CO(C[380]) );
  FA_4001 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n893), .CI(C[380]), .S(S[380]), .CO(C[381]) );
  FA_4000 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n894), .CI(C[381]), .S(S[381]), .CO(C[382]) );
  FA_3999 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n895), .CI(C[382]), .S(S[382]), .CO(C[383]) );
  FA_3998 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n896), .CI(C[383]), .S(S[383]), .CO(C[384]) );
  FA_3997 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n897), .CI(C[384]), .S(S[384]), .CO(C[385]) );
  FA_3996 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n898), .CI(C[385]), .S(S[385]), .CO(C[386]) );
  FA_3995 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n899), .CI(C[386]), .S(S[386]), .CO(C[387]) );
  FA_3994 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n900), .CI(C[387]), .S(S[387]), .CO(C[388]) );
  FA_3993 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n901), .CI(C[388]), .S(S[388]), .CO(C[389]) );
  FA_3992 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n902), .CI(C[389]), .S(S[389]), .CO(C[390]) );
  FA_3991 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n903), .CI(C[390]), .S(S[390]), .CO(C[391]) );
  FA_3990 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n904), .CI(C[391]), .S(S[391]), .CO(C[392]) );
  FA_3989 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n905), .CI(C[392]), .S(S[392]), .CO(C[393]) );
  FA_3988 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n906), .CI(C[393]), .S(S[393]), .CO(C[394]) );
  FA_3987 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n907), .CI(C[394]), .S(S[394]), .CO(C[395]) );
  FA_3986 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n908), .CI(C[395]), .S(S[395]), .CO(C[396]) );
  FA_3985 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n909), .CI(C[396]), .S(S[396]), .CO(C[397]) );
  FA_3984 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n910), .CI(C[397]), .S(S[397]), .CO(C[398]) );
  FA_3983 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n911), .CI(C[398]), .S(S[398]), .CO(C[399]) );
  FA_3982 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n912), .CI(C[399]), .S(S[399]), .CO(C[400]) );
  FA_3981 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n913), .CI(C[400]), .S(S[400]), .CO(C[401]) );
  FA_3980 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n914), .CI(C[401]), .S(S[401]), .CO(C[402]) );
  FA_3979 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n915), .CI(C[402]), .S(S[402]), .CO(C[403]) );
  FA_3978 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n916), .CI(C[403]), .S(S[403]), .CO(C[404]) );
  FA_3977 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n917), .CI(C[404]), .S(S[404]), .CO(C[405]) );
  FA_3976 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n918), .CI(C[405]), .S(S[405]), .CO(C[406]) );
  FA_3975 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n919), .CI(C[406]), .S(S[406]), .CO(C[407]) );
  FA_3974 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n920), .CI(C[407]), .S(S[407]), .CO(C[408]) );
  FA_3973 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n921), .CI(C[408]), .S(S[408]), .CO(C[409]) );
  FA_3972 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n922), .CI(C[409]), .S(S[409]), .CO(C[410]) );
  FA_3971 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n923), .CI(C[410]), .S(S[410]), .CO(C[411]) );
  FA_3970 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n924), .CI(C[411]), .S(S[411]), .CO(C[412]) );
  FA_3969 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n925), .CI(C[412]), .S(S[412]), .CO(C[413]) );
  FA_3968 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n926), .CI(C[413]), .S(S[413]), .CO(C[414]) );
  FA_3967 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n927), .CI(C[414]), .S(S[414]), .CO(C[415]) );
  FA_3966 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n928), .CI(C[415]), .S(S[415]), .CO(C[416]) );
  FA_3965 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n929), .CI(C[416]), .S(S[416]), .CO(C[417]) );
  FA_3964 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n930), .CI(C[417]), .S(S[417]), .CO(C[418]) );
  FA_3963 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n931), .CI(C[418]), .S(S[418]), .CO(C[419]) );
  FA_3962 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n932), .CI(C[419]), .S(S[419]), .CO(C[420]) );
  FA_3961 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n933), .CI(C[420]), .S(S[420]), .CO(C[421]) );
  FA_3960 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n934), .CI(C[421]), .S(S[421]), .CO(C[422]) );
  FA_3959 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n935), .CI(C[422]), .S(S[422]), .CO(C[423]) );
  FA_3958 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n936), .CI(C[423]), .S(S[423]), .CO(C[424]) );
  FA_3957 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n937), .CI(C[424]), .S(S[424]), .CO(C[425]) );
  FA_3956 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n938), .CI(C[425]), .S(S[425]), .CO(C[426]) );
  FA_3955 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n939), .CI(C[426]), .S(S[426]), .CO(C[427]) );
  FA_3954 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n940), .CI(C[427]), .S(S[427]), .CO(C[428]) );
  FA_3953 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n941), .CI(C[428]), .S(S[428]), .CO(C[429]) );
  FA_3952 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n942), .CI(C[429]), .S(S[429]), .CO(C[430]) );
  FA_3951 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n943), .CI(C[430]), .S(S[430]), .CO(C[431]) );
  FA_3950 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n944), .CI(C[431]), .S(S[431]), .CO(C[432]) );
  FA_3949 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n945), .CI(C[432]), .S(S[432]), .CO(C[433]) );
  FA_3948 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n946), .CI(C[433]), .S(S[433]), .CO(C[434]) );
  FA_3947 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n947), .CI(C[434]), .S(S[434]), .CO(C[435]) );
  FA_3946 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n948), .CI(C[435]), .S(S[435]), .CO(C[436]) );
  FA_3945 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n949), .CI(C[436]), .S(S[436]), .CO(C[437]) );
  FA_3944 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n950), .CI(C[437]), .S(S[437]), .CO(C[438]) );
  FA_3943 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n951), .CI(C[438]), .S(S[438]), .CO(C[439]) );
  FA_3942 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n952), .CI(C[439]), .S(S[439]), .CO(C[440]) );
  FA_3941 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n953), .CI(C[440]), .S(S[440]), .CO(C[441]) );
  FA_3940 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n954), .CI(C[441]), .S(S[441]), .CO(C[442]) );
  FA_3939 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n955), .CI(C[442]), .S(S[442]), .CO(C[443]) );
  FA_3938 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n956), .CI(C[443]), .S(S[443]), .CO(C[444]) );
  FA_3937 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n957), .CI(C[444]), .S(S[444]), .CO(C[445]) );
  FA_3936 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n958), .CI(C[445]), .S(S[445]), .CO(C[446]) );
  FA_3935 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n959), .CI(C[446]), .S(S[446]), .CO(C[447]) );
  FA_3934 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n960), .CI(C[447]), .S(S[447]), .CO(C[448]) );
  FA_3933 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n961), .CI(C[448]), .S(S[448]), .CO(C[449]) );
  FA_3932 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n962), .CI(C[449]), .S(S[449]), .CO(C[450]) );
  FA_3931 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n963), .CI(C[450]), .S(S[450]), .CO(C[451]) );
  FA_3930 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n964), .CI(C[451]), .S(S[451]), .CO(C[452]) );
  FA_3929 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n965), .CI(C[452]), .S(S[452]), .CO(C[453]) );
  FA_3928 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n966), .CI(C[453]), .S(S[453]), .CO(C[454]) );
  FA_3927 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n967), .CI(C[454]), .S(S[454]), .CO(C[455]) );
  FA_3926 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n968), .CI(C[455]), .S(S[455]), .CO(C[456]) );
  FA_3925 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n969), .CI(C[456]), .S(S[456]), .CO(C[457]) );
  FA_3924 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n970), .CI(C[457]), .S(S[457]), .CO(C[458]) );
  FA_3923 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n971), .CI(C[458]), .S(S[458]), .CO(C[459]) );
  FA_3922 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n972), .CI(C[459]), .S(S[459]), .CO(C[460]) );
  FA_3921 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n973), .CI(C[460]), .S(S[460]), .CO(C[461]) );
  FA_3920 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n974), .CI(C[461]), .S(S[461]), .CO(C[462]) );
  FA_3919 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n975), .CI(C[462]), .S(S[462]), .CO(C[463]) );
  FA_3918 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n976), .CI(C[463]), .S(S[463]), .CO(C[464]) );
  FA_3917 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n977), .CI(C[464]), .S(S[464]), .CO(C[465]) );
  FA_3916 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n978), .CI(C[465]), .S(S[465]), .CO(C[466]) );
  FA_3915 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n979), .CI(C[466]), .S(S[466]), .CO(C[467]) );
  FA_3914 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n980), .CI(C[467]), .S(S[467]), .CO(C[468]) );
  FA_3913 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n981), .CI(C[468]), .S(S[468]), .CO(C[469]) );
  FA_3912 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n982), .CI(C[469]), .S(S[469]), .CO(C[470]) );
  FA_3911 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n983), .CI(C[470]), .S(S[470]), .CO(C[471]) );
  FA_3910 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n984), .CI(C[471]), .S(S[471]), .CO(C[472]) );
  FA_3909 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n985), .CI(C[472]), .S(S[472]), .CO(C[473]) );
  FA_3908 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n986), .CI(C[473]), .S(S[473]), .CO(C[474]) );
  FA_3907 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n987), .CI(C[474]), .S(S[474]), .CO(C[475]) );
  FA_3906 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n988), .CI(C[475]), .S(S[475]), .CO(C[476]) );
  FA_3905 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n989), .CI(C[476]), .S(S[476]), .CO(C[477]) );
  FA_3904 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n990), .CI(C[477]), .S(S[477]), .CO(C[478]) );
  FA_3903 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n991), .CI(C[478]), .S(S[478]), .CO(C[479]) );
  FA_3902 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n992), .CI(C[479]), .S(S[479]), .CO(C[480]) );
  FA_3901 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n993), .CI(C[480]), .S(S[480]), .CO(C[481]) );
  FA_3900 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n994), .CI(C[481]), .S(S[481]), .CO(C[482]) );
  FA_3899 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n995), .CI(C[482]), .S(S[482]), .CO(C[483]) );
  FA_3898 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n996), .CI(C[483]), .S(S[483]), .CO(C[484]) );
  FA_3897 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n997), .CI(C[484]), .S(S[484]), .CO(C[485]) );
  FA_3896 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n998), .CI(C[485]), .S(S[485]), .CO(C[486]) );
  FA_3895 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n999), .CI(C[486]), .S(S[486]), .CO(C[487]) );
  FA_3894 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n1000), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_3893 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n1001), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_3892 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n1002), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_3891 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n1003), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_3890 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n1004), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_3889 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n1005), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_3888 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n1006), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_3887 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n1007), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_3886 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n1008), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_3885 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n1009), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_3884 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n1010), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_3883 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n1011), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_3882 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n1012), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_3881 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n1013), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_3880 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n1014), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_3879 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n1015), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_3878 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n1016), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_3877 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n1017), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_3876 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n1018), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_3875 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n1019), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_3874 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n1020), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_3873 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n1021), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_3872 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n1022), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_3871 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n1023), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_3870 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n1024), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_3869 \FA_INST_1[512].FA_  ( .A(A[512]), .B(1'b1), .CI(C[512]), .S(S[512])
         );
  IV U2 ( .A(B[415]), .Z(n928) );
  IV U3 ( .A(B[416]), .Z(n929) );
  IV U4 ( .A(B[417]), .Z(n930) );
  IV U5 ( .A(B[418]), .Z(n931) );
  IV U6 ( .A(B[419]), .Z(n932) );
  IV U7 ( .A(B[420]), .Z(n933) );
  IV U8 ( .A(B[421]), .Z(n934) );
  IV U9 ( .A(B[422]), .Z(n935) );
  IV U10 ( .A(B[423]), .Z(n936) );
  IV U11 ( .A(B[424]), .Z(n937) );
  IV U12 ( .A(B[505]), .Z(n1018) );
  IV U13 ( .A(B[425]), .Z(n938) );
  IV U14 ( .A(B[426]), .Z(n939) );
  IV U15 ( .A(B[427]), .Z(n940) );
  IV U16 ( .A(B[428]), .Z(n941) );
  IV U17 ( .A(B[429]), .Z(n942) );
  IV U18 ( .A(B[430]), .Z(n943) );
  IV U19 ( .A(B[431]), .Z(n944) );
  IV U20 ( .A(B[432]), .Z(n945) );
  IV U21 ( .A(B[433]), .Z(n946) );
  IV U22 ( .A(B[434]), .Z(n947) );
  IV U23 ( .A(B[506]), .Z(n1019) );
  IV U24 ( .A(B[435]), .Z(n948) );
  IV U25 ( .A(B[436]), .Z(n949) );
  IV U26 ( .A(B[437]), .Z(n950) );
  IV U27 ( .A(B[438]), .Z(n951) );
  IV U28 ( .A(B[439]), .Z(n952) );
  IV U29 ( .A(B[440]), .Z(n953) );
  IV U30 ( .A(B[441]), .Z(n954) );
  IV U31 ( .A(B[442]), .Z(n955) );
  IV U32 ( .A(B[443]), .Z(n956) );
  IV U33 ( .A(B[444]), .Z(n957) );
  IV U34 ( .A(B[507]), .Z(n1020) );
  IV U35 ( .A(B[445]), .Z(n958) );
  IV U36 ( .A(B[446]), .Z(n959) );
  IV U37 ( .A(B[447]), .Z(n960) );
  IV U38 ( .A(B[448]), .Z(n961) );
  IV U39 ( .A(B[449]), .Z(n962) );
  IV U40 ( .A(B[450]), .Z(n963) );
  IV U41 ( .A(B[451]), .Z(n964) );
  IV U42 ( .A(B[452]), .Z(n965) );
  IV U43 ( .A(B[453]), .Z(n966) );
  IV U44 ( .A(B[454]), .Z(n967) );
  IV U45 ( .A(B[508]), .Z(n1021) );
  IV U46 ( .A(B[455]), .Z(n968) );
  IV U47 ( .A(B[456]), .Z(n969) );
  IV U48 ( .A(B[457]), .Z(n970) );
  IV U49 ( .A(B[458]), .Z(n971) );
  IV U50 ( .A(B[459]), .Z(n972) );
  IV U51 ( .A(B[460]), .Z(n973) );
  IV U52 ( .A(B[461]), .Z(n974) );
  IV U53 ( .A(B[462]), .Z(n975) );
  IV U54 ( .A(B[0]), .Z(n2) );
  IV U55 ( .A(B[1]), .Z(n514) );
  IV U56 ( .A(B[2]), .Z(n515) );
  IV U57 ( .A(B[3]), .Z(n516) );
  IV U58 ( .A(B[4]), .Z(n517) );
  IV U59 ( .A(B[463]), .Z(n976) );
  IV U60 ( .A(B[5]), .Z(n518) );
  IV U61 ( .A(B[6]), .Z(n519) );
  IV U62 ( .A(B[7]), .Z(n520) );
  IV U63 ( .A(B[8]), .Z(n521) );
  IV U64 ( .A(B[9]), .Z(n522) );
  IV U65 ( .A(B[10]), .Z(n523) );
  IV U66 ( .A(B[11]), .Z(n524) );
  IV U67 ( .A(B[12]), .Z(n525) );
  IV U68 ( .A(B[13]), .Z(n526) );
  IV U69 ( .A(B[14]), .Z(n527) );
  IV U70 ( .A(B[464]), .Z(n977) );
  IV U71 ( .A(B[509]), .Z(n1022) );
  IV U72 ( .A(B[15]), .Z(n528) );
  IV U73 ( .A(B[16]), .Z(n529) );
  IV U74 ( .A(B[17]), .Z(n530) );
  IV U75 ( .A(B[18]), .Z(n531) );
  IV U76 ( .A(B[19]), .Z(n532) );
  IV U77 ( .A(B[20]), .Z(n533) );
  IV U78 ( .A(B[21]), .Z(n534) );
  IV U79 ( .A(B[22]), .Z(n535) );
  IV U80 ( .A(B[23]), .Z(n536) );
  IV U81 ( .A(B[24]), .Z(n537) );
  IV U82 ( .A(B[465]), .Z(n978) );
  IV U83 ( .A(B[25]), .Z(n538) );
  IV U84 ( .A(B[26]), .Z(n539) );
  IV U85 ( .A(B[27]), .Z(n540) );
  IV U86 ( .A(B[28]), .Z(n541) );
  IV U87 ( .A(B[29]), .Z(n542) );
  IV U88 ( .A(B[30]), .Z(n543) );
  IV U89 ( .A(B[31]), .Z(n544) );
  IV U90 ( .A(B[32]), .Z(n545) );
  IV U91 ( .A(B[33]), .Z(n546) );
  IV U92 ( .A(B[34]), .Z(n547) );
  IV U93 ( .A(B[466]), .Z(n979) );
  IV U94 ( .A(B[35]), .Z(n548) );
  IV U95 ( .A(B[36]), .Z(n549) );
  IV U96 ( .A(B[37]), .Z(n550) );
  IV U97 ( .A(B[38]), .Z(n551) );
  IV U98 ( .A(B[39]), .Z(n552) );
  IV U99 ( .A(B[40]), .Z(n553) );
  IV U100 ( .A(B[41]), .Z(n554) );
  IV U101 ( .A(B[42]), .Z(n555) );
  IV U102 ( .A(B[43]), .Z(n556) );
  IV U103 ( .A(B[44]), .Z(n557) );
  IV U104 ( .A(B[467]), .Z(n980) );
  IV U105 ( .A(B[45]), .Z(n558) );
  IV U106 ( .A(B[46]), .Z(n559) );
  IV U107 ( .A(B[47]), .Z(n560) );
  IV U108 ( .A(B[48]), .Z(n561) );
  IV U109 ( .A(B[49]), .Z(n562) );
  IV U110 ( .A(B[50]), .Z(n563) );
  IV U111 ( .A(B[51]), .Z(n564) );
  IV U112 ( .A(B[52]), .Z(n565) );
  IV U113 ( .A(B[53]), .Z(n566) );
  IV U114 ( .A(B[54]), .Z(n567) );
  IV U115 ( .A(B[468]), .Z(n981) );
  IV U116 ( .A(B[55]), .Z(n568) );
  IV U117 ( .A(B[56]), .Z(n569) );
  IV U118 ( .A(B[57]), .Z(n570) );
  IV U119 ( .A(B[58]), .Z(n571) );
  IV U120 ( .A(B[59]), .Z(n572) );
  IV U121 ( .A(B[60]), .Z(n573) );
  IV U122 ( .A(B[61]), .Z(n574) );
  IV U123 ( .A(B[62]), .Z(n575) );
  IV U124 ( .A(B[63]), .Z(n576) );
  IV U125 ( .A(B[64]), .Z(n577) );
  IV U126 ( .A(B[469]), .Z(n982) );
  IV U127 ( .A(B[65]), .Z(n578) );
  IV U128 ( .A(B[66]), .Z(n579) );
  IV U129 ( .A(B[67]), .Z(n580) );
  IV U130 ( .A(B[68]), .Z(n581) );
  IV U131 ( .A(B[69]), .Z(n582) );
  IV U132 ( .A(B[70]), .Z(n583) );
  IV U133 ( .A(B[71]), .Z(n584) );
  IV U134 ( .A(B[72]), .Z(n585) );
  IV U135 ( .A(B[73]), .Z(n586) );
  IV U136 ( .A(B[74]), .Z(n587) );
  IV U137 ( .A(B[470]), .Z(n983) );
  IV U138 ( .A(B[75]), .Z(n588) );
  IV U139 ( .A(B[76]), .Z(n589) );
  IV U140 ( .A(B[77]), .Z(n590) );
  IV U141 ( .A(B[78]), .Z(n591) );
  IV U142 ( .A(B[79]), .Z(n592) );
  IV U143 ( .A(B[80]), .Z(n593) );
  IV U144 ( .A(B[81]), .Z(n594) );
  IV U145 ( .A(B[82]), .Z(n595) );
  IV U146 ( .A(B[83]), .Z(n596) );
  IV U147 ( .A(B[84]), .Z(n597) );
  IV U148 ( .A(B[471]), .Z(n984) );
  IV U149 ( .A(B[85]), .Z(n598) );
  IV U150 ( .A(B[86]), .Z(n599) );
  IV U151 ( .A(B[87]), .Z(n600) );
  IV U152 ( .A(B[88]), .Z(n601) );
  IV U153 ( .A(B[89]), .Z(n602) );
  IV U154 ( .A(B[90]), .Z(n603) );
  IV U155 ( .A(B[91]), .Z(n604) );
  IV U156 ( .A(B[92]), .Z(n605) );
  IV U157 ( .A(B[93]), .Z(n606) );
  IV U158 ( .A(B[94]), .Z(n607) );
  IV U159 ( .A(B[472]), .Z(n985) );
  IV U160 ( .A(B[95]), .Z(n608) );
  IV U161 ( .A(B[96]), .Z(n609) );
  IV U162 ( .A(B[97]), .Z(n610) );
  IV U163 ( .A(B[98]), .Z(n611) );
  IV U164 ( .A(B[99]), .Z(n612) );
  IV U165 ( .A(B[100]), .Z(n613) );
  IV U166 ( .A(B[101]), .Z(n614) );
  IV U167 ( .A(B[102]), .Z(n615) );
  IV U168 ( .A(B[103]), .Z(n616) );
  IV U169 ( .A(B[104]), .Z(n617) );
  IV U170 ( .A(B[473]), .Z(n986) );
  IV U171 ( .A(B[105]), .Z(n618) );
  IV U172 ( .A(B[106]), .Z(n619) );
  IV U173 ( .A(B[107]), .Z(n620) );
  IV U174 ( .A(B[108]), .Z(n621) );
  IV U175 ( .A(B[109]), .Z(n622) );
  IV U176 ( .A(B[110]), .Z(n623) );
  IV U177 ( .A(B[111]), .Z(n624) );
  IV U178 ( .A(B[112]), .Z(n625) );
  IV U179 ( .A(B[113]), .Z(n626) );
  IV U180 ( .A(B[114]), .Z(n627) );
  IV U181 ( .A(B[474]), .Z(n987) );
  IV U182 ( .A(B[510]), .Z(n1023) );
  IV U183 ( .A(B[115]), .Z(n628) );
  IV U184 ( .A(B[116]), .Z(n629) );
  IV U185 ( .A(B[117]), .Z(n630) );
  IV U186 ( .A(B[118]), .Z(n631) );
  IV U187 ( .A(B[119]), .Z(n632) );
  IV U188 ( .A(B[120]), .Z(n633) );
  IV U189 ( .A(B[121]), .Z(n634) );
  IV U190 ( .A(B[122]), .Z(n635) );
  IV U191 ( .A(B[123]), .Z(n636) );
  IV U192 ( .A(B[124]), .Z(n637) );
  IV U193 ( .A(B[475]), .Z(n988) );
  IV U194 ( .A(B[125]), .Z(n638) );
  IV U195 ( .A(B[126]), .Z(n639) );
  IV U196 ( .A(B[127]), .Z(n640) );
  IV U197 ( .A(B[128]), .Z(n641) );
  IV U198 ( .A(B[129]), .Z(n642) );
  IV U199 ( .A(B[130]), .Z(n643) );
  IV U200 ( .A(B[131]), .Z(n644) );
  IV U201 ( .A(B[132]), .Z(n645) );
  IV U202 ( .A(B[133]), .Z(n646) );
  IV U203 ( .A(B[134]), .Z(n647) );
  IV U204 ( .A(B[476]), .Z(n989) );
  IV U205 ( .A(B[135]), .Z(n648) );
  IV U206 ( .A(B[136]), .Z(n649) );
  IV U207 ( .A(B[137]), .Z(n650) );
  IV U208 ( .A(B[138]), .Z(n651) );
  IV U209 ( .A(B[139]), .Z(n652) );
  IV U210 ( .A(B[140]), .Z(n653) );
  IV U211 ( .A(B[141]), .Z(n654) );
  IV U212 ( .A(B[142]), .Z(n655) );
  IV U213 ( .A(B[143]), .Z(n656) );
  IV U214 ( .A(B[144]), .Z(n657) );
  IV U215 ( .A(B[477]), .Z(n990) );
  IV U216 ( .A(B[145]), .Z(n658) );
  IV U217 ( .A(B[146]), .Z(n659) );
  IV U218 ( .A(B[147]), .Z(n660) );
  IV U219 ( .A(B[148]), .Z(n661) );
  IV U220 ( .A(B[149]), .Z(n662) );
  IV U221 ( .A(B[150]), .Z(n663) );
  IV U222 ( .A(B[151]), .Z(n664) );
  IV U223 ( .A(B[152]), .Z(n665) );
  IV U224 ( .A(B[153]), .Z(n666) );
  IV U225 ( .A(B[154]), .Z(n667) );
  IV U226 ( .A(B[478]), .Z(n991) );
  IV U227 ( .A(B[155]), .Z(n668) );
  IV U228 ( .A(B[156]), .Z(n669) );
  IV U229 ( .A(B[157]), .Z(n670) );
  IV U230 ( .A(B[158]), .Z(n671) );
  IV U231 ( .A(B[159]), .Z(n672) );
  IV U232 ( .A(B[160]), .Z(n673) );
  IV U233 ( .A(B[161]), .Z(n674) );
  IV U234 ( .A(B[162]), .Z(n675) );
  IV U235 ( .A(B[163]), .Z(n676) );
  IV U236 ( .A(B[164]), .Z(n677) );
  IV U237 ( .A(B[479]), .Z(n992) );
  IV U238 ( .A(B[165]), .Z(n678) );
  IV U239 ( .A(B[166]), .Z(n679) );
  IV U240 ( .A(B[167]), .Z(n680) );
  IV U241 ( .A(B[168]), .Z(n681) );
  IV U242 ( .A(B[169]), .Z(n682) );
  IV U243 ( .A(B[170]), .Z(n683) );
  IV U244 ( .A(B[171]), .Z(n684) );
  IV U245 ( .A(B[172]), .Z(n685) );
  IV U246 ( .A(B[173]), .Z(n686) );
  IV U247 ( .A(B[174]), .Z(n687) );
  IV U248 ( .A(B[480]), .Z(n993) );
  IV U249 ( .A(B[175]), .Z(n688) );
  IV U250 ( .A(B[176]), .Z(n689) );
  IV U251 ( .A(B[177]), .Z(n690) );
  IV U252 ( .A(B[178]), .Z(n691) );
  IV U253 ( .A(B[179]), .Z(n692) );
  IV U254 ( .A(B[180]), .Z(n693) );
  IV U255 ( .A(B[181]), .Z(n694) );
  IV U256 ( .A(B[182]), .Z(n695) );
  IV U257 ( .A(B[183]), .Z(n696) );
  IV U258 ( .A(B[184]), .Z(n697) );
  IV U259 ( .A(B[481]), .Z(n994) );
  IV U260 ( .A(B[185]), .Z(n698) );
  IV U261 ( .A(B[186]), .Z(n699) );
  IV U262 ( .A(B[187]), .Z(n700) );
  IV U263 ( .A(B[188]), .Z(n701) );
  IV U264 ( .A(B[189]), .Z(n702) );
  IV U265 ( .A(B[190]), .Z(n703) );
  IV U266 ( .A(B[191]), .Z(n704) );
  IV U267 ( .A(B[192]), .Z(n705) );
  IV U268 ( .A(B[193]), .Z(n706) );
  IV U269 ( .A(B[194]), .Z(n707) );
  IV U270 ( .A(B[482]), .Z(n995) );
  IV U271 ( .A(B[195]), .Z(n708) );
  IV U272 ( .A(B[196]), .Z(n709) );
  IV U273 ( .A(B[197]), .Z(n710) );
  IV U274 ( .A(B[198]), .Z(n711) );
  IV U275 ( .A(B[199]), .Z(n712) );
  IV U276 ( .A(B[200]), .Z(n713) );
  IV U277 ( .A(B[201]), .Z(n714) );
  IV U278 ( .A(B[202]), .Z(n715) );
  IV U279 ( .A(B[203]), .Z(n716) );
  IV U280 ( .A(B[204]), .Z(n717) );
  IV U281 ( .A(B[483]), .Z(n996) );
  IV U282 ( .A(B[205]), .Z(n718) );
  IV U283 ( .A(B[206]), .Z(n719) );
  IV U284 ( .A(B[207]), .Z(n720) );
  IV U285 ( .A(B[208]), .Z(n721) );
  IV U286 ( .A(B[209]), .Z(n722) );
  IV U287 ( .A(B[210]), .Z(n723) );
  IV U288 ( .A(B[211]), .Z(n724) );
  IV U289 ( .A(B[212]), .Z(n725) );
  IV U290 ( .A(B[213]), .Z(n726) );
  IV U291 ( .A(B[214]), .Z(n727) );
  IV U292 ( .A(B[484]), .Z(n997) );
  IV U293 ( .A(B[511]), .Z(n1024) );
  IV U294 ( .A(B[215]), .Z(n728) );
  IV U295 ( .A(B[216]), .Z(n729) );
  IV U296 ( .A(B[217]), .Z(n730) );
  IV U297 ( .A(B[218]), .Z(n731) );
  IV U298 ( .A(B[219]), .Z(n732) );
  IV U299 ( .A(B[220]), .Z(n733) );
  IV U300 ( .A(B[221]), .Z(n734) );
  IV U301 ( .A(B[222]), .Z(n735) );
  IV U302 ( .A(B[223]), .Z(n736) );
  IV U303 ( .A(B[224]), .Z(n737) );
  IV U304 ( .A(B[485]), .Z(n998) );
  IV U305 ( .A(B[225]), .Z(n738) );
  IV U306 ( .A(B[226]), .Z(n739) );
  IV U307 ( .A(B[227]), .Z(n740) );
  IV U308 ( .A(B[228]), .Z(n741) );
  IV U309 ( .A(B[229]), .Z(n742) );
  IV U310 ( .A(B[230]), .Z(n743) );
  IV U311 ( .A(B[231]), .Z(n744) );
  IV U312 ( .A(B[232]), .Z(n745) );
  IV U313 ( .A(B[233]), .Z(n746) );
  IV U314 ( .A(B[234]), .Z(n747) );
  IV U315 ( .A(B[486]), .Z(n999) );
  IV U316 ( .A(B[235]), .Z(n748) );
  IV U317 ( .A(B[236]), .Z(n749) );
  IV U318 ( .A(B[237]), .Z(n750) );
  IV U319 ( .A(B[238]), .Z(n751) );
  IV U320 ( .A(B[239]), .Z(n752) );
  IV U321 ( .A(B[240]), .Z(n753) );
  IV U322 ( .A(B[241]), .Z(n754) );
  IV U323 ( .A(B[242]), .Z(n755) );
  IV U324 ( .A(B[243]), .Z(n756) );
  IV U325 ( .A(B[244]), .Z(n757) );
  IV U326 ( .A(B[487]), .Z(n1000) );
  IV U327 ( .A(B[245]), .Z(n758) );
  IV U328 ( .A(B[246]), .Z(n759) );
  IV U329 ( .A(B[247]), .Z(n760) );
  IV U330 ( .A(B[248]), .Z(n761) );
  IV U331 ( .A(B[249]), .Z(n762) );
  IV U332 ( .A(B[250]), .Z(n763) );
  IV U333 ( .A(B[251]), .Z(n764) );
  IV U334 ( .A(B[252]), .Z(n765) );
  IV U335 ( .A(B[253]), .Z(n766) );
  IV U336 ( .A(B[254]), .Z(n767) );
  IV U337 ( .A(B[488]), .Z(n1001) );
  IV U338 ( .A(B[255]), .Z(n768) );
  IV U339 ( .A(B[256]), .Z(n769) );
  IV U340 ( .A(B[257]), .Z(n770) );
  IV U341 ( .A(B[258]), .Z(n771) );
  IV U342 ( .A(B[259]), .Z(n772) );
  IV U343 ( .A(B[260]), .Z(n773) );
  IV U344 ( .A(B[261]), .Z(n774) );
  IV U345 ( .A(B[262]), .Z(n775) );
  IV U346 ( .A(B[263]), .Z(n776) );
  IV U347 ( .A(B[264]), .Z(n777) );
  IV U348 ( .A(B[489]), .Z(n1002) );
  IV U349 ( .A(B[265]), .Z(n778) );
  IV U350 ( .A(B[266]), .Z(n779) );
  IV U351 ( .A(B[267]), .Z(n780) );
  IV U352 ( .A(B[268]), .Z(n781) );
  IV U353 ( .A(B[269]), .Z(n782) );
  IV U354 ( .A(B[270]), .Z(n783) );
  IV U355 ( .A(B[271]), .Z(n784) );
  IV U356 ( .A(B[272]), .Z(n785) );
  IV U357 ( .A(B[273]), .Z(n786) );
  IV U358 ( .A(B[274]), .Z(n787) );
  IV U359 ( .A(B[490]), .Z(n1003) );
  IV U360 ( .A(B[275]), .Z(n788) );
  IV U361 ( .A(B[276]), .Z(n789) );
  IV U362 ( .A(B[277]), .Z(n790) );
  IV U363 ( .A(B[278]), .Z(n791) );
  IV U364 ( .A(B[279]), .Z(n792) );
  IV U365 ( .A(B[280]), .Z(n793) );
  IV U366 ( .A(B[281]), .Z(n794) );
  IV U367 ( .A(B[282]), .Z(n795) );
  IV U368 ( .A(B[283]), .Z(n796) );
  IV U369 ( .A(B[284]), .Z(n797) );
  IV U370 ( .A(B[491]), .Z(n1004) );
  IV U371 ( .A(B[285]), .Z(n798) );
  IV U372 ( .A(B[286]), .Z(n799) );
  IV U373 ( .A(B[287]), .Z(n800) );
  IV U374 ( .A(B[288]), .Z(n801) );
  IV U375 ( .A(B[289]), .Z(n802) );
  IV U376 ( .A(B[290]), .Z(n803) );
  IV U377 ( .A(B[291]), .Z(n804) );
  IV U378 ( .A(B[292]), .Z(n805) );
  IV U379 ( .A(B[293]), .Z(n806) );
  IV U380 ( .A(B[294]), .Z(n807) );
  IV U381 ( .A(B[492]), .Z(n1005) );
  IV U382 ( .A(B[295]), .Z(n808) );
  IV U383 ( .A(B[296]), .Z(n809) );
  IV U384 ( .A(B[297]), .Z(n810) );
  IV U385 ( .A(B[298]), .Z(n811) );
  IV U386 ( .A(B[299]), .Z(n812) );
  IV U387 ( .A(B[300]), .Z(n813) );
  IV U388 ( .A(B[301]), .Z(n814) );
  IV U389 ( .A(B[302]), .Z(n815) );
  IV U390 ( .A(B[303]), .Z(n816) );
  IV U391 ( .A(B[304]), .Z(n817) );
  IV U392 ( .A(B[493]), .Z(n1006) );
  IV U393 ( .A(B[305]), .Z(n818) );
  IV U394 ( .A(B[306]), .Z(n819) );
  IV U395 ( .A(B[307]), .Z(n820) );
  IV U396 ( .A(B[308]), .Z(n821) );
  IV U397 ( .A(B[309]), .Z(n822) );
  IV U398 ( .A(B[310]), .Z(n823) );
  IV U399 ( .A(B[311]), .Z(n824) );
  IV U400 ( .A(B[312]), .Z(n825) );
  IV U401 ( .A(B[313]), .Z(n826) );
  IV U402 ( .A(B[314]), .Z(n827) );
  IV U403 ( .A(B[494]), .Z(n1007) );
  IV U404 ( .A(B[315]), .Z(n828) );
  IV U405 ( .A(B[316]), .Z(n829) );
  IV U406 ( .A(B[317]), .Z(n830) );
  IV U407 ( .A(B[318]), .Z(n831) );
  IV U408 ( .A(B[319]), .Z(n832) );
  IV U409 ( .A(B[320]), .Z(n833) );
  IV U410 ( .A(B[321]), .Z(n834) );
  IV U411 ( .A(B[322]), .Z(n835) );
  IV U412 ( .A(B[323]), .Z(n836) );
  IV U413 ( .A(B[324]), .Z(n837) );
  IV U414 ( .A(B[495]), .Z(n1008) );
  IV U415 ( .A(B[325]), .Z(n838) );
  IV U416 ( .A(B[326]), .Z(n839) );
  IV U417 ( .A(B[327]), .Z(n840) );
  IV U418 ( .A(B[328]), .Z(n841) );
  IV U419 ( .A(B[329]), .Z(n842) );
  IV U420 ( .A(B[330]), .Z(n843) );
  IV U421 ( .A(B[331]), .Z(n844) );
  IV U422 ( .A(B[332]), .Z(n845) );
  IV U423 ( .A(B[333]), .Z(n846) );
  IV U424 ( .A(B[334]), .Z(n847) );
  IV U425 ( .A(B[496]), .Z(n1009) );
  IV U426 ( .A(B[335]), .Z(n848) );
  IV U427 ( .A(B[336]), .Z(n849) );
  IV U428 ( .A(B[337]), .Z(n850) );
  IV U429 ( .A(B[338]), .Z(n851) );
  IV U430 ( .A(B[339]), .Z(n852) );
  IV U431 ( .A(B[340]), .Z(n853) );
  IV U432 ( .A(B[341]), .Z(n854) );
  IV U433 ( .A(B[342]), .Z(n855) );
  IV U434 ( .A(B[343]), .Z(n856) );
  IV U435 ( .A(B[344]), .Z(n857) );
  IV U436 ( .A(B[497]), .Z(n1010) );
  IV U437 ( .A(B[345]), .Z(n858) );
  IV U438 ( .A(B[346]), .Z(n859) );
  IV U439 ( .A(B[347]), .Z(n860) );
  IV U440 ( .A(B[348]), .Z(n861) );
  IV U441 ( .A(B[349]), .Z(n862) );
  IV U442 ( .A(B[350]), .Z(n863) );
  IV U443 ( .A(B[351]), .Z(n864) );
  IV U444 ( .A(B[352]), .Z(n865) );
  IV U445 ( .A(B[353]), .Z(n866) );
  IV U446 ( .A(B[354]), .Z(n867) );
  IV U447 ( .A(B[498]), .Z(n1011) );
  IV U448 ( .A(B[355]), .Z(n868) );
  IV U449 ( .A(B[356]), .Z(n869) );
  IV U450 ( .A(B[357]), .Z(n870) );
  IV U451 ( .A(B[358]), .Z(n871) );
  IV U452 ( .A(B[359]), .Z(n872) );
  IV U453 ( .A(B[360]), .Z(n873) );
  IV U454 ( .A(B[361]), .Z(n874) );
  IV U455 ( .A(B[362]), .Z(n875) );
  IV U456 ( .A(B[363]), .Z(n876) );
  IV U457 ( .A(B[364]), .Z(n877) );
  IV U458 ( .A(B[499]), .Z(n1012) );
  IV U459 ( .A(B[365]), .Z(n878) );
  IV U460 ( .A(B[366]), .Z(n879) );
  IV U461 ( .A(B[367]), .Z(n880) );
  IV U462 ( .A(B[368]), .Z(n881) );
  IV U463 ( .A(B[369]), .Z(n882) );
  IV U464 ( .A(B[370]), .Z(n883) );
  IV U465 ( .A(B[371]), .Z(n884) );
  IV U466 ( .A(B[372]), .Z(n885) );
  IV U467 ( .A(B[373]), .Z(n886) );
  IV U468 ( .A(B[374]), .Z(n887) );
  IV U469 ( .A(B[500]), .Z(n1013) );
  IV U470 ( .A(B[375]), .Z(n888) );
  IV U471 ( .A(B[376]), .Z(n889) );
  IV U472 ( .A(B[377]), .Z(n890) );
  IV U473 ( .A(B[378]), .Z(n891) );
  IV U474 ( .A(B[379]), .Z(n892) );
  IV U475 ( .A(B[380]), .Z(n893) );
  IV U476 ( .A(B[381]), .Z(n894) );
  IV U477 ( .A(B[382]), .Z(n895) );
  IV U478 ( .A(B[383]), .Z(n896) );
  IV U479 ( .A(B[384]), .Z(n897) );
  IV U480 ( .A(B[501]), .Z(n1014) );
  IV U481 ( .A(B[385]), .Z(n898) );
  IV U482 ( .A(B[386]), .Z(n899) );
  IV U483 ( .A(B[387]), .Z(n900) );
  IV U484 ( .A(B[388]), .Z(n901) );
  IV U485 ( .A(B[389]), .Z(n902) );
  IV U486 ( .A(B[390]), .Z(n903) );
  IV U487 ( .A(B[391]), .Z(n904) );
  IV U488 ( .A(B[392]), .Z(n905) );
  IV U489 ( .A(B[393]), .Z(n906) );
  IV U490 ( .A(B[394]), .Z(n907) );
  IV U491 ( .A(B[502]), .Z(n1015) );
  IV U492 ( .A(B[395]), .Z(n908) );
  IV U493 ( .A(B[396]), .Z(n909) );
  IV U494 ( .A(B[397]), .Z(n910) );
  IV U495 ( .A(B[398]), .Z(n911) );
  IV U496 ( .A(B[399]), .Z(n912) );
  IV U497 ( .A(B[400]), .Z(n913) );
  IV U498 ( .A(B[401]), .Z(n914) );
  IV U499 ( .A(B[402]), .Z(n915) );
  IV U500 ( .A(B[403]), .Z(n916) );
  IV U501 ( .A(B[404]), .Z(n917) );
  IV U502 ( .A(B[503]), .Z(n1016) );
  IV U503 ( .A(B[405]), .Z(n918) );
  IV U504 ( .A(B[406]), .Z(n919) );
  IV U505 ( .A(B[407]), .Z(n920) );
  IV U506 ( .A(B[408]), .Z(n921) );
  IV U507 ( .A(B[409]), .Z(n922) );
  IV U508 ( .A(B[410]), .Z(n923) );
  IV U509 ( .A(B[411]), .Z(n924) );
  IV U510 ( .A(B[412]), .Z(n925) );
  IV U511 ( .A(B[413]), .Z(n926) );
  IV U512 ( .A(B[414]), .Z(n927) );
  IV U513 ( .A(B[504]), .Z(n1017) );
endmodule


module modmult_step_N512 ( xregN_1, y, n, zin, zout );
  input [511:0] y;
  input [511:0] n;
  input [513:0] zin;
  output [513:0] zout;
  input xregN_1;
  wire   c1, c2, n1;
  wire   [513:0] w1;
  wire   [513:0] w2;
  wire   [513:0] w3;
  wire   [513:0] z2;
  wire   [513:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6;

  MUX_N514_0 MUX_1 ( .A({1'b0, 1'b0, y}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(xregN_1), .O({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, w1[511:0]}) );
  MUX_N514_2 MUX_2 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(c1), .O({SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, w2[511:0]}) );
  MUX_N514_1 MUX_3 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(n1), .O({SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, w3[511:0]}) );
  ADD_N514 ADD_1 ( .A({zin[512:0], 1'b0}), .B({1'b0, 1'b0, w1[511:0]}), .CI(
        1'b0), .S(z2) );
  COMP_N514_0 COMP_1 ( .A(z2), .B({1'b0, 1'b0, n}), .O(c1) );
  SUB_N514_0 SUB_1 ( .A(z2), .B({1'b0, 1'b0, w2[511:0]}), .S(z3) );
  COMP_N514_1 COMP_2 ( .A({1'b0, 1'b0, n}), .B(z3), .O(c2) );
  SUB_N514_1 SUB_2 ( .A({1'b0, z3[512:0]}), .B({1'b0, 1'b0, w3[511:0]}), .S({
        SYNOPSYS_UNCONNECTED__6, zout[512:0]}) );
  IV U2 ( .A(c2), .Z(n1) );
endmodule


module modmult_N512_CC512 ( clk, rst, start, x, y, n, o );
  input [511:0] x;
  input [511:0] y;
  input [511:0] n;
  output [511:0] o;
  input clk, rst, start;
  wire   \zout[0][512] , \zin[0][512] , \zin[0][511] , \zin[0][510] ,
         \zin[0][509] , \zin[0][508] , \zin[0][507] , \zin[0][506] ,
         \zin[0][505] , \zin[0][504] , \zin[0][503] , \zin[0][502] ,
         \zin[0][501] , \zin[0][500] , \zin[0][499] , \zin[0][498] ,
         \zin[0][497] , \zin[0][496] , \zin[0][495] , \zin[0][494] ,
         \zin[0][493] , \zin[0][492] , \zin[0][491] , \zin[0][490] ,
         \zin[0][489] , \zin[0][488] , \zin[0][487] , \zin[0][486] ,
         \zin[0][485] , \zin[0][484] , \zin[0][483] , \zin[0][482] ,
         \zin[0][481] , \zin[0][480] , \zin[0][479] , \zin[0][478] ,
         \zin[0][477] , \zin[0][476] , \zin[0][475] , \zin[0][474] ,
         \zin[0][473] , \zin[0][472] , \zin[0][471] , \zin[0][470] ,
         \zin[0][469] , \zin[0][468] , \zin[0][467] , \zin[0][466] ,
         \zin[0][465] , \zin[0][464] , \zin[0][463] , \zin[0][462] ,
         \zin[0][461] , \zin[0][460] , \zin[0][459] , \zin[0][458] ,
         \zin[0][457] , \zin[0][456] , \zin[0][455] , \zin[0][454] ,
         \zin[0][453] , \zin[0][452] , \zin[0][451] , \zin[0][450] ,
         \zin[0][449] , \zin[0][448] , \zin[0][447] , \zin[0][446] ,
         \zin[0][445] , \zin[0][444] , \zin[0][443] , \zin[0][442] ,
         \zin[0][441] , \zin[0][440] , \zin[0][439] , \zin[0][438] ,
         \zin[0][437] , \zin[0][436] , \zin[0][435] , \zin[0][434] ,
         \zin[0][433] , \zin[0][432] , \zin[0][431] , \zin[0][430] ,
         \zin[0][429] , \zin[0][428] , \zin[0][427] , \zin[0][426] ,
         \zin[0][425] , \zin[0][424] , \zin[0][423] , \zin[0][422] ,
         \zin[0][421] , \zin[0][420] , \zin[0][419] , \zin[0][418] ,
         \zin[0][417] , \zin[0][416] , \zin[0][415] , \zin[0][414] ,
         \zin[0][413] , \zin[0][412] , \zin[0][411] , \zin[0][410] ,
         \zin[0][409] , \zin[0][408] , \zin[0][407] , \zin[0][406] ,
         \zin[0][405] , \zin[0][404] , \zin[0][403] , \zin[0][402] ,
         \zin[0][401] , \zin[0][400] , \zin[0][399] , \zin[0][398] ,
         \zin[0][397] , \zin[0][396] , \zin[0][395] , \zin[0][394] ,
         \zin[0][393] , \zin[0][392] , \zin[0][391] , \zin[0][390] ,
         \zin[0][389] , \zin[0][388] , \zin[0][387] , \zin[0][386] ,
         \zin[0][385] , \zin[0][384] , \zin[0][383] , \zin[0][382] ,
         \zin[0][381] , \zin[0][380] , \zin[0][379] , \zin[0][378] ,
         \zin[0][377] , \zin[0][376] , \zin[0][375] , \zin[0][374] ,
         \zin[0][373] , \zin[0][372] , \zin[0][371] , \zin[0][370] ,
         \zin[0][369] , \zin[0][368] , \zin[0][367] , \zin[0][366] ,
         \zin[0][365] , \zin[0][364] , \zin[0][363] , \zin[0][362] ,
         \zin[0][361] , \zin[0][360] , \zin[0][359] , \zin[0][358] ,
         \zin[0][357] , \zin[0][356] , \zin[0][355] , \zin[0][354] ,
         \zin[0][353] , \zin[0][352] , \zin[0][351] , \zin[0][350] ,
         \zin[0][349] , \zin[0][348] , \zin[0][347] , \zin[0][346] ,
         \zin[0][345] , \zin[0][344] , \zin[0][343] , \zin[0][342] ,
         \zin[0][341] , \zin[0][340] , \zin[0][339] , \zin[0][338] ,
         \zin[0][337] , \zin[0][336] , \zin[0][335] , \zin[0][334] ,
         \zin[0][333] , \zin[0][332] , \zin[0][331] , \zin[0][330] ,
         \zin[0][329] , \zin[0][328] , \zin[0][327] , \zin[0][326] ,
         \zin[0][325] , \zin[0][324] , \zin[0][323] , \zin[0][322] ,
         \zin[0][321] , \zin[0][320] , \zin[0][319] , \zin[0][318] ,
         \zin[0][317] , \zin[0][316] , \zin[0][315] , \zin[0][314] ,
         \zin[0][313] , \zin[0][312] , \zin[0][311] , \zin[0][310] ,
         \zin[0][309] , \zin[0][308] , \zin[0][307] , \zin[0][306] ,
         \zin[0][305] , \zin[0][304] , \zin[0][303] , \zin[0][302] ,
         \zin[0][301] , \zin[0][300] , \zin[0][299] , \zin[0][298] ,
         \zin[0][297] , \zin[0][296] , \zin[0][295] , \zin[0][294] ,
         \zin[0][293] , \zin[0][292] , \zin[0][291] , \zin[0][290] ,
         \zin[0][289] , \zin[0][288] , \zin[0][287] , \zin[0][286] ,
         \zin[0][285] , \zin[0][284] , \zin[0][283] , \zin[0][282] ,
         \zin[0][281] , \zin[0][280] , \zin[0][279] , \zin[0][278] ,
         \zin[0][277] , \zin[0][276] , \zin[0][275] , \zin[0][274] ,
         \zin[0][273] , \zin[0][272] , \zin[0][271] , \zin[0][270] ,
         \zin[0][269] , \zin[0][268] , \zin[0][267] , \zin[0][266] ,
         \zin[0][265] , \zin[0][264] , \zin[0][263] , \zin[0][262] ,
         \zin[0][261] , \zin[0][260] , \zin[0][259] , \zin[0][258] ,
         \zin[0][257] , \zin[0][256] , \zin[0][255] , \zin[0][254] ,
         \zin[0][253] , \zin[0][252] , \zin[0][251] , \zin[0][250] ,
         \zin[0][249] , \zin[0][248] , \zin[0][247] , \zin[0][246] ,
         \zin[0][245] , \zin[0][244] , \zin[0][243] , \zin[0][242] ,
         \zin[0][241] , \zin[0][240] , \zin[0][239] , \zin[0][238] ,
         \zin[0][237] , \zin[0][236] , \zin[0][235] , \zin[0][234] ,
         \zin[0][233] , \zin[0][232] , \zin[0][231] , \zin[0][230] ,
         \zin[0][229] , \zin[0][228] , \zin[0][227] , \zin[0][226] ,
         \zin[0][225] , \zin[0][224] , \zin[0][223] , \zin[0][222] ,
         \zin[0][221] , \zin[0][220] , \zin[0][219] , \zin[0][218] ,
         \zin[0][217] , \zin[0][216] , \zin[0][215] , \zin[0][214] ,
         \zin[0][213] , \zin[0][212] , \zin[0][211] , \zin[0][210] ,
         \zin[0][209] , \zin[0][208] , \zin[0][207] , \zin[0][206] ,
         \zin[0][205] , \zin[0][204] , \zin[0][203] , \zin[0][202] ,
         \zin[0][201] , \zin[0][200] , \zin[0][199] , \zin[0][198] ,
         \zin[0][197] , \zin[0][196] , \zin[0][195] , \zin[0][194] ,
         \zin[0][193] , \zin[0][192] , \zin[0][191] , \zin[0][190] ,
         \zin[0][189] , \zin[0][188] , \zin[0][187] , \zin[0][186] ,
         \zin[0][185] , \zin[0][184] , \zin[0][183] , \zin[0][182] ,
         \zin[0][181] , \zin[0][180] , \zin[0][179] , \zin[0][178] ,
         \zin[0][177] , \zin[0][176] , \zin[0][175] , \zin[0][174] ,
         \zin[0][173] , \zin[0][172] , \zin[0][171] , \zin[0][170] ,
         \zin[0][169] , \zin[0][168] , \zin[0][167] , \zin[0][166] ,
         \zin[0][165] , \zin[0][164] , \zin[0][163] , \zin[0][162] ,
         \zin[0][161] , \zin[0][160] , \zin[0][159] , \zin[0][158] ,
         \zin[0][157] , \zin[0][156] , \zin[0][155] , \zin[0][154] ,
         \zin[0][153] , \zin[0][152] , \zin[0][151] , \zin[0][150] ,
         \zin[0][149] , \zin[0][148] , \zin[0][147] , \zin[0][146] ,
         \zin[0][145] , \zin[0][144] , \zin[0][143] , \zin[0][142] ,
         \zin[0][141] , \zin[0][140] , \zin[0][139] , \zin[0][138] ,
         \zin[0][137] , \zin[0][136] , \zin[0][135] , \zin[0][134] ,
         \zin[0][133] , \zin[0][132] , \zin[0][131] , \zin[0][130] ,
         \zin[0][129] , \zin[0][128] , \zin[0][127] , \zin[0][126] ,
         \zin[0][125] , \zin[0][124] , \zin[0][123] , \zin[0][122] ,
         \zin[0][121] , \zin[0][120] , \zin[0][119] , \zin[0][118] ,
         \zin[0][117] , \zin[0][116] , \zin[0][115] , \zin[0][114] ,
         \zin[0][113] , \zin[0][112] , \zin[0][111] , \zin[0][110] ,
         \zin[0][109] , \zin[0][108] , \zin[0][107] , \zin[0][106] ,
         \zin[0][105] , \zin[0][104] , \zin[0][103] , \zin[0][102] ,
         \zin[0][101] , \zin[0][100] , \zin[0][99] , \zin[0][98] ,
         \zin[0][97] , \zin[0][96] , \zin[0][95] , \zin[0][94] , \zin[0][93] ,
         \zin[0][92] , \zin[0][91] , \zin[0][90] , \zin[0][89] , \zin[0][88] ,
         \zin[0][87] , \zin[0][86] , \zin[0][85] , \zin[0][84] , \zin[0][83] ,
         \zin[0][82] , \zin[0][81] , \zin[0][80] , \zin[0][79] , \zin[0][78] ,
         \zin[0][77] , \zin[0][76] , \zin[0][75] , \zin[0][74] , \zin[0][73] ,
         \zin[0][72] , \zin[0][71] , \zin[0][70] , \zin[0][69] , \zin[0][68] ,
         \zin[0][67] , \zin[0][66] , \zin[0][65] , \zin[0][64] , \zin[0][63] ,
         \zin[0][62] , \zin[0][61] , \zin[0][60] , \zin[0][59] , \zin[0][58] ,
         \zin[0][57] , \zin[0][56] , \zin[0][55] , \zin[0][54] , \zin[0][53] ,
         \zin[0][52] , \zin[0][51] , \zin[0][50] , \zin[0][49] , \zin[0][48] ,
         \zin[0][47] , \zin[0][46] , \zin[0][45] , \zin[0][44] , \zin[0][43] ,
         \zin[0][42] , \zin[0][41] , \zin[0][40] , \zin[0][39] , \zin[0][38] ,
         \zin[0][37] , \zin[0][36] , \zin[0][35] , \zin[0][34] , \zin[0][33] ,
         \zin[0][32] , \zin[0][31] , \zin[0][30] , \zin[0][29] , \zin[0][28] ,
         \zin[0][27] , \zin[0][26] , \zin[0][25] , \zin[0][24] , \zin[0][23] ,
         \zin[0][22] , \zin[0][21] , \zin[0][20] , \zin[0][19] , \zin[0][18] ,
         \zin[0][17] , \zin[0][16] , \zin[0][15] , \zin[0][14] , \zin[0][13] ,
         \zin[0][12] , \zin[0][11] , \zin[0][10] , \zin[0][9] , \zin[0][8] ,
         \zin[0][7] , \zin[0][6] , \zin[0][5] , \zin[0][4] , \zin[0][3] ,
         \zin[0][2] , \zin[0][1] , \zin[0][0] ;
  wire   [511:0] xin;
  wire   SYNOPSYS_UNCONNECTED__0;

  modmult_step_N512 \MODMULT_STEP[0].modmult_step_  ( .xregN_1(xin[511]), .y(y), .n(n), .zin({1'b0, \zin[0][512] , \zin[0][511] , \zin[0][510] , 
        \zin[0][509] , \zin[0][508] , \zin[0][507] , \zin[0][506] , 
        \zin[0][505] , \zin[0][504] , \zin[0][503] , \zin[0][502] , 
        \zin[0][501] , \zin[0][500] , \zin[0][499] , \zin[0][498] , 
        \zin[0][497] , \zin[0][496] , \zin[0][495] , \zin[0][494] , 
        \zin[0][493] , \zin[0][492] , \zin[0][491] , \zin[0][490] , 
        \zin[0][489] , \zin[0][488] , \zin[0][487] , \zin[0][486] , 
        \zin[0][485] , \zin[0][484] , \zin[0][483] , \zin[0][482] , 
        \zin[0][481] , \zin[0][480] , \zin[0][479] , \zin[0][478] , 
        \zin[0][477] , \zin[0][476] , \zin[0][475] , \zin[0][474] , 
        \zin[0][473] , \zin[0][472] , \zin[0][471] , \zin[0][470] , 
        \zin[0][469] , \zin[0][468] , \zin[0][467] , \zin[0][466] , 
        \zin[0][465] , \zin[0][464] , \zin[0][463] , \zin[0][462] , 
        \zin[0][461] , \zin[0][460] , \zin[0][459] , \zin[0][458] , 
        \zin[0][457] , \zin[0][456] , \zin[0][455] , \zin[0][454] , 
        \zin[0][453] , \zin[0][452] , \zin[0][451] , \zin[0][450] , 
        \zin[0][449] , \zin[0][448] , \zin[0][447] , \zin[0][446] , 
        \zin[0][445] , \zin[0][444] , \zin[0][443] , \zin[0][442] , 
        \zin[0][441] , \zin[0][440] , \zin[0][439] , \zin[0][438] , 
        \zin[0][437] , \zin[0][436] , \zin[0][435] , \zin[0][434] , 
        \zin[0][433] , \zin[0][432] , \zin[0][431] , \zin[0][430] , 
        \zin[0][429] , \zin[0][428] , \zin[0][427] , \zin[0][426] , 
        \zin[0][425] , \zin[0][424] , \zin[0][423] , \zin[0][422] , 
        \zin[0][421] , \zin[0][420] , \zin[0][419] , \zin[0][418] , 
        \zin[0][417] , \zin[0][416] , \zin[0][415] , \zin[0][414] , 
        \zin[0][413] , \zin[0][412] , \zin[0][411] , \zin[0][410] , 
        \zin[0][409] , \zin[0][408] , \zin[0][407] , \zin[0][406] , 
        \zin[0][405] , \zin[0][404] , \zin[0][403] , \zin[0][402] , 
        \zin[0][401] , \zin[0][400] , \zin[0][399] , \zin[0][398] , 
        \zin[0][397] , \zin[0][396] , \zin[0][395] , \zin[0][394] , 
        \zin[0][393] , \zin[0][392] , \zin[0][391] , \zin[0][390] , 
        \zin[0][389] , \zin[0][388] , \zin[0][387] , \zin[0][386] , 
        \zin[0][385] , \zin[0][384] , \zin[0][383] , \zin[0][382] , 
        \zin[0][381] , \zin[0][380] , \zin[0][379] , \zin[0][378] , 
        \zin[0][377] , \zin[0][376] , \zin[0][375] , \zin[0][374] , 
        \zin[0][373] , \zin[0][372] , \zin[0][371] , \zin[0][370] , 
        \zin[0][369] , \zin[0][368] , \zin[0][367] , \zin[0][366] , 
        \zin[0][365] , \zin[0][364] , \zin[0][363] , \zin[0][362] , 
        \zin[0][361] , \zin[0][360] , \zin[0][359] , \zin[0][358] , 
        \zin[0][357] , \zin[0][356] , \zin[0][355] , \zin[0][354] , 
        \zin[0][353] , \zin[0][352] , \zin[0][351] , \zin[0][350] , 
        \zin[0][349] , \zin[0][348] , \zin[0][347] , \zin[0][346] , 
        \zin[0][345] , \zin[0][344] , \zin[0][343] , \zin[0][342] , 
        \zin[0][341] , \zin[0][340] , \zin[0][339] , \zin[0][338] , 
        \zin[0][337] , \zin[0][336] , \zin[0][335] , \zin[0][334] , 
        \zin[0][333] , \zin[0][332] , \zin[0][331] , \zin[0][330] , 
        \zin[0][329] , \zin[0][328] , \zin[0][327] , \zin[0][326] , 
        \zin[0][325] , \zin[0][324] , \zin[0][323] , \zin[0][322] , 
        \zin[0][321] , \zin[0][320] , \zin[0][319] , \zin[0][318] , 
        \zin[0][317] , \zin[0][316] , \zin[0][315] , \zin[0][314] , 
        \zin[0][313] , \zin[0][312] , \zin[0][311] , \zin[0][310] , 
        \zin[0][309] , \zin[0][308] , \zin[0][307] , \zin[0][306] , 
        \zin[0][305] , \zin[0][304] , \zin[0][303] , \zin[0][302] , 
        \zin[0][301] , \zin[0][300] , \zin[0][299] , \zin[0][298] , 
        \zin[0][297] , \zin[0][296] , \zin[0][295] , \zin[0][294] , 
        \zin[0][293] , \zin[0][292] , \zin[0][291] , \zin[0][290] , 
        \zin[0][289] , \zin[0][288] , \zin[0][287] , \zin[0][286] , 
        \zin[0][285] , \zin[0][284] , \zin[0][283] , \zin[0][282] , 
        \zin[0][281] , \zin[0][280] , \zin[0][279] , \zin[0][278] , 
        \zin[0][277] , \zin[0][276] , \zin[0][275] , \zin[0][274] , 
        \zin[0][273] , \zin[0][272] , \zin[0][271] , \zin[0][270] , 
        \zin[0][269] , \zin[0][268] , \zin[0][267] , \zin[0][266] , 
        \zin[0][265] , \zin[0][264] , \zin[0][263] , \zin[0][262] , 
        \zin[0][261] , \zin[0][260] , \zin[0][259] , \zin[0][258] , 
        \zin[0][257] , \zin[0][256] , \zin[0][255] , \zin[0][254] , 
        \zin[0][253] , \zin[0][252] , \zin[0][251] , \zin[0][250] , 
        \zin[0][249] , \zin[0][248] , \zin[0][247] , \zin[0][246] , 
        \zin[0][245] , \zin[0][244] , \zin[0][243] , \zin[0][242] , 
        \zin[0][241] , \zin[0][240] , \zin[0][239] , \zin[0][238] , 
        \zin[0][237] , \zin[0][236] , \zin[0][235] , \zin[0][234] , 
        \zin[0][233] , \zin[0][232] , \zin[0][231] , \zin[0][230] , 
        \zin[0][229] , \zin[0][228] , \zin[0][227] , \zin[0][226] , 
        \zin[0][225] , \zin[0][224] , \zin[0][223] , \zin[0][222] , 
        \zin[0][221] , \zin[0][220] , \zin[0][219] , \zin[0][218] , 
        \zin[0][217] , \zin[0][216] , \zin[0][215] , \zin[0][214] , 
        \zin[0][213] , \zin[0][212] , \zin[0][211] , \zin[0][210] , 
        \zin[0][209] , \zin[0][208] , \zin[0][207] , \zin[0][206] , 
        \zin[0][205] , \zin[0][204] , \zin[0][203] , \zin[0][202] , 
        \zin[0][201] , \zin[0][200] , \zin[0][199] , \zin[0][198] , 
        \zin[0][197] , \zin[0][196] , \zin[0][195] , \zin[0][194] , 
        \zin[0][193] , \zin[0][192] , \zin[0][191] , \zin[0][190] , 
        \zin[0][189] , \zin[0][188] , \zin[0][187] , \zin[0][186] , 
        \zin[0][185] , \zin[0][184] , \zin[0][183] , \zin[0][182] , 
        \zin[0][181] , \zin[0][180] , \zin[0][179] , \zin[0][178] , 
        \zin[0][177] , \zin[0][176] , \zin[0][175] , \zin[0][174] , 
        \zin[0][173] , \zin[0][172] , \zin[0][171] , \zin[0][170] , 
        \zin[0][169] , \zin[0][168] , \zin[0][167] , \zin[0][166] , 
        \zin[0][165] , \zin[0][164] , \zin[0][163] , \zin[0][162] , 
        \zin[0][161] , \zin[0][160] , \zin[0][159] , \zin[0][158] , 
        \zin[0][157] , \zin[0][156] , \zin[0][155] , \zin[0][154] , 
        \zin[0][153] , \zin[0][152] , \zin[0][151] , \zin[0][150] , 
        \zin[0][149] , \zin[0][148] , \zin[0][147] , \zin[0][146] , 
        \zin[0][145] , \zin[0][144] , \zin[0][143] , \zin[0][142] , 
        \zin[0][141] , \zin[0][140] , \zin[0][139] , \zin[0][138] , 
        \zin[0][137] , \zin[0][136] , \zin[0][135] , \zin[0][134] , 
        \zin[0][133] , \zin[0][132] , \zin[0][131] , \zin[0][130] , 
        \zin[0][129] , \zin[0][128] , \zin[0][127] , \zin[0][126] , 
        \zin[0][125] , \zin[0][124] , \zin[0][123] , \zin[0][122] , 
        \zin[0][121] , \zin[0][120] , \zin[0][119] , \zin[0][118] , 
        \zin[0][117] , \zin[0][116] , \zin[0][115] , \zin[0][114] , 
        \zin[0][113] , \zin[0][112] , \zin[0][111] , \zin[0][110] , 
        \zin[0][109] , \zin[0][108] , \zin[0][107] , \zin[0][106] , 
        \zin[0][105] , \zin[0][104] , \zin[0][103] , \zin[0][102] , 
        \zin[0][101] , \zin[0][100] , \zin[0][99] , \zin[0][98] , \zin[0][97] , 
        \zin[0][96] , \zin[0][95] , \zin[0][94] , \zin[0][93] , \zin[0][92] , 
        \zin[0][91] , \zin[0][90] , \zin[0][89] , \zin[0][88] , \zin[0][87] , 
        \zin[0][86] , \zin[0][85] , \zin[0][84] , \zin[0][83] , \zin[0][82] , 
        \zin[0][81] , \zin[0][80] , \zin[0][79] , \zin[0][78] , \zin[0][77] , 
        \zin[0][76] , \zin[0][75] , \zin[0][74] , \zin[0][73] , \zin[0][72] , 
        \zin[0][71] , \zin[0][70] , \zin[0][69] , \zin[0][68] , \zin[0][67] , 
        \zin[0][66] , \zin[0][65] , \zin[0][64] , \zin[0][63] , \zin[0][62] , 
        \zin[0][61] , \zin[0][60] , \zin[0][59] , \zin[0][58] , \zin[0][57] , 
        \zin[0][56] , \zin[0][55] , \zin[0][54] , \zin[0][53] , \zin[0][52] , 
        \zin[0][51] , \zin[0][50] , \zin[0][49] , \zin[0][48] , \zin[0][47] , 
        \zin[0][46] , \zin[0][45] , \zin[0][44] , \zin[0][43] , \zin[0][42] , 
        \zin[0][41] , \zin[0][40] , \zin[0][39] , \zin[0][38] , \zin[0][37] , 
        \zin[0][36] , \zin[0][35] , \zin[0][34] , \zin[0][33] , \zin[0][32] , 
        \zin[0][31] , \zin[0][30] , \zin[0][29] , \zin[0][28] , \zin[0][27] , 
        \zin[0][26] , \zin[0][25] , \zin[0][24] , \zin[0][23] , \zin[0][22] , 
        \zin[0][21] , \zin[0][20] , \zin[0][19] , \zin[0][18] , \zin[0][17] , 
        \zin[0][16] , \zin[0][15] , \zin[0][14] , \zin[0][13] , \zin[0][12] , 
        \zin[0][11] , \zin[0][10] , \zin[0][9] , \zin[0][8] , \zin[0][7] , 
        \zin[0][6] , \zin[0][5] , \zin[0][4] , \zin[0][3] , \zin[0][2] , 
        \zin[0][1] , \zin[0][0] }), .zout({SYNOPSYS_UNCONNECTED__0, 
        \zout[0][512] , o}) );
  DFF \xreg_reg[0]  ( .D(1'b0), .CLK(clk), .RST(start), .I(x[0]), .Q(xin[0])
         );
  DFF \xreg_reg[1]  ( .D(xin[0]), .CLK(clk), .RST(start), .I(x[1]), .Q(xin[1])
         );
  DFF \xreg_reg[2]  ( .D(xin[1]), .CLK(clk), .RST(start), .I(x[2]), .Q(xin[2])
         );
  DFF \xreg_reg[3]  ( .D(xin[2]), .CLK(clk), .RST(start), .I(x[3]), .Q(xin[3])
         );
  DFF \xreg_reg[4]  ( .D(xin[3]), .CLK(clk), .RST(start), .I(x[4]), .Q(xin[4])
         );
  DFF \xreg_reg[5]  ( .D(xin[4]), .CLK(clk), .RST(start), .I(x[5]), .Q(xin[5])
         );
  DFF \xreg_reg[6]  ( .D(xin[5]), .CLK(clk), .RST(start), .I(x[6]), .Q(xin[6])
         );
  DFF \xreg_reg[7]  ( .D(xin[6]), .CLK(clk), .RST(start), .I(x[7]), .Q(xin[7])
         );
  DFF \xreg_reg[8]  ( .D(xin[7]), .CLK(clk), .RST(start), .I(x[8]), .Q(xin[8])
         );
  DFF \xreg_reg[9]  ( .D(xin[8]), .CLK(clk), .RST(start), .I(x[9]), .Q(xin[9])
         );
  DFF \xreg_reg[10]  ( .D(xin[9]), .CLK(clk), .RST(start), .I(x[10]), .Q(
        xin[10]) );
  DFF \xreg_reg[11]  ( .D(xin[10]), .CLK(clk), .RST(start), .I(x[11]), .Q(
        xin[11]) );
  DFF \xreg_reg[12]  ( .D(xin[11]), .CLK(clk), .RST(start), .I(x[12]), .Q(
        xin[12]) );
  DFF \xreg_reg[13]  ( .D(xin[12]), .CLK(clk), .RST(start), .I(x[13]), .Q(
        xin[13]) );
  DFF \xreg_reg[14]  ( .D(xin[13]), .CLK(clk), .RST(start), .I(x[14]), .Q(
        xin[14]) );
  DFF \xreg_reg[15]  ( .D(xin[14]), .CLK(clk), .RST(start), .I(x[15]), .Q(
        xin[15]) );
  DFF \xreg_reg[16]  ( .D(xin[15]), .CLK(clk), .RST(start), .I(x[16]), .Q(
        xin[16]) );
  DFF \xreg_reg[17]  ( .D(xin[16]), .CLK(clk), .RST(start), .I(x[17]), .Q(
        xin[17]) );
  DFF \xreg_reg[18]  ( .D(xin[17]), .CLK(clk), .RST(start), .I(x[18]), .Q(
        xin[18]) );
  DFF \xreg_reg[19]  ( .D(xin[18]), .CLK(clk), .RST(start), .I(x[19]), .Q(
        xin[19]) );
  DFF \xreg_reg[20]  ( .D(xin[19]), .CLK(clk), .RST(start), .I(x[20]), .Q(
        xin[20]) );
  DFF \xreg_reg[21]  ( .D(xin[20]), .CLK(clk), .RST(start), .I(x[21]), .Q(
        xin[21]) );
  DFF \xreg_reg[22]  ( .D(xin[21]), .CLK(clk), .RST(start), .I(x[22]), .Q(
        xin[22]) );
  DFF \xreg_reg[23]  ( .D(xin[22]), .CLK(clk), .RST(start), .I(x[23]), .Q(
        xin[23]) );
  DFF \xreg_reg[24]  ( .D(xin[23]), .CLK(clk), .RST(start), .I(x[24]), .Q(
        xin[24]) );
  DFF \xreg_reg[25]  ( .D(xin[24]), .CLK(clk), .RST(start), .I(x[25]), .Q(
        xin[25]) );
  DFF \xreg_reg[26]  ( .D(xin[25]), .CLK(clk), .RST(start), .I(x[26]), .Q(
        xin[26]) );
  DFF \xreg_reg[27]  ( .D(xin[26]), .CLK(clk), .RST(start), .I(x[27]), .Q(
        xin[27]) );
  DFF \xreg_reg[28]  ( .D(xin[27]), .CLK(clk), .RST(start), .I(x[28]), .Q(
        xin[28]) );
  DFF \xreg_reg[29]  ( .D(xin[28]), .CLK(clk), .RST(start), .I(x[29]), .Q(
        xin[29]) );
  DFF \xreg_reg[30]  ( .D(xin[29]), .CLK(clk), .RST(start), .I(x[30]), .Q(
        xin[30]) );
  DFF \xreg_reg[31]  ( .D(xin[30]), .CLK(clk), .RST(start), .I(x[31]), .Q(
        xin[31]) );
  DFF \xreg_reg[32]  ( .D(xin[31]), .CLK(clk), .RST(start), .I(x[32]), .Q(
        xin[32]) );
  DFF \xreg_reg[33]  ( .D(xin[32]), .CLK(clk), .RST(start), .I(x[33]), .Q(
        xin[33]) );
  DFF \xreg_reg[34]  ( .D(xin[33]), .CLK(clk), .RST(start), .I(x[34]), .Q(
        xin[34]) );
  DFF \xreg_reg[35]  ( .D(xin[34]), .CLK(clk), .RST(start), .I(x[35]), .Q(
        xin[35]) );
  DFF \xreg_reg[36]  ( .D(xin[35]), .CLK(clk), .RST(start), .I(x[36]), .Q(
        xin[36]) );
  DFF \xreg_reg[37]  ( .D(xin[36]), .CLK(clk), .RST(start), .I(x[37]), .Q(
        xin[37]) );
  DFF \xreg_reg[38]  ( .D(xin[37]), .CLK(clk), .RST(start), .I(x[38]), .Q(
        xin[38]) );
  DFF \xreg_reg[39]  ( .D(xin[38]), .CLK(clk), .RST(start), .I(x[39]), .Q(
        xin[39]) );
  DFF \xreg_reg[40]  ( .D(xin[39]), .CLK(clk), .RST(start), .I(x[40]), .Q(
        xin[40]) );
  DFF \xreg_reg[41]  ( .D(xin[40]), .CLK(clk), .RST(start), .I(x[41]), .Q(
        xin[41]) );
  DFF \xreg_reg[42]  ( .D(xin[41]), .CLK(clk), .RST(start), .I(x[42]), .Q(
        xin[42]) );
  DFF \xreg_reg[43]  ( .D(xin[42]), .CLK(clk), .RST(start), .I(x[43]), .Q(
        xin[43]) );
  DFF \xreg_reg[44]  ( .D(xin[43]), .CLK(clk), .RST(start), .I(x[44]), .Q(
        xin[44]) );
  DFF \xreg_reg[45]  ( .D(xin[44]), .CLK(clk), .RST(start), .I(x[45]), .Q(
        xin[45]) );
  DFF \xreg_reg[46]  ( .D(xin[45]), .CLK(clk), .RST(start), .I(x[46]), .Q(
        xin[46]) );
  DFF \xreg_reg[47]  ( .D(xin[46]), .CLK(clk), .RST(start), .I(x[47]), .Q(
        xin[47]) );
  DFF \xreg_reg[48]  ( .D(xin[47]), .CLK(clk), .RST(start), .I(x[48]), .Q(
        xin[48]) );
  DFF \xreg_reg[49]  ( .D(xin[48]), .CLK(clk), .RST(start), .I(x[49]), .Q(
        xin[49]) );
  DFF \xreg_reg[50]  ( .D(xin[49]), .CLK(clk), .RST(start), .I(x[50]), .Q(
        xin[50]) );
  DFF \xreg_reg[51]  ( .D(xin[50]), .CLK(clk), .RST(start), .I(x[51]), .Q(
        xin[51]) );
  DFF \xreg_reg[52]  ( .D(xin[51]), .CLK(clk), .RST(start), .I(x[52]), .Q(
        xin[52]) );
  DFF \xreg_reg[53]  ( .D(xin[52]), .CLK(clk), .RST(start), .I(x[53]), .Q(
        xin[53]) );
  DFF \xreg_reg[54]  ( .D(xin[53]), .CLK(clk), .RST(start), .I(x[54]), .Q(
        xin[54]) );
  DFF \xreg_reg[55]  ( .D(xin[54]), .CLK(clk), .RST(start), .I(x[55]), .Q(
        xin[55]) );
  DFF \xreg_reg[56]  ( .D(xin[55]), .CLK(clk), .RST(start), .I(x[56]), .Q(
        xin[56]) );
  DFF \xreg_reg[57]  ( .D(xin[56]), .CLK(clk), .RST(start), .I(x[57]), .Q(
        xin[57]) );
  DFF \xreg_reg[58]  ( .D(xin[57]), .CLK(clk), .RST(start), .I(x[58]), .Q(
        xin[58]) );
  DFF \xreg_reg[59]  ( .D(xin[58]), .CLK(clk), .RST(start), .I(x[59]), .Q(
        xin[59]) );
  DFF \xreg_reg[60]  ( .D(xin[59]), .CLK(clk), .RST(start), .I(x[60]), .Q(
        xin[60]) );
  DFF \xreg_reg[61]  ( .D(xin[60]), .CLK(clk), .RST(start), .I(x[61]), .Q(
        xin[61]) );
  DFF \xreg_reg[62]  ( .D(xin[61]), .CLK(clk), .RST(start), .I(x[62]), .Q(
        xin[62]) );
  DFF \xreg_reg[63]  ( .D(xin[62]), .CLK(clk), .RST(start), .I(x[63]), .Q(
        xin[63]) );
  DFF \xreg_reg[64]  ( .D(xin[63]), .CLK(clk), .RST(start), .I(x[64]), .Q(
        xin[64]) );
  DFF \xreg_reg[65]  ( .D(xin[64]), .CLK(clk), .RST(start), .I(x[65]), .Q(
        xin[65]) );
  DFF \xreg_reg[66]  ( .D(xin[65]), .CLK(clk), .RST(start), .I(x[66]), .Q(
        xin[66]) );
  DFF \xreg_reg[67]  ( .D(xin[66]), .CLK(clk), .RST(start), .I(x[67]), .Q(
        xin[67]) );
  DFF \xreg_reg[68]  ( .D(xin[67]), .CLK(clk), .RST(start), .I(x[68]), .Q(
        xin[68]) );
  DFF \xreg_reg[69]  ( .D(xin[68]), .CLK(clk), .RST(start), .I(x[69]), .Q(
        xin[69]) );
  DFF \xreg_reg[70]  ( .D(xin[69]), .CLK(clk), .RST(start), .I(x[70]), .Q(
        xin[70]) );
  DFF \xreg_reg[71]  ( .D(xin[70]), .CLK(clk), .RST(start), .I(x[71]), .Q(
        xin[71]) );
  DFF \xreg_reg[72]  ( .D(xin[71]), .CLK(clk), .RST(start), .I(x[72]), .Q(
        xin[72]) );
  DFF \xreg_reg[73]  ( .D(xin[72]), .CLK(clk), .RST(start), .I(x[73]), .Q(
        xin[73]) );
  DFF \xreg_reg[74]  ( .D(xin[73]), .CLK(clk), .RST(start), .I(x[74]), .Q(
        xin[74]) );
  DFF \xreg_reg[75]  ( .D(xin[74]), .CLK(clk), .RST(start), .I(x[75]), .Q(
        xin[75]) );
  DFF \xreg_reg[76]  ( .D(xin[75]), .CLK(clk), .RST(start), .I(x[76]), .Q(
        xin[76]) );
  DFF \xreg_reg[77]  ( .D(xin[76]), .CLK(clk), .RST(start), .I(x[77]), .Q(
        xin[77]) );
  DFF \xreg_reg[78]  ( .D(xin[77]), .CLK(clk), .RST(start), .I(x[78]), .Q(
        xin[78]) );
  DFF \xreg_reg[79]  ( .D(xin[78]), .CLK(clk), .RST(start), .I(x[79]), .Q(
        xin[79]) );
  DFF \xreg_reg[80]  ( .D(xin[79]), .CLK(clk), .RST(start), .I(x[80]), .Q(
        xin[80]) );
  DFF \xreg_reg[81]  ( .D(xin[80]), .CLK(clk), .RST(start), .I(x[81]), .Q(
        xin[81]) );
  DFF \xreg_reg[82]  ( .D(xin[81]), .CLK(clk), .RST(start), .I(x[82]), .Q(
        xin[82]) );
  DFF \xreg_reg[83]  ( .D(xin[82]), .CLK(clk), .RST(start), .I(x[83]), .Q(
        xin[83]) );
  DFF \xreg_reg[84]  ( .D(xin[83]), .CLK(clk), .RST(start), .I(x[84]), .Q(
        xin[84]) );
  DFF \xreg_reg[85]  ( .D(xin[84]), .CLK(clk), .RST(start), .I(x[85]), .Q(
        xin[85]) );
  DFF \xreg_reg[86]  ( .D(xin[85]), .CLK(clk), .RST(start), .I(x[86]), .Q(
        xin[86]) );
  DFF \xreg_reg[87]  ( .D(xin[86]), .CLK(clk), .RST(start), .I(x[87]), .Q(
        xin[87]) );
  DFF \xreg_reg[88]  ( .D(xin[87]), .CLK(clk), .RST(start), .I(x[88]), .Q(
        xin[88]) );
  DFF \xreg_reg[89]  ( .D(xin[88]), .CLK(clk), .RST(start), .I(x[89]), .Q(
        xin[89]) );
  DFF \xreg_reg[90]  ( .D(xin[89]), .CLK(clk), .RST(start), .I(x[90]), .Q(
        xin[90]) );
  DFF \xreg_reg[91]  ( .D(xin[90]), .CLK(clk), .RST(start), .I(x[91]), .Q(
        xin[91]) );
  DFF \xreg_reg[92]  ( .D(xin[91]), .CLK(clk), .RST(start), .I(x[92]), .Q(
        xin[92]) );
  DFF \xreg_reg[93]  ( .D(xin[92]), .CLK(clk), .RST(start), .I(x[93]), .Q(
        xin[93]) );
  DFF \xreg_reg[94]  ( .D(xin[93]), .CLK(clk), .RST(start), .I(x[94]), .Q(
        xin[94]) );
  DFF \xreg_reg[95]  ( .D(xin[94]), .CLK(clk), .RST(start), .I(x[95]), .Q(
        xin[95]) );
  DFF \xreg_reg[96]  ( .D(xin[95]), .CLK(clk), .RST(start), .I(x[96]), .Q(
        xin[96]) );
  DFF \xreg_reg[97]  ( .D(xin[96]), .CLK(clk), .RST(start), .I(x[97]), .Q(
        xin[97]) );
  DFF \xreg_reg[98]  ( .D(xin[97]), .CLK(clk), .RST(start), .I(x[98]), .Q(
        xin[98]) );
  DFF \xreg_reg[99]  ( .D(xin[98]), .CLK(clk), .RST(start), .I(x[99]), .Q(
        xin[99]) );
  DFF \xreg_reg[100]  ( .D(xin[99]), .CLK(clk), .RST(start), .I(x[100]), .Q(
        xin[100]) );
  DFF \xreg_reg[101]  ( .D(xin[100]), .CLK(clk), .RST(start), .I(x[101]), .Q(
        xin[101]) );
  DFF \xreg_reg[102]  ( .D(xin[101]), .CLK(clk), .RST(start), .I(x[102]), .Q(
        xin[102]) );
  DFF \xreg_reg[103]  ( .D(xin[102]), .CLK(clk), .RST(start), .I(x[103]), .Q(
        xin[103]) );
  DFF \xreg_reg[104]  ( .D(xin[103]), .CLK(clk), .RST(start), .I(x[104]), .Q(
        xin[104]) );
  DFF \xreg_reg[105]  ( .D(xin[104]), .CLK(clk), .RST(start), .I(x[105]), .Q(
        xin[105]) );
  DFF \xreg_reg[106]  ( .D(xin[105]), .CLK(clk), .RST(start), .I(x[106]), .Q(
        xin[106]) );
  DFF \xreg_reg[107]  ( .D(xin[106]), .CLK(clk), .RST(start), .I(x[107]), .Q(
        xin[107]) );
  DFF \xreg_reg[108]  ( .D(xin[107]), .CLK(clk), .RST(start), .I(x[108]), .Q(
        xin[108]) );
  DFF \xreg_reg[109]  ( .D(xin[108]), .CLK(clk), .RST(start), .I(x[109]), .Q(
        xin[109]) );
  DFF \xreg_reg[110]  ( .D(xin[109]), .CLK(clk), .RST(start), .I(x[110]), .Q(
        xin[110]) );
  DFF \xreg_reg[111]  ( .D(xin[110]), .CLK(clk), .RST(start), .I(x[111]), .Q(
        xin[111]) );
  DFF \xreg_reg[112]  ( .D(xin[111]), .CLK(clk), .RST(start), .I(x[112]), .Q(
        xin[112]) );
  DFF \xreg_reg[113]  ( .D(xin[112]), .CLK(clk), .RST(start), .I(x[113]), .Q(
        xin[113]) );
  DFF \xreg_reg[114]  ( .D(xin[113]), .CLK(clk), .RST(start), .I(x[114]), .Q(
        xin[114]) );
  DFF \xreg_reg[115]  ( .D(xin[114]), .CLK(clk), .RST(start), .I(x[115]), .Q(
        xin[115]) );
  DFF \xreg_reg[116]  ( .D(xin[115]), .CLK(clk), .RST(start), .I(x[116]), .Q(
        xin[116]) );
  DFF \xreg_reg[117]  ( .D(xin[116]), .CLK(clk), .RST(start), .I(x[117]), .Q(
        xin[117]) );
  DFF \xreg_reg[118]  ( .D(xin[117]), .CLK(clk), .RST(start), .I(x[118]), .Q(
        xin[118]) );
  DFF \xreg_reg[119]  ( .D(xin[118]), .CLK(clk), .RST(start), .I(x[119]), .Q(
        xin[119]) );
  DFF \xreg_reg[120]  ( .D(xin[119]), .CLK(clk), .RST(start), .I(x[120]), .Q(
        xin[120]) );
  DFF \xreg_reg[121]  ( .D(xin[120]), .CLK(clk), .RST(start), .I(x[121]), .Q(
        xin[121]) );
  DFF \xreg_reg[122]  ( .D(xin[121]), .CLK(clk), .RST(start), .I(x[122]), .Q(
        xin[122]) );
  DFF \xreg_reg[123]  ( .D(xin[122]), .CLK(clk), .RST(start), .I(x[123]), .Q(
        xin[123]) );
  DFF \xreg_reg[124]  ( .D(xin[123]), .CLK(clk), .RST(start), .I(x[124]), .Q(
        xin[124]) );
  DFF \xreg_reg[125]  ( .D(xin[124]), .CLK(clk), .RST(start), .I(x[125]), .Q(
        xin[125]) );
  DFF \xreg_reg[126]  ( .D(xin[125]), .CLK(clk), .RST(start), .I(x[126]), .Q(
        xin[126]) );
  DFF \xreg_reg[127]  ( .D(xin[126]), .CLK(clk), .RST(start), .I(x[127]), .Q(
        xin[127]) );
  DFF \xreg_reg[128]  ( .D(xin[127]), .CLK(clk), .RST(start), .I(x[128]), .Q(
        xin[128]) );
  DFF \xreg_reg[129]  ( .D(xin[128]), .CLK(clk), .RST(start), .I(x[129]), .Q(
        xin[129]) );
  DFF \xreg_reg[130]  ( .D(xin[129]), .CLK(clk), .RST(start), .I(x[130]), .Q(
        xin[130]) );
  DFF \xreg_reg[131]  ( .D(xin[130]), .CLK(clk), .RST(start), .I(x[131]), .Q(
        xin[131]) );
  DFF \xreg_reg[132]  ( .D(xin[131]), .CLK(clk), .RST(start), .I(x[132]), .Q(
        xin[132]) );
  DFF \xreg_reg[133]  ( .D(xin[132]), .CLK(clk), .RST(start), .I(x[133]), .Q(
        xin[133]) );
  DFF \xreg_reg[134]  ( .D(xin[133]), .CLK(clk), .RST(start), .I(x[134]), .Q(
        xin[134]) );
  DFF \xreg_reg[135]  ( .D(xin[134]), .CLK(clk), .RST(start), .I(x[135]), .Q(
        xin[135]) );
  DFF \xreg_reg[136]  ( .D(xin[135]), .CLK(clk), .RST(start), .I(x[136]), .Q(
        xin[136]) );
  DFF \xreg_reg[137]  ( .D(xin[136]), .CLK(clk), .RST(start), .I(x[137]), .Q(
        xin[137]) );
  DFF \xreg_reg[138]  ( .D(xin[137]), .CLK(clk), .RST(start), .I(x[138]), .Q(
        xin[138]) );
  DFF \xreg_reg[139]  ( .D(xin[138]), .CLK(clk), .RST(start), .I(x[139]), .Q(
        xin[139]) );
  DFF \xreg_reg[140]  ( .D(xin[139]), .CLK(clk), .RST(start), .I(x[140]), .Q(
        xin[140]) );
  DFF \xreg_reg[141]  ( .D(xin[140]), .CLK(clk), .RST(start), .I(x[141]), .Q(
        xin[141]) );
  DFF \xreg_reg[142]  ( .D(xin[141]), .CLK(clk), .RST(start), .I(x[142]), .Q(
        xin[142]) );
  DFF \xreg_reg[143]  ( .D(xin[142]), .CLK(clk), .RST(start), .I(x[143]), .Q(
        xin[143]) );
  DFF \xreg_reg[144]  ( .D(xin[143]), .CLK(clk), .RST(start), .I(x[144]), .Q(
        xin[144]) );
  DFF \xreg_reg[145]  ( .D(xin[144]), .CLK(clk), .RST(start), .I(x[145]), .Q(
        xin[145]) );
  DFF \xreg_reg[146]  ( .D(xin[145]), .CLK(clk), .RST(start), .I(x[146]), .Q(
        xin[146]) );
  DFF \xreg_reg[147]  ( .D(xin[146]), .CLK(clk), .RST(start), .I(x[147]), .Q(
        xin[147]) );
  DFF \xreg_reg[148]  ( .D(xin[147]), .CLK(clk), .RST(start), .I(x[148]), .Q(
        xin[148]) );
  DFF \xreg_reg[149]  ( .D(xin[148]), .CLK(clk), .RST(start), .I(x[149]), .Q(
        xin[149]) );
  DFF \xreg_reg[150]  ( .D(xin[149]), .CLK(clk), .RST(start), .I(x[150]), .Q(
        xin[150]) );
  DFF \xreg_reg[151]  ( .D(xin[150]), .CLK(clk), .RST(start), .I(x[151]), .Q(
        xin[151]) );
  DFF \xreg_reg[152]  ( .D(xin[151]), .CLK(clk), .RST(start), .I(x[152]), .Q(
        xin[152]) );
  DFF \xreg_reg[153]  ( .D(xin[152]), .CLK(clk), .RST(start), .I(x[153]), .Q(
        xin[153]) );
  DFF \xreg_reg[154]  ( .D(xin[153]), .CLK(clk), .RST(start), .I(x[154]), .Q(
        xin[154]) );
  DFF \xreg_reg[155]  ( .D(xin[154]), .CLK(clk), .RST(start), .I(x[155]), .Q(
        xin[155]) );
  DFF \xreg_reg[156]  ( .D(xin[155]), .CLK(clk), .RST(start), .I(x[156]), .Q(
        xin[156]) );
  DFF \xreg_reg[157]  ( .D(xin[156]), .CLK(clk), .RST(start), .I(x[157]), .Q(
        xin[157]) );
  DFF \xreg_reg[158]  ( .D(xin[157]), .CLK(clk), .RST(start), .I(x[158]), .Q(
        xin[158]) );
  DFF \xreg_reg[159]  ( .D(xin[158]), .CLK(clk), .RST(start), .I(x[159]), .Q(
        xin[159]) );
  DFF \xreg_reg[160]  ( .D(xin[159]), .CLK(clk), .RST(start), .I(x[160]), .Q(
        xin[160]) );
  DFF \xreg_reg[161]  ( .D(xin[160]), .CLK(clk), .RST(start), .I(x[161]), .Q(
        xin[161]) );
  DFF \xreg_reg[162]  ( .D(xin[161]), .CLK(clk), .RST(start), .I(x[162]), .Q(
        xin[162]) );
  DFF \xreg_reg[163]  ( .D(xin[162]), .CLK(clk), .RST(start), .I(x[163]), .Q(
        xin[163]) );
  DFF \xreg_reg[164]  ( .D(xin[163]), .CLK(clk), .RST(start), .I(x[164]), .Q(
        xin[164]) );
  DFF \xreg_reg[165]  ( .D(xin[164]), .CLK(clk), .RST(start), .I(x[165]), .Q(
        xin[165]) );
  DFF \xreg_reg[166]  ( .D(xin[165]), .CLK(clk), .RST(start), .I(x[166]), .Q(
        xin[166]) );
  DFF \xreg_reg[167]  ( .D(xin[166]), .CLK(clk), .RST(start), .I(x[167]), .Q(
        xin[167]) );
  DFF \xreg_reg[168]  ( .D(xin[167]), .CLK(clk), .RST(start), .I(x[168]), .Q(
        xin[168]) );
  DFF \xreg_reg[169]  ( .D(xin[168]), .CLK(clk), .RST(start), .I(x[169]), .Q(
        xin[169]) );
  DFF \xreg_reg[170]  ( .D(xin[169]), .CLK(clk), .RST(start), .I(x[170]), .Q(
        xin[170]) );
  DFF \xreg_reg[171]  ( .D(xin[170]), .CLK(clk), .RST(start), .I(x[171]), .Q(
        xin[171]) );
  DFF \xreg_reg[172]  ( .D(xin[171]), .CLK(clk), .RST(start), .I(x[172]), .Q(
        xin[172]) );
  DFF \xreg_reg[173]  ( .D(xin[172]), .CLK(clk), .RST(start), .I(x[173]), .Q(
        xin[173]) );
  DFF \xreg_reg[174]  ( .D(xin[173]), .CLK(clk), .RST(start), .I(x[174]), .Q(
        xin[174]) );
  DFF \xreg_reg[175]  ( .D(xin[174]), .CLK(clk), .RST(start), .I(x[175]), .Q(
        xin[175]) );
  DFF \xreg_reg[176]  ( .D(xin[175]), .CLK(clk), .RST(start), .I(x[176]), .Q(
        xin[176]) );
  DFF \xreg_reg[177]  ( .D(xin[176]), .CLK(clk), .RST(start), .I(x[177]), .Q(
        xin[177]) );
  DFF \xreg_reg[178]  ( .D(xin[177]), .CLK(clk), .RST(start), .I(x[178]), .Q(
        xin[178]) );
  DFF \xreg_reg[179]  ( .D(xin[178]), .CLK(clk), .RST(start), .I(x[179]), .Q(
        xin[179]) );
  DFF \xreg_reg[180]  ( .D(xin[179]), .CLK(clk), .RST(start), .I(x[180]), .Q(
        xin[180]) );
  DFF \xreg_reg[181]  ( .D(xin[180]), .CLK(clk), .RST(start), .I(x[181]), .Q(
        xin[181]) );
  DFF \xreg_reg[182]  ( .D(xin[181]), .CLK(clk), .RST(start), .I(x[182]), .Q(
        xin[182]) );
  DFF \xreg_reg[183]  ( .D(xin[182]), .CLK(clk), .RST(start), .I(x[183]), .Q(
        xin[183]) );
  DFF \xreg_reg[184]  ( .D(xin[183]), .CLK(clk), .RST(start), .I(x[184]), .Q(
        xin[184]) );
  DFF \xreg_reg[185]  ( .D(xin[184]), .CLK(clk), .RST(start), .I(x[185]), .Q(
        xin[185]) );
  DFF \xreg_reg[186]  ( .D(xin[185]), .CLK(clk), .RST(start), .I(x[186]), .Q(
        xin[186]) );
  DFF \xreg_reg[187]  ( .D(xin[186]), .CLK(clk), .RST(start), .I(x[187]), .Q(
        xin[187]) );
  DFF \xreg_reg[188]  ( .D(xin[187]), .CLK(clk), .RST(start), .I(x[188]), .Q(
        xin[188]) );
  DFF \xreg_reg[189]  ( .D(xin[188]), .CLK(clk), .RST(start), .I(x[189]), .Q(
        xin[189]) );
  DFF \xreg_reg[190]  ( .D(xin[189]), .CLK(clk), .RST(start), .I(x[190]), .Q(
        xin[190]) );
  DFF \xreg_reg[191]  ( .D(xin[190]), .CLK(clk), .RST(start), .I(x[191]), .Q(
        xin[191]) );
  DFF \xreg_reg[192]  ( .D(xin[191]), .CLK(clk), .RST(start), .I(x[192]), .Q(
        xin[192]) );
  DFF \xreg_reg[193]  ( .D(xin[192]), .CLK(clk), .RST(start), .I(x[193]), .Q(
        xin[193]) );
  DFF \xreg_reg[194]  ( .D(xin[193]), .CLK(clk), .RST(start), .I(x[194]), .Q(
        xin[194]) );
  DFF \xreg_reg[195]  ( .D(xin[194]), .CLK(clk), .RST(start), .I(x[195]), .Q(
        xin[195]) );
  DFF \xreg_reg[196]  ( .D(xin[195]), .CLK(clk), .RST(start), .I(x[196]), .Q(
        xin[196]) );
  DFF \xreg_reg[197]  ( .D(xin[196]), .CLK(clk), .RST(start), .I(x[197]), .Q(
        xin[197]) );
  DFF \xreg_reg[198]  ( .D(xin[197]), .CLK(clk), .RST(start), .I(x[198]), .Q(
        xin[198]) );
  DFF \xreg_reg[199]  ( .D(xin[198]), .CLK(clk), .RST(start), .I(x[199]), .Q(
        xin[199]) );
  DFF \xreg_reg[200]  ( .D(xin[199]), .CLK(clk), .RST(start), .I(x[200]), .Q(
        xin[200]) );
  DFF \xreg_reg[201]  ( .D(xin[200]), .CLK(clk), .RST(start), .I(x[201]), .Q(
        xin[201]) );
  DFF \xreg_reg[202]  ( .D(xin[201]), .CLK(clk), .RST(start), .I(x[202]), .Q(
        xin[202]) );
  DFF \xreg_reg[203]  ( .D(xin[202]), .CLK(clk), .RST(start), .I(x[203]), .Q(
        xin[203]) );
  DFF \xreg_reg[204]  ( .D(xin[203]), .CLK(clk), .RST(start), .I(x[204]), .Q(
        xin[204]) );
  DFF \xreg_reg[205]  ( .D(xin[204]), .CLK(clk), .RST(start), .I(x[205]), .Q(
        xin[205]) );
  DFF \xreg_reg[206]  ( .D(xin[205]), .CLK(clk), .RST(start), .I(x[206]), .Q(
        xin[206]) );
  DFF \xreg_reg[207]  ( .D(xin[206]), .CLK(clk), .RST(start), .I(x[207]), .Q(
        xin[207]) );
  DFF \xreg_reg[208]  ( .D(xin[207]), .CLK(clk), .RST(start), .I(x[208]), .Q(
        xin[208]) );
  DFF \xreg_reg[209]  ( .D(xin[208]), .CLK(clk), .RST(start), .I(x[209]), .Q(
        xin[209]) );
  DFF \xreg_reg[210]  ( .D(xin[209]), .CLK(clk), .RST(start), .I(x[210]), .Q(
        xin[210]) );
  DFF \xreg_reg[211]  ( .D(xin[210]), .CLK(clk), .RST(start), .I(x[211]), .Q(
        xin[211]) );
  DFF \xreg_reg[212]  ( .D(xin[211]), .CLK(clk), .RST(start), .I(x[212]), .Q(
        xin[212]) );
  DFF \xreg_reg[213]  ( .D(xin[212]), .CLK(clk), .RST(start), .I(x[213]), .Q(
        xin[213]) );
  DFF \xreg_reg[214]  ( .D(xin[213]), .CLK(clk), .RST(start), .I(x[214]), .Q(
        xin[214]) );
  DFF \xreg_reg[215]  ( .D(xin[214]), .CLK(clk), .RST(start), .I(x[215]), .Q(
        xin[215]) );
  DFF \xreg_reg[216]  ( .D(xin[215]), .CLK(clk), .RST(start), .I(x[216]), .Q(
        xin[216]) );
  DFF \xreg_reg[217]  ( .D(xin[216]), .CLK(clk), .RST(start), .I(x[217]), .Q(
        xin[217]) );
  DFF \xreg_reg[218]  ( .D(xin[217]), .CLK(clk), .RST(start), .I(x[218]), .Q(
        xin[218]) );
  DFF \xreg_reg[219]  ( .D(xin[218]), .CLK(clk), .RST(start), .I(x[219]), .Q(
        xin[219]) );
  DFF \xreg_reg[220]  ( .D(xin[219]), .CLK(clk), .RST(start), .I(x[220]), .Q(
        xin[220]) );
  DFF \xreg_reg[221]  ( .D(xin[220]), .CLK(clk), .RST(start), .I(x[221]), .Q(
        xin[221]) );
  DFF \xreg_reg[222]  ( .D(xin[221]), .CLK(clk), .RST(start), .I(x[222]), .Q(
        xin[222]) );
  DFF \xreg_reg[223]  ( .D(xin[222]), .CLK(clk), .RST(start), .I(x[223]), .Q(
        xin[223]) );
  DFF \xreg_reg[224]  ( .D(xin[223]), .CLK(clk), .RST(start), .I(x[224]), .Q(
        xin[224]) );
  DFF \xreg_reg[225]  ( .D(xin[224]), .CLK(clk), .RST(start), .I(x[225]), .Q(
        xin[225]) );
  DFF \xreg_reg[226]  ( .D(xin[225]), .CLK(clk), .RST(start), .I(x[226]), .Q(
        xin[226]) );
  DFF \xreg_reg[227]  ( .D(xin[226]), .CLK(clk), .RST(start), .I(x[227]), .Q(
        xin[227]) );
  DFF \xreg_reg[228]  ( .D(xin[227]), .CLK(clk), .RST(start), .I(x[228]), .Q(
        xin[228]) );
  DFF \xreg_reg[229]  ( .D(xin[228]), .CLK(clk), .RST(start), .I(x[229]), .Q(
        xin[229]) );
  DFF \xreg_reg[230]  ( .D(xin[229]), .CLK(clk), .RST(start), .I(x[230]), .Q(
        xin[230]) );
  DFF \xreg_reg[231]  ( .D(xin[230]), .CLK(clk), .RST(start), .I(x[231]), .Q(
        xin[231]) );
  DFF \xreg_reg[232]  ( .D(xin[231]), .CLK(clk), .RST(start), .I(x[232]), .Q(
        xin[232]) );
  DFF \xreg_reg[233]  ( .D(xin[232]), .CLK(clk), .RST(start), .I(x[233]), .Q(
        xin[233]) );
  DFF \xreg_reg[234]  ( .D(xin[233]), .CLK(clk), .RST(start), .I(x[234]), .Q(
        xin[234]) );
  DFF \xreg_reg[235]  ( .D(xin[234]), .CLK(clk), .RST(start), .I(x[235]), .Q(
        xin[235]) );
  DFF \xreg_reg[236]  ( .D(xin[235]), .CLK(clk), .RST(start), .I(x[236]), .Q(
        xin[236]) );
  DFF \xreg_reg[237]  ( .D(xin[236]), .CLK(clk), .RST(start), .I(x[237]), .Q(
        xin[237]) );
  DFF \xreg_reg[238]  ( .D(xin[237]), .CLK(clk), .RST(start), .I(x[238]), .Q(
        xin[238]) );
  DFF \xreg_reg[239]  ( .D(xin[238]), .CLK(clk), .RST(start), .I(x[239]), .Q(
        xin[239]) );
  DFF \xreg_reg[240]  ( .D(xin[239]), .CLK(clk), .RST(start), .I(x[240]), .Q(
        xin[240]) );
  DFF \xreg_reg[241]  ( .D(xin[240]), .CLK(clk), .RST(start), .I(x[241]), .Q(
        xin[241]) );
  DFF \xreg_reg[242]  ( .D(xin[241]), .CLK(clk), .RST(start), .I(x[242]), .Q(
        xin[242]) );
  DFF \xreg_reg[243]  ( .D(xin[242]), .CLK(clk), .RST(start), .I(x[243]), .Q(
        xin[243]) );
  DFF \xreg_reg[244]  ( .D(xin[243]), .CLK(clk), .RST(start), .I(x[244]), .Q(
        xin[244]) );
  DFF \xreg_reg[245]  ( .D(xin[244]), .CLK(clk), .RST(start), .I(x[245]), .Q(
        xin[245]) );
  DFF \xreg_reg[246]  ( .D(xin[245]), .CLK(clk), .RST(start), .I(x[246]), .Q(
        xin[246]) );
  DFF \xreg_reg[247]  ( .D(xin[246]), .CLK(clk), .RST(start), .I(x[247]), .Q(
        xin[247]) );
  DFF \xreg_reg[248]  ( .D(xin[247]), .CLK(clk), .RST(start), .I(x[248]), .Q(
        xin[248]) );
  DFF \xreg_reg[249]  ( .D(xin[248]), .CLK(clk), .RST(start), .I(x[249]), .Q(
        xin[249]) );
  DFF \xreg_reg[250]  ( .D(xin[249]), .CLK(clk), .RST(start), .I(x[250]), .Q(
        xin[250]) );
  DFF \xreg_reg[251]  ( .D(xin[250]), .CLK(clk), .RST(start), .I(x[251]), .Q(
        xin[251]) );
  DFF \xreg_reg[252]  ( .D(xin[251]), .CLK(clk), .RST(start), .I(x[252]), .Q(
        xin[252]) );
  DFF \xreg_reg[253]  ( .D(xin[252]), .CLK(clk), .RST(start), .I(x[253]), .Q(
        xin[253]) );
  DFF \xreg_reg[254]  ( .D(xin[253]), .CLK(clk), .RST(start), .I(x[254]), .Q(
        xin[254]) );
  DFF \xreg_reg[255]  ( .D(xin[254]), .CLK(clk), .RST(start), .I(x[255]), .Q(
        xin[255]) );
  DFF \xreg_reg[256]  ( .D(xin[255]), .CLK(clk), .RST(start), .I(x[256]), .Q(
        xin[256]) );
  DFF \xreg_reg[257]  ( .D(xin[256]), .CLK(clk), .RST(start), .I(x[257]), .Q(
        xin[257]) );
  DFF \xreg_reg[258]  ( .D(xin[257]), .CLK(clk), .RST(start), .I(x[258]), .Q(
        xin[258]) );
  DFF \xreg_reg[259]  ( .D(xin[258]), .CLK(clk), .RST(start), .I(x[259]), .Q(
        xin[259]) );
  DFF \xreg_reg[260]  ( .D(xin[259]), .CLK(clk), .RST(start), .I(x[260]), .Q(
        xin[260]) );
  DFF \xreg_reg[261]  ( .D(xin[260]), .CLK(clk), .RST(start), .I(x[261]), .Q(
        xin[261]) );
  DFF \xreg_reg[262]  ( .D(xin[261]), .CLK(clk), .RST(start), .I(x[262]), .Q(
        xin[262]) );
  DFF \xreg_reg[263]  ( .D(xin[262]), .CLK(clk), .RST(start), .I(x[263]), .Q(
        xin[263]) );
  DFF \xreg_reg[264]  ( .D(xin[263]), .CLK(clk), .RST(start), .I(x[264]), .Q(
        xin[264]) );
  DFF \xreg_reg[265]  ( .D(xin[264]), .CLK(clk), .RST(start), .I(x[265]), .Q(
        xin[265]) );
  DFF \xreg_reg[266]  ( .D(xin[265]), .CLK(clk), .RST(start), .I(x[266]), .Q(
        xin[266]) );
  DFF \xreg_reg[267]  ( .D(xin[266]), .CLK(clk), .RST(start), .I(x[267]), .Q(
        xin[267]) );
  DFF \xreg_reg[268]  ( .D(xin[267]), .CLK(clk), .RST(start), .I(x[268]), .Q(
        xin[268]) );
  DFF \xreg_reg[269]  ( .D(xin[268]), .CLK(clk), .RST(start), .I(x[269]), .Q(
        xin[269]) );
  DFF \xreg_reg[270]  ( .D(xin[269]), .CLK(clk), .RST(start), .I(x[270]), .Q(
        xin[270]) );
  DFF \xreg_reg[271]  ( .D(xin[270]), .CLK(clk), .RST(start), .I(x[271]), .Q(
        xin[271]) );
  DFF \xreg_reg[272]  ( .D(xin[271]), .CLK(clk), .RST(start), .I(x[272]), .Q(
        xin[272]) );
  DFF \xreg_reg[273]  ( .D(xin[272]), .CLK(clk), .RST(start), .I(x[273]), .Q(
        xin[273]) );
  DFF \xreg_reg[274]  ( .D(xin[273]), .CLK(clk), .RST(start), .I(x[274]), .Q(
        xin[274]) );
  DFF \xreg_reg[275]  ( .D(xin[274]), .CLK(clk), .RST(start), .I(x[275]), .Q(
        xin[275]) );
  DFF \xreg_reg[276]  ( .D(xin[275]), .CLK(clk), .RST(start), .I(x[276]), .Q(
        xin[276]) );
  DFF \xreg_reg[277]  ( .D(xin[276]), .CLK(clk), .RST(start), .I(x[277]), .Q(
        xin[277]) );
  DFF \xreg_reg[278]  ( .D(xin[277]), .CLK(clk), .RST(start), .I(x[278]), .Q(
        xin[278]) );
  DFF \xreg_reg[279]  ( .D(xin[278]), .CLK(clk), .RST(start), .I(x[279]), .Q(
        xin[279]) );
  DFF \xreg_reg[280]  ( .D(xin[279]), .CLK(clk), .RST(start), .I(x[280]), .Q(
        xin[280]) );
  DFF \xreg_reg[281]  ( .D(xin[280]), .CLK(clk), .RST(start), .I(x[281]), .Q(
        xin[281]) );
  DFF \xreg_reg[282]  ( .D(xin[281]), .CLK(clk), .RST(start), .I(x[282]), .Q(
        xin[282]) );
  DFF \xreg_reg[283]  ( .D(xin[282]), .CLK(clk), .RST(start), .I(x[283]), .Q(
        xin[283]) );
  DFF \xreg_reg[284]  ( .D(xin[283]), .CLK(clk), .RST(start), .I(x[284]), .Q(
        xin[284]) );
  DFF \xreg_reg[285]  ( .D(xin[284]), .CLK(clk), .RST(start), .I(x[285]), .Q(
        xin[285]) );
  DFF \xreg_reg[286]  ( .D(xin[285]), .CLK(clk), .RST(start), .I(x[286]), .Q(
        xin[286]) );
  DFF \xreg_reg[287]  ( .D(xin[286]), .CLK(clk), .RST(start), .I(x[287]), .Q(
        xin[287]) );
  DFF \xreg_reg[288]  ( .D(xin[287]), .CLK(clk), .RST(start), .I(x[288]), .Q(
        xin[288]) );
  DFF \xreg_reg[289]  ( .D(xin[288]), .CLK(clk), .RST(start), .I(x[289]), .Q(
        xin[289]) );
  DFF \xreg_reg[290]  ( .D(xin[289]), .CLK(clk), .RST(start), .I(x[290]), .Q(
        xin[290]) );
  DFF \xreg_reg[291]  ( .D(xin[290]), .CLK(clk), .RST(start), .I(x[291]), .Q(
        xin[291]) );
  DFF \xreg_reg[292]  ( .D(xin[291]), .CLK(clk), .RST(start), .I(x[292]), .Q(
        xin[292]) );
  DFF \xreg_reg[293]  ( .D(xin[292]), .CLK(clk), .RST(start), .I(x[293]), .Q(
        xin[293]) );
  DFF \xreg_reg[294]  ( .D(xin[293]), .CLK(clk), .RST(start), .I(x[294]), .Q(
        xin[294]) );
  DFF \xreg_reg[295]  ( .D(xin[294]), .CLK(clk), .RST(start), .I(x[295]), .Q(
        xin[295]) );
  DFF \xreg_reg[296]  ( .D(xin[295]), .CLK(clk), .RST(start), .I(x[296]), .Q(
        xin[296]) );
  DFF \xreg_reg[297]  ( .D(xin[296]), .CLK(clk), .RST(start), .I(x[297]), .Q(
        xin[297]) );
  DFF \xreg_reg[298]  ( .D(xin[297]), .CLK(clk), .RST(start), .I(x[298]), .Q(
        xin[298]) );
  DFF \xreg_reg[299]  ( .D(xin[298]), .CLK(clk), .RST(start), .I(x[299]), .Q(
        xin[299]) );
  DFF \xreg_reg[300]  ( .D(xin[299]), .CLK(clk), .RST(start), .I(x[300]), .Q(
        xin[300]) );
  DFF \xreg_reg[301]  ( .D(xin[300]), .CLK(clk), .RST(start), .I(x[301]), .Q(
        xin[301]) );
  DFF \xreg_reg[302]  ( .D(xin[301]), .CLK(clk), .RST(start), .I(x[302]), .Q(
        xin[302]) );
  DFF \xreg_reg[303]  ( .D(xin[302]), .CLK(clk), .RST(start), .I(x[303]), .Q(
        xin[303]) );
  DFF \xreg_reg[304]  ( .D(xin[303]), .CLK(clk), .RST(start), .I(x[304]), .Q(
        xin[304]) );
  DFF \xreg_reg[305]  ( .D(xin[304]), .CLK(clk), .RST(start), .I(x[305]), .Q(
        xin[305]) );
  DFF \xreg_reg[306]  ( .D(xin[305]), .CLK(clk), .RST(start), .I(x[306]), .Q(
        xin[306]) );
  DFF \xreg_reg[307]  ( .D(xin[306]), .CLK(clk), .RST(start), .I(x[307]), .Q(
        xin[307]) );
  DFF \xreg_reg[308]  ( .D(xin[307]), .CLK(clk), .RST(start), .I(x[308]), .Q(
        xin[308]) );
  DFF \xreg_reg[309]  ( .D(xin[308]), .CLK(clk), .RST(start), .I(x[309]), .Q(
        xin[309]) );
  DFF \xreg_reg[310]  ( .D(xin[309]), .CLK(clk), .RST(start), .I(x[310]), .Q(
        xin[310]) );
  DFF \xreg_reg[311]  ( .D(xin[310]), .CLK(clk), .RST(start), .I(x[311]), .Q(
        xin[311]) );
  DFF \xreg_reg[312]  ( .D(xin[311]), .CLK(clk), .RST(start), .I(x[312]), .Q(
        xin[312]) );
  DFF \xreg_reg[313]  ( .D(xin[312]), .CLK(clk), .RST(start), .I(x[313]), .Q(
        xin[313]) );
  DFF \xreg_reg[314]  ( .D(xin[313]), .CLK(clk), .RST(start), .I(x[314]), .Q(
        xin[314]) );
  DFF \xreg_reg[315]  ( .D(xin[314]), .CLK(clk), .RST(start), .I(x[315]), .Q(
        xin[315]) );
  DFF \xreg_reg[316]  ( .D(xin[315]), .CLK(clk), .RST(start), .I(x[316]), .Q(
        xin[316]) );
  DFF \xreg_reg[317]  ( .D(xin[316]), .CLK(clk), .RST(start), .I(x[317]), .Q(
        xin[317]) );
  DFF \xreg_reg[318]  ( .D(xin[317]), .CLK(clk), .RST(start), .I(x[318]), .Q(
        xin[318]) );
  DFF \xreg_reg[319]  ( .D(xin[318]), .CLK(clk), .RST(start), .I(x[319]), .Q(
        xin[319]) );
  DFF \xreg_reg[320]  ( .D(xin[319]), .CLK(clk), .RST(start), .I(x[320]), .Q(
        xin[320]) );
  DFF \xreg_reg[321]  ( .D(xin[320]), .CLK(clk), .RST(start), .I(x[321]), .Q(
        xin[321]) );
  DFF \xreg_reg[322]  ( .D(xin[321]), .CLK(clk), .RST(start), .I(x[322]), .Q(
        xin[322]) );
  DFF \xreg_reg[323]  ( .D(xin[322]), .CLK(clk), .RST(start), .I(x[323]), .Q(
        xin[323]) );
  DFF \xreg_reg[324]  ( .D(xin[323]), .CLK(clk), .RST(start), .I(x[324]), .Q(
        xin[324]) );
  DFF \xreg_reg[325]  ( .D(xin[324]), .CLK(clk), .RST(start), .I(x[325]), .Q(
        xin[325]) );
  DFF \xreg_reg[326]  ( .D(xin[325]), .CLK(clk), .RST(start), .I(x[326]), .Q(
        xin[326]) );
  DFF \xreg_reg[327]  ( .D(xin[326]), .CLK(clk), .RST(start), .I(x[327]), .Q(
        xin[327]) );
  DFF \xreg_reg[328]  ( .D(xin[327]), .CLK(clk), .RST(start), .I(x[328]), .Q(
        xin[328]) );
  DFF \xreg_reg[329]  ( .D(xin[328]), .CLK(clk), .RST(start), .I(x[329]), .Q(
        xin[329]) );
  DFF \xreg_reg[330]  ( .D(xin[329]), .CLK(clk), .RST(start), .I(x[330]), .Q(
        xin[330]) );
  DFF \xreg_reg[331]  ( .D(xin[330]), .CLK(clk), .RST(start), .I(x[331]), .Q(
        xin[331]) );
  DFF \xreg_reg[332]  ( .D(xin[331]), .CLK(clk), .RST(start), .I(x[332]), .Q(
        xin[332]) );
  DFF \xreg_reg[333]  ( .D(xin[332]), .CLK(clk), .RST(start), .I(x[333]), .Q(
        xin[333]) );
  DFF \xreg_reg[334]  ( .D(xin[333]), .CLK(clk), .RST(start), .I(x[334]), .Q(
        xin[334]) );
  DFF \xreg_reg[335]  ( .D(xin[334]), .CLK(clk), .RST(start), .I(x[335]), .Q(
        xin[335]) );
  DFF \xreg_reg[336]  ( .D(xin[335]), .CLK(clk), .RST(start), .I(x[336]), .Q(
        xin[336]) );
  DFF \xreg_reg[337]  ( .D(xin[336]), .CLK(clk), .RST(start), .I(x[337]), .Q(
        xin[337]) );
  DFF \xreg_reg[338]  ( .D(xin[337]), .CLK(clk), .RST(start), .I(x[338]), .Q(
        xin[338]) );
  DFF \xreg_reg[339]  ( .D(xin[338]), .CLK(clk), .RST(start), .I(x[339]), .Q(
        xin[339]) );
  DFF \xreg_reg[340]  ( .D(xin[339]), .CLK(clk), .RST(start), .I(x[340]), .Q(
        xin[340]) );
  DFF \xreg_reg[341]  ( .D(xin[340]), .CLK(clk), .RST(start), .I(x[341]), .Q(
        xin[341]) );
  DFF \xreg_reg[342]  ( .D(xin[341]), .CLK(clk), .RST(start), .I(x[342]), .Q(
        xin[342]) );
  DFF \xreg_reg[343]  ( .D(xin[342]), .CLK(clk), .RST(start), .I(x[343]), .Q(
        xin[343]) );
  DFF \xreg_reg[344]  ( .D(xin[343]), .CLK(clk), .RST(start), .I(x[344]), .Q(
        xin[344]) );
  DFF \xreg_reg[345]  ( .D(xin[344]), .CLK(clk), .RST(start), .I(x[345]), .Q(
        xin[345]) );
  DFF \xreg_reg[346]  ( .D(xin[345]), .CLK(clk), .RST(start), .I(x[346]), .Q(
        xin[346]) );
  DFF \xreg_reg[347]  ( .D(xin[346]), .CLK(clk), .RST(start), .I(x[347]), .Q(
        xin[347]) );
  DFF \xreg_reg[348]  ( .D(xin[347]), .CLK(clk), .RST(start), .I(x[348]), .Q(
        xin[348]) );
  DFF \xreg_reg[349]  ( .D(xin[348]), .CLK(clk), .RST(start), .I(x[349]), .Q(
        xin[349]) );
  DFF \xreg_reg[350]  ( .D(xin[349]), .CLK(clk), .RST(start), .I(x[350]), .Q(
        xin[350]) );
  DFF \xreg_reg[351]  ( .D(xin[350]), .CLK(clk), .RST(start), .I(x[351]), .Q(
        xin[351]) );
  DFF \xreg_reg[352]  ( .D(xin[351]), .CLK(clk), .RST(start), .I(x[352]), .Q(
        xin[352]) );
  DFF \xreg_reg[353]  ( .D(xin[352]), .CLK(clk), .RST(start), .I(x[353]), .Q(
        xin[353]) );
  DFF \xreg_reg[354]  ( .D(xin[353]), .CLK(clk), .RST(start), .I(x[354]), .Q(
        xin[354]) );
  DFF \xreg_reg[355]  ( .D(xin[354]), .CLK(clk), .RST(start), .I(x[355]), .Q(
        xin[355]) );
  DFF \xreg_reg[356]  ( .D(xin[355]), .CLK(clk), .RST(start), .I(x[356]), .Q(
        xin[356]) );
  DFF \xreg_reg[357]  ( .D(xin[356]), .CLK(clk), .RST(start), .I(x[357]), .Q(
        xin[357]) );
  DFF \xreg_reg[358]  ( .D(xin[357]), .CLK(clk), .RST(start), .I(x[358]), .Q(
        xin[358]) );
  DFF \xreg_reg[359]  ( .D(xin[358]), .CLK(clk), .RST(start), .I(x[359]), .Q(
        xin[359]) );
  DFF \xreg_reg[360]  ( .D(xin[359]), .CLK(clk), .RST(start), .I(x[360]), .Q(
        xin[360]) );
  DFF \xreg_reg[361]  ( .D(xin[360]), .CLK(clk), .RST(start), .I(x[361]), .Q(
        xin[361]) );
  DFF \xreg_reg[362]  ( .D(xin[361]), .CLK(clk), .RST(start), .I(x[362]), .Q(
        xin[362]) );
  DFF \xreg_reg[363]  ( .D(xin[362]), .CLK(clk), .RST(start), .I(x[363]), .Q(
        xin[363]) );
  DFF \xreg_reg[364]  ( .D(xin[363]), .CLK(clk), .RST(start), .I(x[364]), .Q(
        xin[364]) );
  DFF \xreg_reg[365]  ( .D(xin[364]), .CLK(clk), .RST(start), .I(x[365]), .Q(
        xin[365]) );
  DFF \xreg_reg[366]  ( .D(xin[365]), .CLK(clk), .RST(start), .I(x[366]), .Q(
        xin[366]) );
  DFF \xreg_reg[367]  ( .D(xin[366]), .CLK(clk), .RST(start), .I(x[367]), .Q(
        xin[367]) );
  DFF \xreg_reg[368]  ( .D(xin[367]), .CLK(clk), .RST(start), .I(x[368]), .Q(
        xin[368]) );
  DFF \xreg_reg[369]  ( .D(xin[368]), .CLK(clk), .RST(start), .I(x[369]), .Q(
        xin[369]) );
  DFF \xreg_reg[370]  ( .D(xin[369]), .CLK(clk), .RST(start), .I(x[370]), .Q(
        xin[370]) );
  DFF \xreg_reg[371]  ( .D(xin[370]), .CLK(clk), .RST(start), .I(x[371]), .Q(
        xin[371]) );
  DFF \xreg_reg[372]  ( .D(xin[371]), .CLK(clk), .RST(start), .I(x[372]), .Q(
        xin[372]) );
  DFF \xreg_reg[373]  ( .D(xin[372]), .CLK(clk), .RST(start), .I(x[373]), .Q(
        xin[373]) );
  DFF \xreg_reg[374]  ( .D(xin[373]), .CLK(clk), .RST(start), .I(x[374]), .Q(
        xin[374]) );
  DFF \xreg_reg[375]  ( .D(xin[374]), .CLK(clk), .RST(start), .I(x[375]), .Q(
        xin[375]) );
  DFF \xreg_reg[376]  ( .D(xin[375]), .CLK(clk), .RST(start), .I(x[376]), .Q(
        xin[376]) );
  DFF \xreg_reg[377]  ( .D(xin[376]), .CLK(clk), .RST(start), .I(x[377]), .Q(
        xin[377]) );
  DFF \xreg_reg[378]  ( .D(xin[377]), .CLK(clk), .RST(start), .I(x[378]), .Q(
        xin[378]) );
  DFF \xreg_reg[379]  ( .D(xin[378]), .CLK(clk), .RST(start), .I(x[379]), .Q(
        xin[379]) );
  DFF \xreg_reg[380]  ( .D(xin[379]), .CLK(clk), .RST(start), .I(x[380]), .Q(
        xin[380]) );
  DFF \xreg_reg[381]  ( .D(xin[380]), .CLK(clk), .RST(start), .I(x[381]), .Q(
        xin[381]) );
  DFF \xreg_reg[382]  ( .D(xin[381]), .CLK(clk), .RST(start), .I(x[382]), .Q(
        xin[382]) );
  DFF \xreg_reg[383]  ( .D(xin[382]), .CLK(clk), .RST(start), .I(x[383]), .Q(
        xin[383]) );
  DFF \xreg_reg[384]  ( .D(xin[383]), .CLK(clk), .RST(start), .I(x[384]), .Q(
        xin[384]) );
  DFF \xreg_reg[385]  ( .D(xin[384]), .CLK(clk), .RST(start), .I(x[385]), .Q(
        xin[385]) );
  DFF \xreg_reg[386]  ( .D(xin[385]), .CLK(clk), .RST(start), .I(x[386]), .Q(
        xin[386]) );
  DFF \xreg_reg[387]  ( .D(xin[386]), .CLK(clk), .RST(start), .I(x[387]), .Q(
        xin[387]) );
  DFF \xreg_reg[388]  ( .D(xin[387]), .CLK(clk), .RST(start), .I(x[388]), .Q(
        xin[388]) );
  DFF \xreg_reg[389]  ( .D(xin[388]), .CLK(clk), .RST(start), .I(x[389]), .Q(
        xin[389]) );
  DFF \xreg_reg[390]  ( .D(xin[389]), .CLK(clk), .RST(start), .I(x[390]), .Q(
        xin[390]) );
  DFF \xreg_reg[391]  ( .D(xin[390]), .CLK(clk), .RST(start), .I(x[391]), .Q(
        xin[391]) );
  DFF \xreg_reg[392]  ( .D(xin[391]), .CLK(clk), .RST(start), .I(x[392]), .Q(
        xin[392]) );
  DFF \xreg_reg[393]  ( .D(xin[392]), .CLK(clk), .RST(start), .I(x[393]), .Q(
        xin[393]) );
  DFF \xreg_reg[394]  ( .D(xin[393]), .CLK(clk), .RST(start), .I(x[394]), .Q(
        xin[394]) );
  DFF \xreg_reg[395]  ( .D(xin[394]), .CLK(clk), .RST(start), .I(x[395]), .Q(
        xin[395]) );
  DFF \xreg_reg[396]  ( .D(xin[395]), .CLK(clk), .RST(start), .I(x[396]), .Q(
        xin[396]) );
  DFF \xreg_reg[397]  ( .D(xin[396]), .CLK(clk), .RST(start), .I(x[397]), .Q(
        xin[397]) );
  DFF \xreg_reg[398]  ( .D(xin[397]), .CLK(clk), .RST(start), .I(x[398]), .Q(
        xin[398]) );
  DFF \xreg_reg[399]  ( .D(xin[398]), .CLK(clk), .RST(start), .I(x[399]), .Q(
        xin[399]) );
  DFF \xreg_reg[400]  ( .D(xin[399]), .CLK(clk), .RST(start), .I(x[400]), .Q(
        xin[400]) );
  DFF \xreg_reg[401]  ( .D(xin[400]), .CLK(clk), .RST(start), .I(x[401]), .Q(
        xin[401]) );
  DFF \xreg_reg[402]  ( .D(xin[401]), .CLK(clk), .RST(start), .I(x[402]), .Q(
        xin[402]) );
  DFF \xreg_reg[403]  ( .D(xin[402]), .CLK(clk), .RST(start), .I(x[403]), .Q(
        xin[403]) );
  DFF \xreg_reg[404]  ( .D(xin[403]), .CLK(clk), .RST(start), .I(x[404]), .Q(
        xin[404]) );
  DFF \xreg_reg[405]  ( .D(xin[404]), .CLK(clk), .RST(start), .I(x[405]), .Q(
        xin[405]) );
  DFF \xreg_reg[406]  ( .D(xin[405]), .CLK(clk), .RST(start), .I(x[406]), .Q(
        xin[406]) );
  DFF \xreg_reg[407]  ( .D(xin[406]), .CLK(clk), .RST(start), .I(x[407]), .Q(
        xin[407]) );
  DFF \xreg_reg[408]  ( .D(xin[407]), .CLK(clk), .RST(start), .I(x[408]), .Q(
        xin[408]) );
  DFF \xreg_reg[409]  ( .D(xin[408]), .CLK(clk), .RST(start), .I(x[409]), .Q(
        xin[409]) );
  DFF \xreg_reg[410]  ( .D(xin[409]), .CLK(clk), .RST(start), .I(x[410]), .Q(
        xin[410]) );
  DFF \xreg_reg[411]  ( .D(xin[410]), .CLK(clk), .RST(start), .I(x[411]), .Q(
        xin[411]) );
  DFF \xreg_reg[412]  ( .D(xin[411]), .CLK(clk), .RST(start), .I(x[412]), .Q(
        xin[412]) );
  DFF \xreg_reg[413]  ( .D(xin[412]), .CLK(clk), .RST(start), .I(x[413]), .Q(
        xin[413]) );
  DFF \xreg_reg[414]  ( .D(xin[413]), .CLK(clk), .RST(start), .I(x[414]), .Q(
        xin[414]) );
  DFF \xreg_reg[415]  ( .D(xin[414]), .CLK(clk), .RST(start), .I(x[415]), .Q(
        xin[415]) );
  DFF \xreg_reg[416]  ( .D(xin[415]), .CLK(clk), .RST(start), .I(x[416]), .Q(
        xin[416]) );
  DFF \xreg_reg[417]  ( .D(xin[416]), .CLK(clk), .RST(start), .I(x[417]), .Q(
        xin[417]) );
  DFF \xreg_reg[418]  ( .D(xin[417]), .CLK(clk), .RST(start), .I(x[418]), .Q(
        xin[418]) );
  DFF \xreg_reg[419]  ( .D(xin[418]), .CLK(clk), .RST(start), .I(x[419]), .Q(
        xin[419]) );
  DFF \xreg_reg[420]  ( .D(xin[419]), .CLK(clk), .RST(start), .I(x[420]), .Q(
        xin[420]) );
  DFF \xreg_reg[421]  ( .D(xin[420]), .CLK(clk), .RST(start), .I(x[421]), .Q(
        xin[421]) );
  DFF \xreg_reg[422]  ( .D(xin[421]), .CLK(clk), .RST(start), .I(x[422]), .Q(
        xin[422]) );
  DFF \xreg_reg[423]  ( .D(xin[422]), .CLK(clk), .RST(start), .I(x[423]), .Q(
        xin[423]) );
  DFF \xreg_reg[424]  ( .D(xin[423]), .CLK(clk), .RST(start), .I(x[424]), .Q(
        xin[424]) );
  DFF \xreg_reg[425]  ( .D(xin[424]), .CLK(clk), .RST(start), .I(x[425]), .Q(
        xin[425]) );
  DFF \xreg_reg[426]  ( .D(xin[425]), .CLK(clk), .RST(start), .I(x[426]), .Q(
        xin[426]) );
  DFF \xreg_reg[427]  ( .D(xin[426]), .CLK(clk), .RST(start), .I(x[427]), .Q(
        xin[427]) );
  DFF \xreg_reg[428]  ( .D(xin[427]), .CLK(clk), .RST(start), .I(x[428]), .Q(
        xin[428]) );
  DFF \xreg_reg[429]  ( .D(xin[428]), .CLK(clk), .RST(start), .I(x[429]), .Q(
        xin[429]) );
  DFF \xreg_reg[430]  ( .D(xin[429]), .CLK(clk), .RST(start), .I(x[430]), .Q(
        xin[430]) );
  DFF \xreg_reg[431]  ( .D(xin[430]), .CLK(clk), .RST(start), .I(x[431]), .Q(
        xin[431]) );
  DFF \xreg_reg[432]  ( .D(xin[431]), .CLK(clk), .RST(start), .I(x[432]), .Q(
        xin[432]) );
  DFF \xreg_reg[433]  ( .D(xin[432]), .CLK(clk), .RST(start), .I(x[433]), .Q(
        xin[433]) );
  DFF \xreg_reg[434]  ( .D(xin[433]), .CLK(clk), .RST(start), .I(x[434]), .Q(
        xin[434]) );
  DFF \xreg_reg[435]  ( .D(xin[434]), .CLK(clk), .RST(start), .I(x[435]), .Q(
        xin[435]) );
  DFF \xreg_reg[436]  ( .D(xin[435]), .CLK(clk), .RST(start), .I(x[436]), .Q(
        xin[436]) );
  DFF \xreg_reg[437]  ( .D(xin[436]), .CLK(clk), .RST(start), .I(x[437]), .Q(
        xin[437]) );
  DFF \xreg_reg[438]  ( .D(xin[437]), .CLK(clk), .RST(start), .I(x[438]), .Q(
        xin[438]) );
  DFF \xreg_reg[439]  ( .D(xin[438]), .CLK(clk), .RST(start), .I(x[439]), .Q(
        xin[439]) );
  DFF \xreg_reg[440]  ( .D(xin[439]), .CLK(clk), .RST(start), .I(x[440]), .Q(
        xin[440]) );
  DFF \xreg_reg[441]  ( .D(xin[440]), .CLK(clk), .RST(start), .I(x[441]), .Q(
        xin[441]) );
  DFF \xreg_reg[442]  ( .D(xin[441]), .CLK(clk), .RST(start), .I(x[442]), .Q(
        xin[442]) );
  DFF \xreg_reg[443]  ( .D(xin[442]), .CLK(clk), .RST(start), .I(x[443]), .Q(
        xin[443]) );
  DFF \xreg_reg[444]  ( .D(xin[443]), .CLK(clk), .RST(start), .I(x[444]), .Q(
        xin[444]) );
  DFF \xreg_reg[445]  ( .D(xin[444]), .CLK(clk), .RST(start), .I(x[445]), .Q(
        xin[445]) );
  DFF \xreg_reg[446]  ( .D(xin[445]), .CLK(clk), .RST(start), .I(x[446]), .Q(
        xin[446]) );
  DFF \xreg_reg[447]  ( .D(xin[446]), .CLK(clk), .RST(start), .I(x[447]), .Q(
        xin[447]) );
  DFF \xreg_reg[448]  ( .D(xin[447]), .CLK(clk), .RST(start), .I(x[448]), .Q(
        xin[448]) );
  DFF \xreg_reg[449]  ( .D(xin[448]), .CLK(clk), .RST(start), .I(x[449]), .Q(
        xin[449]) );
  DFF \xreg_reg[450]  ( .D(xin[449]), .CLK(clk), .RST(start), .I(x[450]), .Q(
        xin[450]) );
  DFF \xreg_reg[451]  ( .D(xin[450]), .CLK(clk), .RST(start), .I(x[451]), .Q(
        xin[451]) );
  DFF \xreg_reg[452]  ( .D(xin[451]), .CLK(clk), .RST(start), .I(x[452]), .Q(
        xin[452]) );
  DFF \xreg_reg[453]  ( .D(xin[452]), .CLK(clk), .RST(start), .I(x[453]), .Q(
        xin[453]) );
  DFF \xreg_reg[454]  ( .D(xin[453]), .CLK(clk), .RST(start), .I(x[454]), .Q(
        xin[454]) );
  DFF \xreg_reg[455]  ( .D(xin[454]), .CLK(clk), .RST(start), .I(x[455]), .Q(
        xin[455]) );
  DFF \xreg_reg[456]  ( .D(xin[455]), .CLK(clk), .RST(start), .I(x[456]), .Q(
        xin[456]) );
  DFF \xreg_reg[457]  ( .D(xin[456]), .CLK(clk), .RST(start), .I(x[457]), .Q(
        xin[457]) );
  DFF \xreg_reg[458]  ( .D(xin[457]), .CLK(clk), .RST(start), .I(x[458]), .Q(
        xin[458]) );
  DFF \xreg_reg[459]  ( .D(xin[458]), .CLK(clk), .RST(start), .I(x[459]), .Q(
        xin[459]) );
  DFF \xreg_reg[460]  ( .D(xin[459]), .CLK(clk), .RST(start), .I(x[460]), .Q(
        xin[460]) );
  DFF \xreg_reg[461]  ( .D(xin[460]), .CLK(clk), .RST(start), .I(x[461]), .Q(
        xin[461]) );
  DFF \xreg_reg[462]  ( .D(xin[461]), .CLK(clk), .RST(start), .I(x[462]), .Q(
        xin[462]) );
  DFF \xreg_reg[463]  ( .D(xin[462]), .CLK(clk), .RST(start), .I(x[463]), .Q(
        xin[463]) );
  DFF \xreg_reg[464]  ( .D(xin[463]), .CLK(clk), .RST(start), .I(x[464]), .Q(
        xin[464]) );
  DFF \xreg_reg[465]  ( .D(xin[464]), .CLK(clk), .RST(start), .I(x[465]), .Q(
        xin[465]) );
  DFF \xreg_reg[466]  ( .D(xin[465]), .CLK(clk), .RST(start), .I(x[466]), .Q(
        xin[466]) );
  DFF \xreg_reg[467]  ( .D(xin[466]), .CLK(clk), .RST(start), .I(x[467]), .Q(
        xin[467]) );
  DFF \xreg_reg[468]  ( .D(xin[467]), .CLK(clk), .RST(start), .I(x[468]), .Q(
        xin[468]) );
  DFF \xreg_reg[469]  ( .D(xin[468]), .CLK(clk), .RST(start), .I(x[469]), .Q(
        xin[469]) );
  DFF \xreg_reg[470]  ( .D(xin[469]), .CLK(clk), .RST(start), .I(x[470]), .Q(
        xin[470]) );
  DFF \xreg_reg[471]  ( .D(xin[470]), .CLK(clk), .RST(start), .I(x[471]), .Q(
        xin[471]) );
  DFF \xreg_reg[472]  ( .D(xin[471]), .CLK(clk), .RST(start), .I(x[472]), .Q(
        xin[472]) );
  DFF \xreg_reg[473]  ( .D(xin[472]), .CLK(clk), .RST(start), .I(x[473]), .Q(
        xin[473]) );
  DFF \xreg_reg[474]  ( .D(xin[473]), .CLK(clk), .RST(start), .I(x[474]), .Q(
        xin[474]) );
  DFF \xreg_reg[475]  ( .D(xin[474]), .CLK(clk), .RST(start), .I(x[475]), .Q(
        xin[475]) );
  DFF \xreg_reg[476]  ( .D(xin[475]), .CLK(clk), .RST(start), .I(x[476]), .Q(
        xin[476]) );
  DFF \xreg_reg[477]  ( .D(xin[476]), .CLK(clk), .RST(start), .I(x[477]), .Q(
        xin[477]) );
  DFF \xreg_reg[478]  ( .D(xin[477]), .CLK(clk), .RST(start), .I(x[478]), .Q(
        xin[478]) );
  DFF \xreg_reg[479]  ( .D(xin[478]), .CLK(clk), .RST(start), .I(x[479]), .Q(
        xin[479]) );
  DFF \xreg_reg[480]  ( .D(xin[479]), .CLK(clk), .RST(start), .I(x[480]), .Q(
        xin[480]) );
  DFF \xreg_reg[481]  ( .D(xin[480]), .CLK(clk), .RST(start), .I(x[481]), .Q(
        xin[481]) );
  DFF \xreg_reg[482]  ( .D(xin[481]), .CLK(clk), .RST(start), .I(x[482]), .Q(
        xin[482]) );
  DFF \xreg_reg[483]  ( .D(xin[482]), .CLK(clk), .RST(start), .I(x[483]), .Q(
        xin[483]) );
  DFF \xreg_reg[484]  ( .D(xin[483]), .CLK(clk), .RST(start), .I(x[484]), .Q(
        xin[484]) );
  DFF \xreg_reg[485]  ( .D(xin[484]), .CLK(clk), .RST(start), .I(x[485]), .Q(
        xin[485]) );
  DFF \xreg_reg[486]  ( .D(xin[485]), .CLK(clk), .RST(start), .I(x[486]), .Q(
        xin[486]) );
  DFF \xreg_reg[487]  ( .D(xin[486]), .CLK(clk), .RST(start), .I(x[487]), .Q(
        xin[487]) );
  DFF \xreg_reg[488]  ( .D(xin[487]), .CLK(clk), .RST(start), .I(x[488]), .Q(
        xin[488]) );
  DFF \xreg_reg[489]  ( .D(xin[488]), .CLK(clk), .RST(start), .I(x[489]), .Q(
        xin[489]) );
  DFF \xreg_reg[490]  ( .D(xin[489]), .CLK(clk), .RST(start), .I(x[490]), .Q(
        xin[490]) );
  DFF \xreg_reg[491]  ( .D(xin[490]), .CLK(clk), .RST(start), .I(x[491]), .Q(
        xin[491]) );
  DFF \xreg_reg[492]  ( .D(xin[491]), .CLK(clk), .RST(start), .I(x[492]), .Q(
        xin[492]) );
  DFF \xreg_reg[493]  ( .D(xin[492]), .CLK(clk), .RST(start), .I(x[493]), .Q(
        xin[493]) );
  DFF \xreg_reg[494]  ( .D(xin[493]), .CLK(clk), .RST(start), .I(x[494]), .Q(
        xin[494]) );
  DFF \xreg_reg[495]  ( .D(xin[494]), .CLK(clk), .RST(start), .I(x[495]), .Q(
        xin[495]) );
  DFF \xreg_reg[496]  ( .D(xin[495]), .CLK(clk), .RST(start), .I(x[496]), .Q(
        xin[496]) );
  DFF \xreg_reg[497]  ( .D(xin[496]), .CLK(clk), .RST(start), .I(x[497]), .Q(
        xin[497]) );
  DFF \xreg_reg[498]  ( .D(xin[497]), .CLK(clk), .RST(start), .I(x[498]), .Q(
        xin[498]) );
  DFF \xreg_reg[499]  ( .D(xin[498]), .CLK(clk), .RST(start), .I(x[499]), .Q(
        xin[499]) );
  DFF \xreg_reg[500]  ( .D(xin[499]), .CLK(clk), .RST(start), .I(x[500]), .Q(
        xin[500]) );
  DFF \xreg_reg[501]  ( .D(xin[500]), .CLK(clk), .RST(start), .I(x[501]), .Q(
        xin[501]) );
  DFF \xreg_reg[502]  ( .D(xin[501]), .CLK(clk), .RST(start), .I(x[502]), .Q(
        xin[502]) );
  DFF \xreg_reg[503]  ( .D(xin[502]), .CLK(clk), .RST(start), .I(x[503]), .Q(
        xin[503]) );
  DFF \xreg_reg[504]  ( .D(xin[503]), .CLK(clk), .RST(start), .I(x[504]), .Q(
        xin[504]) );
  DFF \xreg_reg[505]  ( .D(xin[504]), .CLK(clk), .RST(start), .I(x[505]), .Q(
        xin[505]) );
  DFF \xreg_reg[506]  ( .D(xin[505]), .CLK(clk), .RST(start), .I(x[506]), .Q(
        xin[506]) );
  DFF \xreg_reg[507]  ( .D(xin[506]), .CLK(clk), .RST(start), .I(x[507]), .Q(
        xin[507]) );
  DFF \xreg_reg[508]  ( .D(xin[507]), .CLK(clk), .RST(start), .I(x[508]), .Q(
        xin[508]) );
  DFF \xreg_reg[509]  ( .D(xin[508]), .CLK(clk), .RST(start), .I(x[509]), .Q(
        xin[509]) );
  DFF \xreg_reg[510]  ( .D(xin[509]), .CLK(clk), .RST(start), .I(x[510]), .Q(
        xin[510]) );
  DFF \xreg_reg[511]  ( .D(xin[510]), .CLK(clk), .RST(start), .I(x[511]), .Q(
        xin[511]) );
  DFF \zreg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][0] ) );
  DFF \zreg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1] ) );
  DFF \zreg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][2] ) );
  DFF \zreg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][3] ) );
  DFF \zreg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][4] ) );
  DFF \zreg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][5] ) );
  DFF \zreg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][6] ) );
  DFF \zreg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][7] ) );
  DFF \zreg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][8] ) );
  DFF \zreg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][9] ) );
  DFF \zreg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][10] ) );
  DFF \zreg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][11] ) );
  DFF \zreg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][12] ) );
  DFF \zreg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][13] ) );
  DFF \zreg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][14] ) );
  DFF \zreg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][15] ) );
  DFF \zreg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][16] ) );
  DFF \zreg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][17] ) );
  DFF \zreg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][18] ) );
  DFF \zreg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][19] ) );
  DFF \zreg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][20] ) );
  DFF \zreg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][21] ) );
  DFF \zreg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][22] ) );
  DFF \zreg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][23] ) );
  DFF \zreg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][24] ) );
  DFF \zreg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][25] ) );
  DFF \zreg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][26] ) );
  DFF \zreg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][27] ) );
  DFF \zreg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][28] ) );
  DFF \zreg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][29] ) );
  DFF \zreg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][30] ) );
  DFF \zreg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][31] ) );
  DFF \zreg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][32] ) );
  DFF \zreg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][33] ) );
  DFF \zreg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][34] ) );
  DFF \zreg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][35] ) );
  DFF \zreg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][36] ) );
  DFF \zreg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][37] ) );
  DFF \zreg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][38] ) );
  DFF \zreg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][39] ) );
  DFF \zreg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][40] ) );
  DFF \zreg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][41] ) );
  DFF \zreg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][42] ) );
  DFF \zreg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][43] ) );
  DFF \zreg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][44] ) );
  DFF \zreg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][45] ) );
  DFF \zreg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][46] ) );
  DFF \zreg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][47] ) );
  DFF \zreg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][48] ) );
  DFF \zreg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][49] ) );
  DFF \zreg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][50] ) );
  DFF \zreg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][51] ) );
  DFF \zreg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][52] ) );
  DFF \zreg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][53] ) );
  DFF \zreg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][54] ) );
  DFF \zreg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][55] ) );
  DFF \zreg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][56] ) );
  DFF \zreg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][57] ) );
  DFF \zreg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][58] ) );
  DFF \zreg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][59] ) );
  DFF \zreg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][60] ) );
  DFF \zreg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][61] ) );
  DFF \zreg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][62] ) );
  DFF \zreg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][63] ) );
  DFF \zreg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][64] ) );
  DFF \zreg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][65] ) );
  DFF \zreg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][66] ) );
  DFF \zreg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][67] ) );
  DFF \zreg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][68] ) );
  DFF \zreg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][69] ) );
  DFF \zreg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][70] ) );
  DFF \zreg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][71] ) );
  DFF \zreg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][72] ) );
  DFF \zreg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][73] ) );
  DFF \zreg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][74] ) );
  DFF \zreg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][75] ) );
  DFF \zreg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][76] ) );
  DFF \zreg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][77] ) );
  DFF \zreg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][78] ) );
  DFF \zreg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][79] ) );
  DFF \zreg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][80] ) );
  DFF \zreg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][81] ) );
  DFF \zreg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][82] ) );
  DFF \zreg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][83] ) );
  DFF \zreg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][84] ) );
  DFF \zreg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][85] ) );
  DFF \zreg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][86] ) );
  DFF \zreg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][87] ) );
  DFF \zreg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][88] ) );
  DFF \zreg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][89] ) );
  DFF \zreg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][90] ) );
  DFF \zreg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][91] ) );
  DFF \zreg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][92] ) );
  DFF \zreg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][93] ) );
  DFF \zreg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][94] ) );
  DFF \zreg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][95] ) );
  DFF \zreg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][96] ) );
  DFF \zreg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][97] ) );
  DFF \zreg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][98] ) );
  DFF \zreg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][99] ) );
  DFF \zreg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][100] ) );
  DFF \zreg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][101] ) );
  DFF \zreg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][102] ) );
  DFF \zreg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][103] ) );
  DFF \zreg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][104] ) );
  DFF \zreg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][105] ) );
  DFF \zreg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][106] ) );
  DFF \zreg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][107] ) );
  DFF \zreg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][108] ) );
  DFF \zreg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][109] ) );
  DFF \zreg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][110] ) );
  DFF \zreg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][111] ) );
  DFF \zreg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][112] ) );
  DFF \zreg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][113] ) );
  DFF \zreg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][114] ) );
  DFF \zreg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][115] ) );
  DFF \zreg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][116] ) );
  DFF \zreg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][117] ) );
  DFF \zreg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][118] ) );
  DFF \zreg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][119] ) );
  DFF \zreg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][120] ) );
  DFF \zreg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][121] ) );
  DFF \zreg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][122] ) );
  DFF \zreg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][123] ) );
  DFF \zreg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][124] ) );
  DFF \zreg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][125] ) );
  DFF \zreg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][126] ) );
  DFF \zreg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][127] ) );
  DFF \zreg_reg[128]  ( .D(o[128]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][128] ) );
  DFF \zreg_reg[129]  ( .D(o[129]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][129] ) );
  DFF \zreg_reg[130]  ( .D(o[130]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][130] ) );
  DFF \zreg_reg[131]  ( .D(o[131]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][131] ) );
  DFF \zreg_reg[132]  ( .D(o[132]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][132] ) );
  DFF \zreg_reg[133]  ( .D(o[133]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][133] ) );
  DFF \zreg_reg[134]  ( .D(o[134]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][134] ) );
  DFF \zreg_reg[135]  ( .D(o[135]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][135] ) );
  DFF \zreg_reg[136]  ( .D(o[136]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][136] ) );
  DFF \zreg_reg[137]  ( .D(o[137]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][137] ) );
  DFF \zreg_reg[138]  ( .D(o[138]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][138] ) );
  DFF \zreg_reg[139]  ( .D(o[139]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][139] ) );
  DFF \zreg_reg[140]  ( .D(o[140]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][140] ) );
  DFF \zreg_reg[141]  ( .D(o[141]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][141] ) );
  DFF \zreg_reg[142]  ( .D(o[142]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][142] ) );
  DFF \zreg_reg[143]  ( .D(o[143]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][143] ) );
  DFF \zreg_reg[144]  ( .D(o[144]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][144] ) );
  DFF \zreg_reg[145]  ( .D(o[145]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][145] ) );
  DFF \zreg_reg[146]  ( .D(o[146]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][146] ) );
  DFF \zreg_reg[147]  ( .D(o[147]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][147] ) );
  DFF \zreg_reg[148]  ( .D(o[148]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][148] ) );
  DFF \zreg_reg[149]  ( .D(o[149]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][149] ) );
  DFF \zreg_reg[150]  ( .D(o[150]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][150] ) );
  DFF \zreg_reg[151]  ( .D(o[151]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][151] ) );
  DFF \zreg_reg[152]  ( .D(o[152]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][152] ) );
  DFF \zreg_reg[153]  ( .D(o[153]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][153] ) );
  DFF \zreg_reg[154]  ( .D(o[154]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][154] ) );
  DFF \zreg_reg[155]  ( .D(o[155]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][155] ) );
  DFF \zreg_reg[156]  ( .D(o[156]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][156] ) );
  DFF \zreg_reg[157]  ( .D(o[157]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][157] ) );
  DFF \zreg_reg[158]  ( .D(o[158]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][158] ) );
  DFF \zreg_reg[159]  ( .D(o[159]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][159] ) );
  DFF \zreg_reg[160]  ( .D(o[160]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][160] ) );
  DFF \zreg_reg[161]  ( .D(o[161]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][161] ) );
  DFF \zreg_reg[162]  ( .D(o[162]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][162] ) );
  DFF \zreg_reg[163]  ( .D(o[163]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][163] ) );
  DFF \zreg_reg[164]  ( .D(o[164]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][164] ) );
  DFF \zreg_reg[165]  ( .D(o[165]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][165] ) );
  DFF \zreg_reg[166]  ( .D(o[166]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][166] ) );
  DFF \zreg_reg[167]  ( .D(o[167]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][167] ) );
  DFF \zreg_reg[168]  ( .D(o[168]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][168] ) );
  DFF \zreg_reg[169]  ( .D(o[169]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][169] ) );
  DFF \zreg_reg[170]  ( .D(o[170]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][170] ) );
  DFF \zreg_reg[171]  ( .D(o[171]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][171] ) );
  DFF \zreg_reg[172]  ( .D(o[172]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][172] ) );
  DFF \zreg_reg[173]  ( .D(o[173]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][173] ) );
  DFF \zreg_reg[174]  ( .D(o[174]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][174] ) );
  DFF \zreg_reg[175]  ( .D(o[175]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][175] ) );
  DFF \zreg_reg[176]  ( .D(o[176]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][176] ) );
  DFF \zreg_reg[177]  ( .D(o[177]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][177] ) );
  DFF \zreg_reg[178]  ( .D(o[178]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][178] ) );
  DFF \zreg_reg[179]  ( .D(o[179]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][179] ) );
  DFF \zreg_reg[180]  ( .D(o[180]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][180] ) );
  DFF \zreg_reg[181]  ( .D(o[181]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][181] ) );
  DFF \zreg_reg[182]  ( .D(o[182]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][182] ) );
  DFF \zreg_reg[183]  ( .D(o[183]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][183] ) );
  DFF \zreg_reg[184]  ( .D(o[184]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][184] ) );
  DFF \zreg_reg[185]  ( .D(o[185]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][185] ) );
  DFF \zreg_reg[186]  ( .D(o[186]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][186] ) );
  DFF \zreg_reg[187]  ( .D(o[187]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][187] ) );
  DFF \zreg_reg[188]  ( .D(o[188]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][188] ) );
  DFF \zreg_reg[189]  ( .D(o[189]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][189] ) );
  DFF \zreg_reg[190]  ( .D(o[190]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][190] ) );
  DFF \zreg_reg[191]  ( .D(o[191]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][191] ) );
  DFF \zreg_reg[192]  ( .D(o[192]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][192] ) );
  DFF \zreg_reg[193]  ( .D(o[193]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][193] ) );
  DFF \zreg_reg[194]  ( .D(o[194]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][194] ) );
  DFF \zreg_reg[195]  ( .D(o[195]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][195] ) );
  DFF \zreg_reg[196]  ( .D(o[196]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][196] ) );
  DFF \zreg_reg[197]  ( .D(o[197]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][197] ) );
  DFF \zreg_reg[198]  ( .D(o[198]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][198] ) );
  DFF \zreg_reg[199]  ( .D(o[199]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][199] ) );
  DFF \zreg_reg[200]  ( .D(o[200]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][200] ) );
  DFF \zreg_reg[201]  ( .D(o[201]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][201] ) );
  DFF \zreg_reg[202]  ( .D(o[202]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][202] ) );
  DFF \zreg_reg[203]  ( .D(o[203]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][203] ) );
  DFF \zreg_reg[204]  ( .D(o[204]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][204] ) );
  DFF \zreg_reg[205]  ( .D(o[205]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][205] ) );
  DFF \zreg_reg[206]  ( .D(o[206]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][206] ) );
  DFF \zreg_reg[207]  ( .D(o[207]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][207] ) );
  DFF \zreg_reg[208]  ( .D(o[208]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][208] ) );
  DFF \zreg_reg[209]  ( .D(o[209]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][209] ) );
  DFF \zreg_reg[210]  ( .D(o[210]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][210] ) );
  DFF \zreg_reg[211]  ( .D(o[211]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][211] ) );
  DFF \zreg_reg[212]  ( .D(o[212]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][212] ) );
  DFF \zreg_reg[213]  ( .D(o[213]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][213] ) );
  DFF \zreg_reg[214]  ( .D(o[214]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][214] ) );
  DFF \zreg_reg[215]  ( .D(o[215]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][215] ) );
  DFF \zreg_reg[216]  ( .D(o[216]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][216] ) );
  DFF \zreg_reg[217]  ( .D(o[217]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][217] ) );
  DFF \zreg_reg[218]  ( .D(o[218]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][218] ) );
  DFF \zreg_reg[219]  ( .D(o[219]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][219] ) );
  DFF \zreg_reg[220]  ( .D(o[220]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][220] ) );
  DFF \zreg_reg[221]  ( .D(o[221]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][221] ) );
  DFF \zreg_reg[222]  ( .D(o[222]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][222] ) );
  DFF \zreg_reg[223]  ( .D(o[223]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][223] ) );
  DFF \zreg_reg[224]  ( .D(o[224]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][224] ) );
  DFF \zreg_reg[225]  ( .D(o[225]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][225] ) );
  DFF \zreg_reg[226]  ( .D(o[226]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][226] ) );
  DFF \zreg_reg[227]  ( .D(o[227]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][227] ) );
  DFF \zreg_reg[228]  ( .D(o[228]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][228] ) );
  DFF \zreg_reg[229]  ( .D(o[229]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][229] ) );
  DFF \zreg_reg[230]  ( .D(o[230]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][230] ) );
  DFF \zreg_reg[231]  ( .D(o[231]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][231] ) );
  DFF \zreg_reg[232]  ( .D(o[232]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][232] ) );
  DFF \zreg_reg[233]  ( .D(o[233]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][233] ) );
  DFF \zreg_reg[234]  ( .D(o[234]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][234] ) );
  DFF \zreg_reg[235]  ( .D(o[235]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][235] ) );
  DFF \zreg_reg[236]  ( .D(o[236]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][236] ) );
  DFF \zreg_reg[237]  ( .D(o[237]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][237] ) );
  DFF \zreg_reg[238]  ( .D(o[238]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][238] ) );
  DFF \zreg_reg[239]  ( .D(o[239]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][239] ) );
  DFF \zreg_reg[240]  ( .D(o[240]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][240] ) );
  DFF \zreg_reg[241]  ( .D(o[241]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][241] ) );
  DFF \zreg_reg[242]  ( .D(o[242]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][242] ) );
  DFF \zreg_reg[243]  ( .D(o[243]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][243] ) );
  DFF \zreg_reg[244]  ( .D(o[244]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][244] ) );
  DFF \zreg_reg[245]  ( .D(o[245]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][245] ) );
  DFF \zreg_reg[246]  ( .D(o[246]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][246] ) );
  DFF \zreg_reg[247]  ( .D(o[247]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][247] ) );
  DFF \zreg_reg[248]  ( .D(o[248]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][248] ) );
  DFF \zreg_reg[249]  ( .D(o[249]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][249] ) );
  DFF \zreg_reg[250]  ( .D(o[250]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][250] ) );
  DFF \zreg_reg[251]  ( .D(o[251]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][251] ) );
  DFF \zreg_reg[252]  ( .D(o[252]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][252] ) );
  DFF \zreg_reg[253]  ( .D(o[253]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][253] ) );
  DFF \zreg_reg[254]  ( .D(o[254]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][254] ) );
  DFF \zreg_reg[255]  ( .D(o[255]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][255] ) );
  DFF \zreg_reg[256]  ( .D(o[256]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][256] ) );
  DFF \zreg_reg[257]  ( .D(o[257]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][257] ) );
  DFF \zreg_reg[258]  ( .D(o[258]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][258] ) );
  DFF \zreg_reg[259]  ( .D(o[259]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][259] ) );
  DFF \zreg_reg[260]  ( .D(o[260]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][260] ) );
  DFF \zreg_reg[261]  ( .D(o[261]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][261] ) );
  DFF \zreg_reg[262]  ( .D(o[262]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][262] ) );
  DFF \zreg_reg[263]  ( .D(o[263]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][263] ) );
  DFF \zreg_reg[264]  ( .D(o[264]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][264] ) );
  DFF \zreg_reg[265]  ( .D(o[265]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][265] ) );
  DFF \zreg_reg[266]  ( .D(o[266]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][266] ) );
  DFF \zreg_reg[267]  ( .D(o[267]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][267] ) );
  DFF \zreg_reg[268]  ( .D(o[268]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][268] ) );
  DFF \zreg_reg[269]  ( .D(o[269]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][269] ) );
  DFF \zreg_reg[270]  ( .D(o[270]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][270] ) );
  DFF \zreg_reg[271]  ( .D(o[271]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][271] ) );
  DFF \zreg_reg[272]  ( .D(o[272]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][272] ) );
  DFF \zreg_reg[273]  ( .D(o[273]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][273] ) );
  DFF \zreg_reg[274]  ( .D(o[274]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][274] ) );
  DFF \zreg_reg[275]  ( .D(o[275]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][275] ) );
  DFF \zreg_reg[276]  ( .D(o[276]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][276] ) );
  DFF \zreg_reg[277]  ( .D(o[277]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][277] ) );
  DFF \zreg_reg[278]  ( .D(o[278]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][278] ) );
  DFF \zreg_reg[279]  ( .D(o[279]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][279] ) );
  DFF \zreg_reg[280]  ( .D(o[280]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][280] ) );
  DFF \zreg_reg[281]  ( .D(o[281]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][281] ) );
  DFF \zreg_reg[282]  ( .D(o[282]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][282] ) );
  DFF \zreg_reg[283]  ( .D(o[283]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][283] ) );
  DFF \zreg_reg[284]  ( .D(o[284]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][284] ) );
  DFF \zreg_reg[285]  ( .D(o[285]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][285] ) );
  DFF \zreg_reg[286]  ( .D(o[286]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][286] ) );
  DFF \zreg_reg[287]  ( .D(o[287]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][287] ) );
  DFF \zreg_reg[288]  ( .D(o[288]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][288] ) );
  DFF \zreg_reg[289]  ( .D(o[289]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][289] ) );
  DFF \zreg_reg[290]  ( .D(o[290]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][290] ) );
  DFF \zreg_reg[291]  ( .D(o[291]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][291] ) );
  DFF \zreg_reg[292]  ( .D(o[292]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][292] ) );
  DFF \zreg_reg[293]  ( .D(o[293]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][293] ) );
  DFF \zreg_reg[294]  ( .D(o[294]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][294] ) );
  DFF \zreg_reg[295]  ( .D(o[295]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][295] ) );
  DFF \zreg_reg[296]  ( .D(o[296]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][296] ) );
  DFF \zreg_reg[297]  ( .D(o[297]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][297] ) );
  DFF \zreg_reg[298]  ( .D(o[298]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][298] ) );
  DFF \zreg_reg[299]  ( .D(o[299]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][299] ) );
  DFF \zreg_reg[300]  ( .D(o[300]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][300] ) );
  DFF \zreg_reg[301]  ( .D(o[301]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][301] ) );
  DFF \zreg_reg[302]  ( .D(o[302]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][302] ) );
  DFF \zreg_reg[303]  ( .D(o[303]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][303] ) );
  DFF \zreg_reg[304]  ( .D(o[304]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][304] ) );
  DFF \zreg_reg[305]  ( .D(o[305]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][305] ) );
  DFF \zreg_reg[306]  ( .D(o[306]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][306] ) );
  DFF \zreg_reg[307]  ( .D(o[307]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][307] ) );
  DFF \zreg_reg[308]  ( .D(o[308]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][308] ) );
  DFF \zreg_reg[309]  ( .D(o[309]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][309] ) );
  DFF \zreg_reg[310]  ( .D(o[310]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][310] ) );
  DFF \zreg_reg[311]  ( .D(o[311]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][311] ) );
  DFF \zreg_reg[312]  ( .D(o[312]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][312] ) );
  DFF \zreg_reg[313]  ( .D(o[313]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][313] ) );
  DFF \zreg_reg[314]  ( .D(o[314]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][314] ) );
  DFF \zreg_reg[315]  ( .D(o[315]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][315] ) );
  DFF \zreg_reg[316]  ( .D(o[316]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][316] ) );
  DFF \zreg_reg[317]  ( .D(o[317]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][317] ) );
  DFF \zreg_reg[318]  ( .D(o[318]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][318] ) );
  DFF \zreg_reg[319]  ( .D(o[319]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][319] ) );
  DFF \zreg_reg[320]  ( .D(o[320]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][320] ) );
  DFF \zreg_reg[321]  ( .D(o[321]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][321] ) );
  DFF \zreg_reg[322]  ( .D(o[322]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][322] ) );
  DFF \zreg_reg[323]  ( .D(o[323]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][323] ) );
  DFF \zreg_reg[324]  ( .D(o[324]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][324] ) );
  DFF \zreg_reg[325]  ( .D(o[325]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][325] ) );
  DFF \zreg_reg[326]  ( .D(o[326]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][326] ) );
  DFF \zreg_reg[327]  ( .D(o[327]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][327] ) );
  DFF \zreg_reg[328]  ( .D(o[328]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][328] ) );
  DFF \zreg_reg[329]  ( .D(o[329]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][329] ) );
  DFF \zreg_reg[330]  ( .D(o[330]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][330] ) );
  DFF \zreg_reg[331]  ( .D(o[331]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][331] ) );
  DFF \zreg_reg[332]  ( .D(o[332]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][332] ) );
  DFF \zreg_reg[333]  ( .D(o[333]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][333] ) );
  DFF \zreg_reg[334]  ( .D(o[334]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][334] ) );
  DFF \zreg_reg[335]  ( .D(o[335]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][335] ) );
  DFF \zreg_reg[336]  ( .D(o[336]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][336] ) );
  DFF \zreg_reg[337]  ( .D(o[337]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][337] ) );
  DFF \zreg_reg[338]  ( .D(o[338]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][338] ) );
  DFF \zreg_reg[339]  ( .D(o[339]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][339] ) );
  DFF \zreg_reg[340]  ( .D(o[340]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][340] ) );
  DFF \zreg_reg[341]  ( .D(o[341]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][341] ) );
  DFF \zreg_reg[342]  ( .D(o[342]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][342] ) );
  DFF \zreg_reg[343]  ( .D(o[343]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][343] ) );
  DFF \zreg_reg[344]  ( .D(o[344]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][344] ) );
  DFF \zreg_reg[345]  ( .D(o[345]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][345] ) );
  DFF \zreg_reg[346]  ( .D(o[346]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][346] ) );
  DFF \zreg_reg[347]  ( .D(o[347]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][347] ) );
  DFF \zreg_reg[348]  ( .D(o[348]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][348] ) );
  DFF \zreg_reg[349]  ( .D(o[349]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][349] ) );
  DFF \zreg_reg[350]  ( .D(o[350]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][350] ) );
  DFF \zreg_reg[351]  ( .D(o[351]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][351] ) );
  DFF \zreg_reg[352]  ( .D(o[352]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][352] ) );
  DFF \zreg_reg[353]  ( .D(o[353]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][353] ) );
  DFF \zreg_reg[354]  ( .D(o[354]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][354] ) );
  DFF \zreg_reg[355]  ( .D(o[355]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][355] ) );
  DFF \zreg_reg[356]  ( .D(o[356]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][356] ) );
  DFF \zreg_reg[357]  ( .D(o[357]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][357] ) );
  DFF \zreg_reg[358]  ( .D(o[358]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][358] ) );
  DFF \zreg_reg[359]  ( .D(o[359]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][359] ) );
  DFF \zreg_reg[360]  ( .D(o[360]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][360] ) );
  DFF \zreg_reg[361]  ( .D(o[361]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][361] ) );
  DFF \zreg_reg[362]  ( .D(o[362]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][362] ) );
  DFF \zreg_reg[363]  ( .D(o[363]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][363] ) );
  DFF \zreg_reg[364]  ( .D(o[364]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][364] ) );
  DFF \zreg_reg[365]  ( .D(o[365]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][365] ) );
  DFF \zreg_reg[366]  ( .D(o[366]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][366] ) );
  DFF \zreg_reg[367]  ( .D(o[367]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][367] ) );
  DFF \zreg_reg[368]  ( .D(o[368]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][368] ) );
  DFF \zreg_reg[369]  ( .D(o[369]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][369] ) );
  DFF \zreg_reg[370]  ( .D(o[370]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][370] ) );
  DFF \zreg_reg[371]  ( .D(o[371]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][371] ) );
  DFF \zreg_reg[372]  ( .D(o[372]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][372] ) );
  DFF \zreg_reg[373]  ( .D(o[373]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][373] ) );
  DFF \zreg_reg[374]  ( .D(o[374]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][374] ) );
  DFF \zreg_reg[375]  ( .D(o[375]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][375] ) );
  DFF \zreg_reg[376]  ( .D(o[376]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][376] ) );
  DFF \zreg_reg[377]  ( .D(o[377]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][377] ) );
  DFF \zreg_reg[378]  ( .D(o[378]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][378] ) );
  DFF \zreg_reg[379]  ( .D(o[379]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][379] ) );
  DFF \zreg_reg[380]  ( .D(o[380]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][380] ) );
  DFF \zreg_reg[381]  ( .D(o[381]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][381] ) );
  DFF \zreg_reg[382]  ( .D(o[382]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][382] ) );
  DFF \zreg_reg[383]  ( .D(o[383]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][383] ) );
  DFF \zreg_reg[384]  ( .D(o[384]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][384] ) );
  DFF \zreg_reg[385]  ( .D(o[385]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][385] ) );
  DFF \zreg_reg[386]  ( .D(o[386]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][386] ) );
  DFF \zreg_reg[387]  ( .D(o[387]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][387] ) );
  DFF \zreg_reg[388]  ( .D(o[388]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][388] ) );
  DFF \zreg_reg[389]  ( .D(o[389]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][389] ) );
  DFF \zreg_reg[390]  ( .D(o[390]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][390] ) );
  DFF \zreg_reg[391]  ( .D(o[391]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][391] ) );
  DFF \zreg_reg[392]  ( .D(o[392]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][392] ) );
  DFF \zreg_reg[393]  ( .D(o[393]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][393] ) );
  DFF \zreg_reg[394]  ( .D(o[394]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][394] ) );
  DFF \zreg_reg[395]  ( .D(o[395]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][395] ) );
  DFF \zreg_reg[396]  ( .D(o[396]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][396] ) );
  DFF \zreg_reg[397]  ( .D(o[397]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][397] ) );
  DFF \zreg_reg[398]  ( .D(o[398]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][398] ) );
  DFF \zreg_reg[399]  ( .D(o[399]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][399] ) );
  DFF \zreg_reg[400]  ( .D(o[400]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][400] ) );
  DFF \zreg_reg[401]  ( .D(o[401]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][401] ) );
  DFF \zreg_reg[402]  ( .D(o[402]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][402] ) );
  DFF \zreg_reg[403]  ( .D(o[403]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][403] ) );
  DFF \zreg_reg[404]  ( .D(o[404]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][404] ) );
  DFF \zreg_reg[405]  ( .D(o[405]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][405] ) );
  DFF \zreg_reg[406]  ( .D(o[406]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][406] ) );
  DFF \zreg_reg[407]  ( .D(o[407]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][407] ) );
  DFF \zreg_reg[408]  ( .D(o[408]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][408] ) );
  DFF \zreg_reg[409]  ( .D(o[409]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][409] ) );
  DFF \zreg_reg[410]  ( .D(o[410]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][410] ) );
  DFF \zreg_reg[411]  ( .D(o[411]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][411] ) );
  DFF \zreg_reg[412]  ( .D(o[412]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][412] ) );
  DFF \zreg_reg[413]  ( .D(o[413]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][413] ) );
  DFF \zreg_reg[414]  ( .D(o[414]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][414] ) );
  DFF \zreg_reg[415]  ( .D(o[415]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][415] ) );
  DFF \zreg_reg[416]  ( .D(o[416]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][416] ) );
  DFF \zreg_reg[417]  ( .D(o[417]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][417] ) );
  DFF \zreg_reg[418]  ( .D(o[418]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][418] ) );
  DFF \zreg_reg[419]  ( .D(o[419]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][419] ) );
  DFF \zreg_reg[420]  ( .D(o[420]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][420] ) );
  DFF \zreg_reg[421]  ( .D(o[421]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][421] ) );
  DFF \zreg_reg[422]  ( .D(o[422]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][422] ) );
  DFF \zreg_reg[423]  ( .D(o[423]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][423] ) );
  DFF \zreg_reg[424]  ( .D(o[424]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][424] ) );
  DFF \zreg_reg[425]  ( .D(o[425]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][425] ) );
  DFF \zreg_reg[426]  ( .D(o[426]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][426] ) );
  DFF \zreg_reg[427]  ( .D(o[427]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][427] ) );
  DFF \zreg_reg[428]  ( .D(o[428]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][428] ) );
  DFF \zreg_reg[429]  ( .D(o[429]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][429] ) );
  DFF \zreg_reg[430]  ( .D(o[430]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][430] ) );
  DFF \zreg_reg[431]  ( .D(o[431]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][431] ) );
  DFF \zreg_reg[432]  ( .D(o[432]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][432] ) );
  DFF \zreg_reg[433]  ( .D(o[433]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][433] ) );
  DFF \zreg_reg[434]  ( .D(o[434]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][434] ) );
  DFF \zreg_reg[435]  ( .D(o[435]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][435] ) );
  DFF \zreg_reg[436]  ( .D(o[436]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][436] ) );
  DFF \zreg_reg[437]  ( .D(o[437]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][437] ) );
  DFF \zreg_reg[438]  ( .D(o[438]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][438] ) );
  DFF \zreg_reg[439]  ( .D(o[439]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][439] ) );
  DFF \zreg_reg[440]  ( .D(o[440]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][440] ) );
  DFF \zreg_reg[441]  ( .D(o[441]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][441] ) );
  DFF \zreg_reg[442]  ( .D(o[442]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][442] ) );
  DFF \zreg_reg[443]  ( .D(o[443]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][443] ) );
  DFF \zreg_reg[444]  ( .D(o[444]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][444] ) );
  DFF \zreg_reg[445]  ( .D(o[445]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][445] ) );
  DFF \zreg_reg[446]  ( .D(o[446]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][446] ) );
  DFF \zreg_reg[447]  ( .D(o[447]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][447] ) );
  DFF \zreg_reg[448]  ( .D(o[448]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][448] ) );
  DFF \zreg_reg[449]  ( .D(o[449]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][449] ) );
  DFF \zreg_reg[450]  ( .D(o[450]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][450] ) );
  DFF \zreg_reg[451]  ( .D(o[451]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][451] ) );
  DFF \zreg_reg[452]  ( .D(o[452]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][452] ) );
  DFF \zreg_reg[453]  ( .D(o[453]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][453] ) );
  DFF \zreg_reg[454]  ( .D(o[454]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][454] ) );
  DFF \zreg_reg[455]  ( .D(o[455]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][455] ) );
  DFF \zreg_reg[456]  ( .D(o[456]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][456] ) );
  DFF \zreg_reg[457]  ( .D(o[457]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][457] ) );
  DFF \zreg_reg[458]  ( .D(o[458]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][458] ) );
  DFF \zreg_reg[459]  ( .D(o[459]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][459] ) );
  DFF \zreg_reg[460]  ( .D(o[460]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][460] ) );
  DFF \zreg_reg[461]  ( .D(o[461]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][461] ) );
  DFF \zreg_reg[462]  ( .D(o[462]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][462] ) );
  DFF \zreg_reg[463]  ( .D(o[463]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][463] ) );
  DFF \zreg_reg[464]  ( .D(o[464]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][464] ) );
  DFF \zreg_reg[465]  ( .D(o[465]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][465] ) );
  DFF \zreg_reg[466]  ( .D(o[466]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][466] ) );
  DFF \zreg_reg[467]  ( .D(o[467]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][467] ) );
  DFF \zreg_reg[468]  ( .D(o[468]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][468] ) );
  DFF \zreg_reg[469]  ( .D(o[469]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][469] ) );
  DFF \zreg_reg[470]  ( .D(o[470]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][470] ) );
  DFF \zreg_reg[471]  ( .D(o[471]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][471] ) );
  DFF \zreg_reg[472]  ( .D(o[472]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][472] ) );
  DFF \zreg_reg[473]  ( .D(o[473]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][473] ) );
  DFF \zreg_reg[474]  ( .D(o[474]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][474] ) );
  DFF \zreg_reg[475]  ( .D(o[475]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][475] ) );
  DFF \zreg_reg[476]  ( .D(o[476]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][476] ) );
  DFF \zreg_reg[477]  ( .D(o[477]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][477] ) );
  DFF \zreg_reg[478]  ( .D(o[478]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][478] ) );
  DFF \zreg_reg[479]  ( .D(o[479]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][479] ) );
  DFF \zreg_reg[480]  ( .D(o[480]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][480] ) );
  DFF \zreg_reg[481]  ( .D(o[481]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][481] ) );
  DFF \zreg_reg[482]  ( .D(o[482]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][482] ) );
  DFF \zreg_reg[483]  ( .D(o[483]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][483] ) );
  DFF \zreg_reg[484]  ( .D(o[484]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][484] ) );
  DFF \zreg_reg[485]  ( .D(o[485]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][485] ) );
  DFF \zreg_reg[486]  ( .D(o[486]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][486] ) );
  DFF \zreg_reg[487]  ( .D(o[487]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][487] ) );
  DFF \zreg_reg[488]  ( .D(o[488]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][488] ) );
  DFF \zreg_reg[489]  ( .D(o[489]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][489] ) );
  DFF \zreg_reg[490]  ( .D(o[490]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][490] ) );
  DFF \zreg_reg[491]  ( .D(o[491]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][491] ) );
  DFF \zreg_reg[492]  ( .D(o[492]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][492] ) );
  DFF \zreg_reg[493]  ( .D(o[493]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][493] ) );
  DFF \zreg_reg[494]  ( .D(o[494]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][494] ) );
  DFF \zreg_reg[495]  ( .D(o[495]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][495] ) );
  DFF \zreg_reg[496]  ( .D(o[496]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][496] ) );
  DFF \zreg_reg[497]  ( .D(o[497]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][497] ) );
  DFF \zreg_reg[498]  ( .D(o[498]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][498] ) );
  DFF \zreg_reg[499]  ( .D(o[499]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][499] ) );
  DFF \zreg_reg[500]  ( .D(o[500]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][500] ) );
  DFF \zreg_reg[501]  ( .D(o[501]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][501] ) );
  DFF \zreg_reg[502]  ( .D(o[502]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][502] ) );
  DFF \zreg_reg[503]  ( .D(o[503]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][503] ) );
  DFF \zreg_reg[504]  ( .D(o[504]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][504] ) );
  DFF \zreg_reg[505]  ( .D(o[505]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][505] ) );
  DFF \zreg_reg[506]  ( .D(o[506]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][506] ) );
  DFF \zreg_reg[507]  ( .D(o[507]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][507] ) );
  DFF \zreg_reg[508]  ( .D(o[508]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][508] ) );
  DFF \zreg_reg[509]  ( .D(o[509]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][509] ) );
  DFF \zreg_reg[510]  ( .D(o[510]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][510] ) );
  DFF \zreg_reg[511]  ( .D(o[511]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][511] ) );
  DFF \zreg_reg[512]  ( .D(\zout[0][512] ), .CLK(clk), .RST(start), .I(1'b0), 
        .Q(\zin[0][512] ) );
endmodule


module MUX_N512_1 ( A, B, S, O );
  input [511:0] A;
  input [511:0] B;
  output [511:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024;

  XOR U1 ( .A(A[9]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U4 ( .A(A[99]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U7 ( .A(A[98]), .B(n5), .Z(O[98]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[98]), .B(A[98]), .Z(n6) );
  XOR U10 ( .A(A[97]), .B(n7), .Z(O[97]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[97]), .B(A[97]), .Z(n8) );
  XOR U13 ( .A(A[96]), .B(n9), .Z(O[96]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[96]), .B(A[96]), .Z(n10) );
  XOR U16 ( .A(A[95]), .B(n11), .Z(O[95]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[95]), .B(A[95]), .Z(n12) );
  XOR U19 ( .A(A[94]), .B(n13), .Z(O[94]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[94]), .B(A[94]), .Z(n14) );
  XOR U22 ( .A(A[93]), .B(n15), .Z(O[93]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[93]), .B(A[93]), .Z(n16) );
  XOR U25 ( .A(A[92]), .B(n17), .Z(O[92]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[92]), .B(A[92]), .Z(n18) );
  XOR U28 ( .A(A[91]), .B(n19), .Z(O[91]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[91]), .B(A[91]), .Z(n20) );
  XOR U31 ( .A(A[90]), .B(n21), .Z(O[90]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[90]), .B(A[90]), .Z(n22) );
  XOR U34 ( .A(A[8]), .B(n23), .Z(O[8]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR U37 ( .A(A[89]), .B(n25), .Z(O[89]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[89]), .B(A[89]), .Z(n26) );
  XOR U40 ( .A(A[88]), .B(n27), .Z(O[88]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[88]), .B(A[88]), .Z(n28) );
  XOR U43 ( .A(A[87]), .B(n29), .Z(O[87]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[87]), .B(A[87]), .Z(n30) );
  XOR U46 ( .A(A[86]), .B(n31), .Z(O[86]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[86]), .B(A[86]), .Z(n32) );
  XOR U49 ( .A(A[85]), .B(n33), .Z(O[85]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[85]), .B(A[85]), .Z(n34) );
  XOR U52 ( .A(A[84]), .B(n35), .Z(O[84]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[84]), .B(A[84]), .Z(n36) );
  XOR U55 ( .A(A[83]), .B(n37), .Z(O[83]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[83]), .B(A[83]), .Z(n38) );
  XOR U58 ( .A(A[82]), .B(n39), .Z(O[82]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[82]), .B(A[82]), .Z(n40) );
  XOR U61 ( .A(A[81]), .B(n41), .Z(O[81]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[81]), .B(A[81]), .Z(n42) );
  XOR U64 ( .A(A[80]), .B(n43), .Z(O[80]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[80]), .B(A[80]), .Z(n44) );
  XOR U67 ( .A(A[7]), .B(n45), .Z(O[7]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[7]), .B(A[7]), .Z(n46) );
  XOR U70 ( .A(A[79]), .B(n47), .Z(O[79]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[79]), .B(A[79]), .Z(n48) );
  XOR U73 ( .A(A[78]), .B(n49), .Z(O[78]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[78]), .B(A[78]), .Z(n50) );
  XOR U76 ( .A(A[77]), .B(n51), .Z(O[77]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[77]), .B(A[77]), .Z(n52) );
  XOR U79 ( .A(A[76]), .B(n53), .Z(O[76]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[76]), .B(A[76]), .Z(n54) );
  XOR U82 ( .A(A[75]), .B(n55), .Z(O[75]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[75]), .B(A[75]), .Z(n56) );
  XOR U85 ( .A(A[74]), .B(n57), .Z(O[74]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[74]), .B(A[74]), .Z(n58) );
  XOR U88 ( .A(A[73]), .B(n59), .Z(O[73]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[73]), .B(A[73]), .Z(n60) );
  XOR U91 ( .A(A[72]), .B(n61), .Z(O[72]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[72]), .B(A[72]), .Z(n62) );
  XOR U94 ( .A(A[71]), .B(n63), .Z(O[71]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[71]), .B(A[71]), .Z(n64) );
  XOR U97 ( .A(A[70]), .B(n65), .Z(O[70]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[70]), .B(A[70]), .Z(n66) );
  XOR U100 ( .A(A[6]), .B(n67), .Z(O[6]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[6]), .B(A[6]), .Z(n68) );
  XOR U103 ( .A(A[69]), .B(n69), .Z(O[69]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[69]), .B(A[69]), .Z(n70) );
  XOR U106 ( .A(A[68]), .B(n71), .Z(O[68]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[68]), .B(A[68]), .Z(n72) );
  XOR U109 ( .A(A[67]), .B(n73), .Z(O[67]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[67]), .B(A[67]), .Z(n74) );
  XOR U112 ( .A(A[66]), .B(n75), .Z(O[66]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[66]), .B(A[66]), .Z(n76) );
  XOR U115 ( .A(A[65]), .B(n77), .Z(O[65]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[65]), .B(A[65]), .Z(n78) );
  XOR U118 ( .A(A[64]), .B(n79), .Z(O[64]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[64]), .B(A[64]), .Z(n80) );
  XOR U121 ( .A(A[63]), .B(n81), .Z(O[63]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[63]), .B(A[63]), .Z(n82) );
  XOR U124 ( .A(A[62]), .B(n83), .Z(O[62]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[62]), .B(A[62]), .Z(n84) );
  XOR U127 ( .A(A[61]), .B(n85), .Z(O[61]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[61]), .B(A[61]), .Z(n86) );
  XOR U130 ( .A(A[60]), .B(n87), .Z(O[60]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[60]), .B(A[60]), .Z(n88) );
  XOR U133 ( .A(A[5]), .B(n89), .Z(O[5]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[5]), .B(A[5]), .Z(n90) );
  XOR U136 ( .A(A[59]), .B(n91), .Z(O[59]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[59]), .B(A[59]), .Z(n92) );
  XOR U139 ( .A(A[58]), .B(n93), .Z(O[58]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[58]), .B(A[58]), .Z(n94) );
  XOR U142 ( .A(A[57]), .B(n95), .Z(O[57]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[57]), .B(A[57]), .Z(n96) );
  XOR U145 ( .A(A[56]), .B(n97), .Z(O[56]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[56]), .B(A[56]), .Z(n98) );
  XOR U148 ( .A(A[55]), .B(n99), .Z(O[55]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[55]), .B(A[55]), .Z(n100) );
  XOR U151 ( .A(A[54]), .B(n101), .Z(O[54]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[54]), .B(A[54]), .Z(n102) );
  XOR U154 ( .A(A[53]), .B(n103), .Z(O[53]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[53]), .B(A[53]), .Z(n104) );
  XOR U157 ( .A(A[52]), .B(n105), .Z(O[52]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[52]), .B(A[52]), .Z(n106) );
  XOR U160 ( .A(A[51]), .B(n107), .Z(O[51]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[51]), .B(A[51]), .Z(n108) );
  XOR U163 ( .A(A[511]), .B(n109), .Z(O[511]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[511]), .B(A[511]), .Z(n110) );
  XOR U166 ( .A(A[510]), .B(n111), .Z(O[510]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[510]), .B(A[510]), .Z(n112) );
  XOR U169 ( .A(A[50]), .B(n113), .Z(O[50]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[50]), .B(A[50]), .Z(n114) );
  XOR U172 ( .A(A[509]), .B(n115), .Z(O[509]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[509]), .B(A[509]), .Z(n116) );
  XOR U175 ( .A(A[508]), .B(n117), .Z(O[508]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[508]), .B(A[508]), .Z(n118) );
  XOR U178 ( .A(A[507]), .B(n119), .Z(O[507]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[507]), .B(A[507]), .Z(n120) );
  XOR U181 ( .A(A[506]), .B(n121), .Z(O[506]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[506]), .B(A[506]), .Z(n122) );
  XOR U184 ( .A(A[505]), .B(n123), .Z(O[505]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[505]), .B(A[505]), .Z(n124) );
  XOR U187 ( .A(A[504]), .B(n125), .Z(O[504]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[504]), .B(A[504]), .Z(n126) );
  XOR U190 ( .A(A[503]), .B(n127), .Z(O[503]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[503]), .B(A[503]), .Z(n128) );
  XOR U193 ( .A(A[502]), .B(n129), .Z(O[502]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[502]), .B(A[502]), .Z(n130) );
  XOR U196 ( .A(A[501]), .B(n131), .Z(O[501]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[501]), .B(A[501]), .Z(n132) );
  XOR U199 ( .A(A[500]), .B(n133), .Z(O[500]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[500]), .B(A[500]), .Z(n134) );
  XOR U202 ( .A(A[4]), .B(n135), .Z(O[4]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[4]), .B(A[4]), .Z(n136) );
  XOR U205 ( .A(A[49]), .B(n137), .Z(O[49]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[49]), .B(A[49]), .Z(n138) );
  XOR U208 ( .A(A[499]), .B(n139), .Z(O[499]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[499]), .B(A[499]), .Z(n140) );
  XOR U211 ( .A(A[498]), .B(n141), .Z(O[498]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[498]), .B(A[498]), .Z(n142) );
  XOR U214 ( .A(A[497]), .B(n143), .Z(O[497]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[497]), .B(A[497]), .Z(n144) );
  XOR U217 ( .A(A[496]), .B(n145), .Z(O[496]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[496]), .B(A[496]), .Z(n146) );
  XOR U220 ( .A(A[495]), .B(n147), .Z(O[495]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[495]), .B(A[495]), .Z(n148) );
  XOR U223 ( .A(A[494]), .B(n149), .Z(O[494]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[494]), .B(A[494]), .Z(n150) );
  XOR U226 ( .A(A[493]), .B(n151), .Z(O[493]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[493]), .B(A[493]), .Z(n152) );
  XOR U229 ( .A(A[492]), .B(n153), .Z(O[492]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[492]), .B(A[492]), .Z(n154) );
  XOR U232 ( .A(A[491]), .B(n155), .Z(O[491]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[491]), .B(A[491]), .Z(n156) );
  XOR U235 ( .A(A[490]), .B(n157), .Z(O[490]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[490]), .B(A[490]), .Z(n158) );
  XOR U238 ( .A(A[48]), .B(n159), .Z(O[48]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[48]), .B(A[48]), .Z(n160) );
  XOR U241 ( .A(A[489]), .B(n161), .Z(O[489]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[489]), .B(A[489]), .Z(n162) );
  XOR U244 ( .A(A[488]), .B(n163), .Z(O[488]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[488]), .B(A[488]), .Z(n164) );
  XOR U247 ( .A(A[487]), .B(n165), .Z(O[487]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[487]), .B(A[487]), .Z(n166) );
  XOR U250 ( .A(A[486]), .B(n167), .Z(O[486]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[486]), .B(A[486]), .Z(n168) );
  XOR U253 ( .A(A[485]), .B(n169), .Z(O[485]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[485]), .B(A[485]), .Z(n170) );
  XOR U256 ( .A(A[484]), .B(n171), .Z(O[484]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[484]), .B(A[484]), .Z(n172) );
  XOR U259 ( .A(A[483]), .B(n173), .Z(O[483]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[483]), .B(A[483]), .Z(n174) );
  XOR U262 ( .A(A[482]), .B(n175), .Z(O[482]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[482]), .B(A[482]), .Z(n176) );
  XOR U265 ( .A(A[481]), .B(n177), .Z(O[481]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[481]), .B(A[481]), .Z(n178) );
  XOR U268 ( .A(A[480]), .B(n179), .Z(O[480]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[480]), .B(A[480]), .Z(n180) );
  XOR U271 ( .A(A[47]), .B(n181), .Z(O[47]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[47]), .B(A[47]), .Z(n182) );
  XOR U274 ( .A(A[479]), .B(n183), .Z(O[479]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[479]), .B(A[479]), .Z(n184) );
  XOR U277 ( .A(A[478]), .B(n185), .Z(O[478]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[478]), .B(A[478]), .Z(n186) );
  XOR U280 ( .A(A[477]), .B(n187), .Z(O[477]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[477]), .B(A[477]), .Z(n188) );
  XOR U283 ( .A(A[476]), .B(n189), .Z(O[476]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[476]), .B(A[476]), .Z(n190) );
  XOR U286 ( .A(A[475]), .B(n191), .Z(O[475]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[475]), .B(A[475]), .Z(n192) );
  XOR U289 ( .A(A[474]), .B(n193), .Z(O[474]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[474]), .B(A[474]), .Z(n194) );
  XOR U292 ( .A(A[473]), .B(n195), .Z(O[473]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[473]), .B(A[473]), .Z(n196) );
  XOR U295 ( .A(A[472]), .B(n197), .Z(O[472]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[472]), .B(A[472]), .Z(n198) );
  XOR U298 ( .A(A[471]), .B(n199), .Z(O[471]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[471]), .B(A[471]), .Z(n200) );
  XOR U301 ( .A(A[470]), .B(n201), .Z(O[470]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[470]), .B(A[470]), .Z(n202) );
  XOR U304 ( .A(A[46]), .B(n203), .Z(O[46]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[46]), .B(A[46]), .Z(n204) );
  XOR U307 ( .A(A[469]), .B(n205), .Z(O[469]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[469]), .B(A[469]), .Z(n206) );
  XOR U310 ( .A(A[468]), .B(n207), .Z(O[468]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[468]), .B(A[468]), .Z(n208) );
  XOR U313 ( .A(A[467]), .B(n209), .Z(O[467]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[467]), .B(A[467]), .Z(n210) );
  XOR U316 ( .A(A[466]), .B(n211), .Z(O[466]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[466]), .B(A[466]), .Z(n212) );
  XOR U319 ( .A(A[465]), .B(n213), .Z(O[465]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[465]), .B(A[465]), .Z(n214) );
  XOR U322 ( .A(A[464]), .B(n215), .Z(O[464]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[464]), .B(A[464]), .Z(n216) );
  XOR U325 ( .A(A[463]), .B(n217), .Z(O[463]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[463]), .B(A[463]), .Z(n218) );
  XOR U328 ( .A(A[462]), .B(n219), .Z(O[462]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[462]), .B(A[462]), .Z(n220) );
  XOR U331 ( .A(A[461]), .B(n221), .Z(O[461]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[461]), .B(A[461]), .Z(n222) );
  XOR U334 ( .A(A[460]), .B(n223), .Z(O[460]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[460]), .B(A[460]), .Z(n224) );
  XOR U337 ( .A(A[45]), .B(n225), .Z(O[45]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[45]), .B(A[45]), .Z(n226) );
  XOR U340 ( .A(A[459]), .B(n227), .Z(O[459]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[459]), .B(A[459]), .Z(n228) );
  XOR U343 ( .A(A[458]), .B(n229), .Z(O[458]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[458]), .B(A[458]), .Z(n230) );
  XOR U346 ( .A(A[457]), .B(n231), .Z(O[457]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[457]), .B(A[457]), .Z(n232) );
  XOR U349 ( .A(A[456]), .B(n233), .Z(O[456]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[456]), .B(A[456]), .Z(n234) );
  XOR U352 ( .A(A[455]), .B(n235), .Z(O[455]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[455]), .B(A[455]), .Z(n236) );
  XOR U355 ( .A(A[454]), .B(n237), .Z(O[454]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[454]), .B(A[454]), .Z(n238) );
  XOR U358 ( .A(A[453]), .B(n239), .Z(O[453]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[453]), .B(A[453]), .Z(n240) );
  XOR U361 ( .A(A[452]), .B(n241), .Z(O[452]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[452]), .B(A[452]), .Z(n242) );
  XOR U364 ( .A(A[451]), .B(n243), .Z(O[451]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[451]), .B(A[451]), .Z(n244) );
  XOR U367 ( .A(A[450]), .B(n245), .Z(O[450]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[450]), .B(A[450]), .Z(n246) );
  XOR U370 ( .A(A[44]), .B(n247), .Z(O[44]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[44]), .B(A[44]), .Z(n248) );
  XOR U373 ( .A(A[449]), .B(n249), .Z(O[449]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[449]), .B(A[449]), .Z(n250) );
  XOR U376 ( .A(A[448]), .B(n251), .Z(O[448]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[448]), .B(A[448]), .Z(n252) );
  XOR U379 ( .A(A[447]), .B(n253), .Z(O[447]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[447]), .B(A[447]), .Z(n254) );
  XOR U382 ( .A(A[446]), .B(n255), .Z(O[446]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[446]), .B(A[446]), .Z(n256) );
  XOR U385 ( .A(A[445]), .B(n257), .Z(O[445]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[445]), .B(A[445]), .Z(n258) );
  XOR U388 ( .A(A[444]), .B(n259), .Z(O[444]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[444]), .B(A[444]), .Z(n260) );
  XOR U391 ( .A(A[443]), .B(n261), .Z(O[443]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[443]), .B(A[443]), .Z(n262) );
  XOR U394 ( .A(A[442]), .B(n263), .Z(O[442]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[442]), .B(A[442]), .Z(n264) );
  XOR U397 ( .A(A[441]), .B(n265), .Z(O[441]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[441]), .B(A[441]), .Z(n266) );
  XOR U400 ( .A(A[440]), .B(n267), .Z(O[440]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[440]), .B(A[440]), .Z(n268) );
  XOR U403 ( .A(A[43]), .B(n269), .Z(O[43]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[43]), .B(A[43]), .Z(n270) );
  XOR U406 ( .A(A[439]), .B(n271), .Z(O[439]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[439]), .B(A[439]), .Z(n272) );
  XOR U409 ( .A(A[438]), .B(n273), .Z(O[438]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[438]), .B(A[438]), .Z(n274) );
  XOR U412 ( .A(A[437]), .B(n275), .Z(O[437]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[437]), .B(A[437]), .Z(n276) );
  XOR U415 ( .A(A[436]), .B(n277), .Z(O[436]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[436]), .B(A[436]), .Z(n278) );
  XOR U418 ( .A(A[435]), .B(n279), .Z(O[435]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[435]), .B(A[435]), .Z(n280) );
  XOR U421 ( .A(A[434]), .B(n281), .Z(O[434]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[434]), .B(A[434]), .Z(n282) );
  XOR U424 ( .A(A[433]), .B(n283), .Z(O[433]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[433]), .B(A[433]), .Z(n284) );
  XOR U427 ( .A(A[432]), .B(n285), .Z(O[432]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[432]), .B(A[432]), .Z(n286) );
  XOR U430 ( .A(A[431]), .B(n287), .Z(O[431]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[431]), .B(A[431]), .Z(n288) );
  XOR U433 ( .A(A[430]), .B(n289), .Z(O[430]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[430]), .B(A[430]), .Z(n290) );
  XOR U436 ( .A(A[42]), .B(n291), .Z(O[42]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[42]), .B(A[42]), .Z(n292) );
  XOR U439 ( .A(A[429]), .B(n293), .Z(O[429]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[429]), .B(A[429]), .Z(n294) );
  XOR U442 ( .A(A[428]), .B(n295), .Z(O[428]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[428]), .B(A[428]), .Z(n296) );
  XOR U445 ( .A(A[427]), .B(n297), .Z(O[427]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[427]), .B(A[427]), .Z(n298) );
  XOR U448 ( .A(A[426]), .B(n299), .Z(O[426]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[426]), .B(A[426]), .Z(n300) );
  XOR U451 ( .A(A[425]), .B(n301), .Z(O[425]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[425]), .B(A[425]), .Z(n302) );
  XOR U454 ( .A(A[424]), .B(n303), .Z(O[424]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[424]), .B(A[424]), .Z(n304) );
  XOR U457 ( .A(A[423]), .B(n305), .Z(O[423]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[423]), .B(A[423]), .Z(n306) );
  XOR U460 ( .A(A[422]), .B(n307), .Z(O[422]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[422]), .B(A[422]), .Z(n308) );
  XOR U463 ( .A(A[421]), .B(n309), .Z(O[421]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[421]), .B(A[421]), .Z(n310) );
  XOR U466 ( .A(A[420]), .B(n311), .Z(O[420]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[420]), .B(A[420]), .Z(n312) );
  XOR U469 ( .A(A[41]), .B(n313), .Z(O[41]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[41]), .B(A[41]), .Z(n314) );
  XOR U472 ( .A(A[419]), .B(n315), .Z(O[419]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[419]), .B(A[419]), .Z(n316) );
  XOR U475 ( .A(A[418]), .B(n317), .Z(O[418]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[418]), .B(A[418]), .Z(n318) );
  XOR U478 ( .A(A[417]), .B(n319), .Z(O[417]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[417]), .B(A[417]), .Z(n320) );
  XOR U481 ( .A(A[416]), .B(n321), .Z(O[416]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[416]), .B(A[416]), .Z(n322) );
  XOR U484 ( .A(A[415]), .B(n323), .Z(O[415]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[415]), .B(A[415]), .Z(n324) );
  XOR U487 ( .A(A[414]), .B(n325), .Z(O[414]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[414]), .B(A[414]), .Z(n326) );
  XOR U490 ( .A(A[413]), .B(n327), .Z(O[413]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[413]), .B(A[413]), .Z(n328) );
  XOR U493 ( .A(A[412]), .B(n329), .Z(O[412]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[412]), .B(A[412]), .Z(n330) );
  XOR U496 ( .A(A[411]), .B(n331), .Z(O[411]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[411]), .B(A[411]), .Z(n332) );
  XOR U499 ( .A(A[410]), .B(n333), .Z(O[410]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[410]), .B(A[410]), .Z(n334) );
  XOR U502 ( .A(A[40]), .B(n335), .Z(O[40]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[40]), .B(A[40]), .Z(n336) );
  XOR U505 ( .A(A[409]), .B(n337), .Z(O[409]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[409]), .B(A[409]), .Z(n338) );
  XOR U508 ( .A(A[408]), .B(n339), .Z(O[408]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[408]), .B(A[408]), .Z(n340) );
  XOR U511 ( .A(A[407]), .B(n341), .Z(O[407]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[407]), .B(A[407]), .Z(n342) );
  XOR U514 ( .A(A[406]), .B(n343), .Z(O[406]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[406]), .B(A[406]), .Z(n344) );
  XOR U517 ( .A(A[405]), .B(n345), .Z(O[405]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[405]), .B(A[405]), .Z(n346) );
  XOR U520 ( .A(A[404]), .B(n347), .Z(O[404]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[404]), .B(A[404]), .Z(n348) );
  XOR U523 ( .A(A[403]), .B(n349), .Z(O[403]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[403]), .B(A[403]), .Z(n350) );
  XOR U526 ( .A(A[402]), .B(n351), .Z(O[402]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[402]), .B(A[402]), .Z(n352) );
  XOR U529 ( .A(A[401]), .B(n353), .Z(O[401]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[401]), .B(A[401]), .Z(n354) );
  XOR U532 ( .A(A[400]), .B(n355), .Z(O[400]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[400]), .B(A[400]), .Z(n356) );
  XOR U535 ( .A(A[3]), .B(n357), .Z(O[3]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[3]), .B(A[3]), .Z(n358) );
  XOR U538 ( .A(A[39]), .B(n359), .Z(O[39]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[39]), .B(A[39]), .Z(n360) );
  XOR U541 ( .A(A[399]), .B(n361), .Z(O[399]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[399]), .B(A[399]), .Z(n362) );
  XOR U544 ( .A(A[398]), .B(n363), .Z(O[398]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[398]), .B(A[398]), .Z(n364) );
  XOR U547 ( .A(A[397]), .B(n365), .Z(O[397]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[397]), .B(A[397]), .Z(n366) );
  XOR U550 ( .A(A[396]), .B(n367), .Z(O[396]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[396]), .B(A[396]), .Z(n368) );
  XOR U553 ( .A(A[395]), .B(n369), .Z(O[395]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[395]), .B(A[395]), .Z(n370) );
  XOR U556 ( .A(A[394]), .B(n371), .Z(O[394]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[394]), .B(A[394]), .Z(n372) );
  XOR U559 ( .A(A[393]), .B(n373), .Z(O[393]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[393]), .B(A[393]), .Z(n374) );
  XOR U562 ( .A(A[392]), .B(n375), .Z(O[392]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[392]), .B(A[392]), .Z(n376) );
  XOR U565 ( .A(A[391]), .B(n377), .Z(O[391]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[391]), .B(A[391]), .Z(n378) );
  XOR U568 ( .A(A[390]), .B(n379), .Z(O[390]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[390]), .B(A[390]), .Z(n380) );
  XOR U571 ( .A(A[38]), .B(n381), .Z(O[38]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[38]), .B(A[38]), .Z(n382) );
  XOR U574 ( .A(A[389]), .B(n383), .Z(O[389]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[389]), .B(A[389]), .Z(n384) );
  XOR U577 ( .A(A[388]), .B(n385), .Z(O[388]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[388]), .B(A[388]), .Z(n386) );
  XOR U580 ( .A(A[387]), .B(n387), .Z(O[387]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[387]), .B(A[387]), .Z(n388) );
  XOR U583 ( .A(A[386]), .B(n389), .Z(O[386]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[386]), .B(A[386]), .Z(n390) );
  XOR U586 ( .A(A[385]), .B(n391), .Z(O[385]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[385]), .B(A[385]), .Z(n392) );
  XOR U589 ( .A(A[384]), .B(n393), .Z(O[384]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[384]), .B(A[384]), .Z(n394) );
  XOR U592 ( .A(A[383]), .B(n395), .Z(O[383]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[383]), .B(A[383]), .Z(n396) );
  XOR U595 ( .A(A[382]), .B(n397), .Z(O[382]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[382]), .B(A[382]), .Z(n398) );
  XOR U598 ( .A(A[381]), .B(n399), .Z(O[381]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[381]), .B(A[381]), .Z(n400) );
  XOR U601 ( .A(A[380]), .B(n401), .Z(O[380]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[380]), .B(A[380]), .Z(n402) );
  XOR U604 ( .A(A[37]), .B(n403), .Z(O[37]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[37]), .B(A[37]), .Z(n404) );
  XOR U607 ( .A(A[379]), .B(n405), .Z(O[379]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[379]), .B(A[379]), .Z(n406) );
  XOR U610 ( .A(A[378]), .B(n407), .Z(O[378]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[378]), .B(A[378]), .Z(n408) );
  XOR U613 ( .A(A[377]), .B(n409), .Z(O[377]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[377]), .B(A[377]), .Z(n410) );
  XOR U616 ( .A(A[376]), .B(n411), .Z(O[376]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[376]), .B(A[376]), .Z(n412) );
  XOR U619 ( .A(A[375]), .B(n413), .Z(O[375]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[375]), .B(A[375]), .Z(n414) );
  XOR U622 ( .A(A[374]), .B(n415), .Z(O[374]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[374]), .B(A[374]), .Z(n416) );
  XOR U625 ( .A(A[373]), .B(n417), .Z(O[373]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[373]), .B(A[373]), .Z(n418) );
  XOR U628 ( .A(A[372]), .B(n419), .Z(O[372]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[372]), .B(A[372]), .Z(n420) );
  XOR U631 ( .A(A[371]), .B(n421), .Z(O[371]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[371]), .B(A[371]), .Z(n422) );
  XOR U634 ( .A(A[370]), .B(n423), .Z(O[370]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[370]), .B(A[370]), .Z(n424) );
  XOR U637 ( .A(A[36]), .B(n425), .Z(O[36]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[36]), .B(A[36]), .Z(n426) );
  XOR U640 ( .A(A[369]), .B(n427), .Z(O[369]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[369]), .B(A[369]), .Z(n428) );
  XOR U643 ( .A(A[368]), .B(n429), .Z(O[368]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[368]), .B(A[368]), .Z(n430) );
  XOR U646 ( .A(A[367]), .B(n431), .Z(O[367]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[367]), .B(A[367]), .Z(n432) );
  XOR U649 ( .A(A[366]), .B(n433), .Z(O[366]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[366]), .B(A[366]), .Z(n434) );
  XOR U652 ( .A(A[365]), .B(n435), .Z(O[365]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[365]), .B(A[365]), .Z(n436) );
  XOR U655 ( .A(A[364]), .B(n437), .Z(O[364]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[364]), .B(A[364]), .Z(n438) );
  XOR U658 ( .A(A[363]), .B(n439), .Z(O[363]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[363]), .B(A[363]), .Z(n440) );
  XOR U661 ( .A(A[362]), .B(n441), .Z(O[362]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[362]), .B(A[362]), .Z(n442) );
  XOR U664 ( .A(A[361]), .B(n443), .Z(O[361]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[361]), .B(A[361]), .Z(n444) );
  XOR U667 ( .A(A[360]), .B(n445), .Z(O[360]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[360]), .B(A[360]), .Z(n446) );
  XOR U670 ( .A(A[35]), .B(n447), .Z(O[35]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[35]), .B(A[35]), .Z(n448) );
  XOR U673 ( .A(A[359]), .B(n449), .Z(O[359]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[359]), .B(A[359]), .Z(n450) );
  XOR U676 ( .A(A[358]), .B(n451), .Z(O[358]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[358]), .B(A[358]), .Z(n452) );
  XOR U679 ( .A(A[357]), .B(n453), .Z(O[357]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[357]), .B(A[357]), .Z(n454) );
  XOR U682 ( .A(A[356]), .B(n455), .Z(O[356]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[356]), .B(A[356]), .Z(n456) );
  XOR U685 ( .A(A[355]), .B(n457), .Z(O[355]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[355]), .B(A[355]), .Z(n458) );
  XOR U688 ( .A(A[354]), .B(n459), .Z(O[354]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[354]), .B(A[354]), .Z(n460) );
  XOR U691 ( .A(A[353]), .B(n461), .Z(O[353]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[353]), .B(A[353]), .Z(n462) );
  XOR U694 ( .A(A[352]), .B(n463), .Z(O[352]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[352]), .B(A[352]), .Z(n464) );
  XOR U697 ( .A(A[351]), .B(n465), .Z(O[351]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[351]), .B(A[351]), .Z(n466) );
  XOR U700 ( .A(A[350]), .B(n467), .Z(O[350]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[350]), .B(A[350]), .Z(n468) );
  XOR U703 ( .A(A[34]), .B(n469), .Z(O[34]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[34]), .B(A[34]), .Z(n470) );
  XOR U706 ( .A(A[349]), .B(n471), .Z(O[349]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[349]), .B(A[349]), .Z(n472) );
  XOR U709 ( .A(A[348]), .B(n473), .Z(O[348]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[348]), .B(A[348]), .Z(n474) );
  XOR U712 ( .A(A[347]), .B(n475), .Z(O[347]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[347]), .B(A[347]), .Z(n476) );
  XOR U715 ( .A(A[346]), .B(n477), .Z(O[346]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[346]), .B(A[346]), .Z(n478) );
  XOR U718 ( .A(A[345]), .B(n479), .Z(O[345]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[345]), .B(A[345]), .Z(n480) );
  XOR U721 ( .A(A[344]), .B(n481), .Z(O[344]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[344]), .B(A[344]), .Z(n482) );
  XOR U724 ( .A(A[343]), .B(n483), .Z(O[343]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[343]), .B(A[343]), .Z(n484) );
  XOR U727 ( .A(A[342]), .B(n485), .Z(O[342]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[342]), .B(A[342]), .Z(n486) );
  XOR U730 ( .A(A[341]), .B(n487), .Z(O[341]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[341]), .B(A[341]), .Z(n488) );
  XOR U733 ( .A(A[340]), .B(n489), .Z(O[340]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[340]), .B(A[340]), .Z(n490) );
  XOR U736 ( .A(A[33]), .B(n491), .Z(O[33]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[33]), .B(A[33]), .Z(n492) );
  XOR U739 ( .A(A[339]), .B(n493), .Z(O[339]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[339]), .B(A[339]), .Z(n494) );
  XOR U742 ( .A(A[338]), .B(n495), .Z(O[338]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[338]), .B(A[338]), .Z(n496) );
  XOR U745 ( .A(A[337]), .B(n497), .Z(O[337]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[337]), .B(A[337]), .Z(n498) );
  XOR U748 ( .A(A[336]), .B(n499), .Z(O[336]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[336]), .B(A[336]), .Z(n500) );
  XOR U751 ( .A(A[335]), .B(n501), .Z(O[335]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[335]), .B(A[335]), .Z(n502) );
  XOR U754 ( .A(A[334]), .B(n503), .Z(O[334]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[334]), .B(A[334]), .Z(n504) );
  XOR U757 ( .A(A[333]), .B(n505), .Z(O[333]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[333]), .B(A[333]), .Z(n506) );
  XOR U760 ( .A(A[332]), .B(n507), .Z(O[332]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[332]), .B(A[332]), .Z(n508) );
  XOR U763 ( .A(A[331]), .B(n509), .Z(O[331]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[331]), .B(A[331]), .Z(n510) );
  XOR U766 ( .A(A[330]), .B(n511), .Z(O[330]) );
  AND U767 ( .A(S), .B(n512), .Z(n511) );
  XOR U768 ( .A(B[330]), .B(A[330]), .Z(n512) );
  XOR U769 ( .A(A[32]), .B(n513), .Z(O[32]) );
  AND U770 ( .A(S), .B(n514), .Z(n513) );
  XOR U771 ( .A(B[32]), .B(A[32]), .Z(n514) );
  XOR U772 ( .A(A[329]), .B(n515), .Z(O[329]) );
  AND U773 ( .A(S), .B(n516), .Z(n515) );
  XOR U774 ( .A(B[329]), .B(A[329]), .Z(n516) );
  XOR U775 ( .A(A[328]), .B(n517), .Z(O[328]) );
  AND U776 ( .A(S), .B(n518), .Z(n517) );
  XOR U777 ( .A(B[328]), .B(A[328]), .Z(n518) );
  XOR U778 ( .A(A[327]), .B(n519), .Z(O[327]) );
  AND U779 ( .A(S), .B(n520), .Z(n519) );
  XOR U780 ( .A(B[327]), .B(A[327]), .Z(n520) );
  XOR U781 ( .A(A[326]), .B(n521), .Z(O[326]) );
  AND U782 ( .A(S), .B(n522), .Z(n521) );
  XOR U783 ( .A(B[326]), .B(A[326]), .Z(n522) );
  XOR U784 ( .A(A[325]), .B(n523), .Z(O[325]) );
  AND U785 ( .A(S), .B(n524), .Z(n523) );
  XOR U786 ( .A(B[325]), .B(A[325]), .Z(n524) );
  XOR U787 ( .A(A[324]), .B(n525), .Z(O[324]) );
  AND U788 ( .A(S), .B(n526), .Z(n525) );
  XOR U789 ( .A(B[324]), .B(A[324]), .Z(n526) );
  XOR U790 ( .A(A[323]), .B(n527), .Z(O[323]) );
  AND U791 ( .A(S), .B(n528), .Z(n527) );
  XOR U792 ( .A(B[323]), .B(A[323]), .Z(n528) );
  XOR U793 ( .A(A[322]), .B(n529), .Z(O[322]) );
  AND U794 ( .A(S), .B(n530), .Z(n529) );
  XOR U795 ( .A(B[322]), .B(A[322]), .Z(n530) );
  XOR U796 ( .A(A[321]), .B(n531), .Z(O[321]) );
  AND U797 ( .A(S), .B(n532), .Z(n531) );
  XOR U798 ( .A(B[321]), .B(A[321]), .Z(n532) );
  XOR U799 ( .A(A[320]), .B(n533), .Z(O[320]) );
  AND U800 ( .A(S), .B(n534), .Z(n533) );
  XOR U801 ( .A(B[320]), .B(A[320]), .Z(n534) );
  XOR U802 ( .A(A[31]), .B(n535), .Z(O[31]) );
  AND U803 ( .A(S), .B(n536), .Z(n535) );
  XOR U804 ( .A(B[31]), .B(A[31]), .Z(n536) );
  XOR U805 ( .A(A[319]), .B(n537), .Z(O[319]) );
  AND U806 ( .A(S), .B(n538), .Z(n537) );
  XOR U807 ( .A(B[319]), .B(A[319]), .Z(n538) );
  XOR U808 ( .A(A[318]), .B(n539), .Z(O[318]) );
  AND U809 ( .A(S), .B(n540), .Z(n539) );
  XOR U810 ( .A(B[318]), .B(A[318]), .Z(n540) );
  XOR U811 ( .A(A[317]), .B(n541), .Z(O[317]) );
  AND U812 ( .A(S), .B(n542), .Z(n541) );
  XOR U813 ( .A(B[317]), .B(A[317]), .Z(n542) );
  XOR U814 ( .A(A[316]), .B(n543), .Z(O[316]) );
  AND U815 ( .A(S), .B(n544), .Z(n543) );
  XOR U816 ( .A(B[316]), .B(A[316]), .Z(n544) );
  XOR U817 ( .A(A[315]), .B(n545), .Z(O[315]) );
  AND U818 ( .A(S), .B(n546), .Z(n545) );
  XOR U819 ( .A(B[315]), .B(A[315]), .Z(n546) );
  XOR U820 ( .A(A[314]), .B(n547), .Z(O[314]) );
  AND U821 ( .A(S), .B(n548), .Z(n547) );
  XOR U822 ( .A(B[314]), .B(A[314]), .Z(n548) );
  XOR U823 ( .A(A[313]), .B(n549), .Z(O[313]) );
  AND U824 ( .A(S), .B(n550), .Z(n549) );
  XOR U825 ( .A(B[313]), .B(A[313]), .Z(n550) );
  XOR U826 ( .A(A[312]), .B(n551), .Z(O[312]) );
  AND U827 ( .A(S), .B(n552), .Z(n551) );
  XOR U828 ( .A(B[312]), .B(A[312]), .Z(n552) );
  XOR U829 ( .A(A[311]), .B(n553), .Z(O[311]) );
  AND U830 ( .A(S), .B(n554), .Z(n553) );
  XOR U831 ( .A(B[311]), .B(A[311]), .Z(n554) );
  XOR U832 ( .A(A[310]), .B(n555), .Z(O[310]) );
  AND U833 ( .A(S), .B(n556), .Z(n555) );
  XOR U834 ( .A(B[310]), .B(A[310]), .Z(n556) );
  XOR U835 ( .A(A[30]), .B(n557), .Z(O[30]) );
  AND U836 ( .A(S), .B(n558), .Z(n557) );
  XOR U837 ( .A(B[30]), .B(A[30]), .Z(n558) );
  XOR U838 ( .A(A[309]), .B(n559), .Z(O[309]) );
  AND U839 ( .A(S), .B(n560), .Z(n559) );
  XOR U840 ( .A(B[309]), .B(A[309]), .Z(n560) );
  XOR U841 ( .A(A[308]), .B(n561), .Z(O[308]) );
  AND U842 ( .A(S), .B(n562), .Z(n561) );
  XOR U843 ( .A(B[308]), .B(A[308]), .Z(n562) );
  XOR U844 ( .A(A[307]), .B(n563), .Z(O[307]) );
  AND U845 ( .A(S), .B(n564), .Z(n563) );
  XOR U846 ( .A(B[307]), .B(A[307]), .Z(n564) );
  XOR U847 ( .A(A[306]), .B(n565), .Z(O[306]) );
  AND U848 ( .A(S), .B(n566), .Z(n565) );
  XOR U849 ( .A(B[306]), .B(A[306]), .Z(n566) );
  XOR U850 ( .A(A[305]), .B(n567), .Z(O[305]) );
  AND U851 ( .A(S), .B(n568), .Z(n567) );
  XOR U852 ( .A(B[305]), .B(A[305]), .Z(n568) );
  XOR U853 ( .A(A[304]), .B(n569), .Z(O[304]) );
  AND U854 ( .A(S), .B(n570), .Z(n569) );
  XOR U855 ( .A(B[304]), .B(A[304]), .Z(n570) );
  XOR U856 ( .A(A[303]), .B(n571), .Z(O[303]) );
  AND U857 ( .A(S), .B(n572), .Z(n571) );
  XOR U858 ( .A(B[303]), .B(A[303]), .Z(n572) );
  XOR U859 ( .A(A[302]), .B(n573), .Z(O[302]) );
  AND U860 ( .A(S), .B(n574), .Z(n573) );
  XOR U861 ( .A(B[302]), .B(A[302]), .Z(n574) );
  XOR U862 ( .A(A[301]), .B(n575), .Z(O[301]) );
  AND U863 ( .A(S), .B(n576), .Z(n575) );
  XOR U864 ( .A(B[301]), .B(A[301]), .Z(n576) );
  XOR U865 ( .A(A[300]), .B(n577), .Z(O[300]) );
  AND U866 ( .A(S), .B(n578), .Z(n577) );
  XOR U867 ( .A(B[300]), .B(A[300]), .Z(n578) );
  XOR U868 ( .A(A[2]), .B(n579), .Z(O[2]) );
  AND U869 ( .A(S), .B(n580), .Z(n579) );
  XOR U870 ( .A(B[2]), .B(A[2]), .Z(n580) );
  XOR U871 ( .A(A[29]), .B(n581), .Z(O[29]) );
  AND U872 ( .A(S), .B(n582), .Z(n581) );
  XOR U873 ( .A(B[29]), .B(A[29]), .Z(n582) );
  XOR U874 ( .A(A[299]), .B(n583), .Z(O[299]) );
  AND U875 ( .A(S), .B(n584), .Z(n583) );
  XOR U876 ( .A(B[299]), .B(A[299]), .Z(n584) );
  XOR U877 ( .A(A[298]), .B(n585), .Z(O[298]) );
  AND U878 ( .A(S), .B(n586), .Z(n585) );
  XOR U879 ( .A(B[298]), .B(A[298]), .Z(n586) );
  XOR U880 ( .A(A[297]), .B(n587), .Z(O[297]) );
  AND U881 ( .A(S), .B(n588), .Z(n587) );
  XOR U882 ( .A(B[297]), .B(A[297]), .Z(n588) );
  XOR U883 ( .A(A[296]), .B(n589), .Z(O[296]) );
  AND U884 ( .A(S), .B(n590), .Z(n589) );
  XOR U885 ( .A(B[296]), .B(A[296]), .Z(n590) );
  XOR U886 ( .A(A[295]), .B(n591), .Z(O[295]) );
  AND U887 ( .A(S), .B(n592), .Z(n591) );
  XOR U888 ( .A(B[295]), .B(A[295]), .Z(n592) );
  XOR U889 ( .A(A[294]), .B(n593), .Z(O[294]) );
  AND U890 ( .A(S), .B(n594), .Z(n593) );
  XOR U891 ( .A(B[294]), .B(A[294]), .Z(n594) );
  XOR U892 ( .A(A[293]), .B(n595), .Z(O[293]) );
  AND U893 ( .A(S), .B(n596), .Z(n595) );
  XOR U894 ( .A(B[293]), .B(A[293]), .Z(n596) );
  XOR U895 ( .A(A[292]), .B(n597), .Z(O[292]) );
  AND U896 ( .A(S), .B(n598), .Z(n597) );
  XOR U897 ( .A(B[292]), .B(A[292]), .Z(n598) );
  XOR U898 ( .A(A[291]), .B(n599), .Z(O[291]) );
  AND U899 ( .A(S), .B(n600), .Z(n599) );
  XOR U900 ( .A(B[291]), .B(A[291]), .Z(n600) );
  XOR U901 ( .A(A[290]), .B(n601), .Z(O[290]) );
  AND U902 ( .A(S), .B(n602), .Z(n601) );
  XOR U903 ( .A(B[290]), .B(A[290]), .Z(n602) );
  XOR U904 ( .A(A[28]), .B(n603), .Z(O[28]) );
  AND U905 ( .A(S), .B(n604), .Z(n603) );
  XOR U906 ( .A(B[28]), .B(A[28]), .Z(n604) );
  XOR U907 ( .A(A[289]), .B(n605), .Z(O[289]) );
  AND U908 ( .A(S), .B(n606), .Z(n605) );
  XOR U909 ( .A(B[289]), .B(A[289]), .Z(n606) );
  XOR U910 ( .A(A[288]), .B(n607), .Z(O[288]) );
  AND U911 ( .A(S), .B(n608), .Z(n607) );
  XOR U912 ( .A(B[288]), .B(A[288]), .Z(n608) );
  XOR U913 ( .A(A[287]), .B(n609), .Z(O[287]) );
  AND U914 ( .A(S), .B(n610), .Z(n609) );
  XOR U915 ( .A(B[287]), .B(A[287]), .Z(n610) );
  XOR U916 ( .A(A[286]), .B(n611), .Z(O[286]) );
  AND U917 ( .A(S), .B(n612), .Z(n611) );
  XOR U918 ( .A(B[286]), .B(A[286]), .Z(n612) );
  XOR U919 ( .A(A[285]), .B(n613), .Z(O[285]) );
  AND U920 ( .A(S), .B(n614), .Z(n613) );
  XOR U921 ( .A(B[285]), .B(A[285]), .Z(n614) );
  XOR U922 ( .A(A[284]), .B(n615), .Z(O[284]) );
  AND U923 ( .A(S), .B(n616), .Z(n615) );
  XOR U924 ( .A(B[284]), .B(A[284]), .Z(n616) );
  XOR U925 ( .A(A[283]), .B(n617), .Z(O[283]) );
  AND U926 ( .A(S), .B(n618), .Z(n617) );
  XOR U927 ( .A(B[283]), .B(A[283]), .Z(n618) );
  XOR U928 ( .A(A[282]), .B(n619), .Z(O[282]) );
  AND U929 ( .A(S), .B(n620), .Z(n619) );
  XOR U930 ( .A(B[282]), .B(A[282]), .Z(n620) );
  XOR U931 ( .A(A[281]), .B(n621), .Z(O[281]) );
  AND U932 ( .A(S), .B(n622), .Z(n621) );
  XOR U933 ( .A(B[281]), .B(A[281]), .Z(n622) );
  XOR U934 ( .A(A[280]), .B(n623), .Z(O[280]) );
  AND U935 ( .A(S), .B(n624), .Z(n623) );
  XOR U936 ( .A(B[280]), .B(A[280]), .Z(n624) );
  XOR U937 ( .A(A[27]), .B(n625), .Z(O[27]) );
  AND U938 ( .A(S), .B(n626), .Z(n625) );
  XOR U939 ( .A(B[27]), .B(A[27]), .Z(n626) );
  XOR U940 ( .A(A[279]), .B(n627), .Z(O[279]) );
  AND U941 ( .A(S), .B(n628), .Z(n627) );
  XOR U942 ( .A(B[279]), .B(A[279]), .Z(n628) );
  XOR U943 ( .A(A[278]), .B(n629), .Z(O[278]) );
  AND U944 ( .A(S), .B(n630), .Z(n629) );
  XOR U945 ( .A(B[278]), .B(A[278]), .Z(n630) );
  XOR U946 ( .A(A[277]), .B(n631), .Z(O[277]) );
  AND U947 ( .A(S), .B(n632), .Z(n631) );
  XOR U948 ( .A(B[277]), .B(A[277]), .Z(n632) );
  XOR U949 ( .A(A[276]), .B(n633), .Z(O[276]) );
  AND U950 ( .A(S), .B(n634), .Z(n633) );
  XOR U951 ( .A(B[276]), .B(A[276]), .Z(n634) );
  XOR U952 ( .A(A[275]), .B(n635), .Z(O[275]) );
  AND U953 ( .A(S), .B(n636), .Z(n635) );
  XOR U954 ( .A(B[275]), .B(A[275]), .Z(n636) );
  XOR U955 ( .A(A[274]), .B(n637), .Z(O[274]) );
  AND U956 ( .A(S), .B(n638), .Z(n637) );
  XOR U957 ( .A(B[274]), .B(A[274]), .Z(n638) );
  XOR U958 ( .A(A[273]), .B(n639), .Z(O[273]) );
  AND U959 ( .A(S), .B(n640), .Z(n639) );
  XOR U960 ( .A(B[273]), .B(A[273]), .Z(n640) );
  XOR U961 ( .A(A[272]), .B(n641), .Z(O[272]) );
  AND U962 ( .A(S), .B(n642), .Z(n641) );
  XOR U963 ( .A(B[272]), .B(A[272]), .Z(n642) );
  XOR U964 ( .A(A[271]), .B(n643), .Z(O[271]) );
  AND U965 ( .A(S), .B(n644), .Z(n643) );
  XOR U966 ( .A(B[271]), .B(A[271]), .Z(n644) );
  XOR U967 ( .A(A[270]), .B(n645), .Z(O[270]) );
  AND U968 ( .A(S), .B(n646), .Z(n645) );
  XOR U969 ( .A(B[270]), .B(A[270]), .Z(n646) );
  XOR U970 ( .A(A[26]), .B(n647), .Z(O[26]) );
  AND U971 ( .A(S), .B(n648), .Z(n647) );
  XOR U972 ( .A(B[26]), .B(A[26]), .Z(n648) );
  XOR U973 ( .A(A[269]), .B(n649), .Z(O[269]) );
  AND U974 ( .A(S), .B(n650), .Z(n649) );
  XOR U975 ( .A(B[269]), .B(A[269]), .Z(n650) );
  XOR U976 ( .A(A[268]), .B(n651), .Z(O[268]) );
  AND U977 ( .A(S), .B(n652), .Z(n651) );
  XOR U978 ( .A(B[268]), .B(A[268]), .Z(n652) );
  XOR U979 ( .A(A[267]), .B(n653), .Z(O[267]) );
  AND U980 ( .A(S), .B(n654), .Z(n653) );
  XOR U981 ( .A(B[267]), .B(A[267]), .Z(n654) );
  XOR U982 ( .A(A[266]), .B(n655), .Z(O[266]) );
  AND U983 ( .A(S), .B(n656), .Z(n655) );
  XOR U984 ( .A(B[266]), .B(A[266]), .Z(n656) );
  XOR U985 ( .A(A[265]), .B(n657), .Z(O[265]) );
  AND U986 ( .A(S), .B(n658), .Z(n657) );
  XOR U987 ( .A(B[265]), .B(A[265]), .Z(n658) );
  XOR U988 ( .A(A[264]), .B(n659), .Z(O[264]) );
  AND U989 ( .A(S), .B(n660), .Z(n659) );
  XOR U990 ( .A(B[264]), .B(A[264]), .Z(n660) );
  XOR U991 ( .A(A[263]), .B(n661), .Z(O[263]) );
  AND U992 ( .A(S), .B(n662), .Z(n661) );
  XOR U993 ( .A(B[263]), .B(A[263]), .Z(n662) );
  XOR U994 ( .A(A[262]), .B(n663), .Z(O[262]) );
  AND U995 ( .A(S), .B(n664), .Z(n663) );
  XOR U996 ( .A(B[262]), .B(A[262]), .Z(n664) );
  XOR U997 ( .A(A[261]), .B(n665), .Z(O[261]) );
  AND U998 ( .A(S), .B(n666), .Z(n665) );
  XOR U999 ( .A(B[261]), .B(A[261]), .Z(n666) );
  XOR U1000 ( .A(A[260]), .B(n667), .Z(O[260]) );
  AND U1001 ( .A(S), .B(n668), .Z(n667) );
  XOR U1002 ( .A(B[260]), .B(A[260]), .Z(n668) );
  XOR U1003 ( .A(A[25]), .B(n669), .Z(O[25]) );
  AND U1004 ( .A(S), .B(n670), .Z(n669) );
  XOR U1005 ( .A(B[25]), .B(A[25]), .Z(n670) );
  XOR U1006 ( .A(A[259]), .B(n671), .Z(O[259]) );
  AND U1007 ( .A(S), .B(n672), .Z(n671) );
  XOR U1008 ( .A(B[259]), .B(A[259]), .Z(n672) );
  XOR U1009 ( .A(A[258]), .B(n673), .Z(O[258]) );
  AND U1010 ( .A(S), .B(n674), .Z(n673) );
  XOR U1011 ( .A(B[258]), .B(A[258]), .Z(n674) );
  XOR U1012 ( .A(A[257]), .B(n675), .Z(O[257]) );
  AND U1013 ( .A(S), .B(n676), .Z(n675) );
  XOR U1014 ( .A(B[257]), .B(A[257]), .Z(n676) );
  XOR U1015 ( .A(A[256]), .B(n677), .Z(O[256]) );
  AND U1016 ( .A(S), .B(n678), .Z(n677) );
  XOR U1017 ( .A(B[256]), .B(A[256]), .Z(n678) );
  XOR U1018 ( .A(A[255]), .B(n679), .Z(O[255]) );
  AND U1019 ( .A(S), .B(n680), .Z(n679) );
  XOR U1020 ( .A(B[255]), .B(A[255]), .Z(n680) );
  XOR U1021 ( .A(A[254]), .B(n681), .Z(O[254]) );
  AND U1022 ( .A(S), .B(n682), .Z(n681) );
  XOR U1023 ( .A(B[254]), .B(A[254]), .Z(n682) );
  XOR U1024 ( .A(A[253]), .B(n683), .Z(O[253]) );
  AND U1025 ( .A(S), .B(n684), .Z(n683) );
  XOR U1026 ( .A(B[253]), .B(A[253]), .Z(n684) );
  XOR U1027 ( .A(A[252]), .B(n685), .Z(O[252]) );
  AND U1028 ( .A(S), .B(n686), .Z(n685) );
  XOR U1029 ( .A(B[252]), .B(A[252]), .Z(n686) );
  XOR U1030 ( .A(A[251]), .B(n687), .Z(O[251]) );
  AND U1031 ( .A(S), .B(n688), .Z(n687) );
  XOR U1032 ( .A(B[251]), .B(A[251]), .Z(n688) );
  XOR U1033 ( .A(A[250]), .B(n689), .Z(O[250]) );
  AND U1034 ( .A(S), .B(n690), .Z(n689) );
  XOR U1035 ( .A(B[250]), .B(A[250]), .Z(n690) );
  XOR U1036 ( .A(A[24]), .B(n691), .Z(O[24]) );
  AND U1037 ( .A(S), .B(n692), .Z(n691) );
  XOR U1038 ( .A(B[24]), .B(A[24]), .Z(n692) );
  XOR U1039 ( .A(A[249]), .B(n693), .Z(O[249]) );
  AND U1040 ( .A(S), .B(n694), .Z(n693) );
  XOR U1041 ( .A(B[249]), .B(A[249]), .Z(n694) );
  XOR U1042 ( .A(A[248]), .B(n695), .Z(O[248]) );
  AND U1043 ( .A(S), .B(n696), .Z(n695) );
  XOR U1044 ( .A(B[248]), .B(A[248]), .Z(n696) );
  XOR U1045 ( .A(A[247]), .B(n697), .Z(O[247]) );
  AND U1046 ( .A(S), .B(n698), .Z(n697) );
  XOR U1047 ( .A(B[247]), .B(A[247]), .Z(n698) );
  XOR U1048 ( .A(A[246]), .B(n699), .Z(O[246]) );
  AND U1049 ( .A(S), .B(n700), .Z(n699) );
  XOR U1050 ( .A(B[246]), .B(A[246]), .Z(n700) );
  XOR U1051 ( .A(A[245]), .B(n701), .Z(O[245]) );
  AND U1052 ( .A(S), .B(n702), .Z(n701) );
  XOR U1053 ( .A(B[245]), .B(A[245]), .Z(n702) );
  XOR U1054 ( .A(A[244]), .B(n703), .Z(O[244]) );
  AND U1055 ( .A(S), .B(n704), .Z(n703) );
  XOR U1056 ( .A(B[244]), .B(A[244]), .Z(n704) );
  XOR U1057 ( .A(A[243]), .B(n705), .Z(O[243]) );
  AND U1058 ( .A(S), .B(n706), .Z(n705) );
  XOR U1059 ( .A(B[243]), .B(A[243]), .Z(n706) );
  XOR U1060 ( .A(A[242]), .B(n707), .Z(O[242]) );
  AND U1061 ( .A(S), .B(n708), .Z(n707) );
  XOR U1062 ( .A(B[242]), .B(A[242]), .Z(n708) );
  XOR U1063 ( .A(A[241]), .B(n709), .Z(O[241]) );
  AND U1064 ( .A(S), .B(n710), .Z(n709) );
  XOR U1065 ( .A(B[241]), .B(A[241]), .Z(n710) );
  XOR U1066 ( .A(A[240]), .B(n711), .Z(O[240]) );
  AND U1067 ( .A(S), .B(n712), .Z(n711) );
  XOR U1068 ( .A(B[240]), .B(A[240]), .Z(n712) );
  XOR U1069 ( .A(A[23]), .B(n713), .Z(O[23]) );
  AND U1070 ( .A(S), .B(n714), .Z(n713) );
  XOR U1071 ( .A(B[23]), .B(A[23]), .Z(n714) );
  XOR U1072 ( .A(A[239]), .B(n715), .Z(O[239]) );
  AND U1073 ( .A(S), .B(n716), .Z(n715) );
  XOR U1074 ( .A(B[239]), .B(A[239]), .Z(n716) );
  XOR U1075 ( .A(A[238]), .B(n717), .Z(O[238]) );
  AND U1076 ( .A(S), .B(n718), .Z(n717) );
  XOR U1077 ( .A(B[238]), .B(A[238]), .Z(n718) );
  XOR U1078 ( .A(A[237]), .B(n719), .Z(O[237]) );
  AND U1079 ( .A(S), .B(n720), .Z(n719) );
  XOR U1080 ( .A(B[237]), .B(A[237]), .Z(n720) );
  XOR U1081 ( .A(A[236]), .B(n721), .Z(O[236]) );
  AND U1082 ( .A(S), .B(n722), .Z(n721) );
  XOR U1083 ( .A(B[236]), .B(A[236]), .Z(n722) );
  XOR U1084 ( .A(A[235]), .B(n723), .Z(O[235]) );
  AND U1085 ( .A(S), .B(n724), .Z(n723) );
  XOR U1086 ( .A(B[235]), .B(A[235]), .Z(n724) );
  XOR U1087 ( .A(A[234]), .B(n725), .Z(O[234]) );
  AND U1088 ( .A(S), .B(n726), .Z(n725) );
  XOR U1089 ( .A(B[234]), .B(A[234]), .Z(n726) );
  XOR U1090 ( .A(A[233]), .B(n727), .Z(O[233]) );
  AND U1091 ( .A(S), .B(n728), .Z(n727) );
  XOR U1092 ( .A(B[233]), .B(A[233]), .Z(n728) );
  XOR U1093 ( .A(A[232]), .B(n729), .Z(O[232]) );
  AND U1094 ( .A(S), .B(n730), .Z(n729) );
  XOR U1095 ( .A(B[232]), .B(A[232]), .Z(n730) );
  XOR U1096 ( .A(A[231]), .B(n731), .Z(O[231]) );
  AND U1097 ( .A(S), .B(n732), .Z(n731) );
  XOR U1098 ( .A(B[231]), .B(A[231]), .Z(n732) );
  XOR U1099 ( .A(A[230]), .B(n733), .Z(O[230]) );
  AND U1100 ( .A(S), .B(n734), .Z(n733) );
  XOR U1101 ( .A(B[230]), .B(A[230]), .Z(n734) );
  XOR U1102 ( .A(A[22]), .B(n735), .Z(O[22]) );
  AND U1103 ( .A(S), .B(n736), .Z(n735) );
  XOR U1104 ( .A(B[22]), .B(A[22]), .Z(n736) );
  XOR U1105 ( .A(A[229]), .B(n737), .Z(O[229]) );
  AND U1106 ( .A(S), .B(n738), .Z(n737) );
  XOR U1107 ( .A(B[229]), .B(A[229]), .Z(n738) );
  XOR U1108 ( .A(A[228]), .B(n739), .Z(O[228]) );
  AND U1109 ( .A(S), .B(n740), .Z(n739) );
  XOR U1110 ( .A(B[228]), .B(A[228]), .Z(n740) );
  XOR U1111 ( .A(A[227]), .B(n741), .Z(O[227]) );
  AND U1112 ( .A(S), .B(n742), .Z(n741) );
  XOR U1113 ( .A(B[227]), .B(A[227]), .Z(n742) );
  XOR U1114 ( .A(A[226]), .B(n743), .Z(O[226]) );
  AND U1115 ( .A(S), .B(n744), .Z(n743) );
  XOR U1116 ( .A(B[226]), .B(A[226]), .Z(n744) );
  XOR U1117 ( .A(A[225]), .B(n745), .Z(O[225]) );
  AND U1118 ( .A(S), .B(n746), .Z(n745) );
  XOR U1119 ( .A(B[225]), .B(A[225]), .Z(n746) );
  XOR U1120 ( .A(A[224]), .B(n747), .Z(O[224]) );
  AND U1121 ( .A(S), .B(n748), .Z(n747) );
  XOR U1122 ( .A(B[224]), .B(A[224]), .Z(n748) );
  XOR U1123 ( .A(A[223]), .B(n749), .Z(O[223]) );
  AND U1124 ( .A(S), .B(n750), .Z(n749) );
  XOR U1125 ( .A(B[223]), .B(A[223]), .Z(n750) );
  XOR U1126 ( .A(A[222]), .B(n751), .Z(O[222]) );
  AND U1127 ( .A(S), .B(n752), .Z(n751) );
  XOR U1128 ( .A(B[222]), .B(A[222]), .Z(n752) );
  XOR U1129 ( .A(A[221]), .B(n753), .Z(O[221]) );
  AND U1130 ( .A(S), .B(n754), .Z(n753) );
  XOR U1131 ( .A(B[221]), .B(A[221]), .Z(n754) );
  XOR U1132 ( .A(A[220]), .B(n755), .Z(O[220]) );
  AND U1133 ( .A(S), .B(n756), .Z(n755) );
  XOR U1134 ( .A(B[220]), .B(A[220]), .Z(n756) );
  XOR U1135 ( .A(A[21]), .B(n757), .Z(O[21]) );
  AND U1136 ( .A(S), .B(n758), .Z(n757) );
  XOR U1137 ( .A(B[21]), .B(A[21]), .Z(n758) );
  XOR U1138 ( .A(A[219]), .B(n759), .Z(O[219]) );
  AND U1139 ( .A(S), .B(n760), .Z(n759) );
  XOR U1140 ( .A(B[219]), .B(A[219]), .Z(n760) );
  XOR U1141 ( .A(A[218]), .B(n761), .Z(O[218]) );
  AND U1142 ( .A(S), .B(n762), .Z(n761) );
  XOR U1143 ( .A(B[218]), .B(A[218]), .Z(n762) );
  XOR U1144 ( .A(A[217]), .B(n763), .Z(O[217]) );
  AND U1145 ( .A(S), .B(n764), .Z(n763) );
  XOR U1146 ( .A(B[217]), .B(A[217]), .Z(n764) );
  XOR U1147 ( .A(A[216]), .B(n765), .Z(O[216]) );
  AND U1148 ( .A(S), .B(n766), .Z(n765) );
  XOR U1149 ( .A(B[216]), .B(A[216]), .Z(n766) );
  XOR U1150 ( .A(A[215]), .B(n767), .Z(O[215]) );
  AND U1151 ( .A(S), .B(n768), .Z(n767) );
  XOR U1152 ( .A(B[215]), .B(A[215]), .Z(n768) );
  XOR U1153 ( .A(A[214]), .B(n769), .Z(O[214]) );
  AND U1154 ( .A(S), .B(n770), .Z(n769) );
  XOR U1155 ( .A(B[214]), .B(A[214]), .Z(n770) );
  XOR U1156 ( .A(A[213]), .B(n771), .Z(O[213]) );
  AND U1157 ( .A(S), .B(n772), .Z(n771) );
  XOR U1158 ( .A(B[213]), .B(A[213]), .Z(n772) );
  XOR U1159 ( .A(A[212]), .B(n773), .Z(O[212]) );
  AND U1160 ( .A(S), .B(n774), .Z(n773) );
  XOR U1161 ( .A(B[212]), .B(A[212]), .Z(n774) );
  XOR U1162 ( .A(A[211]), .B(n775), .Z(O[211]) );
  AND U1163 ( .A(S), .B(n776), .Z(n775) );
  XOR U1164 ( .A(B[211]), .B(A[211]), .Z(n776) );
  XOR U1165 ( .A(A[210]), .B(n777), .Z(O[210]) );
  AND U1166 ( .A(S), .B(n778), .Z(n777) );
  XOR U1167 ( .A(B[210]), .B(A[210]), .Z(n778) );
  XOR U1168 ( .A(A[20]), .B(n779), .Z(O[20]) );
  AND U1169 ( .A(S), .B(n780), .Z(n779) );
  XOR U1170 ( .A(B[20]), .B(A[20]), .Z(n780) );
  XOR U1171 ( .A(A[209]), .B(n781), .Z(O[209]) );
  AND U1172 ( .A(S), .B(n782), .Z(n781) );
  XOR U1173 ( .A(B[209]), .B(A[209]), .Z(n782) );
  XOR U1174 ( .A(A[208]), .B(n783), .Z(O[208]) );
  AND U1175 ( .A(S), .B(n784), .Z(n783) );
  XOR U1176 ( .A(B[208]), .B(A[208]), .Z(n784) );
  XOR U1177 ( .A(A[207]), .B(n785), .Z(O[207]) );
  AND U1178 ( .A(S), .B(n786), .Z(n785) );
  XOR U1179 ( .A(B[207]), .B(A[207]), .Z(n786) );
  XOR U1180 ( .A(A[206]), .B(n787), .Z(O[206]) );
  AND U1181 ( .A(S), .B(n788), .Z(n787) );
  XOR U1182 ( .A(B[206]), .B(A[206]), .Z(n788) );
  XOR U1183 ( .A(A[205]), .B(n789), .Z(O[205]) );
  AND U1184 ( .A(S), .B(n790), .Z(n789) );
  XOR U1185 ( .A(B[205]), .B(A[205]), .Z(n790) );
  XOR U1186 ( .A(A[204]), .B(n791), .Z(O[204]) );
  AND U1187 ( .A(S), .B(n792), .Z(n791) );
  XOR U1188 ( .A(B[204]), .B(A[204]), .Z(n792) );
  XOR U1189 ( .A(A[203]), .B(n793), .Z(O[203]) );
  AND U1190 ( .A(S), .B(n794), .Z(n793) );
  XOR U1191 ( .A(B[203]), .B(A[203]), .Z(n794) );
  XOR U1192 ( .A(A[202]), .B(n795), .Z(O[202]) );
  AND U1193 ( .A(S), .B(n796), .Z(n795) );
  XOR U1194 ( .A(B[202]), .B(A[202]), .Z(n796) );
  XOR U1195 ( .A(A[201]), .B(n797), .Z(O[201]) );
  AND U1196 ( .A(S), .B(n798), .Z(n797) );
  XOR U1197 ( .A(B[201]), .B(A[201]), .Z(n798) );
  XOR U1198 ( .A(A[200]), .B(n799), .Z(O[200]) );
  AND U1199 ( .A(S), .B(n800), .Z(n799) );
  XOR U1200 ( .A(B[200]), .B(A[200]), .Z(n800) );
  XOR U1201 ( .A(A[1]), .B(n801), .Z(O[1]) );
  AND U1202 ( .A(S), .B(n802), .Z(n801) );
  XOR U1203 ( .A(B[1]), .B(A[1]), .Z(n802) );
  XOR U1204 ( .A(A[19]), .B(n803), .Z(O[19]) );
  AND U1205 ( .A(S), .B(n804), .Z(n803) );
  XOR U1206 ( .A(B[19]), .B(A[19]), .Z(n804) );
  XOR U1207 ( .A(A[199]), .B(n805), .Z(O[199]) );
  AND U1208 ( .A(S), .B(n806), .Z(n805) );
  XOR U1209 ( .A(B[199]), .B(A[199]), .Z(n806) );
  XOR U1210 ( .A(A[198]), .B(n807), .Z(O[198]) );
  AND U1211 ( .A(S), .B(n808), .Z(n807) );
  XOR U1212 ( .A(B[198]), .B(A[198]), .Z(n808) );
  XOR U1213 ( .A(A[197]), .B(n809), .Z(O[197]) );
  AND U1214 ( .A(S), .B(n810), .Z(n809) );
  XOR U1215 ( .A(B[197]), .B(A[197]), .Z(n810) );
  XOR U1216 ( .A(A[196]), .B(n811), .Z(O[196]) );
  AND U1217 ( .A(S), .B(n812), .Z(n811) );
  XOR U1218 ( .A(B[196]), .B(A[196]), .Z(n812) );
  XOR U1219 ( .A(A[195]), .B(n813), .Z(O[195]) );
  AND U1220 ( .A(S), .B(n814), .Z(n813) );
  XOR U1221 ( .A(B[195]), .B(A[195]), .Z(n814) );
  XOR U1222 ( .A(A[194]), .B(n815), .Z(O[194]) );
  AND U1223 ( .A(S), .B(n816), .Z(n815) );
  XOR U1224 ( .A(B[194]), .B(A[194]), .Z(n816) );
  XOR U1225 ( .A(A[193]), .B(n817), .Z(O[193]) );
  AND U1226 ( .A(S), .B(n818), .Z(n817) );
  XOR U1227 ( .A(B[193]), .B(A[193]), .Z(n818) );
  XOR U1228 ( .A(A[192]), .B(n819), .Z(O[192]) );
  AND U1229 ( .A(S), .B(n820), .Z(n819) );
  XOR U1230 ( .A(B[192]), .B(A[192]), .Z(n820) );
  XOR U1231 ( .A(A[191]), .B(n821), .Z(O[191]) );
  AND U1232 ( .A(S), .B(n822), .Z(n821) );
  XOR U1233 ( .A(B[191]), .B(A[191]), .Z(n822) );
  XOR U1234 ( .A(A[190]), .B(n823), .Z(O[190]) );
  AND U1235 ( .A(S), .B(n824), .Z(n823) );
  XOR U1236 ( .A(B[190]), .B(A[190]), .Z(n824) );
  XOR U1237 ( .A(A[18]), .B(n825), .Z(O[18]) );
  AND U1238 ( .A(S), .B(n826), .Z(n825) );
  XOR U1239 ( .A(B[18]), .B(A[18]), .Z(n826) );
  XOR U1240 ( .A(A[189]), .B(n827), .Z(O[189]) );
  AND U1241 ( .A(S), .B(n828), .Z(n827) );
  XOR U1242 ( .A(B[189]), .B(A[189]), .Z(n828) );
  XOR U1243 ( .A(A[188]), .B(n829), .Z(O[188]) );
  AND U1244 ( .A(S), .B(n830), .Z(n829) );
  XOR U1245 ( .A(B[188]), .B(A[188]), .Z(n830) );
  XOR U1246 ( .A(A[187]), .B(n831), .Z(O[187]) );
  AND U1247 ( .A(S), .B(n832), .Z(n831) );
  XOR U1248 ( .A(B[187]), .B(A[187]), .Z(n832) );
  XOR U1249 ( .A(A[186]), .B(n833), .Z(O[186]) );
  AND U1250 ( .A(S), .B(n834), .Z(n833) );
  XOR U1251 ( .A(B[186]), .B(A[186]), .Z(n834) );
  XOR U1252 ( .A(A[185]), .B(n835), .Z(O[185]) );
  AND U1253 ( .A(S), .B(n836), .Z(n835) );
  XOR U1254 ( .A(B[185]), .B(A[185]), .Z(n836) );
  XOR U1255 ( .A(A[184]), .B(n837), .Z(O[184]) );
  AND U1256 ( .A(S), .B(n838), .Z(n837) );
  XOR U1257 ( .A(B[184]), .B(A[184]), .Z(n838) );
  XOR U1258 ( .A(A[183]), .B(n839), .Z(O[183]) );
  AND U1259 ( .A(S), .B(n840), .Z(n839) );
  XOR U1260 ( .A(B[183]), .B(A[183]), .Z(n840) );
  XOR U1261 ( .A(A[182]), .B(n841), .Z(O[182]) );
  AND U1262 ( .A(S), .B(n842), .Z(n841) );
  XOR U1263 ( .A(B[182]), .B(A[182]), .Z(n842) );
  XOR U1264 ( .A(A[181]), .B(n843), .Z(O[181]) );
  AND U1265 ( .A(S), .B(n844), .Z(n843) );
  XOR U1266 ( .A(B[181]), .B(A[181]), .Z(n844) );
  XOR U1267 ( .A(A[180]), .B(n845), .Z(O[180]) );
  AND U1268 ( .A(S), .B(n846), .Z(n845) );
  XOR U1269 ( .A(B[180]), .B(A[180]), .Z(n846) );
  XOR U1270 ( .A(A[17]), .B(n847), .Z(O[17]) );
  AND U1271 ( .A(S), .B(n848), .Z(n847) );
  XOR U1272 ( .A(B[17]), .B(A[17]), .Z(n848) );
  XOR U1273 ( .A(A[179]), .B(n849), .Z(O[179]) );
  AND U1274 ( .A(S), .B(n850), .Z(n849) );
  XOR U1275 ( .A(B[179]), .B(A[179]), .Z(n850) );
  XOR U1276 ( .A(A[178]), .B(n851), .Z(O[178]) );
  AND U1277 ( .A(S), .B(n852), .Z(n851) );
  XOR U1278 ( .A(B[178]), .B(A[178]), .Z(n852) );
  XOR U1279 ( .A(A[177]), .B(n853), .Z(O[177]) );
  AND U1280 ( .A(S), .B(n854), .Z(n853) );
  XOR U1281 ( .A(B[177]), .B(A[177]), .Z(n854) );
  XOR U1282 ( .A(A[176]), .B(n855), .Z(O[176]) );
  AND U1283 ( .A(S), .B(n856), .Z(n855) );
  XOR U1284 ( .A(B[176]), .B(A[176]), .Z(n856) );
  XOR U1285 ( .A(A[175]), .B(n857), .Z(O[175]) );
  AND U1286 ( .A(S), .B(n858), .Z(n857) );
  XOR U1287 ( .A(B[175]), .B(A[175]), .Z(n858) );
  XOR U1288 ( .A(A[174]), .B(n859), .Z(O[174]) );
  AND U1289 ( .A(S), .B(n860), .Z(n859) );
  XOR U1290 ( .A(B[174]), .B(A[174]), .Z(n860) );
  XOR U1291 ( .A(A[173]), .B(n861), .Z(O[173]) );
  AND U1292 ( .A(S), .B(n862), .Z(n861) );
  XOR U1293 ( .A(B[173]), .B(A[173]), .Z(n862) );
  XOR U1294 ( .A(A[172]), .B(n863), .Z(O[172]) );
  AND U1295 ( .A(S), .B(n864), .Z(n863) );
  XOR U1296 ( .A(B[172]), .B(A[172]), .Z(n864) );
  XOR U1297 ( .A(A[171]), .B(n865), .Z(O[171]) );
  AND U1298 ( .A(S), .B(n866), .Z(n865) );
  XOR U1299 ( .A(B[171]), .B(A[171]), .Z(n866) );
  XOR U1300 ( .A(A[170]), .B(n867), .Z(O[170]) );
  AND U1301 ( .A(S), .B(n868), .Z(n867) );
  XOR U1302 ( .A(B[170]), .B(A[170]), .Z(n868) );
  XOR U1303 ( .A(A[16]), .B(n869), .Z(O[16]) );
  AND U1304 ( .A(S), .B(n870), .Z(n869) );
  XOR U1305 ( .A(B[16]), .B(A[16]), .Z(n870) );
  XOR U1306 ( .A(A[169]), .B(n871), .Z(O[169]) );
  AND U1307 ( .A(S), .B(n872), .Z(n871) );
  XOR U1308 ( .A(B[169]), .B(A[169]), .Z(n872) );
  XOR U1309 ( .A(A[168]), .B(n873), .Z(O[168]) );
  AND U1310 ( .A(S), .B(n874), .Z(n873) );
  XOR U1311 ( .A(B[168]), .B(A[168]), .Z(n874) );
  XOR U1312 ( .A(A[167]), .B(n875), .Z(O[167]) );
  AND U1313 ( .A(S), .B(n876), .Z(n875) );
  XOR U1314 ( .A(B[167]), .B(A[167]), .Z(n876) );
  XOR U1315 ( .A(A[166]), .B(n877), .Z(O[166]) );
  AND U1316 ( .A(S), .B(n878), .Z(n877) );
  XOR U1317 ( .A(B[166]), .B(A[166]), .Z(n878) );
  XOR U1318 ( .A(A[165]), .B(n879), .Z(O[165]) );
  AND U1319 ( .A(S), .B(n880), .Z(n879) );
  XOR U1320 ( .A(B[165]), .B(A[165]), .Z(n880) );
  XOR U1321 ( .A(A[164]), .B(n881), .Z(O[164]) );
  AND U1322 ( .A(S), .B(n882), .Z(n881) );
  XOR U1323 ( .A(B[164]), .B(A[164]), .Z(n882) );
  XOR U1324 ( .A(A[163]), .B(n883), .Z(O[163]) );
  AND U1325 ( .A(S), .B(n884), .Z(n883) );
  XOR U1326 ( .A(B[163]), .B(A[163]), .Z(n884) );
  XOR U1327 ( .A(A[162]), .B(n885), .Z(O[162]) );
  AND U1328 ( .A(S), .B(n886), .Z(n885) );
  XOR U1329 ( .A(B[162]), .B(A[162]), .Z(n886) );
  XOR U1330 ( .A(A[161]), .B(n887), .Z(O[161]) );
  AND U1331 ( .A(S), .B(n888), .Z(n887) );
  XOR U1332 ( .A(B[161]), .B(A[161]), .Z(n888) );
  XOR U1333 ( .A(A[160]), .B(n889), .Z(O[160]) );
  AND U1334 ( .A(S), .B(n890), .Z(n889) );
  XOR U1335 ( .A(B[160]), .B(A[160]), .Z(n890) );
  XOR U1336 ( .A(A[15]), .B(n891), .Z(O[15]) );
  AND U1337 ( .A(S), .B(n892), .Z(n891) );
  XOR U1338 ( .A(B[15]), .B(A[15]), .Z(n892) );
  XOR U1339 ( .A(A[159]), .B(n893), .Z(O[159]) );
  AND U1340 ( .A(S), .B(n894), .Z(n893) );
  XOR U1341 ( .A(B[159]), .B(A[159]), .Z(n894) );
  XOR U1342 ( .A(A[158]), .B(n895), .Z(O[158]) );
  AND U1343 ( .A(S), .B(n896), .Z(n895) );
  XOR U1344 ( .A(B[158]), .B(A[158]), .Z(n896) );
  XOR U1345 ( .A(A[157]), .B(n897), .Z(O[157]) );
  AND U1346 ( .A(S), .B(n898), .Z(n897) );
  XOR U1347 ( .A(B[157]), .B(A[157]), .Z(n898) );
  XOR U1348 ( .A(A[156]), .B(n899), .Z(O[156]) );
  AND U1349 ( .A(S), .B(n900), .Z(n899) );
  XOR U1350 ( .A(B[156]), .B(A[156]), .Z(n900) );
  XOR U1351 ( .A(A[155]), .B(n901), .Z(O[155]) );
  AND U1352 ( .A(S), .B(n902), .Z(n901) );
  XOR U1353 ( .A(B[155]), .B(A[155]), .Z(n902) );
  XOR U1354 ( .A(A[154]), .B(n903), .Z(O[154]) );
  AND U1355 ( .A(S), .B(n904), .Z(n903) );
  XOR U1356 ( .A(B[154]), .B(A[154]), .Z(n904) );
  XOR U1357 ( .A(A[153]), .B(n905), .Z(O[153]) );
  AND U1358 ( .A(S), .B(n906), .Z(n905) );
  XOR U1359 ( .A(B[153]), .B(A[153]), .Z(n906) );
  XOR U1360 ( .A(A[152]), .B(n907), .Z(O[152]) );
  AND U1361 ( .A(S), .B(n908), .Z(n907) );
  XOR U1362 ( .A(B[152]), .B(A[152]), .Z(n908) );
  XOR U1363 ( .A(A[151]), .B(n909), .Z(O[151]) );
  AND U1364 ( .A(S), .B(n910), .Z(n909) );
  XOR U1365 ( .A(B[151]), .B(A[151]), .Z(n910) );
  XOR U1366 ( .A(A[150]), .B(n911), .Z(O[150]) );
  AND U1367 ( .A(S), .B(n912), .Z(n911) );
  XOR U1368 ( .A(B[150]), .B(A[150]), .Z(n912) );
  XOR U1369 ( .A(A[14]), .B(n913), .Z(O[14]) );
  AND U1370 ( .A(S), .B(n914), .Z(n913) );
  XOR U1371 ( .A(B[14]), .B(A[14]), .Z(n914) );
  XOR U1372 ( .A(A[149]), .B(n915), .Z(O[149]) );
  AND U1373 ( .A(S), .B(n916), .Z(n915) );
  XOR U1374 ( .A(B[149]), .B(A[149]), .Z(n916) );
  XOR U1375 ( .A(A[148]), .B(n917), .Z(O[148]) );
  AND U1376 ( .A(S), .B(n918), .Z(n917) );
  XOR U1377 ( .A(B[148]), .B(A[148]), .Z(n918) );
  XOR U1378 ( .A(A[147]), .B(n919), .Z(O[147]) );
  AND U1379 ( .A(S), .B(n920), .Z(n919) );
  XOR U1380 ( .A(B[147]), .B(A[147]), .Z(n920) );
  XOR U1381 ( .A(A[146]), .B(n921), .Z(O[146]) );
  AND U1382 ( .A(S), .B(n922), .Z(n921) );
  XOR U1383 ( .A(B[146]), .B(A[146]), .Z(n922) );
  XOR U1384 ( .A(A[145]), .B(n923), .Z(O[145]) );
  AND U1385 ( .A(S), .B(n924), .Z(n923) );
  XOR U1386 ( .A(B[145]), .B(A[145]), .Z(n924) );
  XOR U1387 ( .A(A[144]), .B(n925), .Z(O[144]) );
  AND U1388 ( .A(S), .B(n926), .Z(n925) );
  XOR U1389 ( .A(B[144]), .B(A[144]), .Z(n926) );
  XOR U1390 ( .A(A[143]), .B(n927), .Z(O[143]) );
  AND U1391 ( .A(S), .B(n928), .Z(n927) );
  XOR U1392 ( .A(B[143]), .B(A[143]), .Z(n928) );
  XOR U1393 ( .A(A[142]), .B(n929), .Z(O[142]) );
  AND U1394 ( .A(S), .B(n930), .Z(n929) );
  XOR U1395 ( .A(B[142]), .B(A[142]), .Z(n930) );
  XOR U1396 ( .A(A[141]), .B(n931), .Z(O[141]) );
  AND U1397 ( .A(S), .B(n932), .Z(n931) );
  XOR U1398 ( .A(B[141]), .B(A[141]), .Z(n932) );
  XOR U1399 ( .A(A[140]), .B(n933), .Z(O[140]) );
  AND U1400 ( .A(S), .B(n934), .Z(n933) );
  XOR U1401 ( .A(B[140]), .B(A[140]), .Z(n934) );
  XOR U1402 ( .A(A[13]), .B(n935), .Z(O[13]) );
  AND U1403 ( .A(S), .B(n936), .Z(n935) );
  XOR U1404 ( .A(B[13]), .B(A[13]), .Z(n936) );
  XOR U1405 ( .A(A[139]), .B(n937), .Z(O[139]) );
  AND U1406 ( .A(S), .B(n938), .Z(n937) );
  XOR U1407 ( .A(B[139]), .B(A[139]), .Z(n938) );
  XOR U1408 ( .A(A[138]), .B(n939), .Z(O[138]) );
  AND U1409 ( .A(S), .B(n940), .Z(n939) );
  XOR U1410 ( .A(B[138]), .B(A[138]), .Z(n940) );
  XOR U1411 ( .A(A[137]), .B(n941), .Z(O[137]) );
  AND U1412 ( .A(S), .B(n942), .Z(n941) );
  XOR U1413 ( .A(B[137]), .B(A[137]), .Z(n942) );
  XOR U1414 ( .A(A[136]), .B(n943), .Z(O[136]) );
  AND U1415 ( .A(S), .B(n944), .Z(n943) );
  XOR U1416 ( .A(B[136]), .B(A[136]), .Z(n944) );
  XOR U1417 ( .A(A[135]), .B(n945), .Z(O[135]) );
  AND U1418 ( .A(S), .B(n946), .Z(n945) );
  XOR U1419 ( .A(B[135]), .B(A[135]), .Z(n946) );
  XOR U1420 ( .A(A[134]), .B(n947), .Z(O[134]) );
  AND U1421 ( .A(S), .B(n948), .Z(n947) );
  XOR U1422 ( .A(B[134]), .B(A[134]), .Z(n948) );
  XOR U1423 ( .A(A[133]), .B(n949), .Z(O[133]) );
  AND U1424 ( .A(S), .B(n950), .Z(n949) );
  XOR U1425 ( .A(B[133]), .B(A[133]), .Z(n950) );
  XOR U1426 ( .A(A[132]), .B(n951), .Z(O[132]) );
  AND U1427 ( .A(S), .B(n952), .Z(n951) );
  XOR U1428 ( .A(B[132]), .B(A[132]), .Z(n952) );
  XOR U1429 ( .A(A[131]), .B(n953), .Z(O[131]) );
  AND U1430 ( .A(S), .B(n954), .Z(n953) );
  XOR U1431 ( .A(B[131]), .B(A[131]), .Z(n954) );
  XOR U1432 ( .A(A[130]), .B(n955), .Z(O[130]) );
  AND U1433 ( .A(S), .B(n956), .Z(n955) );
  XOR U1434 ( .A(B[130]), .B(A[130]), .Z(n956) );
  XOR U1435 ( .A(A[12]), .B(n957), .Z(O[12]) );
  AND U1436 ( .A(S), .B(n958), .Z(n957) );
  XOR U1437 ( .A(B[12]), .B(A[12]), .Z(n958) );
  XOR U1438 ( .A(A[129]), .B(n959), .Z(O[129]) );
  AND U1439 ( .A(S), .B(n960), .Z(n959) );
  XOR U1440 ( .A(B[129]), .B(A[129]), .Z(n960) );
  XOR U1441 ( .A(A[128]), .B(n961), .Z(O[128]) );
  AND U1442 ( .A(S), .B(n962), .Z(n961) );
  XOR U1443 ( .A(B[128]), .B(A[128]), .Z(n962) );
  XOR U1444 ( .A(A[127]), .B(n963), .Z(O[127]) );
  AND U1445 ( .A(S), .B(n964), .Z(n963) );
  XOR U1446 ( .A(B[127]), .B(A[127]), .Z(n964) );
  XOR U1447 ( .A(A[126]), .B(n965), .Z(O[126]) );
  AND U1448 ( .A(S), .B(n966), .Z(n965) );
  XOR U1449 ( .A(B[126]), .B(A[126]), .Z(n966) );
  XOR U1450 ( .A(A[125]), .B(n967), .Z(O[125]) );
  AND U1451 ( .A(S), .B(n968), .Z(n967) );
  XOR U1452 ( .A(B[125]), .B(A[125]), .Z(n968) );
  XOR U1453 ( .A(A[124]), .B(n969), .Z(O[124]) );
  AND U1454 ( .A(S), .B(n970), .Z(n969) );
  XOR U1455 ( .A(B[124]), .B(A[124]), .Z(n970) );
  XOR U1456 ( .A(A[123]), .B(n971), .Z(O[123]) );
  AND U1457 ( .A(S), .B(n972), .Z(n971) );
  XOR U1458 ( .A(B[123]), .B(A[123]), .Z(n972) );
  XOR U1459 ( .A(A[122]), .B(n973), .Z(O[122]) );
  AND U1460 ( .A(S), .B(n974), .Z(n973) );
  XOR U1461 ( .A(B[122]), .B(A[122]), .Z(n974) );
  XOR U1462 ( .A(A[121]), .B(n975), .Z(O[121]) );
  AND U1463 ( .A(S), .B(n976), .Z(n975) );
  XOR U1464 ( .A(B[121]), .B(A[121]), .Z(n976) );
  XOR U1465 ( .A(A[120]), .B(n977), .Z(O[120]) );
  AND U1466 ( .A(S), .B(n978), .Z(n977) );
  XOR U1467 ( .A(B[120]), .B(A[120]), .Z(n978) );
  XOR U1468 ( .A(A[11]), .B(n979), .Z(O[11]) );
  AND U1469 ( .A(S), .B(n980), .Z(n979) );
  XOR U1470 ( .A(B[11]), .B(A[11]), .Z(n980) );
  XOR U1471 ( .A(A[119]), .B(n981), .Z(O[119]) );
  AND U1472 ( .A(S), .B(n982), .Z(n981) );
  XOR U1473 ( .A(B[119]), .B(A[119]), .Z(n982) );
  XOR U1474 ( .A(A[118]), .B(n983), .Z(O[118]) );
  AND U1475 ( .A(S), .B(n984), .Z(n983) );
  XOR U1476 ( .A(B[118]), .B(A[118]), .Z(n984) );
  XOR U1477 ( .A(A[117]), .B(n985), .Z(O[117]) );
  AND U1478 ( .A(S), .B(n986), .Z(n985) );
  XOR U1479 ( .A(B[117]), .B(A[117]), .Z(n986) );
  XOR U1480 ( .A(A[116]), .B(n987), .Z(O[116]) );
  AND U1481 ( .A(S), .B(n988), .Z(n987) );
  XOR U1482 ( .A(B[116]), .B(A[116]), .Z(n988) );
  XOR U1483 ( .A(A[115]), .B(n989), .Z(O[115]) );
  AND U1484 ( .A(S), .B(n990), .Z(n989) );
  XOR U1485 ( .A(B[115]), .B(A[115]), .Z(n990) );
  XOR U1486 ( .A(A[114]), .B(n991), .Z(O[114]) );
  AND U1487 ( .A(S), .B(n992), .Z(n991) );
  XOR U1488 ( .A(B[114]), .B(A[114]), .Z(n992) );
  XOR U1489 ( .A(A[113]), .B(n993), .Z(O[113]) );
  AND U1490 ( .A(S), .B(n994), .Z(n993) );
  XOR U1491 ( .A(B[113]), .B(A[113]), .Z(n994) );
  XOR U1492 ( .A(A[112]), .B(n995), .Z(O[112]) );
  AND U1493 ( .A(S), .B(n996), .Z(n995) );
  XOR U1494 ( .A(B[112]), .B(A[112]), .Z(n996) );
  XOR U1495 ( .A(A[111]), .B(n997), .Z(O[111]) );
  AND U1496 ( .A(S), .B(n998), .Z(n997) );
  XOR U1497 ( .A(B[111]), .B(A[111]), .Z(n998) );
  XOR U1498 ( .A(A[110]), .B(n999), .Z(O[110]) );
  AND U1499 ( .A(S), .B(n1000), .Z(n999) );
  XOR U1500 ( .A(B[110]), .B(A[110]), .Z(n1000) );
  XOR U1501 ( .A(A[10]), .B(n1001), .Z(O[10]) );
  AND U1502 ( .A(S), .B(n1002), .Z(n1001) );
  XOR U1503 ( .A(B[10]), .B(A[10]), .Z(n1002) );
  XOR U1504 ( .A(A[109]), .B(n1003), .Z(O[109]) );
  AND U1505 ( .A(S), .B(n1004), .Z(n1003) );
  XOR U1506 ( .A(B[109]), .B(A[109]), .Z(n1004) );
  XOR U1507 ( .A(A[108]), .B(n1005), .Z(O[108]) );
  AND U1508 ( .A(S), .B(n1006), .Z(n1005) );
  XOR U1509 ( .A(B[108]), .B(A[108]), .Z(n1006) );
  XOR U1510 ( .A(A[107]), .B(n1007), .Z(O[107]) );
  AND U1511 ( .A(S), .B(n1008), .Z(n1007) );
  XOR U1512 ( .A(B[107]), .B(A[107]), .Z(n1008) );
  XOR U1513 ( .A(A[106]), .B(n1009), .Z(O[106]) );
  AND U1514 ( .A(S), .B(n1010), .Z(n1009) );
  XOR U1515 ( .A(B[106]), .B(A[106]), .Z(n1010) );
  XOR U1516 ( .A(A[105]), .B(n1011), .Z(O[105]) );
  AND U1517 ( .A(S), .B(n1012), .Z(n1011) );
  XOR U1518 ( .A(B[105]), .B(A[105]), .Z(n1012) );
  XOR U1519 ( .A(A[104]), .B(n1013), .Z(O[104]) );
  AND U1520 ( .A(S), .B(n1014), .Z(n1013) );
  XOR U1521 ( .A(B[104]), .B(A[104]), .Z(n1014) );
  XOR U1522 ( .A(A[103]), .B(n1015), .Z(O[103]) );
  AND U1523 ( .A(S), .B(n1016), .Z(n1015) );
  XOR U1524 ( .A(B[103]), .B(A[103]), .Z(n1016) );
  XOR U1525 ( .A(A[102]), .B(n1017), .Z(O[102]) );
  AND U1526 ( .A(S), .B(n1018), .Z(n1017) );
  XOR U1527 ( .A(B[102]), .B(A[102]), .Z(n1018) );
  XOR U1528 ( .A(A[101]), .B(n1019), .Z(O[101]) );
  AND U1529 ( .A(S), .B(n1020), .Z(n1019) );
  XOR U1530 ( .A(B[101]), .B(A[101]), .Z(n1020) );
  XOR U1531 ( .A(A[100]), .B(n1021), .Z(O[100]) );
  AND U1532 ( .A(S), .B(n1022), .Z(n1021) );
  XOR U1533 ( .A(B[100]), .B(A[100]), .Z(n1022) );
  XOR U1534 ( .A(A[0]), .B(n1023), .Z(O[0]) );
  AND U1535 ( .A(S), .B(n1024), .Z(n1023) );
  XOR U1536 ( .A(B[0]), .B(A[0]), .Z(n1024) );
endmodule


module MUX_N512_2 ( A, B, S, O );
  input [511:0] A;
  input [511:0] B;
  output [511:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;

  XOR U1 ( .A(B[8]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(B[8]), .Z(n2) );
  XOR U4 ( .A(B[98]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(B[98]), .Z(n4) );
  XOR U7 ( .A(B[97]), .B(n5), .Z(O[98]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[98]), .B(B[97]), .Z(n6) );
  XOR U10 ( .A(B[96]), .B(n7), .Z(O[97]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[97]), .B(B[96]), .Z(n8) );
  XOR U13 ( .A(B[95]), .B(n9), .Z(O[96]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[96]), .B(B[95]), .Z(n10) );
  XOR U16 ( .A(B[94]), .B(n11), .Z(O[95]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[95]), .B(B[94]), .Z(n12) );
  XOR U19 ( .A(B[93]), .B(n13), .Z(O[94]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[94]), .B(B[93]), .Z(n14) );
  XOR U22 ( .A(B[92]), .B(n15), .Z(O[93]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[93]), .B(B[92]), .Z(n16) );
  XOR U25 ( .A(B[91]), .B(n17), .Z(O[92]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[92]), .B(B[91]), .Z(n18) );
  XOR U28 ( .A(B[90]), .B(n19), .Z(O[91]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[91]), .B(B[90]), .Z(n20) );
  XOR U31 ( .A(B[89]), .B(n21), .Z(O[90]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[90]), .B(B[89]), .Z(n22) );
  XOR U34 ( .A(B[7]), .B(n23), .Z(O[8]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[8]), .B(B[7]), .Z(n24) );
  XOR U37 ( .A(B[88]), .B(n25), .Z(O[89]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[89]), .B(B[88]), .Z(n26) );
  XOR U40 ( .A(B[87]), .B(n27), .Z(O[88]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[88]), .B(B[87]), .Z(n28) );
  XOR U43 ( .A(B[86]), .B(n29), .Z(O[87]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[87]), .B(B[86]), .Z(n30) );
  XOR U46 ( .A(B[85]), .B(n31), .Z(O[86]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[86]), .B(B[85]), .Z(n32) );
  XOR U49 ( .A(B[84]), .B(n33), .Z(O[85]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[85]), .B(B[84]), .Z(n34) );
  XOR U52 ( .A(B[83]), .B(n35), .Z(O[84]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[84]), .B(B[83]), .Z(n36) );
  XOR U55 ( .A(B[82]), .B(n37), .Z(O[83]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[83]), .B(B[82]), .Z(n38) );
  XOR U58 ( .A(B[81]), .B(n39), .Z(O[82]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[82]), .B(B[81]), .Z(n40) );
  XOR U61 ( .A(B[80]), .B(n41), .Z(O[81]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[81]), .B(B[80]), .Z(n42) );
  XOR U64 ( .A(B[79]), .B(n43), .Z(O[80]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[80]), .B(B[79]), .Z(n44) );
  XOR U67 ( .A(B[6]), .B(n45), .Z(O[7]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[7]), .B(B[6]), .Z(n46) );
  XOR U70 ( .A(B[78]), .B(n47), .Z(O[79]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[79]), .B(B[78]), .Z(n48) );
  XOR U73 ( .A(B[77]), .B(n49), .Z(O[78]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[78]), .B(B[77]), .Z(n50) );
  XOR U76 ( .A(B[76]), .B(n51), .Z(O[77]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[77]), .B(B[76]), .Z(n52) );
  XOR U79 ( .A(B[75]), .B(n53), .Z(O[76]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[76]), .B(B[75]), .Z(n54) );
  XOR U82 ( .A(B[74]), .B(n55), .Z(O[75]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[75]), .B(B[74]), .Z(n56) );
  XOR U85 ( .A(B[73]), .B(n57), .Z(O[74]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[74]), .B(B[73]), .Z(n58) );
  XOR U88 ( .A(B[72]), .B(n59), .Z(O[73]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[73]), .B(B[72]), .Z(n60) );
  XOR U91 ( .A(B[71]), .B(n61), .Z(O[72]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[72]), .B(B[71]), .Z(n62) );
  XOR U94 ( .A(B[70]), .B(n63), .Z(O[71]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[71]), .B(B[70]), .Z(n64) );
  XOR U97 ( .A(B[69]), .B(n65), .Z(O[70]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[70]), .B(B[69]), .Z(n66) );
  XOR U100 ( .A(B[5]), .B(n67), .Z(O[6]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[6]), .B(B[5]), .Z(n68) );
  XOR U103 ( .A(B[68]), .B(n69), .Z(O[69]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[69]), .B(B[68]), .Z(n70) );
  XOR U106 ( .A(B[67]), .B(n71), .Z(O[68]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[68]), .B(B[67]), .Z(n72) );
  XOR U109 ( .A(B[66]), .B(n73), .Z(O[67]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[67]), .B(B[66]), .Z(n74) );
  XOR U112 ( .A(B[65]), .B(n75), .Z(O[66]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[66]), .B(B[65]), .Z(n76) );
  XOR U115 ( .A(B[64]), .B(n77), .Z(O[65]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[65]), .B(B[64]), .Z(n78) );
  XOR U118 ( .A(B[63]), .B(n79), .Z(O[64]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[64]), .B(B[63]), .Z(n80) );
  XOR U121 ( .A(B[62]), .B(n81), .Z(O[63]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[63]), .B(B[62]), .Z(n82) );
  XOR U124 ( .A(B[61]), .B(n83), .Z(O[62]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[62]), .B(B[61]), .Z(n84) );
  XOR U127 ( .A(B[60]), .B(n85), .Z(O[61]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[61]), .B(B[60]), .Z(n86) );
  XOR U130 ( .A(B[59]), .B(n87), .Z(O[60]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[60]), .B(B[59]), .Z(n88) );
  XOR U133 ( .A(B[4]), .B(n89), .Z(O[5]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[5]), .B(B[4]), .Z(n90) );
  XOR U136 ( .A(B[58]), .B(n91), .Z(O[59]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[59]), .B(B[58]), .Z(n92) );
  XOR U139 ( .A(B[57]), .B(n93), .Z(O[58]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[58]), .B(B[57]), .Z(n94) );
  XOR U142 ( .A(B[56]), .B(n95), .Z(O[57]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[57]), .B(B[56]), .Z(n96) );
  XOR U145 ( .A(B[55]), .B(n97), .Z(O[56]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[56]), .B(B[55]), .Z(n98) );
  XOR U148 ( .A(B[54]), .B(n99), .Z(O[55]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[55]), .B(B[54]), .Z(n100) );
  XOR U151 ( .A(B[53]), .B(n101), .Z(O[54]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[54]), .B(B[53]), .Z(n102) );
  XOR U154 ( .A(B[52]), .B(n103), .Z(O[53]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[53]), .B(B[52]), .Z(n104) );
  XOR U157 ( .A(B[51]), .B(n105), .Z(O[52]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[52]), .B(B[51]), .Z(n106) );
  XOR U160 ( .A(B[50]), .B(n107), .Z(O[51]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[51]), .B(B[50]), .Z(n108) );
  XOR U163 ( .A(B[510]), .B(n109), .Z(O[511]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[511]), .B(B[510]), .Z(n110) );
  XOR U166 ( .A(B[509]), .B(n111), .Z(O[510]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[510]), .B(B[509]), .Z(n112) );
  XOR U169 ( .A(B[49]), .B(n113), .Z(O[50]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[50]), .B(B[49]), .Z(n114) );
  XOR U172 ( .A(B[508]), .B(n115), .Z(O[509]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[509]), .B(B[508]), .Z(n116) );
  XOR U175 ( .A(B[507]), .B(n117), .Z(O[508]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[508]), .B(B[507]), .Z(n118) );
  XOR U178 ( .A(B[506]), .B(n119), .Z(O[507]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[507]), .B(B[506]), .Z(n120) );
  XOR U181 ( .A(B[505]), .B(n121), .Z(O[506]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[506]), .B(B[505]), .Z(n122) );
  XOR U184 ( .A(B[504]), .B(n123), .Z(O[505]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[505]), .B(B[504]), .Z(n124) );
  XOR U187 ( .A(B[503]), .B(n125), .Z(O[504]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[504]), .B(B[503]), .Z(n126) );
  XOR U190 ( .A(B[502]), .B(n127), .Z(O[503]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[503]), .B(B[502]), .Z(n128) );
  XOR U193 ( .A(B[501]), .B(n129), .Z(O[502]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[502]), .B(B[501]), .Z(n130) );
  XOR U196 ( .A(B[500]), .B(n131), .Z(O[501]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[501]), .B(B[500]), .Z(n132) );
  XOR U199 ( .A(B[499]), .B(n133), .Z(O[500]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[500]), .B(B[499]), .Z(n134) );
  XOR U202 ( .A(B[3]), .B(n135), .Z(O[4]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[4]), .B(B[3]), .Z(n136) );
  XOR U205 ( .A(B[48]), .B(n137), .Z(O[49]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[49]), .B(B[48]), .Z(n138) );
  XOR U208 ( .A(B[498]), .B(n139), .Z(O[499]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[499]), .B(B[498]), .Z(n140) );
  XOR U211 ( .A(B[497]), .B(n141), .Z(O[498]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[498]), .B(B[497]), .Z(n142) );
  XOR U214 ( .A(B[496]), .B(n143), .Z(O[497]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[497]), .B(B[496]), .Z(n144) );
  XOR U217 ( .A(B[495]), .B(n145), .Z(O[496]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[496]), .B(B[495]), .Z(n146) );
  XOR U220 ( .A(B[494]), .B(n147), .Z(O[495]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[495]), .B(B[494]), .Z(n148) );
  XOR U223 ( .A(B[493]), .B(n149), .Z(O[494]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[494]), .B(B[493]), .Z(n150) );
  XOR U226 ( .A(B[492]), .B(n151), .Z(O[493]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[493]), .B(B[492]), .Z(n152) );
  XOR U229 ( .A(B[491]), .B(n153), .Z(O[492]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[492]), .B(B[491]), .Z(n154) );
  XOR U232 ( .A(B[490]), .B(n155), .Z(O[491]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[491]), .B(B[490]), .Z(n156) );
  XOR U235 ( .A(B[489]), .B(n157), .Z(O[490]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[490]), .B(B[489]), .Z(n158) );
  XOR U238 ( .A(B[47]), .B(n159), .Z(O[48]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[48]), .B(B[47]), .Z(n160) );
  XOR U241 ( .A(B[488]), .B(n161), .Z(O[489]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[489]), .B(B[488]), .Z(n162) );
  XOR U244 ( .A(B[487]), .B(n163), .Z(O[488]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[488]), .B(B[487]), .Z(n164) );
  XOR U247 ( .A(B[486]), .B(n165), .Z(O[487]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[487]), .B(B[486]), .Z(n166) );
  XOR U250 ( .A(B[485]), .B(n167), .Z(O[486]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[486]), .B(B[485]), .Z(n168) );
  XOR U253 ( .A(B[484]), .B(n169), .Z(O[485]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[485]), .B(B[484]), .Z(n170) );
  XOR U256 ( .A(B[483]), .B(n171), .Z(O[484]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[484]), .B(B[483]), .Z(n172) );
  XOR U259 ( .A(B[482]), .B(n173), .Z(O[483]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[483]), .B(B[482]), .Z(n174) );
  XOR U262 ( .A(B[481]), .B(n175), .Z(O[482]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[482]), .B(B[481]), .Z(n176) );
  XOR U265 ( .A(B[480]), .B(n177), .Z(O[481]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[481]), .B(B[480]), .Z(n178) );
  XOR U268 ( .A(B[479]), .B(n179), .Z(O[480]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[480]), .B(B[479]), .Z(n180) );
  XOR U271 ( .A(B[46]), .B(n181), .Z(O[47]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[47]), .B(B[46]), .Z(n182) );
  XOR U274 ( .A(B[478]), .B(n183), .Z(O[479]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[479]), .B(B[478]), .Z(n184) );
  XOR U277 ( .A(B[477]), .B(n185), .Z(O[478]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[478]), .B(B[477]), .Z(n186) );
  XOR U280 ( .A(B[476]), .B(n187), .Z(O[477]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[477]), .B(B[476]), .Z(n188) );
  XOR U283 ( .A(B[475]), .B(n189), .Z(O[476]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[476]), .B(B[475]), .Z(n190) );
  XOR U286 ( .A(B[474]), .B(n191), .Z(O[475]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[475]), .B(B[474]), .Z(n192) );
  XOR U289 ( .A(B[473]), .B(n193), .Z(O[474]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[474]), .B(B[473]), .Z(n194) );
  XOR U292 ( .A(B[472]), .B(n195), .Z(O[473]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[473]), .B(B[472]), .Z(n196) );
  XOR U295 ( .A(B[471]), .B(n197), .Z(O[472]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[472]), .B(B[471]), .Z(n198) );
  XOR U298 ( .A(B[470]), .B(n199), .Z(O[471]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[471]), .B(B[470]), .Z(n200) );
  XOR U301 ( .A(B[469]), .B(n201), .Z(O[470]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[470]), .B(B[469]), .Z(n202) );
  XOR U304 ( .A(B[45]), .B(n203), .Z(O[46]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[46]), .B(B[45]), .Z(n204) );
  XOR U307 ( .A(B[468]), .B(n205), .Z(O[469]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[469]), .B(B[468]), .Z(n206) );
  XOR U310 ( .A(B[467]), .B(n207), .Z(O[468]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[468]), .B(B[467]), .Z(n208) );
  XOR U313 ( .A(B[466]), .B(n209), .Z(O[467]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[467]), .B(B[466]), .Z(n210) );
  XOR U316 ( .A(B[465]), .B(n211), .Z(O[466]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[466]), .B(B[465]), .Z(n212) );
  XOR U319 ( .A(B[464]), .B(n213), .Z(O[465]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[465]), .B(B[464]), .Z(n214) );
  XOR U322 ( .A(B[463]), .B(n215), .Z(O[464]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[464]), .B(B[463]), .Z(n216) );
  XOR U325 ( .A(B[462]), .B(n217), .Z(O[463]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[463]), .B(B[462]), .Z(n218) );
  XOR U328 ( .A(B[461]), .B(n219), .Z(O[462]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[462]), .B(B[461]), .Z(n220) );
  XOR U331 ( .A(B[460]), .B(n221), .Z(O[461]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[461]), .B(B[460]), .Z(n222) );
  XOR U334 ( .A(B[459]), .B(n223), .Z(O[460]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[460]), .B(B[459]), .Z(n224) );
  XOR U337 ( .A(B[44]), .B(n225), .Z(O[45]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[45]), .B(B[44]), .Z(n226) );
  XOR U340 ( .A(B[458]), .B(n227), .Z(O[459]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[459]), .B(B[458]), .Z(n228) );
  XOR U343 ( .A(B[457]), .B(n229), .Z(O[458]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[458]), .B(B[457]), .Z(n230) );
  XOR U346 ( .A(B[456]), .B(n231), .Z(O[457]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[457]), .B(B[456]), .Z(n232) );
  XOR U349 ( .A(B[455]), .B(n233), .Z(O[456]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[456]), .B(B[455]), .Z(n234) );
  XOR U352 ( .A(B[454]), .B(n235), .Z(O[455]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[455]), .B(B[454]), .Z(n236) );
  XOR U355 ( .A(B[453]), .B(n237), .Z(O[454]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[454]), .B(B[453]), .Z(n238) );
  XOR U358 ( .A(B[452]), .B(n239), .Z(O[453]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[453]), .B(B[452]), .Z(n240) );
  XOR U361 ( .A(B[451]), .B(n241), .Z(O[452]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[452]), .B(B[451]), .Z(n242) );
  XOR U364 ( .A(B[450]), .B(n243), .Z(O[451]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[451]), .B(B[450]), .Z(n244) );
  XOR U367 ( .A(B[449]), .B(n245), .Z(O[450]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[450]), .B(B[449]), .Z(n246) );
  XOR U370 ( .A(B[43]), .B(n247), .Z(O[44]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[44]), .B(B[43]), .Z(n248) );
  XOR U373 ( .A(B[448]), .B(n249), .Z(O[449]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[449]), .B(B[448]), .Z(n250) );
  XOR U376 ( .A(B[447]), .B(n251), .Z(O[448]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[448]), .B(B[447]), .Z(n252) );
  XOR U379 ( .A(B[446]), .B(n253), .Z(O[447]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[447]), .B(B[446]), .Z(n254) );
  XOR U382 ( .A(B[445]), .B(n255), .Z(O[446]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[446]), .B(B[445]), .Z(n256) );
  XOR U385 ( .A(B[444]), .B(n257), .Z(O[445]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[445]), .B(B[444]), .Z(n258) );
  XOR U388 ( .A(B[443]), .B(n259), .Z(O[444]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[444]), .B(B[443]), .Z(n260) );
  XOR U391 ( .A(B[442]), .B(n261), .Z(O[443]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[443]), .B(B[442]), .Z(n262) );
  XOR U394 ( .A(B[441]), .B(n263), .Z(O[442]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[442]), .B(B[441]), .Z(n264) );
  XOR U397 ( .A(B[440]), .B(n265), .Z(O[441]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[441]), .B(B[440]), .Z(n266) );
  XOR U400 ( .A(B[439]), .B(n267), .Z(O[440]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[440]), .B(B[439]), .Z(n268) );
  XOR U403 ( .A(B[42]), .B(n269), .Z(O[43]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[43]), .B(B[42]), .Z(n270) );
  XOR U406 ( .A(B[438]), .B(n271), .Z(O[439]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[439]), .B(B[438]), .Z(n272) );
  XOR U409 ( .A(B[437]), .B(n273), .Z(O[438]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[438]), .B(B[437]), .Z(n274) );
  XOR U412 ( .A(B[436]), .B(n275), .Z(O[437]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[437]), .B(B[436]), .Z(n276) );
  XOR U415 ( .A(B[435]), .B(n277), .Z(O[436]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[436]), .B(B[435]), .Z(n278) );
  XOR U418 ( .A(B[434]), .B(n279), .Z(O[435]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[435]), .B(B[434]), .Z(n280) );
  XOR U421 ( .A(B[433]), .B(n281), .Z(O[434]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[434]), .B(B[433]), .Z(n282) );
  XOR U424 ( .A(B[432]), .B(n283), .Z(O[433]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[433]), .B(B[432]), .Z(n284) );
  XOR U427 ( .A(B[431]), .B(n285), .Z(O[432]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[432]), .B(B[431]), .Z(n286) );
  XOR U430 ( .A(B[430]), .B(n287), .Z(O[431]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[431]), .B(B[430]), .Z(n288) );
  XOR U433 ( .A(B[429]), .B(n289), .Z(O[430]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[430]), .B(B[429]), .Z(n290) );
  XOR U436 ( .A(B[41]), .B(n291), .Z(O[42]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[42]), .B(B[41]), .Z(n292) );
  XOR U439 ( .A(B[428]), .B(n293), .Z(O[429]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[429]), .B(B[428]), .Z(n294) );
  XOR U442 ( .A(B[427]), .B(n295), .Z(O[428]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[428]), .B(B[427]), .Z(n296) );
  XOR U445 ( .A(B[426]), .B(n297), .Z(O[427]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[427]), .B(B[426]), .Z(n298) );
  XOR U448 ( .A(B[425]), .B(n299), .Z(O[426]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[426]), .B(B[425]), .Z(n300) );
  XOR U451 ( .A(B[424]), .B(n301), .Z(O[425]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[425]), .B(B[424]), .Z(n302) );
  XOR U454 ( .A(B[423]), .B(n303), .Z(O[424]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[424]), .B(B[423]), .Z(n304) );
  XOR U457 ( .A(B[422]), .B(n305), .Z(O[423]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[423]), .B(B[422]), .Z(n306) );
  XOR U460 ( .A(B[421]), .B(n307), .Z(O[422]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[422]), .B(B[421]), .Z(n308) );
  XOR U463 ( .A(B[420]), .B(n309), .Z(O[421]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[421]), .B(B[420]), .Z(n310) );
  XOR U466 ( .A(B[419]), .B(n311), .Z(O[420]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[420]), .B(B[419]), .Z(n312) );
  XOR U469 ( .A(B[40]), .B(n313), .Z(O[41]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[41]), .B(B[40]), .Z(n314) );
  XOR U472 ( .A(B[418]), .B(n315), .Z(O[419]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[419]), .B(B[418]), .Z(n316) );
  XOR U475 ( .A(B[417]), .B(n317), .Z(O[418]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[418]), .B(B[417]), .Z(n318) );
  XOR U478 ( .A(B[416]), .B(n319), .Z(O[417]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[417]), .B(B[416]), .Z(n320) );
  XOR U481 ( .A(B[415]), .B(n321), .Z(O[416]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[416]), .B(B[415]), .Z(n322) );
  XOR U484 ( .A(B[414]), .B(n323), .Z(O[415]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[415]), .B(B[414]), .Z(n324) );
  XOR U487 ( .A(B[413]), .B(n325), .Z(O[414]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[414]), .B(B[413]), .Z(n326) );
  XOR U490 ( .A(B[412]), .B(n327), .Z(O[413]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[413]), .B(B[412]), .Z(n328) );
  XOR U493 ( .A(B[411]), .B(n329), .Z(O[412]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[412]), .B(B[411]), .Z(n330) );
  XOR U496 ( .A(B[410]), .B(n331), .Z(O[411]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[411]), .B(B[410]), .Z(n332) );
  XOR U499 ( .A(B[409]), .B(n333), .Z(O[410]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[410]), .B(B[409]), .Z(n334) );
  XOR U502 ( .A(B[39]), .B(n335), .Z(O[40]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[40]), .B(B[39]), .Z(n336) );
  XOR U505 ( .A(B[408]), .B(n337), .Z(O[409]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[409]), .B(B[408]), .Z(n338) );
  XOR U508 ( .A(B[407]), .B(n339), .Z(O[408]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[408]), .B(B[407]), .Z(n340) );
  XOR U511 ( .A(B[406]), .B(n341), .Z(O[407]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[407]), .B(B[406]), .Z(n342) );
  XOR U514 ( .A(B[405]), .B(n343), .Z(O[406]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[406]), .B(B[405]), .Z(n344) );
  XOR U517 ( .A(B[404]), .B(n345), .Z(O[405]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[405]), .B(B[404]), .Z(n346) );
  XOR U520 ( .A(B[403]), .B(n347), .Z(O[404]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[404]), .B(B[403]), .Z(n348) );
  XOR U523 ( .A(B[402]), .B(n349), .Z(O[403]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[403]), .B(B[402]), .Z(n350) );
  XOR U526 ( .A(B[401]), .B(n351), .Z(O[402]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[402]), .B(B[401]), .Z(n352) );
  XOR U529 ( .A(B[400]), .B(n353), .Z(O[401]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[401]), .B(B[400]), .Z(n354) );
  XOR U532 ( .A(B[399]), .B(n355), .Z(O[400]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[400]), .B(B[399]), .Z(n356) );
  XOR U535 ( .A(B[2]), .B(n357), .Z(O[3]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[3]), .B(B[2]), .Z(n358) );
  XOR U538 ( .A(B[38]), .B(n359), .Z(O[39]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[39]), .B(B[38]), .Z(n360) );
  XOR U541 ( .A(B[398]), .B(n361), .Z(O[399]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[399]), .B(B[398]), .Z(n362) );
  XOR U544 ( .A(B[397]), .B(n363), .Z(O[398]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[398]), .B(B[397]), .Z(n364) );
  XOR U547 ( .A(B[396]), .B(n365), .Z(O[397]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[397]), .B(B[396]), .Z(n366) );
  XOR U550 ( .A(B[395]), .B(n367), .Z(O[396]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[396]), .B(B[395]), .Z(n368) );
  XOR U553 ( .A(B[394]), .B(n369), .Z(O[395]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[395]), .B(B[394]), .Z(n370) );
  XOR U556 ( .A(B[393]), .B(n371), .Z(O[394]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[394]), .B(B[393]), .Z(n372) );
  XOR U559 ( .A(B[392]), .B(n373), .Z(O[393]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[393]), .B(B[392]), .Z(n374) );
  XOR U562 ( .A(B[391]), .B(n375), .Z(O[392]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[392]), .B(B[391]), .Z(n376) );
  XOR U565 ( .A(B[390]), .B(n377), .Z(O[391]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[391]), .B(B[390]), .Z(n378) );
  XOR U568 ( .A(B[389]), .B(n379), .Z(O[390]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[390]), .B(B[389]), .Z(n380) );
  XOR U571 ( .A(B[37]), .B(n381), .Z(O[38]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[38]), .B(B[37]), .Z(n382) );
  XOR U574 ( .A(B[388]), .B(n383), .Z(O[389]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[389]), .B(B[388]), .Z(n384) );
  XOR U577 ( .A(B[387]), .B(n385), .Z(O[388]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[388]), .B(B[387]), .Z(n386) );
  XOR U580 ( .A(B[386]), .B(n387), .Z(O[387]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[387]), .B(B[386]), .Z(n388) );
  XOR U583 ( .A(B[385]), .B(n389), .Z(O[386]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[386]), .B(B[385]), .Z(n390) );
  XOR U586 ( .A(B[384]), .B(n391), .Z(O[385]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[385]), .B(B[384]), .Z(n392) );
  XOR U589 ( .A(B[383]), .B(n393), .Z(O[384]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[384]), .B(B[383]), .Z(n394) );
  XOR U592 ( .A(B[382]), .B(n395), .Z(O[383]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[383]), .B(B[382]), .Z(n396) );
  XOR U595 ( .A(B[381]), .B(n397), .Z(O[382]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[382]), .B(B[381]), .Z(n398) );
  XOR U598 ( .A(B[380]), .B(n399), .Z(O[381]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[381]), .B(B[380]), .Z(n400) );
  XOR U601 ( .A(B[379]), .B(n401), .Z(O[380]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[380]), .B(B[379]), .Z(n402) );
  XOR U604 ( .A(B[36]), .B(n403), .Z(O[37]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[37]), .B(B[36]), .Z(n404) );
  XOR U607 ( .A(B[378]), .B(n405), .Z(O[379]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[379]), .B(B[378]), .Z(n406) );
  XOR U610 ( .A(B[377]), .B(n407), .Z(O[378]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[378]), .B(B[377]), .Z(n408) );
  XOR U613 ( .A(B[376]), .B(n409), .Z(O[377]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[377]), .B(B[376]), .Z(n410) );
  XOR U616 ( .A(B[375]), .B(n411), .Z(O[376]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[376]), .B(B[375]), .Z(n412) );
  XOR U619 ( .A(B[374]), .B(n413), .Z(O[375]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[375]), .B(B[374]), .Z(n414) );
  XOR U622 ( .A(B[373]), .B(n415), .Z(O[374]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[374]), .B(B[373]), .Z(n416) );
  XOR U625 ( .A(B[372]), .B(n417), .Z(O[373]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[373]), .B(B[372]), .Z(n418) );
  XOR U628 ( .A(B[371]), .B(n419), .Z(O[372]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[372]), .B(B[371]), .Z(n420) );
  XOR U631 ( .A(B[370]), .B(n421), .Z(O[371]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[371]), .B(B[370]), .Z(n422) );
  XOR U634 ( .A(B[369]), .B(n423), .Z(O[370]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[370]), .B(B[369]), .Z(n424) );
  XOR U637 ( .A(B[35]), .B(n425), .Z(O[36]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[36]), .B(B[35]), .Z(n426) );
  XOR U640 ( .A(B[368]), .B(n427), .Z(O[369]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[369]), .B(B[368]), .Z(n428) );
  XOR U643 ( .A(B[367]), .B(n429), .Z(O[368]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[368]), .B(B[367]), .Z(n430) );
  XOR U646 ( .A(B[366]), .B(n431), .Z(O[367]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[367]), .B(B[366]), .Z(n432) );
  XOR U649 ( .A(B[365]), .B(n433), .Z(O[366]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[366]), .B(B[365]), .Z(n434) );
  XOR U652 ( .A(B[364]), .B(n435), .Z(O[365]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[365]), .B(B[364]), .Z(n436) );
  XOR U655 ( .A(B[363]), .B(n437), .Z(O[364]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[364]), .B(B[363]), .Z(n438) );
  XOR U658 ( .A(B[362]), .B(n439), .Z(O[363]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[363]), .B(B[362]), .Z(n440) );
  XOR U661 ( .A(B[361]), .B(n441), .Z(O[362]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[362]), .B(B[361]), .Z(n442) );
  XOR U664 ( .A(B[360]), .B(n443), .Z(O[361]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[361]), .B(B[360]), .Z(n444) );
  XOR U667 ( .A(B[359]), .B(n445), .Z(O[360]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[360]), .B(B[359]), .Z(n446) );
  XOR U670 ( .A(B[34]), .B(n447), .Z(O[35]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[35]), .B(B[34]), .Z(n448) );
  XOR U673 ( .A(B[358]), .B(n449), .Z(O[359]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[359]), .B(B[358]), .Z(n450) );
  XOR U676 ( .A(B[357]), .B(n451), .Z(O[358]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[358]), .B(B[357]), .Z(n452) );
  XOR U679 ( .A(B[356]), .B(n453), .Z(O[357]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[357]), .B(B[356]), .Z(n454) );
  XOR U682 ( .A(B[355]), .B(n455), .Z(O[356]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[356]), .B(B[355]), .Z(n456) );
  XOR U685 ( .A(B[354]), .B(n457), .Z(O[355]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[355]), .B(B[354]), .Z(n458) );
  XOR U688 ( .A(B[353]), .B(n459), .Z(O[354]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[354]), .B(B[353]), .Z(n460) );
  XOR U691 ( .A(B[352]), .B(n461), .Z(O[353]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[353]), .B(B[352]), .Z(n462) );
  XOR U694 ( .A(B[351]), .B(n463), .Z(O[352]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[352]), .B(B[351]), .Z(n464) );
  XOR U697 ( .A(B[350]), .B(n465), .Z(O[351]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[351]), .B(B[350]), .Z(n466) );
  XOR U700 ( .A(B[349]), .B(n467), .Z(O[350]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[350]), .B(B[349]), .Z(n468) );
  XOR U703 ( .A(B[33]), .B(n469), .Z(O[34]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[34]), .B(B[33]), .Z(n470) );
  XOR U706 ( .A(B[348]), .B(n471), .Z(O[349]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[349]), .B(B[348]), .Z(n472) );
  XOR U709 ( .A(B[347]), .B(n473), .Z(O[348]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[348]), .B(B[347]), .Z(n474) );
  XOR U712 ( .A(B[346]), .B(n475), .Z(O[347]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[347]), .B(B[346]), .Z(n476) );
  XOR U715 ( .A(B[345]), .B(n477), .Z(O[346]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[346]), .B(B[345]), .Z(n478) );
  XOR U718 ( .A(B[344]), .B(n479), .Z(O[345]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[345]), .B(B[344]), .Z(n480) );
  XOR U721 ( .A(B[343]), .B(n481), .Z(O[344]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[344]), .B(B[343]), .Z(n482) );
  XOR U724 ( .A(B[342]), .B(n483), .Z(O[343]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[343]), .B(B[342]), .Z(n484) );
  XOR U727 ( .A(B[341]), .B(n485), .Z(O[342]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[342]), .B(B[341]), .Z(n486) );
  XOR U730 ( .A(B[340]), .B(n487), .Z(O[341]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[341]), .B(B[340]), .Z(n488) );
  XOR U733 ( .A(B[339]), .B(n489), .Z(O[340]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[340]), .B(B[339]), .Z(n490) );
  XOR U736 ( .A(B[32]), .B(n491), .Z(O[33]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[33]), .B(B[32]), .Z(n492) );
  XOR U739 ( .A(B[338]), .B(n493), .Z(O[339]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[339]), .B(B[338]), .Z(n494) );
  XOR U742 ( .A(B[337]), .B(n495), .Z(O[338]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[338]), .B(B[337]), .Z(n496) );
  XOR U745 ( .A(B[336]), .B(n497), .Z(O[337]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[337]), .B(B[336]), .Z(n498) );
  XOR U748 ( .A(B[335]), .B(n499), .Z(O[336]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[336]), .B(B[335]), .Z(n500) );
  XOR U751 ( .A(B[334]), .B(n501), .Z(O[335]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[335]), .B(B[334]), .Z(n502) );
  XOR U754 ( .A(B[333]), .B(n503), .Z(O[334]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[334]), .B(B[333]), .Z(n504) );
  XOR U757 ( .A(B[332]), .B(n505), .Z(O[333]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[333]), .B(B[332]), .Z(n506) );
  XOR U760 ( .A(B[331]), .B(n507), .Z(O[332]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[332]), .B(B[331]), .Z(n508) );
  XOR U763 ( .A(B[330]), .B(n509), .Z(O[331]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[331]), .B(B[330]), .Z(n510) );
  XOR U766 ( .A(B[329]), .B(n511), .Z(O[330]) );
  AND U767 ( .A(S), .B(n512), .Z(n511) );
  XOR U768 ( .A(B[330]), .B(B[329]), .Z(n512) );
  XOR U769 ( .A(B[31]), .B(n513), .Z(O[32]) );
  AND U770 ( .A(S), .B(n514), .Z(n513) );
  XOR U771 ( .A(B[32]), .B(B[31]), .Z(n514) );
  XOR U772 ( .A(B[328]), .B(n515), .Z(O[329]) );
  AND U773 ( .A(S), .B(n516), .Z(n515) );
  XOR U774 ( .A(B[329]), .B(B[328]), .Z(n516) );
  XOR U775 ( .A(B[327]), .B(n517), .Z(O[328]) );
  AND U776 ( .A(S), .B(n518), .Z(n517) );
  XOR U777 ( .A(B[328]), .B(B[327]), .Z(n518) );
  XOR U778 ( .A(B[326]), .B(n519), .Z(O[327]) );
  AND U779 ( .A(S), .B(n520), .Z(n519) );
  XOR U780 ( .A(B[327]), .B(B[326]), .Z(n520) );
  XOR U781 ( .A(B[325]), .B(n521), .Z(O[326]) );
  AND U782 ( .A(S), .B(n522), .Z(n521) );
  XOR U783 ( .A(B[326]), .B(B[325]), .Z(n522) );
  XOR U784 ( .A(B[324]), .B(n523), .Z(O[325]) );
  AND U785 ( .A(S), .B(n524), .Z(n523) );
  XOR U786 ( .A(B[325]), .B(B[324]), .Z(n524) );
  XOR U787 ( .A(B[323]), .B(n525), .Z(O[324]) );
  AND U788 ( .A(S), .B(n526), .Z(n525) );
  XOR U789 ( .A(B[324]), .B(B[323]), .Z(n526) );
  XOR U790 ( .A(B[322]), .B(n527), .Z(O[323]) );
  AND U791 ( .A(S), .B(n528), .Z(n527) );
  XOR U792 ( .A(B[323]), .B(B[322]), .Z(n528) );
  XOR U793 ( .A(B[321]), .B(n529), .Z(O[322]) );
  AND U794 ( .A(S), .B(n530), .Z(n529) );
  XOR U795 ( .A(B[322]), .B(B[321]), .Z(n530) );
  XOR U796 ( .A(B[320]), .B(n531), .Z(O[321]) );
  AND U797 ( .A(S), .B(n532), .Z(n531) );
  XOR U798 ( .A(B[321]), .B(B[320]), .Z(n532) );
  XOR U799 ( .A(B[319]), .B(n533), .Z(O[320]) );
  AND U800 ( .A(S), .B(n534), .Z(n533) );
  XOR U801 ( .A(B[320]), .B(B[319]), .Z(n534) );
  XOR U802 ( .A(B[30]), .B(n535), .Z(O[31]) );
  AND U803 ( .A(S), .B(n536), .Z(n535) );
  XOR U804 ( .A(B[31]), .B(B[30]), .Z(n536) );
  XOR U805 ( .A(B[318]), .B(n537), .Z(O[319]) );
  AND U806 ( .A(S), .B(n538), .Z(n537) );
  XOR U807 ( .A(B[319]), .B(B[318]), .Z(n538) );
  XOR U808 ( .A(B[317]), .B(n539), .Z(O[318]) );
  AND U809 ( .A(S), .B(n540), .Z(n539) );
  XOR U810 ( .A(B[318]), .B(B[317]), .Z(n540) );
  XOR U811 ( .A(B[316]), .B(n541), .Z(O[317]) );
  AND U812 ( .A(S), .B(n542), .Z(n541) );
  XOR U813 ( .A(B[317]), .B(B[316]), .Z(n542) );
  XOR U814 ( .A(B[315]), .B(n543), .Z(O[316]) );
  AND U815 ( .A(S), .B(n544), .Z(n543) );
  XOR U816 ( .A(B[316]), .B(B[315]), .Z(n544) );
  XOR U817 ( .A(B[314]), .B(n545), .Z(O[315]) );
  AND U818 ( .A(S), .B(n546), .Z(n545) );
  XOR U819 ( .A(B[315]), .B(B[314]), .Z(n546) );
  XOR U820 ( .A(B[313]), .B(n547), .Z(O[314]) );
  AND U821 ( .A(S), .B(n548), .Z(n547) );
  XOR U822 ( .A(B[314]), .B(B[313]), .Z(n548) );
  XOR U823 ( .A(B[312]), .B(n549), .Z(O[313]) );
  AND U824 ( .A(S), .B(n550), .Z(n549) );
  XOR U825 ( .A(B[313]), .B(B[312]), .Z(n550) );
  XOR U826 ( .A(B[311]), .B(n551), .Z(O[312]) );
  AND U827 ( .A(S), .B(n552), .Z(n551) );
  XOR U828 ( .A(B[312]), .B(B[311]), .Z(n552) );
  XOR U829 ( .A(B[310]), .B(n553), .Z(O[311]) );
  AND U830 ( .A(S), .B(n554), .Z(n553) );
  XOR U831 ( .A(B[311]), .B(B[310]), .Z(n554) );
  XOR U832 ( .A(B[309]), .B(n555), .Z(O[310]) );
  AND U833 ( .A(S), .B(n556), .Z(n555) );
  XOR U834 ( .A(B[310]), .B(B[309]), .Z(n556) );
  XOR U835 ( .A(B[29]), .B(n557), .Z(O[30]) );
  AND U836 ( .A(S), .B(n558), .Z(n557) );
  XOR U837 ( .A(B[30]), .B(B[29]), .Z(n558) );
  XOR U838 ( .A(B[308]), .B(n559), .Z(O[309]) );
  AND U839 ( .A(S), .B(n560), .Z(n559) );
  XOR U840 ( .A(B[309]), .B(B[308]), .Z(n560) );
  XOR U841 ( .A(B[307]), .B(n561), .Z(O[308]) );
  AND U842 ( .A(S), .B(n562), .Z(n561) );
  XOR U843 ( .A(B[308]), .B(B[307]), .Z(n562) );
  XOR U844 ( .A(B[306]), .B(n563), .Z(O[307]) );
  AND U845 ( .A(S), .B(n564), .Z(n563) );
  XOR U846 ( .A(B[307]), .B(B[306]), .Z(n564) );
  XOR U847 ( .A(B[305]), .B(n565), .Z(O[306]) );
  AND U848 ( .A(S), .B(n566), .Z(n565) );
  XOR U849 ( .A(B[306]), .B(B[305]), .Z(n566) );
  XOR U850 ( .A(B[304]), .B(n567), .Z(O[305]) );
  AND U851 ( .A(S), .B(n568), .Z(n567) );
  XOR U852 ( .A(B[305]), .B(B[304]), .Z(n568) );
  XOR U853 ( .A(B[303]), .B(n569), .Z(O[304]) );
  AND U854 ( .A(S), .B(n570), .Z(n569) );
  XOR U855 ( .A(B[304]), .B(B[303]), .Z(n570) );
  XOR U856 ( .A(B[302]), .B(n571), .Z(O[303]) );
  AND U857 ( .A(S), .B(n572), .Z(n571) );
  XOR U858 ( .A(B[303]), .B(B[302]), .Z(n572) );
  XOR U859 ( .A(B[301]), .B(n573), .Z(O[302]) );
  AND U860 ( .A(S), .B(n574), .Z(n573) );
  XOR U861 ( .A(B[302]), .B(B[301]), .Z(n574) );
  XOR U862 ( .A(B[300]), .B(n575), .Z(O[301]) );
  AND U863 ( .A(S), .B(n576), .Z(n575) );
  XOR U864 ( .A(B[301]), .B(B[300]), .Z(n576) );
  XOR U865 ( .A(B[299]), .B(n577), .Z(O[300]) );
  AND U866 ( .A(S), .B(n578), .Z(n577) );
  XOR U867 ( .A(B[300]), .B(B[299]), .Z(n578) );
  XOR U868 ( .A(B[1]), .B(n579), .Z(O[2]) );
  AND U869 ( .A(S), .B(n580), .Z(n579) );
  XOR U870 ( .A(B[2]), .B(B[1]), .Z(n580) );
  XOR U871 ( .A(B[28]), .B(n581), .Z(O[29]) );
  AND U872 ( .A(S), .B(n582), .Z(n581) );
  XOR U873 ( .A(B[29]), .B(B[28]), .Z(n582) );
  XOR U874 ( .A(B[298]), .B(n583), .Z(O[299]) );
  AND U875 ( .A(S), .B(n584), .Z(n583) );
  XOR U876 ( .A(B[299]), .B(B[298]), .Z(n584) );
  XOR U877 ( .A(B[297]), .B(n585), .Z(O[298]) );
  AND U878 ( .A(S), .B(n586), .Z(n585) );
  XOR U879 ( .A(B[298]), .B(B[297]), .Z(n586) );
  XOR U880 ( .A(B[296]), .B(n587), .Z(O[297]) );
  AND U881 ( .A(S), .B(n588), .Z(n587) );
  XOR U882 ( .A(B[297]), .B(B[296]), .Z(n588) );
  XOR U883 ( .A(B[295]), .B(n589), .Z(O[296]) );
  AND U884 ( .A(S), .B(n590), .Z(n589) );
  XOR U885 ( .A(B[296]), .B(B[295]), .Z(n590) );
  XOR U886 ( .A(B[294]), .B(n591), .Z(O[295]) );
  AND U887 ( .A(S), .B(n592), .Z(n591) );
  XOR U888 ( .A(B[295]), .B(B[294]), .Z(n592) );
  XOR U889 ( .A(B[293]), .B(n593), .Z(O[294]) );
  AND U890 ( .A(S), .B(n594), .Z(n593) );
  XOR U891 ( .A(B[294]), .B(B[293]), .Z(n594) );
  XOR U892 ( .A(B[292]), .B(n595), .Z(O[293]) );
  AND U893 ( .A(S), .B(n596), .Z(n595) );
  XOR U894 ( .A(B[293]), .B(B[292]), .Z(n596) );
  XOR U895 ( .A(B[291]), .B(n597), .Z(O[292]) );
  AND U896 ( .A(S), .B(n598), .Z(n597) );
  XOR U897 ( .A(B[292]), .B(B[291]), .Z(n598) );
  XOR U898 ( .A(B[290]), .B(n599), .Z(O[291]) );
  AND U899 ( .A(S), .B(n600), .Z(n599) );
  XOR U900 ( .A(B[291]), .B(B[290]), .Z(n600) );
  XOR U901 ( .A(B[289]), .B(n601), .Z(O[290]) );
  AND U902 ( .A(S), .B(n602), .Z(n601) );
  XOR U903 ( .A(B[290]), .B(B[289]), .Z(n602) );
  XOR U904 ( .A(B[27]), .B(n603), .Z(O[28]) );
  AND U905 ( .A(S), .B(n604), .Z(n603) );
  XOR U906 ( .A(B[28]), .B(B[27]), .Z(n604) );
  XOR U907 ( .A(B[288]), .B(n605), .Z(O[289]) );
  AND U908 ( .A(S), .B(n606), .Z(n605) );
  XOR U909 ( .A(B[289]), .B(B[288]), .Z(n606) );
  XOR U910 ( .A(B[287]), .B(n607), .Z(O[288]) );
  AND U911 ( .A(S), .B(n608), .Z(n607) );
  XOR U912 ( .A(B[288]), .B(B[287]), .Z(n608) );
  XOR U913 ( .A(B[286]), .B(n609), .Z(O[287]) );
  AND U914 ( .A(S), .B(n610), .Z(n609) );
  XOR U915 ( .A(B[287]), .B(B[286]), .Z(n610) );
  XOR U916 ( .A(B[285]), .B(n611), .Z(O[286]) );
  AND U917 ( .A(S), .B(n612), .Z(n611) );
  XOR U918 ( .A(B[286]), .B(B[285]), .Z(n612) );
  XOR U919 ( .A(B[284]), .B(n613), .Z(O[285]) );
  AND U920 ( .A(S), .B(n614), .Z(n613) );
  XOR U921 ( .A(B[285]), .B(B[284]), .Z(n614) );
  XOR U922 ( .A(B[283]), .B(n615), .Z(O[284]) );
  AND U923 ( .A(S), .B(n616), .Z(n615) );
  XOR U924 ( .A(B[284]), .B(B[283]), .Z(n616) );
  XOR U925 ( .A(B[282]), .B(n617), .Z(O[283]) );
  AND U926 ( .A(S), .B(n618), .Z(n617) );
  XOR U927 ( .A(B[283]), .B(B[282]), .Z(n618) );
  XOR U928 ( .A(B[281]), .B(n619), .Z(O[282]) );
  AND U929 ( .A(S), .B(n620), .Z(n619) );
  XOR U930 ( .A(B[282]), .B(B[281]), .Z(n620) );
  XOR U931 ( .A(B[280]), .B(n621), .Z(O[281]) );
  AND U932 ( .A(S), .B(n622), .Z(n621) );
  XOR U933 ( .A(B[281]), .B(B[280]), .Z(n622) );
  XOR U934 ( .A(B[279]), .B(n623), .Z(O[280]) );
  AND U935 ( .A(S), .B(n624), .Z(n623) );
  XOR U936 ( .A(B[280]), .B(B[279]), .Z(n624) );
  XOR U937 ( .A(B[26]), .B(n625), .Z(O[27]) );
  AND U938 ( .A(S), .B(n626), .Z(n625) );
  XOR U939 ( .A(B[27]), .B(B[26]), .Z(n626) );
  XOR U940 ( .A(B[278]), .B(n627), .Z(O[279]) );
  AND U941 ( .A(S), .B(n628), .Z(n627) );
  XOR U942 ( .A(B[279]), .B(B[278]), .Z(n628) );
  XOR U943 ( .A(B[277]), .B(n629), .Z(O[278]) );
  AND U944 ( .A(S), .B(n630), .Z(n629) );
  XOR U945 ( .A(B[278]), .B(B[277]), .Z(n630) );
  XOR U946 ( .A(B[276]), .B(n631), .Z(O[277]) );
  AND U947 ( .A(S), .B(n632), .Z(n631) );
  XOR U948 ( .A(B[277]), .B(B[276]), .Z(n632) );
  XOR U949 ( .A(B[275]), .B(n633), .Z(O[276]) );
  AND U950 ( .A(S), .B(n634), .Z(n633) );
  XOR U951 ( .A(B[276]), .B(B[275]), .Z(n634) );
  XOR U952 ( .A(B[274]), .B(n635), .Z(O[275]) );
  AND U953 ( .A(S), .B(n636), .Z(n635) );
  XOR U954 ( .A(B[275]), .B(B[274]), .Z(n636) );
  XOR U955 ( .A(B[273]), .B(n637), .Z(O[274]) );
  AND U956 ( .A(S), .B(n638), .Z(n637) );
  XOR U957 ( .A(B[274]), .B(B[273]), .Z(n638) );
  XOR U958 ( .A(B[272]), .B(n639), .Z(O[273]) );
  AND U959 ( .A(S), .B(n640), .Z(n639) );
  XOR U960 ( .A(B[273]), .B(B[272]), .Z(n640) );
  XOR U961 ( .A(B[271]), .B(n641), .Z(O[272]) );
  AND U962 ( .A(S), .B(n642), .Z(n641) );
  XOR U963 ( .A(B[272]), .B(B[271]), .Z(n642) );
  XOR U964 ( .A(B[270]), .B(n643), .Z(O[271]) );
  AND U965 ( .A(S), .B(n644), .Z(n643) );
  XOR U966 ( .A(B[271]), .B(B[270]), .Z(n644) );
  XOR U967 ( .A(B[269]), .B(n645), .Z(O[270]) );
  AND U968 ( .A(S), .B(n646), .Z(n645) );
  XOR U969 ( .A(B[270]), .B(B[269]), .Z(n646) );
  XOR U970 ( .A(B[25]), .B(n647), .Z(O[26]) );
  AND U971 ( .A(S), .B(n648), .Z(n647) );
  XOR U972 ( .A(B[26]), .B(B[25]), .Z(n648) );
  XOR U973 ( .A(B[268]), .B(n649), .Z(O[269]) );
  AND U974 ( .A(S), .B(n650), .Z(n649) );
  XOR U975 ( .A(B[269]), .B(B[268]), .Z(n650) );
  XOR U976 ( .A(B[267]), .B(n651), .Z(O[268]) );
  AND U977 ( .A(S), .B(n652), .Z(n651) );
  XOR U978 ( .A(B[268]), .B(B[267]), .Z(n652) );
  XOR U979 ( .A(B[266]), .B(n653), .Z(O[267]) );
  AND U980 ( .A(S), .B(n654), .Z(n653) );
  XOR U981 ( .A(B[267]), .B(B[266]), .Z(n654) );
  XOR U982 ( .A(B[265]), .B(n655), .Z(O[266]) );
  AND U983 ( .A(S), .B(n656), .Z(n655) );
  XOR U984 ( .A(B[266]), .B(B[265]), .Z(n656) );
  XOR U985 ( .A(B[264]), .B(n657), .Z(O[265]) );
  AND U986 ( .A(S), .B(n658), .Z(n657) );
  XOR U987 ( .A(B[265]), .B(B[264]), .Z(n658) );
  XOR U988 ( .A(B[263]), .B(n659), .Z(O[264]) );
  AND U989 ( .A(S), .B(n660), .Z(n659) );
  XOR U990 ( .A(B[264]), .B(B[263]), .Z(n660) );
  XOR U991 ( .A(B[262]), .B(n661), .Z(O[263]) );
  AND U992 ( .A(S), .B(n662), .Z(n661) );
  XOR U993 ( .A(B[263]), .B(B[262]), .Z(n662) );
  XOR U994 ( .A(B[261]), .B(n663), .Z(O[262]) );
  AND U995 ( .A(S), .B(n664), .Z(n663) );
  XOR U996 ( .A(B[262]), .B(B[261]), .Z(n664) );
  XOR U997 ( .A(B[260]), .B(n665), .Z(O[261]) );
  AND U998 ( .A(S), .B(n666), .Z(n665) );
  XOR U999 ( .A(B[261]), .B(B[260]), .Z(n666) );
  XOR U1000 ( .A(B[259]), .B(n667), .Z(O[260]) );
  AND U1001 ( .A(S), .B(n668), .Z(n667) );
  XOR U1002 ( .A(B[260]), .B(B[259]), .Z(n668) );
  XOR U1003 ( .A(B[24]), .B(n669), .Z(O[25]) );
  AND U1004 ( .A(S), .B(n670), .Z(n669) );
  XOR U1005 ( .A(B[25]), .B(B[24]), .Z(n670) );
  XOR U1006 ( .A(B[258]), .B(n671), .Z(O[259]) );
  AND U1007 ( .A(S), .B(n672), .Z(n671) );
  XOR U1008 ( .A(B[259]), .B(B[258]), .Z(n672) );
  XOR U1009 ( .A(B[257]), .B(n673), .Z(O[258]) );
  AND U1010 ( .A(S), .B(n674), .Z(n673) );
  XOR U1011 ( .A(B[258]), .B(B[257]), .Z(n674) );
  XOR U1012 ( .A(B[256]), .B(n675), .Z(O[257]) );
  AND U1013 ( .A(S), .B(n676), .Z(n675) );
  XOR U1014 ( .A(B[257]), .B(B[256]), .Z(n676) );
  XOR U1015 ( .A(B[255]), .B(n677), .Z(O[256]) );
  AND U1016 ( .A(S), .B(n678), .Z(n677) );
  XOR U1017 ( .A(B[256]), .B(B[255]), .Z(n678) );
  XOR U1018 ( .A(B[254]), .B(n679), .Z(O[255]) );
  AND U1019 ( .A(S), .B(n680), .Z(n679) );
  XOR U1020 ( .A(B[255]), .B(B[254]), .Z(n680) );
  XOR U1021 ( .A(B[253]), .B(n681), .Z(O[254]) );
  AND U1022 ( .A(S), .B(n682), .Z(n681) );
  XOR U1023 ( .A(B[254]), .B(B[253]), .Z(n682) );
  XOR U1024 ( .A(B[252]), .B(n683), .Z(O[253]) );
  AND U1025 ( .A(S), .B(n684), .Z(n683) );
  XOR U1026 ( .A(B[253]), .B(B[252]), .Z(n684) );
  XOR U1027 ( .A(B[251]), .B(n685), .Z(O[252]) );
  AND U1028 ( .A(S), .B(n686), .Z(n685) );
  XOR U1029 ( .A(B[252]), .B(B[251]), .Z(n686) );
  XOR U1030 ( .A(B[250]), .B(n687), .Z(O[251]) );
  AND U1031 ( .A(S), .B(n688), .Z(n687) );
  XOR U1032 ( .A(B[251]), .B(B[250]), .Z(n688) );
  XOR U1033 ( .A(B[249]), .B(n689), .Z(O[250]) );
  AND U1034 ( .A(S), .B(n690), .Z(n689) );
  XOR U1035 ( .A(B[250]), .B(B[249]), .Z(n690) );
  XOR U1036 ( .A(B[23]), .B(n691), .Z(O[24]) );
  AND U1037 ( .A(S), .B(n692), .Z(n691) );
  XOR U1038 ( .A(B[24]), .B(B[23]), .Z(n692) );
  XOR U1039 ( .A(B[248]), .B(n693), .Z(O[249]) );
  AND U1040 ( .A(S), .B(n694), .Z(n693) );
  XOR U1041 ( .A(B[249]), .B(B[248]), .Z(n694) );
  XOR U1042 ( .A(B[247]), .B(n695), .Z(O[248]) );
  AND U1043 ( .A(S), .B(n696), .Z(n695) );
  XOR U1044 ( .A(B[248]), .B(B[247]), .Z(n696) );
  XOR U1045 ( .A(B[246]), .B(n697), .Z(O[247]) );
  AND U1046 ( .A(S), .B(n698), .Z(n697) );
  XOR U1047 ( .A(B[247]), .B(B[246]), .Z(n698) );
  XOR U1048 ( .A(B[245]), .B(n699), .Z(O[246]) );
  AND U1049 ( .A(S), .B(n700), .Z(n699) );
  XOR U1050 ( .A(B[246]), .B(B[245]), .Z(n700) );
  XOR U1051 ( .A(B[244]), .B(n701), .Z(O[245]) );
  AND U1052 ( .A(S), .B(n702), .Z(n701) );
  XOR U1053 ( .A(B[245]), .B(B[244]), .Z(n702) );
  XOR U1054 ( .A(B[243]), .B(n703), .Z(O[244]) );
  AND U1055 ( .A(S), .B(n704), .Z(n703) );
  XOR U1056 ( .A(B[244]), .B(B[243]), .Z(n704) );
  XOR U1057 ( .A(B[242]), .B(n705), .Z(O[243]) );
  AND U1058 ( .A(S), .B(n706), .Z(n705) );
  XOR U1059 ( .A(B[243]), .B(B[242]), .Z(n706) );
  XOR U1060 ( .A(B[241]), .B(n707), .Z(O[242]) );
  AND U1061 ( .A(S), .B(n708), .Z(n707) );
  XOR U1062 ( .A(B[242]), .B(B[241]), .Z(n708) );
  XOR U1063 ( .A(B[240]), .B(n709), .Z(O[241]) );
  AND U1064 ( .A(S), .B(n710), .Z(n709) );
  XOR U1065 ( .A(B[241]), .B(B[240]), .Z(n710) );
  XOR U1066 ( .A(B[239]), .B(n711), .Z(O[240]) );
  AND U1067 ( .A(S), .B(n712), .Z(n711) );
  XOR U1068 ( .A(B[240]), .B(B[239]), .Z(n712) );
  XOR U1069 ( .A(B[22]), .B(n713), .Z(O[23]) );
  AND U1070 ( .A(S), .B(n714), .Z(n713) );
  XOR U1071 ( .A(B[23]), .B(B[22]), .Z(n714) );
  XOR U1072 ( .A(B[238]), .B(n715), .Z(O[239]) );
  AND U1073 ( .A(S), .B(n716), .Z(n715) );
  XOR U1074 ( .A(B[239]), .B(B[238]), .Z(n716) );
  XOR U1075 ( .A(B[237]), .B(n717), .Z(O[238]) );
  AND U1076 ( .A(S), .B(n718), .Z(n717) );
  XOR U1077 ( .A(B[238]), .B(B[237]), .Z(n718) );
  XOR U1078 ( .A(B[236]), .B(n719), .Z(O[237]) );
  AND U1079 ( .A(S), .B(n720), .Z(n719) );
  XOR U1080 ( .A(B[237]), .B(B[236]), .Z(n720) );
  XOR U1081 ( .A(B[235]), .B(n721), .Z(O[236]) );
  AND U1082 ( .A(S), .B(n722), .Z(n721) );
  XOR U1083 ( .A(B[236]), .B(B[235]), .Z(n722) );
  XOR U1084 ( .A(B[234]), .B(n723), .Z(O[235]) );
  AND U1085 ( .A(S), .B(n724), .Z(n723) );
  XOR U1086 ( .A(B[235]), .B(B[234]), .Z(n724) );
  XOR U1087 ( .A(B[233]), .B(n725), .Z(O[234]) );
  AND U1088 ( .A(S), .B(n726), .Z(n725) );
  XOR U1089 ( .A(B[234]), .B(B[233]), .Z(n726) );
  XOR U1090 ( .A(B[232]), .B(n727), .Z(O[233]) );
  AND U1091 ( .A(S), .B(n728), .Z(n727) );
  XOR U1092 ( .A(B[233]), .B(B[232]), .Z(n728) );
  XOR U1093 ( .A(B[231]), .B(n729), .Z(O[232]) );
  AND U1094 ( .A(S), .B(n730), .Z(n729) );
  XOR U1095 ( .A(B[232]), .B(B[231]), .Z(n730) );
  XOR U1096 ( .A(B[230]), .B(n731), .Z(O[231]) );
  AND U1097 ( .A(S), .B(n732), .Z(n731) );
  XOR U1098 ( .A(B[231]), .B(B[230]), .Z(n732) );
  XOR U1099 ( .A(B[229]), .B(n733), .Z(O[230]) );
  AND U1100 ( .A(S), .B(n734), .Z(n733) );
  XOR U1101 ( .A(B[230]), .B(B[229]), .Z(n734) );
  XOR U1102 ( .A(B[21]), .B(n735), .Z(O[22]) );
  AND U1103 ( .A(S), .B(n736), .Z(n735) );
  XOR U1104 ( .A(B[22]), .B(B[21]), .Z(n736) );
  XOR U1105 ( .A(B[228]), .B(n737), .Z(O[229]) );
  AND U1106 ( .A(S), .B(n738), .Z(n737) );
  XOR U1107 ( .A(B[229]), .B(B[228]), .Z(n738) );
  XOR U1108 ( .A(B[227]), .B(n739), .Z(O[228]) );
  AND U1109 ( .A(S), .B(n740), .Z(n739) );
  XOR U1110 ( .A(B[228]), .B(B[227]), .Z(n740) );
  XOR U1111 ( .A(B[226]), .B(n741), .Z(O[227]) );
  AND U1112 ( .A(S), .B(n742), .Z(n741) );
  XOR U1113 ( .A(B[227]), .B(B[226]), .Z(n742) );
  XOR U1114 ( .A(B[225]), .B(n743), .Z(O[226]) );
  AND U1115 ( .A(S), .B(n744), .Z(n743) );
  XOR U1116 ( .A(B[226]), .B(B[225]), .Z(n744) );
  XOR U1117 ( .A(B[224]), .B(n745), .Z(O[225]) );
  AND U1118 ( .A(S), .B(n746), .Z(n745) );
  XOR U1119 ( .A(B[225]), .B(B[224]), .Z(n746) );
  XOR U1120 ( .A(B[223]), .B(n747), .Z(O[224]) );
  AND U1121 ( .A(S), .B(n748), .Z(n747) );
  XOR U1122 ( .A(B[224]), .B(B[223]), .Z(n748) );
  XOR U1123 ( .A(B[222]), .B(n749), .Z(O[223]) );
  AND U1124 ( .A(S), .B(n750), .Z(n749) );
  XOR U1125 ( .A(B[223]), .B(B[222]), .Z(n750) );
  XOR U1126 ( .A(B[221]), .B(n751), .Z(O[222]) );
  AND U1127 ( .A(S), .B(n752), .Z(n751) );
  XOR U1128 ( .A(B[222]), .B(B[221]), .Z(n752) );
  XOR U1129 ( .A(B[220]), .B(n753), .Z(O[221]) );
  AND U1130 ( .A(S), .B(n754), .Z(n753) );
  XOR U1131 ( .A(B[221]), .B(B[220]), .Z(n754) );
  XOR U1132 ( .A(B[219]), .B(n755), .Z(O[220]) );
  AND U1133 ( .A(S), .B(n756), .Z(n755) );
  XOR U1134 ( .A(B[220]), .B(B[219]), .Z(n756) );
  XOR U1135 ( .A(B[20]), .B(n757), .Z(O[21]) );
  AND U1136 ( .A(S), .B(n758), .Z(n757) );
  XOR U1137 ( .A(B[21]), .B(B[20]), .Z(n758) );
  XOR U1138 ( .A(B[218]), .B(n759), .Z(O[219]) );
  AND U1139 ( .A(S), .B(n760), .Z(n759) );
  XOR U1140 ( .A(B[219]), .B(B[218]), .Z(n760) );
  XOR U1141 ( .A(B[217]), .B(n761), .Z(O[218]) );
  AND U1142 ( .A(S), .B(n762), .Z(n761) );
  XOR U1143 ( .A(B[218]), .B(B[217]), .Z(n762) );
  XOR U1144 ( .A(B[216]), .B(n763), .Z(O[217]) );
  AND U1145 ( .A(S), .B(n764), .Z(n763) );
  XOR U1146 ( .A(B[217]), .B(B[216]), .Z(n764) );
  XOR U1147 ( .A(B[215]), .B(n765), .Z(O[216]) );
  AND U1148 ( .A(S), .B(n766), .Z(n765) );
  XOR U1149 ( .A(B[216]), .B(B[215]), .Z(n766) );
  XOR U1150 ( .A(B[214]), .B(n767), .Z(O[215]) );
  AND U1151 ( .A(S), .B(n768), .Z(n767) );
  XOR U1152 ( .A(B[215]), .B(B[214]), .Z(n768) );
  XOR U1153 ( .A(B[213]), .B(n769), .Z(O[214]) );
  AND U1154 ( .A(S), .B(n770), .Z(n769) );
  XOR U1155 ( .A(B[214]), .B(B[213]), .Z(n770) );
  XOR U1156 ( .A(B[212]), .B(n771), .Z(O[213]) );
  AND U1157 ( .A(S), .B(n772), .Z(n771) );
  XOR U1158 ( .A(B[213]), .B(B[212]), .Z(n772) );
  XOR U1159 ( .A(B[211]), .B(n773), .Z(O[212]) );
  AND U1160 ( .A(S), .B(n774), .Z(n773) );
  XOR U1161 ( .A(B[212]), .B(B[211]), .Z(n774) );
  XOR U1162 ( .A(B[210]), .B(n775), .Z(O[211]) );
  AND U1163 ( .A(S), .B(n776), .Z(n775) );
  XOR U1164 ( .A(B[211]), .B(B[210]), .Z(n776) );
  XOR U1165 ( .A(B[209]), .B(n777), .Z(O[210]) );
  AND U1166 ( .A(S), .B(n778), .Z(n777) );
  XOR U1167 ( .A(B[210]), .B(B[209]), .Z(n778) );
  XOR U1168 ( .A(B[19]), .B(n779), .Z(O[20]) );
  AND U1169 ( .A(S), .B(n780), .Z(n779) );
  XOR U1170 ( .A(B[20]), .B(B[19]), .Z(n780) );
  XOR U1171 ( .A(B[208]), .B(n781), .Z(O[209]) );
  AND U1172 ( .A(S), .B(n782), .Z(n781) );
  XOR U1173 ( .A(B[209]), .B(B[208]), .Z(n782) );
  XOR U1174 ( .A(B[207]), .B(n783), .Z(O[208]) );
  AND U1175 ( .A(S), .B(n784), .Z(n783) );
  XOR U1176 ( .A(B[208]), .B(B[207]), .Z(n784) );
  XOR U1177 ( .A(B[206]), .B(n785), .Z(O[207]) );
  AND U1178 ( .A(S), .B(n786), .Z(n785) );
  XOR U1179 ( .A(B[207]), .B(B[206]), .Z(n786) );
  XOR U1180 ( .A(B[205]), .B(n787), .Z(O[206]) );
  AND U1181 ( .A(S), .B(n788), .Z(n787) );
  XOR U1182 ( .A(B[206]), .B(B[205]), .Z(n788) );
  XOR U1183 ( .A(B[204]), .B(n789), .Z(O[205]) );
  AND U1184 ( .A(S), .B(n790), .Z(n789) );
  XOR U1185 ( .A(B[205]), .B(B[204]), .Z(n790) );
  XOR U1186 ( .A(B[203]), .B(n791), .Z(O[204]) );
  AND U1187 ( .A(S), .B(n792), .Z(n791) );
  XOR U1188 ( .A(B[204]), .B(B[203]), .Z(n792) );
  XOR U1189 ( .A(B[202]), .B(n793), .Z(O[203]) );
  AND U1190 ( .A(S), .B(n794), .Z(n793) );
  XOR U1191 ( .A(B[203]), .B(B[202]), .Z(n794) );
  XOR U1192 ( .A(B[201]), .B(n795), .Z(O[202]) );
  AND U1193 ( .A(S), .B(n796), .Z(n795) );
  XOR U1194 ( .A(B[202]), .B(B[201]), .Z(n796) );
  XOR U1195 ( .A(B[200]), .B(n797), .Z(O[201]) );
  AND U1196 ( .A(S), .B(n798), .Z(n797) );
  XOR U1197 ( .A(B[201]), .B(B[200]), .Z(n798) );
  XOR U1198 ( .A(B[199]), .B(n799), .Z(O[200]) );
  AND U1199 ( .A(S), .B(n800), .Z(n799) );
  XOR U1200 ( .A(B[200]), .B(B[199]), .Z(n800) );
  XOR U1201 ( .A(B[0]), .B(n801), .Z(O[1]) );
  AND U1202 ( .A(S), .B(n802), .Z(n801) );
  XOR U1203 ( .A(B[1]), .B(B[0]), .Z(n802) );
  XOR U1204 ( .A(B[18]), .B(n803), .Z(O[19]) );
  AND U1205 ( .A(S), .B(n804), .Z(n803) );
  XOR U1206 ( .A(B[19]), .B(B[18]), .Z(n804) );
  XOR U1207 ( .A(B[198]), .B(n805), .Z(O[199]) );
  AND U1208 ( .A(S), .B(n806), .Z(n805) );
  XOR U1209 ( .A(B[199]), .B(B[198]), .Z(n806) );
  XOR U1210 ( .A(B[197]), .B(n807), .Z(O[198]) );
  AND U1211 ( .A(S), .B(n808), .Z(n807) );
  XOR U1212 ( .A(B[198]), .B(B[197]), .Z(n808) );
  XOR U1213 ( .A(B[196]), .B(n809), .Z(O[197]) );
  AND U1214 ( .A(S), .B(n810), .Z(n809) );
  XOR U1215 ( .A(B[197]), .B(B[196]), .Z(n810) );
  XOR U1216 ( .A(B[195]), .B(n811), .Z(O[196]) );
  AND U1217 ( .A(S), .B(n812), .Z(n811) );
  XOR U1218 ( .A(B[196]), .B(B[195]), .Z(n812) );
  XOR U1219 ( .A(B[194]), .B(n813), .Z(O[195]) );
  AND U1220 ( .A(S), .B(n814), .Z(n813) );
  XOR U1221 ( .A(B[195]), .B(B[194]), .Z(n814) );
  XOR U1222 ( .A(B[193]), .B(n815), .Z(O[194]) );
  AND U1223 ( .A(S), .B(n816), .Z(n815) );
  XOR U1224 ( .A(B[194]), .B(B[193]), .Z(n816) );
  XOR U1225 ( .A(B[192]), .B(n817), .Z(O[193]) );
  AND U1226 ( .A(S), .B(n818), .Z(n817) );
  XOR U1227 ( .A(B[193]), .B(B[192]), .Z(n818) );
  XOR U1228 ( .A(B[191]), .B(n819), .Z(O[192]) );
  AND U1229 ( .A(S), .B(n820), .Z(n819) );
  XOR U1230 ( .A(B[192]), .B(B[191]), .Z(n820) );
  XOR U1231 ( .A(B[190]), .B(n821), .Z(O[191]) );
  AND U1232 ( .A(S), .B(n822), .Z(n821) );
  XOR U1233 ( .A(B[191]), .B(B[190]), .Z(n822) );
  XOR U1234 ( .A(B[189]), .B(n823), .Z(O[190]) );
  AND U1235 ( .A(S), .B(n824), .Z(n823) );
  XOR U1236 ( .A(B[190]), .B(B[189]), .Z(n824) );
  XOR U1237 ( .A(B[17]), .B(n825), .Z(O[18]) );
  AND U1238 ( .A(S), .B(n826), .Z(n825) );
  XOR U1239 ( .A(B[18]), .B(B[17]), .Z(n826) );
  XOR U1240 ( .A(B[188]), .B(n827), .Z(O[189]) );
  AND U1241 ( .A(S), .B(n828), .Z(n827) );
  XOR U1242 ( .A(B[189]), .B(B[188]), .Z(n828) );
  XOR U1243 ( .A(B[187]), .B(n829), .Z(O[188]) );
  AND U1244 ( .A(S), .B(n830), .Z(n829) );
  XOR U1245 ( .A(B[188]), .B(B[187]), .Z(n830) );
  XOR U1246 ( .A(B[186]), .B(n831), .Z(O[187]) );
  AND U1247 ( .A(S), .B(n832), .Z(n831) );
  XOR U1248 ( .A(B[187]), .B(B[186]), .Z(n832) );
  XOR U1249 ( .A(B[185]), .B(n833), .Z(O[186]) );
  AND U1250 ( .A(S), .B(n834), .Z(n833) );
  XOR U1251 ( .A(B[186]), .B(B[185]), .Z(n834) );
  XOR U1252 ( .A(B[184]), .B(n835), .Z(O[185]) );
  AND U1253 ( .A(S), .B(n836), .Z(n835) );
  XOR U1254 ( .A(B[185]), .B(B[184]), .Z(n836) );
  XOR U1255 ( .A(B[183]), .B(n837), .Z(O[184]) );
  AND U1256 ( .A(S), .B(n838), .Z(n837) );
  XOR U1257 ( .A(B[184]), .B(B[183]), .Z(n838) );
  XOR U1258 ( .A(B[182]), .B(n839), .Z(O[183]) );
  AND U1259 ( .A(S), .B(n840), .Z(n839) );
  XOR U1260 ( .A(B[183]), .B(B[182]), .Z(n840) );
  XOR U1261 ( .A(B[181]), .B(n841), .Z(O[182]) );
  AND U1262 ( .A(S), .B(n842), .Z(n841) );
  XOR U1263 ( .A(B[182]), .B(B[181]), .Z(n842) );
  XOR U1264 ( .A(B[180]), .B(n843), .Z(O[181]) );
  AND U1265 ( .A(S), .B(n844), .Z(n843) );
  XOR U1266 ( .A(B[181]), .B(B[180]), .Z(n844) );
  XOR U1267 ( .A(B[179]), .B(n845), .Z(O[180]) );
  AND U1268 ( .A(S), .B(n846), .Z(n845) );
  XOR U1269 ( .A(B[180]), .B(B[179]), .Z(n846) );
  XOR U1270 ( .A(B[16]), .B(n847), .Z(O[17]) );
  AND U1271 ( .A(S), .B(n848), .Z(n847) );
  XOR U1272 ( .A(B[17]), .B(B[16]), .Z(n848) );
  XOR U1273 ( .A(B[178]), .B(n849), .Z(O[179]) );
  AND U1274 ( .A(S), .B(n850), .Z(n849) );
  XOR U1275 ( .A(B[179]), .B(B[178]), .Z(n850) );
  XOR U1276 ( .A(B[177]), .B(n851), .Z(O[178]) );
  AND U1277 ( .A(S), .B(n852), .Z(n851) );
  XOR U1278 ( .A(B[178]), .B(B[177]), .Z(n852) );
  XOR U1279 ( .A(B[176]), .B(n853), .Z(O[177]) );
  AND U1280 ( .A(S), .B(n854), .Z(n853) );
  XOR U1281 ( .A(B[177]), .B(B[176]), .Z(n854) );
  XOR U1282 ( .A(B[175]), .B(n855), .Z(O[176]) );
  AND U1283 ( .A(S), .B(n856), .Z(n855) );
  XOR U1284 ( .A(B[176]), .B(B[175]), .Z(n856) );
  XOR U1285 ( .A(B[174]), .B(n857), .Z(O[175]) );
  AND U1286 ( .A(S), .B(n858), .Z(n857) );
  XOR U1287 ( .A(B[175]), .B(B[174]), .Z(n858) );
  XOR U1288 ( .A(B[173]), .B(n859), .Z(O[174]) );
  AND U1289 ( .A(S), .B(n860), .Z(n859) );
  XOR U1290 ( .A(B[174]), .B(B[173]), .Z(n860) );
  XOR U1291 ( .A(B[172]), .B(n861), .Z(O[173]) );
  AND U1292 ( .A(S), .B(n862), .Z(n861) );
  XOR U1293 ( .A(B[173]), .B(B[172]), .Z(n862) );
  XOR U1294 ( .A(B[171]), .B(n863), .Z(O[172]) );
  AND U1295 ( .A(S), .B(n864), .Z(n863) );
  XOR U1296 ( .A(B[172]), .B(B[171]), .Z(n864) );
  XOR U1297 ( .A(B[170]), .B(n865), .Z(O[171]) );
  AND U1298 ( .A(S), .B(n866), .Z(n865) );
  XOR U1299 ( .A(B[171]), .B(B[170]), .Z(n866) );
  XOR U1300 ( .A(B[169]), .B(n867), .Z(O[170]) );
  AND U1301 ( .A(S), .B(n868), .Z(n867) );
  XOR U1302 ( .A(B[170]), .B(B[169]), .Z(n868) );
  XOR U1303 ( .A(B[15]), .B(n869), .Z(O[16]) );
  AND U1304 ( .A(S), .B(n870), .Z(n869) );
  XOR U1305 ( .A(B[16]), .B(B[15]), .Z(n870) );
  XOR U1306 ( .A(B[168]), .B(n871), .Z(O[169]) );
  AND U1307 ( .A(S), .B(n872), .Z(n871) );
  XOR U1308 ( .A(B[169]), .B(B[168]), .Z(n872) );
  XOR U1309 ( .A(B[167]), .B(n873), .Z(O[168]) );
  AND U1310 ( .A(S), .B(n874), .Z(n873) );
  XOR U1311 ( .A(B[168]), .B(B[167]), .Z(n874) );
  XOR U1312 ( .A(B[166]), .B(n875), .Z(O[167]) );
  AND U1313 ( .A(S), .B(n876), .Z(n875) );
  XOR U1314 ( .A(B[167]), .B(B[166]), .Z(n876) );
  XOR U1315 ( .A(B[165]), .B(n877), .Z(O[166]) );
  AND U1316 ( .A(S), .B(n878), .Z(n877) );
  XOR U1317 ( .A(B[166]), .B(B[165]), .Z(n878) );
  XOR U1318 ( .A(B[164]), .B(n879), .Z(O[165]) );
  AND U1319 ( .A(S), .B(n880), .Z(n879) );
  XOR U1320 ( .A(B[165]), .B(B[164]), .Z(n880) );
  XOR U1321 ( .A(B[163]), .B(n881), .Z(O[164]) );
  AND U1322 ( .A(S), .B(n882), .Z(n881) );
  XOR U1323 ( .A(B[164]), .B(B[163]), .Z(n882) );
  XOR U1324 ( .A(B[162]), .B(n883), .Z(O[163]) );
  AND U1325 ( .A(S), .B(n884), .Z(n883) );
  XOR U1326 ( .A(B[163]), .B(B[162]), .Z(n884) );
  XOR U1327 ( .A(B[161]), .B(n885), .Z(O[162]) );
  AND U1328 ( .A(S), .B(n886), .Z(n885) );
  XOR U1329 ( .A(B[162]), .B(B[161]), .Z(n886) );
  XOR U1330 ( .A(B[160]), .B(n887), .Z(O[161]) );
  AND U1331 ( .A(S), .B(n888), .Z(n887) );
  XOR U1332 ( .A(B[161]), .B(B[160]), .Z(n888) );
  XOR U1333 ( .A(B[159]), .B(n889), .Z(O[160]) );
  AND U1334 ( .A(S), .B(n890), .Z(n889) );
  XOR U1335 ( .A(B[160]), .B(B[159]), .Z(n890) );
  XOR U1336 ( .A(B[14]), .B(n891), .Z(O[15]) );
  AND U1337 ( .A(S), .B(n892), .Z(n891) );
  XOR U1338 ( .A(B[15]), .B(B[14]), .Z(n892) );
  XOR U1339 ( .A(B[158]), .B(n893), .Z(O[159]) );
  AND U1340 ( .A(S), .B(n894), .Z(n893) );
  XOR U1341 ( .A(B[159]), .B(B[158]), .Z(n894) );
  XOR U1342 ( .A(B[157]), .B(n895), .Z(O[158]) );
  AND U1343 ( .A(S), .B(n896), .Z(n895) );
  XOR U1344 ( .A(B[158]), .B(B[157]), .Z(n896) );
  XOR U1345 ( .A(B[156]), .B(n897), .Z(O[157]) );
  AND U1346 ( .A(S), .B(n898), .Z(n897) );
  XOR U1347 ( .A(B[157]), .B(B[156]), .Z(n898) );
  XOR U1348 ( .A(B[155]), .B(n899), .Z(O[156]) );
  AND U1349 ( .A(S), .B(n900), .Z(n899) );
  XOR U1350 ( .A(B[156]), .B(B[155]), .Z(n900) );
  XOR U1351 ( .A(B[154]), .B(n901), .Z(O[155]) );
  AND U1352 ( .A(S), .B(n902), .Z(n901) );
  XOR U1353 ( .A(B[155]), .B(B[154]), .Z(n902) );
  XOR U1354 ( .A(B[153]), .B(n903), .Z(O[154]) );
  AND U1355 ( .A(S), .B(n904), .Z(n903) );
  XOR U1356 ( .A(B[154]), .B(B[153]), .Z(n904) );
  XOR U1357 ( .A(B[152]), .B(n905), .Z(O[153]) );
  AND U1358 ( .A(S), .B(n906), .Z(n905) );
  XOR U1359 ( .A(B[153]), .B(B[152]), .Z(n906) );
  XOR U1360 ( .A(B[151]), .B(n907), .Z(O[152]) );
  AND U1361 ( .A(S), .B(n908), .Z(n907) );
  XOR U1362 ( .A(B[152]), .B(B[151]), .Z(n908) );
  XOR U1363 ( .A(B[150]), .B(n909), .Z(O[151]) );
  AND U1364 ( .A(S), .B(n910), .Z(n909) );
  XOR U1365 ( .A(B[151]), .B(B[150]), .Z(n910) );
  XOR U1366 ( .A(B[149]), .B(n911), .Z(O[150]) );
  AND U1367 ( .A(S), .B(n912), .Z(n911) );
  XOR U1368 ( .A(B[150]), .B(B[149]), .Z(n912) );
  XOR U1369 ( .A(B[13]), .B(n913), .Z(O[14]) );
  AND U1370 ( .A(S), .B(n914), .Z(n913) );
  XOR U1371 ( .A(B[14]), .B(B[13]), .Z(n914) );
  XOR U1372 ( .A(B[148]), .B(n915), .Z(O[149]) );
  AND U1373 ( .A(S), .B(n916), .Z(n915) );
  XOR U1374 ( .A(B[149]), .B(B[148]), .Z(n916) );
  XOR U1375 ( .A(B[147]), .B(n917), .Z(O[148]) );
  AND U1376 ( .A(S), .B(n918), .Z(n917) );
  XOR U1377 ( .A(B[148]), .B(B[147]), .Z(n918) );
  XOR U1378 ( .A(B[146]), .B(n919), .Z(O[147]) );
  AND U1379 ( .A(S), .B(n920), .Z(n919) );
  XOR U1380 ( .A(B[147]), .B(B[146]), .Z(n920) );
  XOR U1381 ( .A(B[145]), .B(n921), .Z(O[146]) );
  AND U1382 ( .A(S), .B(n922), .Z(n921) );
  XOR U1383 ( .A(B[146]), .B(B[145]), .Z(n922) );
  XOR U1384 ( .A(B[144]), .B(n923), .Z(O[145]) );
  AND U1385 ( .A(S), .B(n924), .Z(n923) );
  XOR U1386 ( .A(B[145]), .B(B[144]), .Z(n924) );
  XOR U1387 ( .A(B[143]), .B(n925), .Z(O[144]) );
  AND U1388 ( .A(S), .B(n926), .Z(n925) );
  XOR U1389 ( .A(B[144]), .B(B[143]), .Z(n926) );
  XOR U1390 ( .A(B[142]), .B(n927), .Z(O[143]) );
  AND U1391 ( .A(S), .B(n928), .Z(n927) );
  XOR U1392 ( .A(B[143]), .B(B[142]), .Z(n928) );
  XOR U1393 ( .A(B[141]), .B(n929), .Z(O[142]) );
  AND U1394 ( .A(S), .B(n930), .Z(n929) );
  XOR U1395 ( .A(B[142]), .B(B[141]), .Z(n930) );
  XOR U1396 ( .A(B[140]), .B(n931), .Z(O[141]) );
  AND U1397 ( .A(S), .B(n932), .Z(n931) );
  XOR U1398 ( .A(B[141]), .B(B[140]), .Z(n932) );
  XOR U1399 ( .A(B[139]), .B(n933), .Z(O[140]) );
  AND U1400 ( .A(S), .B(n934), .Z(n933) );
  XOR U1401 ( .A(B[140]), .B(B[139]), .Z(n934) );
  XOR U1402 ( .A(B[12]), .B(n935), .Z(O[13]) );
  AND U1403 ( .A(S), .B(n936), .Z(n935) );
  XOR U1404 ( .A(B[13]), .B(B[12]), .Z(n936) );
  XOR U1405 ( .A(B[138]), .B(n937), .Z(O[139]) );
  AND U1406 ( .A(S), .B(n938), .Z(n937) );
  XOR U1407 ( .A(B[139]), .B(B[138]), .Z(n938) );
  XOR U1408 ( .A(B[137]), .B(n939), .Z(O[138]) );
  AND U1409 ( .A(S), .B(n940), .Z(n939) );
  XOR U1410 ( .A(B[138]), .B(B[137]), .Z(n940) );
  XOR U1411 ( .A(B[136]), .B(n941), .Z(O[137]) );
  AND U1412 ( .A(S), .B(n942), .Z(n941) );
  XOR U1413 ( .A(B[137]), .B(B[136]), .Z(n942) );
  XOR U1414 ( .A(B[135]), .B(n943), .Z(O[136]) );
  AND U1415 ( .A(S), .B(n944), .Z(n943) );
  XOR U1416 ( .A(B[136]), .B(B[135]), .Z(n944) );
  XOR U1417 ( .A(B[134]), .B(n945), .Z(O[135]) );
  AND U1418 ( .A(S), .B(n946), .Z(n945) );
  XOR U1419 ( .A(B[135]), .B(B[134]), .Z(n946) );
  XOR U1420 ( .A(B[133]), .B(n947), .Z(O[134]) );
  AND U1421 ( .A(S), .B(n948), .Z(n947) );
  XOR U1422 ( .A(B[134]), .B(B[133]), .Z(n948) );
  XOR U1423 ( .A(B[132]), .B(n949), .Z(O[133]) );
  AND U1424 ( .A(S), .B(n950), .Z(n949) );
  XOR U1425 ( .A(B[133]), .B(B[132]), .Z(n950) );
  XOR U1426 ( .A(B[131]), .B(n951), .Z(O[132]) );
  AND U1427 ( .A(S), .B(n952), .Z(n951) );
  XOR U1428 ( .A(B[132]), .B(B[131]), .Z(n952) );
  XOR U1429 ( .A(B[130]), .B(n953), .Z(O[131]) );
  AND U1430 ( .A(S), .B(n954), .Z(n953) );
  XOR U1431 ( .A(B[131]), .B(B[130]), .Z(n954) );
  XOR U1432 ( .A(B[129]), .B(n955), .Z(O[130]) );
  AND U1433 ( .A(S), .B(n956), .Z(n955) );
  XOR U1434 ( .A(B[130]), .B(B[129]), .Z(n956) );
  XOR U1435 ( .A(B[11]), .B(n957), .Z(O[12]) );
  AND U1436 ( .A(S), .B(n958), .Z(n957) );
  XOR U1437 ( .A(B[12]), .B(B[11]), .Z(n958) );
  XOR U1438 ( .A(B[128]), .B(n959), .Z(O[129]) );
  AND U1439 ( .A(S), .B(n960), .Z(n959) );
  XOR U1440 ( .A(B[129]), .B(B[128]), .Z(n960) );
  XOR U1441 ( .A(B[127]), .B(n961), .Z(O[128]) );
  AND U1442 ( .A(S), .B(n962), .Z(n961) );
  XOR U1443 ( .A(B[128]), .B(B[127]), .Z(n962) );
  XOR U1444 ( .A(B[126]), .B(n963), .Z(O[127]) );
  AND U1445 ( .A(S), .B(n964), .Z(n963) );
  XOR U1446 ( .A(B[127]), .B(B[126]), .Z(n964) );
  XOR U1447 ( .A(B[125]), .B(n965), .Z(O[126]) );
  AND U1448 ( .A(S), .B(n966), .Z(n965) );
  XOR U1449 ( .A(B[126]), .B(B[125]), .Z(n966) );
  XOR U1450 ( .A(B[124]), .B(n967), .Z(O[125]) );
  AND U1451 ( .A(S), .B(n968), .Z(n967) );
  XOR U1452 ( .A(B[125]), .B(B[124]), .Z(n968) );
  XOR U1453 ( .A(B[123]), .B(n969), .Z(O[124]) );
  AND U1454 ( .A(S), .B(n970), .Z(n969) );
  XOR U1455 ( .A(B[124]), .B(B[123]), .Z(n970) );
  XOR U1456 ( .A(B[122]), .B(n971), .Z(O[123]) );
  AND U1457 ( .A(S), .B(n972), .Z(n971) );
  XOR U1458 ( .A(B[123]), .B(B[122]), .Z(n972) );
  XOR U1459 ( .A(B[121]), .B(n973), .Z(O[122]) );
  AND U1460 ( .A(S), .B(n974), .Z(n973) );
  XOR U1461 ( .A(B[122]), .B(B[121]), .Z(n974) );
  XOR U1462 ( .A(B[120]), .B(n975), .Z(O[121]) );
  AND U1463 ( .A(S), .B(n976), .Z(n975) );
  XOR U1464 ( .A(B[121]), .B(B[120]), .Z(n976) );
  XOR U1465 ( .A(B[119]), .B(n977), .Z(O[120]) );
  AND U1466 ( .A(S), .B(n978), .Z(n977) );
  XOR U1467 ( .A(B[120]), .B(B[119]), .Z(n978) );
  XOR U1468 ( .A(B[10]), .B(n979), .Z(O[11]) );
  AND U1469 ( .A(S), .B(n980), .Z(n979) );
  XOR U1470 ( .A(B[11]), .B(B[10]), .Z(n980) );
  XOR U1471 ( .A(B[118]), .B(n981), .Z(O[119]) );
  AND U1472 ( .A(S), .B(n982), .Z(n981) );
  XOR U1473 ( .A(B[119]), .B(B[118]), .Z(n982) );
  XOR U1474 ( .A(B[117]), .B(n983), .Z(O[118]) );
  AND U1475 ( .A(S), .B(n984), .Z(n983) );
  XOR U1476 ( .A(B[118]), .B(B[117]), .Z(n984) );
  XOR U1477 ( .A(B[116]), .B(n985), .Z(O[117]) );
  AND U1478 ( .A(S), .B(n986), .Z(n985) );
  XOR U1479 ( .A(B[117]), .B(B[116]), .Z(n986) );
  XOR U1480 ( .A(B[115]), .B(n987), .Z(O[116]) );
  AND U1481 ( .A(S), .B(n988), .Z(n987) );
  XOR U1482 ( .A(B[116]), .B(B[115]), .Z(n988) );
  XOR U1483 ( .A(B[114]), .B(n989), .Z(O[115]) );
  AND U1484 ( .A(S), .B(n990), .Z(n989) );
  XOR U1485 ( .A(B[115]), .B(B[114]), .Z(n990) );
  XOR U1486 ( .A(B[113]), .B(n991), .Z(O[114]) );
  AND U1487 ( .A(S), .B(n992), .Z(n991) );
  XOR U1488 ( .A(B[114]), .B(B[113]), .Z(n992) );
  XOR U1489 ( .A(B[112]), .B(n993), .Z(O[113]) );
  AND U1490 ( .A(S), .B(n994), .Z(n993) );
  XOR U1491 ( .A(B[113]), .B(B[112]), .Z(n994) );
  XOR U1492 ( .A(B[111]), .B(n995), .Z(O[112]) );
  AND U1493 ( .A(S), .B(n996), .Z(n995) );
  XOR U1494 ( .A(B[112]), .B(B[111]), .Z(n996) );
  XOR U1495 ( .A(B[110]), .B(n997), .Z(O[111]) );
  AND U1496 ( .A(S), .B(n998), .Z(n997) );
  XOR U1497 ( .A(B[111]), .B(B[110]), .Z(n998) );
  XOR U1498 ( .A(B[109]), .B(n999), .Z(O[110]) );
  AND U1499 ( .A(S), .B(n1000), .Z(n999) );
  XOR U1500 ( .A(B[110]), .B(B[109]), .Z(n1000) );
  XOR U1501 ( .A(B[9]), .B(n1001), .Z(O[10]) );
  AND U1502 ( .A(S), .B(n1002), .Z(n1001) );
  XOR U1503 ( .A(B[9]), .B(B[10]), .Z(n1002) );
  XOR U1504 ( .A(B[108]), .B(n1003), .Z(O[109]) );
  AND U1505 ( .A(S), .B(n1004), .Z(n1003) );
  XOR U1506 ( .A(B[109]), .B(B[108]), .Z(n1004) );
  XOR U1507 ( .A(B[107]), .B(n1005), .Z(O[108]) );
  AND U1508 ( .A(S), .B(n1006), .Z(n1005) );
  XOR U1509 ( .A(B[108]), .B(B[107]), .Z(n1006) );
  XOR U1510 ( .A(B[106]), .B(n1007), .Z(O[107]) );
  AND U1511 ( .A(S), .B(n1008), .Z(n1007) );
  XOR U1512 ( .A(B[107]), .B(B[106]), .Z(n1008) );
  XOR U1513 ( .A(B[105]), .B(n1009), .Z(O[106]) );
  AND U1514 ( .A(S), .B(n1010), .Z(n1009) );
  XOR U1515 ( .A(B[106]), .B(B[105]), .Z(n1010) );
  XOR U1516 ( .A(B[104]), .B(n1011), .Z(O[105]) );
  AND U1517 ( .A(S), .B(n1012), .Z(n1011) );
  XOR U1518 ( .A(B[105]), .B(B[104]), .Z(n1012) );
  XOR U1519 ( .A(B[103]), .B(n1013), .Z(O[104]) );
  AND U1520 ( .A(S), .B(n1014), .Z(n1013) );
  XOR U1521 ( .A(B[104]), .B(B[103]), .Z(n1014) );
  XOR U1522 ( .A(B[102]), .B(n1015), .Z(O[103]) );
  AND U1523 ( .A(S), .B(n1016), .Z(n1015) );
  XOR U1524 ( .A(B[103]), .B(B[102]), .Z(n1016) );
  XOR U1525 ( .A(B[101]), .B(n1017), .Z(O[102]) );
  AND U1526 ( .A(S), .B(n1018), .Z(n1017) );
  XOR U1527 ( .A(B[102]), .B(B[101]), .Z(n1018) );
  XOR U1528 ( .A(B[100]), .B(n1019), .Z(O[101]) );
  AND U1529 ( .A(S), .B(n1020), .Z(n1019) );
  XOR U1530 ( .A(B[101]), .B(B[100]), .Z(n1020) );
  XOR U1531 ( .A(B[99]), .B(n1021), .Z(O[100]) );
  AND U1532 ( .A(S), .B(n1022), .Z(n1021) );
  XOR U1533 ( .A(B[99]), .B(B[100]), .Z(n1022) );
  AND U1534 ( .A(B[0]), .B(S), .Z(O[0]) );
endmodule


module modexp_2N_NN_N512_CC524288 ( clk, rst, m, e, n, c );
  input [511:0] m;
  input [511:0] e;
  input [511:0] n;
  output [511:0] c;
  input clk, rst;
  wire   _0_net_, first_one, mul_pow, n6, n8, n521, n522, n523, n524;
  wire   [511:0] start_in;
  wire   [511:0] ein;
  wire   [511:0] creg_next;
  wire   [511:0] o;
  wire   [511:0] ereg_next;
  wire   [511:0] y;

  MUX_N512_0 MUX_4 ( .A(o), .B(c), .S(_0_net_), .O(creg_next) );
  MUX_N512_2 MUX_6 ( .A({ein[510:0], 1'b0}), .B(ein), .S(mul_pow), .O(
        ereg_next) );
  MUX_N512_1 MUX_9 ( .A(m), .B(c), .S(mul_pow), .O(y) );
  modmult_N512_CC512 modmult_1 ( .clk(clk), .rst(1'b0), .start(start_in[0]), 
        .x(c), .y(y), .n(n), .o(o) );
  DFF \start_reg_reg[0]  ( .D(start_in[511]), .CLK(clk), .RST(rst), .I(1'b1), 
        .Q(start_in[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[127]) );
  DFF \start_reg_reg[128]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[128]) );
  DFF \start_reg_reg[129]  ( .D(start_in[128]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[129]) );
  DFF \start_reg_reg[130]  ( .D(start_in[129]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[130]) );
  DFF \start_reg_reg[131]  ( .D(start_in[130]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[131]) );
  DFF \start_reg_reg[132]  ( .D(start_in[131]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[132]) );
  DFF \start_reg_reg[133]  ( .D(start_in[132]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[133]) );
  DFF \start_reg_reg[134]  ( .D(start_in[133]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[134]) );
  DFF \start_reg_reg[135]  ( .D(start_in[134]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[135]) );
  DFF \start_reg_reg[136]  ( .D(start_in[135]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[136]) );
  DFF \start_reg_reg[137]  ( .D(start_in[136]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[137]) );
  DFF \start_reg_reg[138]  ( .D(start_in[137]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[138]) );
  DFF \start_reg_reg[139]  ( .D(start_in[138]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[139]) );
  DFF \start_reg_reg[140]  ( .D(start_in[139]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[140]) );
  DFF \start_reg_reg[141]  ( .D(start_in[140]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[141]) );
  DFF \start_reg_reg[142]  ( .D(start_in[141]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[142]) );
  DFF \start_reg_reg[143]  ( .D(start_in[142]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[143]) );
  DFF \start_reg_reg[144]  ( .D(start_in[143]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[144]) );
  DFF \start_reg_reg[145]  ( .D(start_in[144]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[145]) );
  DFF \start_reg_reg[146]  ( .D(start_in[145]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[146]) );
  DFF \start_reg_reg[147]  ( .D(start_in[146]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[147]) );
  DFF \start_reg_reg[148]  ( .D(start_in[147]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[148]) );
  DFF \start_reg_reg[149]  ( .D(start_in[148]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[149]) );
  DFF \start_reg_reg[150]  ( .D(start_in[149]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[150]) );
  DFF \start_reg_reg[151]  ( .D(start_in[150]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[151]) );
  DFF \start_reg_reg[152]  ( .D(start_in[151]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[152]) );
  DFF \start_reg_reg[153]  ( .D(start_in[152]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[153]) );
  DFF \start_reg_reg[154]  ( .D(start_in[153]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[154]) );
  DFF \start_reg_reg[155]  ( .D(start_in[154]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[155]) );
  DFF \start_reg_reg[156]  ( .D(start_in[155]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[156]) );
  DFF \start_reg_reg[157]  ( .D(start_in[156]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[157]) );
  DFF \start_reg_reg[158]  ( .D(start_in[157]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[158]) );
  DFF \start_reg_reg[159]  ( .D(start_in[158]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[159]) );
  DFF \start_reg_reg[160]  ( .D(start_in[159]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[160]) );
  DFF \start_reg_reg[161]  ( .D(start_in[160]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[161]) );
  DFF \start_reg_reg[162]  ( .D(start_in[161]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[162]) );
  DFF \start_reg_reg[163]  ( .D(start_in[162]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[163]) );
  DFF \start_reg_reg[164]  ( .D(start_in[163]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[164]) );
  DFF \start_reg_reg[165]  ( .D(start_in[164]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[165]) );
  DFF \start_reg_reg[166]  ( .D(start_in[165]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[166]) );
  DFF \start_reg_reg[167]  ( .D(start_in[166]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[167]) );
  DFF \start_reg_reg[168]  ( .D(start_in[167]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[168]) );
  DFF \start_reg_reg[169]  ( .D(start_in[168]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[169]) );
  DFF \start_reg_reg[170]  ( .D(start_in[169]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[170]) );
  DFF \start_reg_reg[171]  ( .D(start_in[170]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[171]) );
  DFF \start_reg_reg[172]  ( .D(start_in[171]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[172]) );
  DFF \start_reg_reg[173]  ( .D(start_in[172]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[173]) );
  DFF \start_reg_reg[174]  ( .D(start_in[173]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[174]) );
  DFF \start_reg_reg[175]  ( .D(start_in[174]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[175]) );
  DFF \start_reg_reg[176]  ( .D(start_in[175]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[176]) );
  DFF \start_reg_reg[177]  ( .D(start_in[176]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[177]) );
  DFF \start_reg_reg[178]  ( .D(start_in[177]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[178]) );
  DFF \start_reg_reg[179]  ( .D(start_in[178]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[179]) );
  DFF \start_reg_reg[180]  ( .D(start_in[179]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[180]) );
  DFF \start_reg_reg[181]  ( .D(start_in[180]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[181]) );
  DFF \start_reg_reg[182]  ( .D(start_in[181]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[182]) );
  DFF \start_reg_reg[183]  ( .D(start_in[182]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[183]) );
  DFF \start_reg_reg[184]  ( .D(start_in[183]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[184]) );
  DFF \start_reg_reg[185]  ( .D(start_in[184]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[185]) );
  DFF \start_reg_reg[186]  ( .D(start_in[185]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[186]) );
  DFF \start_reg_reg[187]  ( .D(start_in[186]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[187]) );
  DFF \start_reg_reg[188]  ( .D(start_in[187]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[188]) );
  DFF \start_reg_reg[189]  ( .D(start_in[188]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[189]) );
  DFF \start_reg_reg[190]  ( .D(start_in[189]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[190]) );
  DFF \start_reg_reg[191]  ( .D(start_in[190]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[191]) );
  DFF \start_reg_reg[192]  ( .D(start_in[191]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[192]) );
  DFF \start_reg_reg[193]  ( .D(start_in[192]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[193]) );
  DFF \start_reg_reg[194]  ( .D(start_in[193]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[194]) );
  DFF \start_reg_reg[195]  ( .D(start_in[194]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[195]) );
  DFF \start_reg_reg[196]  ( .D(start_in[195]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[196]) );
  DFF \start_reg_reg[197]  ( .D(start_in[196]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[197]) );
  DFF \start_reg_reg[198]  ( .D(start_in[197]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[198]) );
  DFF \start_reg_reg[199]  ( .D(start_in[198]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[199]) );
  DFF \start_reg_reg[200]  ( .D(start_in[199]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[200]) );
  DFF \start_reg_reg[201]  ( .D(start_in[200]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[201]) );
  DFF \start_reg_reg[202]  ( .D(start_in[201]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[202]) );
  DFF \start_reg_reg[203]  ( .D(start_in[202]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[203]) );
  DFF \start_reg_reg[204]  ( .D(start_in[203]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[204]) );
  DFF \start_reg_reg[205]  ( .D(start_in[204]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[205]) );
  DFF \start_reg_reg[206]  ( .D(start_in[205]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[206]) );
  DFF \start_reg_reg[207]  ( .D(start_in[206]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[207]) );
  DFF \start_reg_reg[208]  ( .D(start_in[207]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[208]) );
  DFF \start_reg_reg[209]  ( .D(start_in[208]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[209]) );
  DFF \start_reg_reg[210]  ( .D(start_in[209]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[210]) );
  DFF \start_reg_reg[211]  ( .D(start_in[210]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[211]) );
  DFF \start_reg_reg[212]  ( .D(start_in[211]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[212]) );
  DFF \start_reg_reg[213]  ( .D(start_in[212]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[213]) );
  DFF \start_reg_reg[214]  ( .D(start_in[213]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[214]) );
  DFF \start_reg_reg[215]  ( .D(start_in[214]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[215]) );
  DFF \start_reg_reg[216]  ( .D(start_in[215]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[216]) );
  DFF \start_reg_reg[217]  ( .D(start_in[216]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[217]) );
  DFF \start_reg_reg[218]  ( .D(start_in[217]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[218]) );
  DFF \start_reg_reg[219]  ( .D(start_in[218]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[219]) );
  DFF \start_reg_reg[220]  ( .D(start_in[219]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[220]) );
  DFF \start_reg_reg[221]  ( .D(start_in[220]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[221]) );
  DFF \start_reg_reg[222]  ( .D(start_in[221]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[222]) );
  DFF \start_reg_reg[223]  ( .D(start_in[222]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[223]) );
  DFF \start_reg_reg[224]  ( .D(start_in[223]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[224]) );
  DFF \start_reg_reg[225]  ( .D(start_in[224]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[225]) );
  DFF \start_reg_reg[226]  ( .D(start_in[225]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[226]) );
  DFF \start_reg_reg[227]  ( .D(start_in[226]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[227]) );
  DFF \start_reg_reg[228]  ( .D(start_in[227]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[228]) );
  DFF \start_reg_reg[229]  ( .D(start_in[228]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[229]) );
  DFF \start_reg_reg[230]  ( .D(start_in[229]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[230]) );
  DFF \start_reg_reg[231]  ( .D(start_in[230]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[231]) );
  DFF \start_reg_reg[232]  ( .D(start_in[231]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[232]) );
  DFF \start_reg_reg[233]  ( .D(start_in[232]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[233]) );
  DFF \start_reg_reg[234]  ( .D(start_in[233]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[234]) );
  DFF \start_reg_reg[235]  ( .D(start_in[234]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[235]) );
  DFF \start_reg_reg[236]  ( .D(start_in[235]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[236]) );
  DFF \start_reg_reg[237]  ( .D(start_in[236]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[237]) );
  DFF \start_reg_reg[238]  ( .D(start_in[237]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[238]) );
  DFF \start_reg_reg[239]  ( .D(start_in[238]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[239]) );
  DFF \start_reg_reg[240]  ( .D(start_in[239]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[240]) );
  DFF \start_reg_reg[241]  ( .D(start_in[240]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[241]) );
  DFF \start_reg_reg[242]  ( .D(start_in[241]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[242]) );
  DFF \start_reg_reg[243]  ( .D(start_in[242]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[243]) );
  DFF \start_reg_reg[244]  ( .D(start_in[243]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[244]) );
  DFF \start_reg_reg[245]  ( .D(start_in[244]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[245]) );
  DFF \start_reg_reg[246]  ( .D(start_in[245]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[246]) );
  DFF \start_reg_reg[247]  ( .D(start_in[246]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[247]) );
  DFF \start_reg_reg[248]  ( .D(start_in[247]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[248]) );
  DFF \start_reg_reg[249]  ( .D(start_in[248]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[249]) );
  DFF \start_reg_reg[250]  ( .D(start_in[249]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[250]) );
  DFF \start_reg_reg[251]  ( .D(start_in[250]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[251]) );
  DFF \start_reg_reg[252]  ( .D(start_in[251]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[252]) );
  DFF \start_reg_reg[253]  ( .D(start_in[252]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[253]) );
  DFF \start_reg_reg[254]  ( .D(start_in[253]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[254]) );
  DFF \start_reg_reg[255]  ( .D(start_in[254]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[255]) );
  DFF \start_reg_reg[256]  ( .D(start_in[255]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[256]) );
  DFF \start_reg_reg[257]  ( .D(start_in[256]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[257]) );
  DFF \start_reg_reg[258]  ( .D(start_in[257]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[258]) );
  DFF \start_reg_reg[259]  ( .D(start_in[258]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[259]) );
  DFF \start_reg_reg[260]  ( .D(start_in[259]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[260]) );
  DFF \start_reg_reg[261]  ( .D(start_in[260]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[261]) );
  DFF \start_reg_reg[262]  ( .D(start_in[261]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[262]) );
  DFF \start_reg_reg[263]  ( .D(start_in[262]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[263]) );
  DFF \start_reg_reg[264]  ( .D(start_in[263]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[264]) );
  DFF \start_reg_reg[265]  ( .D(start_in[264]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[265]) );
  DFF \start_reg_reg[266]  ( .D(start_in[265]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[266]) );
  DFF \start_reg_reg[267]  ( .D(start_in[266]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[267]) );
  DFF \start_reg_reg[268]  ( .D(start_in[267]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[268]) );
  DFF \start_reg_reg[269]  ( .D(start_in[268]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[269]) );
  DFF \start_reg_reg[270]  ( .D(start_in[269]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[270]) );
  DFF \start_reg_reg[271]  ( .D(start_in[270]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[271]) );
  DFF \start_reg_reg[272]  ( .D(start_in[271]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[272]) );
  DFF \start_reg_reg[273]  ( .D(start_in[272]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[273]) );
  DFF \start_reg_reg[274]  ( .D(start_in[273]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[274]) );
  DFF \start_reg_reg[275]  ( .D(start_in[274]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[275]) );
  DFF \start_reg_reg[276]  ( .D(start_in[275]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[276]) );
  DFF \start_reg_reg[277]  ( .D(start_in[276]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[277]) );
  DFF \start_reg_reg[278]  ( .D(start_in[277]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[278]) );
  DFF \start_reg_reg[279]  ( .D(start_in[278]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[279]) );
  DFF \start_reg_reg[280]  ( .D(start_in[279]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[280]) );
  DFF \start_reg_reg[281]  ( .D(start_in[280]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[281]) );
  DFF \start_reg_reg[282]  ( .D(start_in[281]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[282]) );
  DFF \start_reg_reg[283]  ( .D(start_in[282]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[283]) );
  DFF \start_reg_reg[284]  ( .D(start_in[283]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[284]) );
  DFF \start_reg_reg[285]  ( .D(start_in[284]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[285]) );
  DFF \start_reg_reg[286]  ( .D(start_in[285]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[286]) );
  DFF \start_reg_reg[287]  ( .D(start_in[286]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[287]) );
  DFF \start_reg_reg[288]  ( .D(start_in[287]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[288]) );
  DFF \start_reg_reg[289]  ( .D(start_in[288]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[289]) );
  DFF \start_reg_reg[290]  ( .D(start_in[289]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[290]) );
  DFF \start_reg_reg[291]  ( .D(start_in[290]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[291]) );
  DFF \start_reg_reg[292]  ( .D(start_in[291]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[292]) );
  DFF \start_reg_reg[293]  ( .D(start_in[292]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[293]) );
  DFF \start_reg_reg[294]  ( .D(start_in[293]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[294]) );
  DFF \start_reg_reg[295]  ( .D(start_in[294]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[295]) );
  DFF \start_reg_reg[296]  ( .D(start_in[295]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[296]) );
  DFF \start_reg_reg[297]  ( .D(start_in[296]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[297]) );
  DFF \start_reg_reg[298]  ( .D(start_in[297]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[298]) );
  DFF \start_reg_reg[299]  ( .D(start_in[298]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[299]) );
  DFF \start_reg_reg[300]  ( .D(start_in[299]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[300]) );
  DFF \start_reg_reg[301]  ( .D(start_in[300]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[301]) );
  DFF \start_reg_reg[302]  ( .D(start_in[301]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[302]) );
  DFF \start_reg_reg[303]  ( .D(start_in[302]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[303]) );
  DFF \start_reg_reg[304]  ( .D(start_in[303]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[304]) );
  DFF \start_reg_reg[305]  ( .D(start_in[304]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[305]) );
  DFF \start_reg_reg[306]  ( .D(start_in[305]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[306]) );
  DFF \start_reg_reg[307]  ( .D(start_in[306]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[307]) );
  DFF \start_reg_reg[308]  ( .D(start_in[307]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[308]) );
  DFF \start_reg_reg[309]  ( .D(start_in[308]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[309]) );
  DFF \start_reg_reg[310]  ( .D(start_in[309]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[310]) );
  DFF \start_reg_reg[311]  ( .D(start_in[310]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[311]) );
  DFF \start_reg_reg[312]  ( .D(start_in[311]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[312]) );
  DFF \start_reg_reg[313]  ( .D(start_in[312]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[313]) );
  DFF \start_reg_reg[314]  ( .D(start_in[313]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[314]) );
  DFF \start_reg_reg[315]  ( .D(start_in[314]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[315]) );
  DFF \start_reg_reg[316]  ( .D(start_in[315]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[316]) );
  DFF \start_reg_reg[317]  ( .D(start_in[316]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[317]) );
  DFF \start_reg_reg[318]  ( .D(start_in[317]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[318]) );
  DFF \start_reg_reg[319]  ( .D(start_in[318]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[319]) );
  DFF \start_reg_reg[320]  ( .D(start_in[319]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[320]) );
  DFF \start_reg_reg[321]  ( .D(start_in[320]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[321]) );
  DFF \start_reg_reg[322]  ( .D(start_in[321]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[322]) );
  DFF \start_reg_reg[323]  ( .D(start_in[322]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[323]) );
  DFF \start_reg_reg[324]  ( .D(start_in[323]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[324]) );
  DFF \start_reg_reg[325]  ( .D(start_in[324]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[325]) );
  DFF \start_reg_reg[326]  ( .D(start_in[325]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[326]) );
  DFF \start_reg_reg[327]  ( .D(start_in[326]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[327]) );
  DFF \start_reg_reg[328]  ( .D(start_in[327]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[328]) );
  DFF \start_reg_reg[329]  ( .D(start_in[328]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[329]) );
  DFF \start_reg_reg[330]  ( .D(start_in[329]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[330]) );
  DFF \start_reg_reg[331]  ( .D(start_in[330]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[331]) );
  DFF \start_reg_reg[332]  ( .D(start_in[331]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[332]) );
  DFF \start_reg_reg[333]  ( .D(start_in[332]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[333]) );
  DFF \start_reg_reg[334]  ( .D(start_in[333]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[334]) );
  DFF \start_reg_reg[335]  ( .D(start_in[334]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[335]) );
  DFF \start_reg_reg[336]  ( .D(start_in[335]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[336]) );
  DFF \start_reg_reg[337]  ( .D(start_in[336]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[337]) );
  DFF \start_reg_reg[338]  ( .D(start_in[337]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[338]) );
  DFF \start_reg_reg[339]  ( .D(start_in[338]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[339]) );
  DFF \start_reg_reg[340]  ( .D(start_in[339]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[340]) );
  DFF \start_reg_reg[341]  ( .D(start_in[340]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[341]) );
  DFF \start_reg_reg[342]  ( .D(start_in[341]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[342]) );
  DFF \start_reg_reg[343]  ( .D(start_in[342]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[343]) );
  DFF \start_reg_reg[344]  ( .D(start_in[343]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[344]) );
  DFF \start_reg_reg[345]  ( .D(start_in[344]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[345]) );
  DFF \start_reg_reg[346]  ( .D(start_in[345]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[346]) );
  DFF \start_reg_reg[347]  ( .D(start_in[346]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[347]) );
  DFF \start_reg_reg[348]  ( .D(start_in[347]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[348]) );
  DFF \start_reg_reg[349]  ( .D(start_in[348]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[349]) );
  DFF \start_reg_reg[350]  ( .D(start_in[349]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[350]) );
  DFF \start_reg_reg[351]  ( .D(start_in[350]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[351]) );
  DFF \start_reg_reg[352]  ( .D(start_in[351]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[352]) );
  DFF \start_reg_reg[353]  ( .D(start_in[352]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[353]) );
  DFF \start_reg_reg[354]  ( .D(start_in[353]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[354]) );
  DFF \start_reg_reg[355]  ( .D(start_in[354]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[355]) );
  DFF \start_reg_reg[356]  ( .D(start_in[355]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[356]) );
  DFF \start_reg_reg[357]  ( .D(start_in[356]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[357]) );
  DFF \start_reg_reg[358]  ( .D(start_in[357]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[358]) );
  DFF \start_reg_reg[359]  ( .D(start_in[358]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[359]) );
  DFF \start_reg_reg[360]  ( .D(start_in[359]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[360]) );
  DFF \start_reg_reg[361]  ( .D(start_in[360]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[361]) );
  DFF \start_reg_reg[362]  ( .D(start_in[361]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[362]) );
  DFF \start_reg_reg[363]  ( .D(start_in[362]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[363]) );
  DFF \start_reg_reg[364]  ( .D(start_in[363]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[364]) );
  DFF \start_reg_reg[365]  ( .D(start_in[364]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[365]) );
  DFF \start_reg_reg[366]  ( .D(start_in[365]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[366]) );
  DFF \start_reg_reg[367]  ( .D(start_in[366]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[367]) );
  DFF \start_reg_reg[368]  ( .D(start_in[367]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[368]) );
  DFF \start_reg_reg[369]  ( .D(start_in[368]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[369]) );
  DFF \start_reg_reg[370]  ( .D(start_in[369]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[370]) );
  DFF \start_reg_reg[371]  ( .D(start_in[370]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[371]) );
  DFF \start_reg_reg[372]  ( .D(start_in[371]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[372]) );
  DFF \start_reg_reg[373]  ( .D(start_in[372]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[373]) );
  DFF \start_reg_reg[374]  ( .D(start_in[373]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[374]) );
  DFF \start_reg_reg[375]  ( .D(start_in[374]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[375]) );
  DFF \start_reg_reg[376]  ( .D(start_in[375]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[376]) );
  DFF \start_reg_reg[377]  ( .D(start_in[376]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[377]) );
  DFF \start_reg_reg[378]  ( .D(start_in[377]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[378]) );
  DFF \start_reg_reg[379]  ( .D(start_in[378]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[379]) );
  DFF \start_reg_reg[380]  ( .D(start_in[379]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[380]) );
  DFF \start_reg_reg[381]  ( .D(start_in[380]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[381]) );
  DFF \start_reg_reg[382]  ( .D(start_in[381]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[382]) );
  DFF \start_reg_reg[383]  ( .D(start_in[382]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[383]) );
  DFF \start_reg_reg[384]  ( .D(start_in[383]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[384]) );
  DFF \start_reg_reg[385]  ( .D(start_in[384]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[385]) );
  DFF \start_reg_reg[386]  ( .D(start_in[385]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[386]) );
  DFF \start_reg_reg[387]  ( .D(start_in[386]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[387]) );
  DFF \start_reg_reg[388]  ( .D(start_in[387]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[388]) );
  DFF \start_reg_reg[389]  ( .D(start_in[388]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[389]) );
  DFF \start_reg_reg[390]  ( .D(start_in[389]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[390]) );
  DFF \start_reg_reg[391]  ( .D(start_in[390]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[391]) );
  DFF \start_reg_reg[392]  ( .D(start_in[391]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[392]) );
  DFF \start_reg_reg[393]  ( .D(start_in[392]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[393]) );
  DFF \start_reg_reg[394]  ( .D(start_in[393]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[394]) );
  DFF \start_reg_reg[395]  ( .D(start_in[394]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[395]) );
  DFF \start_reg_reg[396]  ( .D(start_in[395]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[396]) );
  DFF \start_reg_reg[397]  ( .D(start_in[396]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[397]) );
  DFF \start_reg_reg[398]  ( .D(start_in[397]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[398]) );
  DFF \start_reg_reg[399]  ( .D(start_in[398]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[399]) );
  DFF \start_reg_reg[400]  ( .D(start_in[399]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[400]) );
  DFF \start_reg_reg[401]  ( .D(start_in[400]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[401]) );
  DFF \start_reg_reg[402]  ( .D(start_in[401]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[402]) );
  DFF \start_reg_reg[403]  ( .D(start_in[402]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[403]) );
  DFF \start_reg_reg[404]  ( .D(start_in[403]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[404]) );
  DFF \start_reg_reg[405]  ( .D(start_in[404]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[405]) );
  DFF \start_reg_reg[406]  ( .D(start_in[405]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[406]) );
  DFF \start_reg_reg[407]  ( .D(start_in[406]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[407]) );
  DFF \start_reg_reg[408]  ( .D(start_in[407]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[408]) );
  DFF \start_reg_reg[409]  ( .D(start_in[408]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[409]) );
  DFF \start_reg_reg[410]  ( .D(start_in[409]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[410]) );
  DFF \start_reg_reg[411]  ( .D(start_in[410]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[411]) );
  DFF \start_reg_reg[412]  ( .D(start_in[411]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[412]) );
  DFF \start_reg_reg[413]  ( .D(start_in[412]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[413]) );
  DFF \start_reg_reg[414]  ( .D(start_in[413]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[414]) );
  DFF \start_reg_reg[415]  ( .D(start_in[414]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[415]) );
  DFF \start_reg_reg[416]  ( .D(start_in[415]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[416]) );
  DFF \start_reg_reg[417]  ( .D(start_in[416]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[417]) );
  DFF \start_reg_reg[418]  ( .D(start_in[417]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[418]) );
  DFF \start_reg_reg[419]  ( .D(start_in[418]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[419]) );
  DFF \start_reg_reg[420]  ( .D(start_in[419]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[420]) );
  DFF \start_reg_reg[421]  ( .D(start_in[420]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[421]) );
  DFF \start_reg_reg[422]  ( .D(start_in[421]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[422]) );
  DFF \start_reg_reg[423]  ( .D(start_in[422]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[423]) );
  DFF \start_reg_reg[424]  ( .D(start_in[423]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[424]) );
  DFF \start_reg_reg[425]  ( .D(start_in[424]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[425]) );
  DFF \start_reg_reg[426]  ( .D(start_in[425]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[426]) );
  DFF \start_reg_reg[427]  ( .D(start_in[426]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[427]) );
  DFF \start_reg_reg[428]  ( .D(start_in[427]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[428]) );
  DFF \start_reg_reg[429]  ( .D(start_in[428]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[429]) );
  DFF \start_reg_reg[430]  ( .D(start_in[429]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[430]) );
  DFF \start_reg_reg[431]  ( .D(start_in[430]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[431]) );
  DFF \start_reg_reg[432]  ( .D(start_in[431]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[432]) );
  DFF \start_reg_reg[433]  ( .D(start_in[432]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[433]) );
  DFF \start_reg_reg[434]  ( .D(start_in[433]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[434]) );
  DFF \start_reg_reg[435]  ( .D(start_in[434]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[435]) );
  DFF \start_reg_reg[436]  ( .D(start_in[435]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[436]) );
  DFF \start_reg_reg[437]  ( .D(start_in[436]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[437]) );
  DFF \start_reg_reg[438]  ( .D(start_in[437]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[438]) );
  DFF \start_reg_reg[439]  ( .D(start_in[438]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[439]) );
  DFF \start_reg_reg[440]  ( .D(start_in[439]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[440]) );
  DFF \start_reg_reg[441]  ( .D(start_in[440]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[441]) );
  DFF \start_reg_reg[442]  ( .D(start_in[441]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[442]) );
  DFF \start_reg_reg[443]  ( .D(start_in[442]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[443]) );
  DFF \start_reg_reg[444]  ( .D(start_in[443]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[444]) );
  DFF \start_reg_reg[445]  ( .D(start_in[444]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[445]) );
  DFF \start_reg_reg[446]  ( .D(start_in[445]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[446]) );
  DFF \start_reg_reg[447]  ( .D(start_in[446]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[447]) );
  DFF \start_reg_reg[448]  ( .D(start_in[447]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[448]) );
  DFF \start_reg_reg[449]  ( .D(start_in[448]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[449]) );
  DFF \start_reg_reg[450]  ( .D(start_in[449]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[450]) );
  DFF \start_reg_reg[451]  ( .D(start_in[450]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[451]) );
  DFF \start_reg_reg[452]  ( .D(start_in[451]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[452]) );
  DFF \start_reg_reg[453]  ( .D(start_in[452]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[453]) );
  DFF \start_reg_reg[454]  ( .D(start_in[453]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[454]) );
  DFF \start_reg_reg[455]  ( .D(start_in[454]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[455]) );
  DFF \start_reg_reg[456]  ( .D(start_in[455]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[456]) );
  DFF \start_reg_reg[457]  ( .D(start_in[456]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[457]) );
  DFF \start_reg_reg[458]  ( .D(start_in[457]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[458]) );
  DFF \start_reg_reg[459]  ( .D(start_in[458]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[459]) );
  DFF \start_reg_reg[460]  ( .D(start_in[459]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[460]) );
  DFF \start_reg_reg[461]  ( .D(start_in[460]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[461]) );
  DFF \start_reg_reg[462]  ( .D(start_in[461]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[462]) );
  DFF \start_reg_reg[463]  ( .D(start_in[462]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[463]) );
  DFF \start_reg_reg[464]  ( .D(start_in[463]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[464]) );
  DFF \start_reg_reg[465]  ( .D(start_in[464]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[465]) );
  DFF \start_reg_reg[466]  ( .D(start_in[465]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[466]) );
  DFF \start_reg_reg[467]  ( .D(start_in[466]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[467]) );
  DFF \start_reg_reg[468]  ( .D(start_in[467]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[468]) );
  DFF \start_reg_reg[469]  ( .D(start_in[468]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[469]) );
  DFF \start_reg_reg[470]  ( .D(start_in[469]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[470]) );
  DFF \start_reg_reg[471]  ( .D(start_in[470]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[471]) );
  DFF \start_reg_reg[472]  ( .D(start_in[471]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[472]) );
  DFF \start_reg_reg[473]  ( .D(start_in[472]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[473]) );
  DFF \start_reg_reg[474]  ( .D(start_in[473]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[474]) );
  DFF \start_reg_reg[475]  ( .D(start_in[474]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[475]) );
  DFF \start_reg_reg[476]  ( .D(start_in[475]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[476]) );
  DFF \start_reg_reg[477]  ( .D(start_in[476]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[477]) );
  DFF \start_reg_reg[478]  ( .D(start_in[477]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[478]) );
  DFF \start_reg_reg[479]  ( .D(start_in[478]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[479]) );
  DFF \start_reg_reg[480]  ( .D(start_in[479]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[480]) );
  DFF \start_reg_reg[481]  ( .D(start_in[480]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[481]) );
  DFF \start_reg_reg[482]  ( .D(start_in[481]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[482]) );
  DFF \start_reg_reg[483]  ( .D(start_in[482]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[483]) );
  DFF \start_reg_reg[484]  ( .D(start_in[483]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[484]) );
  DFF \start_reg_reg[485]  ( .D(start_in[484]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[485]) );
  DFF \start_reg_reg[486]  ( .D(start_in[485]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[486]) );
  DFF \start_reg_reg[487]  ( .D(start_in[486]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[487]) );
  DFF \start_reg_reg[488]  ( .D(start_in[487]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[488]) );
  DFF \start_reg_reg[489]  ( .D(start_in[488]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[489]) );
  DFF \start_reg_reg[490]  ( .D(start_in[489]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[490]) );
  DFF \start_reg_reg[491]  ( .D(start_in[490]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[491]) );
  DFF \start_reg_reg[492]  ( .D(start_in[491]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[492]) );
  DFF \start_reg_reg[493]  ( .D(start_in[492]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[493]) );
  DFF \start_reg_reg[494]  ( .D(start_in[493]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[494]) );
  DFF \start_reg_reg[495]  ( .D(start_in[494]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[495]) );
  DFF \start_reg_reg[496]  ( .D(start_in[495]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[496]) );
  DFF \start_reg_reg[497]  ( .D(start_in[496]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[497]) );
  DFF \start_reg_reg[498]  ( .D(start_in[497]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[498]) );
  DFF \start_reg_reg[499]  ( .D(start_in[498]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[499]) );
  DFF \start_reg_reg[500]  ( .D(start_in[499]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[500]) );
  DFF \start_reg_reg[501]  ( .D(start_in[500]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[501]) );
  DFF \start_reg_reg[502]  ( .D(start_in[501]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[502]) );
  DFF \start_reg_reg[503]  ( .D(start_in[502]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[503]) );
  DFF \start_reg_reg[504]  ( .D(start_in[503]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[504]) );
  DFF \start_reg_reg[505]  ( .D(start_in[504]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[505]) );
  DFF \start_reg_reg[506]  ( .D(start_in[505]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[506]) );
  DFF \start_reg_reg[507]  ( .D(start_in[506]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[507]) );
  DFF \start_reg_reg[508]  ( .D(start_in[507]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[508]) );
  DFF \start_reg_reg[509]  ( .D(start_in[508]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[509]) );
  DFF \start_reg_reg[510]  ( .D(start_in[509]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[510]) );
  DFF \start_reg_reg[511]  ( .D(start_in[510]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[511]) );
  DFF mul_pow_reg ( .D(n8), .CLK(clk), .RST(rst), .I(1'b0), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(ereg_next[0]), .CLK(clk), .RST(rst), .I(e[0]), .Q(
        ein[0]) );
  DFF \ereg_reg[1]  ( .D(ereg_next[1]), .CLK(clk), .RST(rst), .I(e[1]), .Q(
        ein[1]) );
  DFF \ereg_reg[2]  ( .D(ereg_next[2]), .CLK(clk), .RST(rst), .I(e[2]), .Q(
        ein[2]) );
  DFF \ereg_reg[3]  ( .D(ereg_next[3]), .CLK(clk), .RST(rst), .I(e[3]), .Q(
        ein[3]) );
  DFF \ereg_reg[4]  ( .D(ereg_next[4]), .CLK(clk), .RST(rst), .I(e[4]), .Q(
        ein[4]) );
  DFF \ereg_reg[5]  ( .D(ereg_next[5]), .CLK(clk), .RST(rst), .I(e[5]), .Q(
        ein[5]) );
  DFF \ereg_reg[6]  ( .D(ereg_next[6]), .CLK(clk), .RST(rst), .I(e[6]), .Q(
        ein[6]) );
  DFF \ereg_reg[7]  ( .D(ereg_next[7]), .CLK(clk), .RST(rst), .I(e[7]), .Q(
        ein[7]) );
  DFF \ereg_reg[8]  ( .D(ereg_next[8]), .CLK(clk), .RST(rst), .I(e[8]), .Q(
        ein[8]) );
  DFF \ereg_reg[9]  ( .D(ereg_next[9]), .CLK(clk), .RST(rst), .I(e[9]), .Q(
        ein[9]) );
  DFF \ereg_reg[10]  ( .D(ereg_next[10]), .CLK(clk), .RST(rst), .I(e[10]), .Q(
        ein[10]) );
  DFF \ereg_reg[11]  ( .D(ereg_next[11]), .CLK(clk), .RST(rst), .I(e[11]), .Q(
        ein[11]) );
  DFF \ereg_reg[12]  ( .D(ereg_next[12]), .CLK(clk), .RST(rst), .I(e[12]), .Q(
        ein[12]) );
  DFF \ereg_reg[13]  ( .D(ereg_next[13]), .CLK(clk), .RST(rst), .I(e[13]), .Q(
        ein[13]) );
  DFF \ereg_reg[14]  ( .D(ereg_next[14]), .CLK(clk), .RST(rst), .I(e[14]), .Q(
        ein[14]) );
  DFF \ereg_reg[15]  ( .D(ereg_next[15]), .CLK(clk), .RST(rst), .I(e[15]), .Q(
        ein[15]) );
  DFF \ereg_reg[16]  ( .D(ereg_next[16]), .CLK(clk), .RST(rst), .I(e[16]), .Q(
        ein[16]) );
  DFF \ereg_reg[17]  ( .D(ereg_next[17]), .CLK(clk), .RST(rst), .I(e[17]), .Q(
        ein[17]) );
  DFF \ereg_reg[18]  ( .D(ereg_next[18]), .CLK(clk), .RST(rst), .I(e[18]), .Q(
        ein[18]) );
  DFF \ereg_reg[19]  ( .D(ereg_next[19]), .CLK(clk), .RST(rst), .I(e[19]), .Q(
        ein[19]) );
  DFF \ereg_reg[20]  ( .D(ereg_next[20]), .CLK(clk), .RST(rst), .I(e[20]), .Q(
        ein[20]) );
  DFF \ereg_reg[21]  ( .D(ereg_next[21]), .CLK(clk), .RST(rst), .I(e[21]), .Q(
        ein[21]) );
  DFF \ereg_reg[22]  ( .D(ereg_next[22]), .CLK(clk), .RST(rst), .I(e[22]), .Q(
        ein[22]) );
  DFF \ereg_reg[23]  ( .D(ereg_next[23]), .CLK(clk), .RST(rst), .I(e[23]), .Q(
        ein[23]) );
  DFF \ereg_reg[24]  ( .D(ereg_next[24]), .CLK(clk), .RST(rst), .I(e[24]), .Q(
        ein[24]) );
  DFF \ereg_reg[25]  ( .D(ereg_next[25]), .CLK(clk), .RST(rst), .I(e[25]), .Q(
        ein[25]) );
  DFF \ereg_reg[26]  ( .D(ereg_next[26]), .CLK(clk), .RST(rst), .I(e[26]), .Q(
        ein[26]) );
  DFF \ereg_reg[27]  ( .D(ereg_next[27]), .CLK(clk), .RST(rst), .I(e[27]), .Q(
        ein[27]) );
  DFF \ereg_reg[28]  ( .D(ereg_next[28]), .CLK(clk), .RST(rst), .I(e[28]), .Q(
        ein[28]) );
  DFF \ereg_reg[29]  ( .D(ereg_next[29]), .CLK(clk), .RST(rst), .I(e[29]), .Q(
        ein[29]) );
  DFF \ereg_reg[30]  ( .D(ereg_next[30]), .CLK(clk), .RST(rst), .I(e[30]), .Q(
        ein[30]) );
  DFF \ereg_reg[31]  ( .D(ereg_next[31]), .CLK(clk), .RST(rst), .I(e[31]), .Q(
        ein[31]) );
  DFF \ereg_reg[32]  ( .D(ereg_next[32]), .CLK(clk), .RST(rst), .I(e[32]), .Q(
        ein[32]) );
  DFF \ereg_reg[33]  ( .D(ereg_next[33]), .CLK(clk), .RST(rst), .I(e[33]), .Q(
        ein[33]) );
  DFF \ereg_reg[34]  ( .D(ereg_next[34]), .CLK(clk), .RST(rst), .I(e[34]), .Q(
        ein[34]) );
  DFF \ereg_reg[35]  ( .D(ereg_next[35]), .CLK(clk), .RST(rst), .I(e[35]), .Q(
        ein[35]) );
  DFF \ereg_reg[36]  ( .D(ereg_next[36]), .CLK(clk), .RST(rst), .I(e[36]), .Q(
        ein[36]) );
  DFF \ereg_reg[37]  ( .D(ereg_next[37]), .CLK(clk), .RST(rst), .I(e[37]), .Q(
        ein[37]) );
  DFF \ereg_reg[38]  ( .D(ereg_next[38]), .CLK(clk), .RST(rst), .I(e[38]), .Q(
        ein[38]) );
  DFF \ereg_reg[39]  ( .D(ereg_next[39]), .CLK(clk), .RST(rst), .I(e[39]), .Q(
        ein[39]) );
  DFF \ereg_reg[40]  ( .D(ereg_next[40]), .CLK(clk), .RST(rst), .I(e[40]), .Q(
        ein[40]) );
  DFF \ereg_reg[41]  ( .D(ereg_next[41]), .CLK(clk), .RST(rst), .I(e[41]), .Q(
        ein[41]) );
  DFF \ereg_reg[42]  ( .D(ereg_next[42]), .CLK(clk), .RST(rst), .I(e[42]), .Q(
        ein[42]) );
  DFF \ereg_reg[43]  ( .D(ereg_next[43]), .CLK(clk), .RST(rst), .I(e[43]), .Q(
        ein[43]) );
  DFF \ereg_reg[44]  ( .D(ereg_next[44]), .CLK(clk), .RST(rst), .I(e[44]), .Q(
        ein[44]) );
  DFF \ereg_reg[45]  ( .D(ereg_next[45]), .CLK(clk), .RST(rst), .I(e[45]), .Q(
        ein[45]) );
  DFF \ereg_reg[46]  ( .D(ereg_next[46]), .CLK(clk), .RST(rst), .I(e[46]), .Q(
        ein[46]) );
  DFF \ereg_reg[47]  ( .D(ereg_next[47]), .CLK(clk), .RST(rst), .I(e[47]), .Q(
        ein[47]) );
  DFF \ereg_reg[48]  ( .D(ereg_next[48]), .CLK(clk), .RST(rst), .I(e[48]), .Q(
        ein[48]) );
  DFF \ereg_reg[49]  ( .D(ereg_next[49]), .CLK(clk), .RST(rst), .I(e[49]), .Q(
        ein[49]) );
  DFF \ereg_reg[50]  ( .D(ereg_next[50]), .CLK(clk), .RST(rst), .I(e[50]), .Q(
        ein[50]) );
  DFF \ereg_reg[51]  ( .D(ereg_next[51]), .CLK(clk), .RST(rst), .I(e[51]), .Q(
        ein[51]) );
  DFF \ereg_reg[52]  ( .D(ereg_next[52]), .CLK(clk), .RST(rst), .I(e[52]), .Q(
        ein[52]) );
  DFF \ereg_reg[53]  ( .D(ereg_next[53]), .CLK(clk), .RST(rst), .I(e[53]), .Q(
        ein[53]) );
  DFF \ereg_reg[54]  ( .D(ereg_next[54]), .CLK(clk), .RST(rst), .I(e[54]), .Q(
        ein[54]) );
  DFF \ereg_reg[55]  ( .D(ereg_next[55]), .CLK(clk), .RST(rst), .I(e[55]), .Q(
        ein[55]) );
  DFF \ereg_reg[56]  ( .D(ereg_next[56]), .CLK(clk), .RST(rst), .I(e[56]), .Q(
        ein[56]) );
  DFF \ereg_reg[57]  ( .D(ereg_next[57]), .CLK(clk), .RST(rst), .I(e[57]), .Q(
        ein[57]) );
  DFF \ereg_reg[58]  ( .D(ereg_next[58]), .CLK(clk), .RST(rst), .I(e[58]), .Q(
        ein[58]) );
  DFF \ereg_reg[59]  ( .D(ereg_next[59]), .CLK(clk), .RST(rst), .I(e[59]), .Q(
        ein[59]) );
  DFF \ereg_reg[60]  ( .D(ereg_next[60]), .CLK(clk), .RST(rst), .I(e[60]), .Q(
        ein[60]) );
  DFF \ereg_reg[61]  ( .D(ereg_next[61]), .CLK(clk), .RST(rst), .I(e[61]), .Q(
        ein[61]) );
  DFF \ereg_reg[62]  ( .D(ereg_next[62]), .CLK(clk), .RST(rst), .I(e[62]), .Q(
        ein[62]) );
  DFF \ereg_reg[63]  ( .D(ereg_next[63]), .CLK(clk), .RST(rst), .I(e[63]), .Q(
        ein[63]) );
  DFF \ereg_reg[64]  ( .D(ereg_next[64]), .CLK(clk), .RST(rst), .I(e[64]), .Q(
        ein[64]) );
  DFF \ereg_reg[65]  ( .D(ereg_next[65]), .CLK(clk), .RST(rst), .I(e[65]), .Q(
        ein[65]) );
  DFF \ereg_reg[66]  ( .D(ereg_next[66]), .CLK(clk), .RST(rst), .I(e[66]), .Q(
        ein[66]) );
  DFF \ereg_reg[67]  ( .D(ereg_next[67]), .CLK(clk), .RST(rst), .I(e[67]), .Q(
        ein[67]) );
  DFF \ereg_reg[68]  ( .D(ereg_next[68]), .CLK(clk), .RST(rst), .I(e[68]), .Q(
        ein[68]) );
  DFF \ereg_reg[69]  ( .D(ereg_next[69]), .CLK(clk), .RST(rst), .I(e[69]), .Q(
        ein[69]) );
  DFF \ereg_reg[70]  ( .D(ereg_next[70]), .CLK(clk), .RST(rst), .I(e[70]), .Q(
        ein[70]) );
  DFF \ereg_reg[71]  ( .D(ereg_next[71]), .CLK(clk), .RST(rst), .I(e[71]), .Q(
        ein[71]) );
  DFF \ereg_reg[72]  ( .D(ereg_next[72]), .CLK(clk), .RST(rst), .I(e[72]), .Q(
        ein[72]) );
  DFF \ereg_reg[73]  ( .D(ereg_next[73]), .CLK(clk), .RST(rst), .I(e[73]), .Q(
        ein[73]) );
  DFF \ereg_reg[74]  ( .D(ereg_next[74]), .CLK(clk), .RST(rst), .I(e[74]), .Q(
        ein[74]) );
  DFF \ereg_reg[75]  ( .D(ereg_next[75]), .CLK(clk), .RST(rst), .I(e[75]), .Q(
        ein[75]) );
  DFF \ereg_reg[76]  ( .D(ereg_next[76]), .CLK(clk), .RST(rst), .I(e[76]), .Q(
        ein[76]) );
  DFF \ereg_reg[77]  ( .D(ereg_next[77]), .CLK(clk), .RST(rst), .I(e[77]), .Q(
        ein[77]) );
  DFF \ereg_reg[78]  ( .D(ereg_next[78]), .CLK(clk), .RST(rst), .I(e[78]), .Q(
        ein[78]) );
  DFF \ereg_reg[79]  ( .D(ereg_next[79]), .CLK(clk), .RST(rst), .I(e[79]), .Q(
        ein[79]) );
  DFF \ereg_reg[80]  ( .D(ereg_next[80]), .CLK(clk), .RST(rst), .I(e[80]), .Q(
        ein[80]) );
  DFF \ereg_reg[81]  ( .D(ereg_next[81]), .CLK(clk), .RST(rst), .I(e[81]), .Q(
        ein[81]) );
  DFF \ereg_reg[82]  ( .D(ereg_next[82]), .CLK(clk), .RST(rst), .I(e[82]), .Q(
        ein[82]) );
  DFF \ereg_reg[83]  ( .D(ereg_next[83]), .CLK(clk), .RST(rst), .I(e[83]), .Q(
        ein[83]) );
  DFF \ereg_reg[84]  ( .D(ereg_next[84]), .CLK(clk), .RST(rst), .I(e[84]), .Q(
        ein[84]) );
  DFF \ereg_reg[85]  ( .D(ereg_next[85]), .CLK(clk), .RST(rst), .I(e[85]), .Q(
        ein[85]) );
  DFF \ereg_reg[86]  ( .D(ereg_next[86]), .CLK(clk), .RST(rst), .I(e[86]), .Q(
        ein[86]) );
  DFF \ereg_reg[87]  ( .D(ereg_next[87]), .CLK(clk), .RST(rst), .I(e[87]), .Q(
        ein[87]) );
  DFF \ereg_reg[88]  ( .D(ereg_next[88]), .CLK(clk), .RST(rst), .I(e[88]), .Q(
        ein[88]) );
  DFF \ereg_reg[89]  ( .D(ereg_next[89]), .CLK(clk), .RST(rst), .I(e[89]), .Q(
        ein[89]) );
  DFF \ereg_reg[90]  ( .D(ereg_next[90]), .CLK(clk), .RST(rst), .I(e[90]), .Q(
        ein[90]) );
  DFF \ereg_reg[91]  ( .D(ereg_next[91]), .CLK(clk), .RST(rst), .I(e[91]), .Q(
        ein[91]) );
  DFF \ereg_reg[92]  ( .D(ereg_next[92]), .CLK(clk), .RST(rst), .I(e[92]), .Q(
        ein[92]) );
  DFF \ereg_reg[93]  ( .D(ereg_next[93]), .CLK(clk), .RST(rst), .I(e[93]), .Q(
        ein[93]) );
  DFF \ereg_reg[94]  ( .D(ereg_next[94]), .CLK(clk), .RST(rst), .I(e[94]), .Q(
        ein[94]) );
  DFF \ereg_reg[95]  ( .D(ereg_next[95]), .CLK(clk), .RST(rst), .I(e[95]), .Q(
        ein[95]) );
  DFF \ereg_reg[96]  ( .D(ereg_next[96]), .CLK(clk), .RST(rst), .I(e[96]), .Q(
        ein[96]) );
  DFF \ereg_reg[97]  ( .D(ereg_next[97]), .CLK(clk), .RST(rst), .I(e[97]), .Q(
        ein[97]) );
  DFF \ereg_reg[98]  ( .D(ereg_next[98]), .CLK(clk), .RST(rst), .I(e[98]), .Q(
        ein[98]) );
  DFF \ereg_reg[99]  ( .D(ereg_next[99]), .CLK(clk), .RST(rst), .I(e[99]), .Q(
        ein[99]) );
  DFF \ereg_reg[100]  ( .D(ereg_next[100]), .CLK(clk), .RST(rst), .I(e[100]), 
        .Q(ein[100]) );
  DFF \ereg_reg[101]  ( .D(ereg_next[101]), .CLK(clk), .RST(rst), .I(e[101]), 
        .Q(ein[101]) );
  DFF \ereg_reg[102]  ( .D(ereg_next[102]), .CLK(clk), .RST(rst), .I(e[102]), 
        .Q(ein[102]) );
  DFF \ereg_reg[103]  ( .D(ereg_next[103]), .CLK(clk), .RST(rst), .I(e[103]), 
        .Q(ein[103]) );
  DFF \ereg_reg[104]  ( .D(ereg_next[104]), .CLK(clk), .RST(rst), .I(e[104]), 
        .Q(ein[104]) );
  DFF \ereg_reg[105]  ( .D(ereg_next[105]), .CLK(clk), .RST(rst), .I(e[105]), 
        .Q(ein[105]) );
  DFF \ereg_reg[106]  ( .D(ereg_next[106]), .CLK(clk), .RST(rst), .I(e[106]), 
        .Q(ein[106]) );
  DFF \ereg_reg[107]  ( .D(ereg_next[107]), .CLK(clk), .RST(rst), .I(e[107]), 
        .Q(ein[107]) );
  DFF \ereg_reg[108]  ( .D(ereg_next[108]), .CLK(clk), .RST(rst), .I(e[108]), 
        .Q(ein[108]) );
  DFF \ereg_reg[109]  ( .D(ereg_next[109]), .CLK(clk), .RST(rst), .I(e[109]), 
        .Q(ein[109]) );
  DFF \ereg_reg[110]  ( .D(ereg_next[110]), .CLK(clk), .RST(rst), .I(e[110]), 
        .Q(ein[110]) );
  DFF \ereg_reg[111]  ( .D(ereg_next[111]), .CLK(clk), .RST(rst), .I(e[111]), 
        .Q(ein[111]) );
  DFF \ereg_reg[112]  ( .D(ereg_next[112]), .CLK(clk), .RST(rst), .I(e[112]), 
        .Q(ein[112]) );
  DFF \ereg_reg[113]  ( .D(ereg_next[113]), .CLK(clk), .RST(rst), .I(e[113]), 
        .Q(ein[113]) );
  DFF \ereg_reg[114]  ( .D(ereg_next[114]), .CLK(clk), .RST(rst), .I(e[114]), 
        .Q(ein[114]) );
  DFF \ereg_reg[115]  ( .D(ereg_next[115]), .CLK(clk), .RST(rst), .I(e[115]), 
        .Q(ein[115]) );
  DFF \ereg_reg[116]  ( .D(ereg_next[116]), .CLK(clk), .RST(rst), .I(e[116]), 
        .Q(ein[116]) );
  DFF \ereg_reg[117]  ( .D(ereg_next[117]), .CLK(clk), .RST(rst), .I(e[117]), 
        .Q(ein[117]) );
  DFF \ereg_reg[118]  ( .D(ereg_next[118]), .CLK(clk), .RST(rst), .I(e[118]), 
        .Q(ein[118]) );
  DFF \ereg_reg[119]  ( .D(ereg_next[119]), .CLK(clk), .RST(rst), .I(e[119]), 
        .Q(ein[119]) );
  DFF \ereg_reg[120]  ( .D(ereg_next[120]), .CLK(clk), .RST(rst), .I(e[120]), 
        .Q(ein[120]) );
  DFF \ereg_reg[121]  ( .D(ereg_next[121]), .CLK(clk), .RST(rst), .I(e[121]), 
        .Q(ein[121]) );
  DFF \ereg_reg[122]  ( .D(ereg_next[122]), .CLK(clk), .RST(rst), .I(e[122]), 
        .Q(ein[122]) );
  DFF \ereg_reg[123]  ( .D(ereg_next[123]), .CLK(clk), .RST(rst), .I(e[123]), 
        .Q(ein[123]) );
  DFF \ereg_reg[124]  ( .D(ereg_next[124]), .CLK(clk), .RST(rst), .I(e[124]), 
        .Q(ein[124]) );
  DFF \ereg_reg[125]  ( .D(ereg_next[125]), .CLK(clk), .RST(rst), .I(e[125]), 
        .Q(ein[125]) );
  DFF \ereg_reg[126]  ( .D(ereg_next[126]), .CLK(clk), .RST(rst), .I(e[126]), 
        .Q(ein[126]) );
  DFF \ereg_reg[127]  ( .D(ereg_next[127]), .CLK(clk), .RST(rst), .I(e[127]), 
        .Q(ein[127]) );
  DFF \ereg_reg[128]  ( .D(ereg_next[128]), .CLK(clk), .RST(rst), .I(e[128]), 
        .Q(ein[128]) );
  DFF \ereg_reg[129]  ( .D(ereg_next[129]), .CLK(clk), .RST(rst), .I(e[129]), 
        .Q(ein[129]) );
  DFF \ereg_reg[130]  ( .D(ereg_next[130]), .CLK(clk), .RST(rst), .I(e[130]), 
        .Q(ein[130]) );
  DFF \ereg_reg[131]  ( .D(ereg_next[131]), .CLK(clk), .RST(rst), .I(e[131]), 
        .Q(ein[131]) );
  DFF \ereg_reg[132]  ( .D(ereg_next[132]), .CLK(clk), .RST(rst), .I(e[132]), 
        .Q(ein[132]) );
  DFF \ereg_reg[133]  ( .D(ereg_next[133]), .CLK(clk), .RST(rst), .I(e[133]), 
        .Q(ein[133]) );
  DFF \ereg_reg[134]  ( .D(ereg_next[134]), .CLK(clk), .RST(rst), .I(e[134]), 
        .Q(ein[134]) );
  DFF \ereg_reg[135]  ( .D(ereg_next[135]), .CLK(clk), .RST(rst), .I(e[135]), 
        .Q(ein[135]) );
  DFF \ereg_reg[136]  ( .D(ereg_next[136]), .CLK(clk), .RST(rst), .I(e[136]), 
        .Q(ein[136]) );
  DFF \ereg_reg[137]  ( .D(ereg_next[137]), .CLK(clk), .RST(rst), .I(e[137]), 
        .Q(ein[137]) );
  DFF \ereg_reg[138]  ( .D(ereg_next[138]), .CLK(clk), .RST(rst), .I(e[138]), 
        .Q(ein[138]) );
  DFF \ereg_reg[139]  ( .D(ereg_next[139]), .CLK(clk), .RST(rst), .I(e[139]), 
        .Q(ein[139]) );
  DFF \ereg_reg[140]  ( .D(ereg_next[140]), .CLK(clk), .RST(rst), .I(e[140]), 
        .Q(ein[140]) );
  DFF \ereg_reg[141]  ( .D(ereg_next[141]), .CLK(clk), .RST(rst), .I(e[141]), 
        .Q(ein[141]) );
  DFF \ereg_reg[142]  ( .D(ereg_next[142]), .CLK(clk), .RST(rst), .I(e[142]), 
        .Q(ein[142]) );
  DFF \ereg_reg[143]  ( .D(ereg_next[143]), .CLK(clk), .RST(rst), .I(e[143]), 
        .Q(ein[143]) );
  DFF \ereg_reg[144]  ( .D(ereg_next[144]), .CLK(clk), .RST(rst), .I(e[144]), 
        .Q(ein[144]) );
  DFF \ereg_reg[145]  ( .D(ereg_next[145]), .CLK(clk), .RST(rst), .I(e[145]), 
        .Q(ein[145]) );
  DFF \ereg_reg[146]  ( .D(ereg_next[146]), .CLK(clk), .RST(rst), .I(e[146]), 
        .Q(ein[146]) );
  DFF \ereg_reg[147]  ( .D(ereg_next[147]), .CLK(clk), .RST(rst), .I(e[147]), 
        .Q(ein[147]) );
  DFF \ereg_reg[148]  ( .D(ereg_next[148]), .CLK(clk), .RST(rst), .I(e[148]), 
        .Q(ein[148]) );
  DFF \ereg_reg[149]  ( .D(ereg_next[149]), .CLK(clk), .RST(rst), .I(e[149]), 
        .Q(ein[149]) );
  DFF \ereg_reg[150]  ( .D(ereg_next[150]), .CLK(clk), .RST(rst), .I(e[150]), 
        .Q(ein[150]) );
  DFF \ereg_reg[151]  ( .D(ereg_next[151]), .CLK(clk), .RST(rst), .I(e[151]), 
        .Q(ein[151]) );
  DFF \ereg_reg[152]  ( .D(ereg_next[152]), .CLK(clk), .RST(rst), .I(e[152]), 
        .Q(ein[152]) );
  DFF \ereg_reg[153]  ( .D(ereg_next[153]), .CLK(clk), .RST(rst), .I(e[153]), 
        .Q(ein[153]) );
  DFF \ereg_reg[154]  ( .D(ereg_next[154]), .CLK(clk), .RST(rst), .I(e[154]), 
        .Q(ein[154]) );
  DFF \ereg_reg[155]  ( .D(ereg_next[155]), .CLK(clk), .RST(rst), .I(e[155]), 
        .Q(ein[155]) );
  DFF \ereg_reg[156]  ( .D(ereg_next[156]), .CLK(clk), .RST(rst), .I(e[156]), 
        .Q(ein[156]) );
  DFF \ereg_reg[157]  ( .D(ereg_next[157]), .CLK(clk), .RST(rst), .I(e[157]), 
        .Q(ein[157]) );
  DFF \ereg_reg[158]  ( .D(ereg_next[158]), .CLK(clk), .RST(rst), .I(e[158]), 
        .Q(ein[158]) );
  DFF \ereg_reg[159]  ( .D(ereg_next[159]), .CLK(clk), .RST(rst), .I(e[159]), 
        .Q(ein[159]) );
  DFF \ereg_reg[160]  ( .D(ereg_next[160]), .CLK(clk), .RST(rst), .I(e[160]), 
        .Q(ein[160]) );
  DFF \ereg_reg[161]  ( .D(ereg_next[161]), .CLK(clk), .RST(rst), .I(e[161]), 
        .Q(ein[161]) );
  DFF \ereg_reg[162]  ( .D(ereg_next[162]), .CLK(clk), .RST(rst), .I(e[162]), 
        .Q(ein[162]) );
  DFF \ereg_reg[163]  ( .D(ereg_next[163]), .CLK(clk), .RST(rst), .I(e[163]), 
        .Q(ein[163]) );
  DFF \ereg_reg[164]  ( .D(ereg_next[164]), .CLK(clk), .RST(rst), .I(e[164]), 
        .Q(ein[164]) );
  DFF \ereg_reg[165]  ( .D(ereg_next[165]), .CLK(clk), .RST(rst), .I(e[165]), 
        .Q(ein[165]) );
  DFF \ereg_reg[166]  ( .D(ereg_next[166]), .CLK(clk), .RST(rst), .I(e[166]), 
        .Q(ein[166]) );
  DFF \ereg_reg[167]  ( .D(ereg_next[167]), .CLK(clk), .RST(rst), .I(e[167]), 
        .Q(ein[167]) );
  DFF \ereg_reg[168]  ( .D(ereg_next[168]), .CLK(clk), .RST(rst), .I(e[168]), 
        .Q(ein[168]) );
  DFF \ereg_reg[169]  ( .D(ereg_next[169]), .CLK(clk), .RST(rst), .I(e[169]), 
        .Q(ein[169]) );
  DFF \ereg_reg[170]  ( .D(ereg_next[170]), .CLK(clk), .RST(rst), .I(e[170]), 
        .Q(ein[170]) );
  DFF \ereg_reg[171]  ( .D(ereg_next[171]), .CLK(clk), .RST(rst), .I(e[171]), 
        .Q(ein[171]) );
  DFF \ereg_reg[172]  ( .D(ereg_next[172]), .CLK(clk), .RST(rst), .I(e[172]), 
        .Q(ein[172]) );
  DFF \ereg_reg[173]  ( .D(ereg_next[173]), .CLK(clk), .RST(rst), .I(e[173]), 
        .Q(ein[173]) );
  DFF \ereg_reg[174]  ( .D(ereg_next[174]), .CLK(clk), .RST(rst), .I(e[174]), 
        .Q(ein[174]) );
  DFF \ereg_reg[175]  ( .D(ereg_next[175]), .CLK(clk), .RST(rst), .I(e[175]), 
        .Q(ein[175]) );
  DFF \ereg_reg[176]  ( .D(ereg_next[176]), .CLK(clk), .RST(rst), .I(e[176]), 
        .Q(ein[176]) );
  DFF \ereg_reg[177]  ( .D(ereg_next[177]), .CLK(clk), .RST(rst), .I(e[177]), 
        .Q(ein[177]) );
  DFF \ereg_reg[178]  ( .D(ereg_next[178]), .CLK(clk), .RST(rst), .I(e[178]), 
        .Q(ein[178]) );
  DFF \ereg_reg[179]  ( .D(ereg_next[179]), .CLK(clk), .RST(rst), .I(e[179]), 
        .Q(ein[179]) );
  DFF \ereg_reg[180]  ( .D(ereg_next[180]), .CLK(clk), .RST(rst), .I(e[180]), 
        .Q(ein[180]) );
  DFF \ereg_reg[181]  ( .D(ereg_next[181]), .CLK(clk), .RST(rst), .I(e[181]), 
        .Q(ein[181]) );
  DFF \ereg_reg[182]  ( .D(ereg_next[182]), .CLK(clk), .RST(rst), .I(e[182]), 
        .Q(ein[182]) );
  DFF \ereg_reg[183]  ( .D(ereg_next[183]), .CLK(clk), .RST(rst), .I(e[183]), 
        .Q(ein[183]) );
  DFF \ereg_reg[184]  ( .D(ereg_next[184]), .CLK(clk), .RST(rst), .I(e[184]), 
        .Q(ein[184]) );
  DFF \ereg_reg[185]  ( .D(ereg_next[185]), .CLK(clk), .RST(rst), .I(e[185]), 
        .Q(ein[185]) );
  DFF \ereg_reg[186]  ( .D(ereg_next[186]), .CLK(clk), .RST(rst), .I(e[186]), 
        .Q(ein[186]) );
  DFF \ereg_reg[187]  ( .D(ereg_next[187]), .CLK(clk), .RST(rst), .I(e[187]), 
        .Q(ein[187]) );
  DFF \ereg_reg[188]  ( .D(ereg_next[188]), .CLK(clk), .RST(rst), .I(e[188]), 
        .Q(ein[188]) );
  DFF \ereg_reg[189]  ( .D(ereg_next[189]), .CLK(clk), .RST(rst), .I(e[189]), 
        .Q(ein[189]) );
  DFF \ereg_reg[190]  ( .D(ereg_next[190]), .CLK(clk), .RST(rst), .I(e[190]), 
        .Q(ein[190]) );
  DFF \ereg_reg[191]  ( .D(ereg_next[191]), .CLK(clk), .RST(rst), .I(e[191]), 
        .Q(ein[191]) );
  DFF \ereg_reg[192]  ( .D(ereg_next[192]), .CLK(clk), .RST(rst), .I(e[192]), 
        .Q(ein[192]) );
  DFF \ereg_reg[193]  ( .D(ereg_next[193]), .CLK(clk), .RST(rst), .I(e[193]), 
        .Q(ein[193]) );
  DFF \ereg_reg[194]  ( .D(ereg_next[194]), .CLK(clk), .RST(rst), .I(e[194]), 
        .Q(ein[194]) );
  DFF \ereg_reg[195]  ( .D(ereg_next[195]), .CLK(clk), .RST(rst), .I(e[195]), 
        .Q(ein[195]) );
  DFF \ereg_reg[196]  ( .D(ereg_next[196]), .CLK(clk), .RST(rst), .I(e[196]), 
        .Q(ein[196]) );
  DFF \ereg_reg[197]  ( .D(ereg_next[197]), .CLK(clk), .RST(rst), .I(e[197]), 
        .Q(ein[197]) );
  DFF \ereg_reg[198]  ( .D(ereg_next[198]), .CLK(clk), .RST(rst), .I(e[198]), 
        .Q(ein[198]) );
  DFF \ereg_reg[199]  ( .D(ereg_next[199]), .CLK(clk), .RST(rst), .I(e[199]), 
        .Q(ein[199]) );
  DFF \ereg_reg[200]  ( .D(ereg_next[200]), .CLK(clk), .RST(rst), .I(e[200]), 
        .Q(ein[200]) );
  DFF \ereg_reg[201]  ( .D(ereg_next[201]), .CLK(clk), .RST(rst), .I(e[201]), 
        .Q(ein[201]) );
  DFF \ereg_reg[202]  ( .D(ereg_next[202]), .CLK(clk), .RST(rst), .I(e[202]), 
        .Q(ein[202]) );
  DFF \ereg_reg[203]  ( .D(ereg_next[203]), .CLK(clk), .RST(rst), .I(e[203]), 
        .Q(ein[203]) );
  DFF \ereg_reg[204]  ( .D(ereg_next[204]), .CLK(clk), .RST(rst), .I(e[204]), 
        .Q(ein[204]) );
  DFF \ereg_reg[205]  ( .D(ereg_next[205]), .CLK(clk), .RST(rst), .I(e[205]), 
        .Q(ein[205]) );
  DFF \ereg_reg[206]  ( .D(ereg_next[206]), .CLK(clk), .RST(rst), .I(e[206]), 
        .Q(ein[206]) );
  DFF \ereg_reg[207]  ( .D(ereg_next[207]), .CLK(clk), .RST(rst), .I(e[207]), 
        .Q(ein[207]) );
  DFF \ereg_reg[208]  ( .D(ereg_next[208]), .CLK(clk), .RST(rst), .I(e[208]), 
        .Q(ein[208]) );
  DFF \ereg_reg[209]  ( .D(ereg_next[209]), .CLK(clk), .RST(rst), .I(e[209]), 
        .Q(ein[209]) );
  DFF \ereg_reg[210]  ( .D(ereg_next[210]), .CLK(clk), .RST(rst), .I(e[210]), 
        .Q(ein[210]) );
  DFF \ereg_reg[211]  ( .D(ereg_next[211]), .CLK(clk), .RST(rst), .I(e[211]), 
        .Q(ein[211]) );
  DFF \ereg_reg[212]  ( .D(ereg_next[212]), .CLK(clk), .RST(rst), .I(e[212]), 
        .Q(ein[212]) );
  DFF \ereg_reg[213]  ( .D(ereg_next[213]), .CLK(clk), .RST(rst), .I(e[213]), 
        .Q(ein[213]) );
  DFF \ereg_reg[214]  ( .D(ereg_next[214]), .CLK(clk), .RST(rst), .I(e[214]), 
        .Q(ein[214]) );
  DFF \ereg_reg[215]  ( .D(ereg_next[215]), .CLK(clk), .RST(rst), .I(e[215]), 
        .Q(ein[215]) );
  DFF \ereg_reg[216]  ( .D(ereg_next[216]), .CLK(clk), .RST(rst), .I(e[216]), 
        .Q(ein[216]) );
  DFF \ereg_reg[217]  ( .D(ereg_next[217]), .CLK(clk), .RST(rst), .I(e[217]), 
        .Q(ein[217]) );
  DFF \ereg_reg[218]  ( .D(ereg_next[218]), .CLK(clk), .RST(rst), .I(e[218]), 
        .Q(ein[218]) );
  DFF \ereg_reg[219]  ( .D(ereg_next[219]), .CLK(clk), .RST(rst), .I(e[219]), 
        .Q(ein[219]) );
  DFF \ereg_reg[220]  ( .D(ereg_next[220]), .CLK(clk), .RST(rst), .I(e[220]), 
        .Q(ein[220]) );
  DFF \ereg_reg[221]  ( .D(ereg_next[221]), .CLK(clk), .RST(rst), .I(e[221]), 
        .Q(ein[221]) );
  DFF \ereg_reg[222]  ( .D(ereg_next[222]), .CLK(clk), .RST(rst), .I(e[222]), 
        .Q(ein[222]) );
  DFF \ereg_reg[223]  ( .D(ereg_next[223]), .CLK(clk), .RST(rst), .I(e[223]), 
        .Q(ein[223]) );
  DFF \ereg_reg[224]  ( .D(ereg_next[224]), .CLK(clk), .RST(rst), .I(e[224]), 
        .Q(ein[224]) );
  DFF \ereg_reg[225]  ( .D(ereg_next[225]), .CLK(clk), .RST(rst), .I(e[225]), 
        .Q(ein[225]) );
  DFF \ereg_reg[226]  ( .D(ereg_next[226]), .CLK(clk), .RST(rst), .I(e[226]), 
        .Q(ein[226]) );
  DFF \ereg_reg[227]  ( .D(ereg_next[227]), .CLK(clk), .RST(rst), .I(e[227]), 
        .Q(ein[227]) );
  DFF \ereg_reg[228]  ( .D(ereg_next[228]), .CLK(clk), .RST(rst), .I(e[228]), 
        .Q(ein[228]) );
  DFF \ereg_reg[229]  ( .D(ereg_next[229]), .CLK(clk), .RST(rst), .I(e[229]), 
        .Q(ein[229]) );
  DFF \ereg_reg[230]  ( .D(ereg_next[230]), .CLK(clk), .RST(rst), .I(e[230]), 
        .Q(ein[230]) );
  DFF \ereg_reg[231]  ( .D(ereg_next[231]), .CLK(clk), .RST(rst), .I(e[231]), 
        .Q(ein[231]) );
  DFF \ereg_reg[232]  ( .D(ereg_next[232]), .CLK(clk), .RST(rst), .I(e[232]), 
        .Q(ein[232]) );
  DFF \ereg_reg[233]  ( .D(ereg_next[233]), .CLK(clk), .RST(rst), .I(e[233]), 
        .Q(ein[233]) );
  DFF \ereg_reg[234]  ( .D(ereg_next[234]), .CLK(clk), .RST(rst), .I(e[234]), 
        .Q(ein[234]) );
  DFF \ereg_reg[235]  ( .D(ereg_next[235]), .CLK(clk), .RST(rst), .I(e[235]), 
        .Q(ein[235]) );
  DFF \ereg_reg[236]  ( .D(ereg_next[236]), .CLK(clk), .RST(rst), .I(e[236]), 
        .Q(ein[236]) );
  DFF \ereg_reg[237]  ( .D(ereg_next[237]), .CLK(clk), .RST(rst), .I(e[237]), 
        .Q(ein[237]) );
  DFF \ereg_reg[238]  ( .D(ereg_next[238]), .CLK(clk), .RST(rst), .I(e[238]), 
        .Q(ein[238]) );
  DFF \ereg_reg[239]  ( .D(ereg_next[239]), .CLK(clk), .RST(rst), .I(e[239]), 
        .Q(ein[239]) );
  DFF \ereg_reg[240]  ( .D(ereg_next[240]), .CLK(clk), .RST(rst), .I(e[240]), 
        .Q(ein[240]) );
  DFF \ereg_reg[241]  ( .D(ereg_next[241]), .CLK(clk), .RST(rst), .I(e[241]), 
        .Q(ein[241]) );
  DFF \ereg_reg[242]  ( .D(ereg_next[242]), .CLK(clk), .RST(rst), .I(e[242]), 
        .Q(ein[242]) );
  DFF \ereg_reg[243]  ( .D(ereg_next[243]), .CLK(clk), .RST(rst), .I(e[243]), 
        .Q(ein[243]) );
  DFF \ereg_reg[244]  ( .D(ereg_next[244]), .CLK(clk), .RST(rst), .I(e[244]), 
        .Q(ein[244]) );
  DFF \ereg_reg[245]  ( .D(ereg_next[245]), .CLK(clk), .RST(rst), .I(e[245]), 
        .Q(ein[245]) );
  DFF \ereg_reg[246]  ( .D(ereg_next[246]), .CLK(clk), .RST(rst), .I(e[246]), 
        .Q(ein[246]) );
  DFF \ereg_reg[247]  ( .D(ereg_next[247]), .CLK(clk), .RST(rst), .I(e[247]), 
        .Q(ein[247]) );
  DFF \ereg_reg[248]  ( .D(ereg_next[248]), .CLK(clk), .RST(rst), .I(e[248]), 
        .Q(ein[248]) );
  DFF \ereg_reg[249]  ( .D(ereg_next[249]), .CLK(clk), .RST(rst), .I(e[249]), 
        .Q(ein[249]) );
  DFF \ereg_reg[250]  ( .D(ereg_next[250]), .CLK(clk), .RST(rst), .I(e[250]), 
        .Q(ein[250]) );
  DFF \ereg_reg[251]  ( .D(ereg_next[251]), .CLK(clk), .RST(rst), .I(e[251]), 
        .Q(ein[251]) );
  DFF \ereg_reg[252]  ( .D(ereg_next[252]), .CLK(clk), .RST(rst), .I(e[252]), 
        .Q(ein[252]) );
  DFF \ereg_reg[253]  ( .D(ereg_next[253]), .CLK(clk), .RST(rst), .I(e[253]), 
        .Q(ein[253]) );
  DFF \ereg_reg[254]  ( .D(ereg_next[254]), .CLK(clk), .RST(rst), .I(e[254]), 
        .Q(ein[254]) );
  DFF \ereg_reg[255]  ( .D(ereg_next[255]), .CLK(clk), .RST(rst), .I(e[255]), 
        .Q(ein[255]) );
  DFF \ereg_reg[256]  ( .D(ereg_next[256]), .CLK(clk), .RST(rst), .I(e[256]), 
        .Q(ein[256]) );
  DFF \ereg_reg[257]  ( .D(ereg_next[257]), .CLK(clk), .RST(rst), .I(e[257]), 
        .Q(ein[257]) );
  DFF \ereg_reg[258]  ( .D(ereg_next[258]), .CLK(clk), .RST(rst), .I(e[258]), 
        .Q(ein[258]) );
  DFF \ereg_reg[259]  ( .D(ereg_next[259]), .CLK(clk), .RST(rst), .I(e[259]), 
        .Q(ein[259]) );
  DFF \ereg_reg[260]  ( .D(ereg_next[260]), .CLK(clk), .RST(rst), .I(e[260]), 
        .Q(ein[260]) );
  DFF \ereg_reg[261]  ( .D(ereg_next[261]), .CLK(clk), .RST(rst), .I(e[261]), 
        .Q(ein[261]) );
  DFF \ereg_reg[262]  ( .D(ereg_next[262]), .CLK(clk), .RST(rst), .I(e[262]), 
        .Q(ein[262]) );
  DFF \ereg_reg[263]  ( .D(ereg_next[263]), .CLK(clk), .RST(rst), .I(e[263]), 
        .Q(ein[263]) );
  DFF \ereg_reg[264]  ( .D(ereg_next[264]), .CLK(clk), .RST(rst), .I(e[264]), 
        .Q(ein[264]) );
  DFF \ereg_reg[265]  ( .D(ereg_next[265]), .CLK(clk), .RST(rst), .I(e[265]), 
        .Q(ein[265]) );
  DFF \ereg_reg[266]  ( .D(ereg_next[266]), .CLK(clk), .RST(rst), .I(e[266]), 
        .Q(ein[266]) );
  DFF \ereg_reg[267]  ( .D(ereg_next[267]), .CLK(clk), .RST(rst), .I(e[267]), 
        .Q(ein[267]) );
  DFF \ereg_reg[268]  ( .D(ereg_next[268]), .CLK(clk), .RST(rst), .I(e[268]), 
        .Q(ein[268]) );
  DFF \ereg_reg[269]  ( .D(ereg_next[269]), .CLK(clk), .RST(rst), .I(e[269]), 
        .Q(ein[269]) );
  DFF \ereg_reg[270]  ( .D(ereg_next[270]), .CLK(clk), .RST(rst), .I(e[270]), 
        .Q(ein[270]) );
  DFF \ereg_reg[271]  ( .D(ereg_next[271]), .CLK(clk), .RST(rst), .I(e[271]), 
        .Q(ein[271]) );
  DFF \ereg_reg[272]  ( .D(ereg_next[272]), .CLK(clk), .RST(rst), .I(e[272]), 
        .Q(ein[272]) );
  DFF \ereg_reg[273]  ( .D(ereg_next[273]), .CLK(clk), .RST(rst), .I(e[273]), 
        .Q(ein[273]) );
  DFF \ereg_reg[274]  ( .D(ereg_next[274]), .CLK(clk), .RST(rst), .I(e[274]), 
        .Q(ein[274]) );
  DFF \ereg_reg[275]  ( .D(ereg_next[275]), .CLK(clk), .RST(rst), .I(e[275]), 
        .Q(ein[275]) );
  DFF \ereg_reg[276]  ( .D(ereg_next[276]), .CLK(clk), .RST(rst), .I(e[276]), 
        .Q(ein[276]) );
  DFF \ereg_reg[277]  ( .D(ereg_next[277]), .CLK(clk), .RST(rst), .I(e[277]), 
        .Q(ein[277]) );
  DFF \ereg_reg[278]  ( .D(ereg_next[278]), .CLK(clk), .RST(rst), .I(e[278]), 
        .Q(ein[278]) );
  DFF \ereg_reg[279]  ( .D(ereg_next[279]), .CLK(clk), .RST(rst), .I(e[279]), 
        .Q(ein[279]) );
  DFF \ereg_reg[280]  ( .D(ereg_next[280]), .CLK(clk), .RST(rst), .I(e[280]), 
        .Q(ein[280]) );
  DFF \ereg_reg[281]  ( .D(ereg_next[281]), .CLK(clk), .RST(rst), .I(e[281]), 
        .Q(ein[281]) );
  DFF \ereg_reg[282]  ( .D(ereg_next[282]), .CLK(clk), .RST(rst), .I(e[282]), 
        .Q(ein[282]) );
  DFF \ereg_reg[283]  ( .D(ereg_next[283]), .CLK(clk), .RST(rst), .I(e[283]), 
        .Q(ein[283]) );
  DFF \ereg_reg[284]  ( .D(ereg_next[284]), .CLK(clk), .RST(rst), .I(e[284]), 
        .Q(ein[284]) );
  DFF \ereg_reg[285]  ( .D(ereg_next[285]), .CLK(clk), .RST(rst), .I(e[285]), 
        .Q(ein[285]) );
  DFF \ereg_reg[286]  ( .D(ereg_next[286]), .CLK(clk), .RST(rst), .I(e[286]), 
        .Q(ein[286]) );
  DFF \ereg_reg[287]  ( .D(ereg_next[287]), .CLK(clk), .RST(rst), .I(e[287]), 
        .Q(ein[287]) );
  DFF \ereg_reg[288]  ( .D(ereg_next[288]), .CLK(clk), .RST(rst), .I(e[288]), 
        .Q(ein[288]) );
  DFF \ereg_reg[289]  ( .D(ereg_next[289]), .CLK(clk), .RST(rst), .I(e[289]), 
        .Q(ein[289]) );
  DFF \ereg_reg[290]  ( .D(ereg_next[290]), .CLK(clk), .RST(rst), .I(e[290]), 
        .Q(ein[290]) );
  DFF \ereg_reg[291]  ( .D(ereg_next[291]), .CLK(clk), .RST(rst), .I(e[291]), 
        .Q(ein[291]) );
  DFF \ereg_reg[292]  ( .D(ereg_next[292]), .CLK(clk), .RST(rst), .I(e[292]), 
        .Q(ein[292]) );
  DFF \ereg_reg[293]  ( .D(ereg_next[293]), .CLK(clk), .RST(rst), .I(e[293]), 
        .Q(ein[293]) );
  DFF \ereg_reg[294]  ( .D(ereg_next[294]), .CLK(clk), .RST(rst), .I(e[294]), 
        .Q(ein[294]) );
  DFF \ereg_reg[295]  ( .D(ereg_next[295]), .CLK(clk), .RST(rst), .I(e[295]), 
        .Q(ein[295]) );
  DFF \ereg_reg[296]  ( .D(ereg_next[296]), .CLK(clk), .RST(rst), .I(e[296]), 
        .Q(ein[296]) );
  DFF \ereg_reg[297]  ( .D(ereg_next[297]), .CLK(clk), .RST(rst), .I(e[297]), 
        .Q(ein[297]) );
  DFF \ereg_reg[298]  ( .D(ereg_next[298]), .CLK(clk), .RST(rst), .I(e[298]), 
        .Q(ein[298]) );
  DFF \ereg_reg[299]  ( .D(ereg_next[299]), .CLK(clk), .RST(rst), .I(e[299]), 
        .Q(ein[299]) );
  DFF \ereg_reg[300]  ( .D(ereg_next[300]), .CLK(clk), .RST(rst), .I(e[300]), 
        .Q(ein[300]) );
  DFF \ereg_reg[301]  ( .D(ereg_next[301]), .CLK(clk), .RST(rst), .I(e[301]), 
        .Q(ein[301]) );
  DFF \ereg_reg[302]  ( .D(ereg_next[302]), .CLK(clk), .RST(rst), .I(e[302]), 
        .Q(ein[302]) );
  DFF \ereg_reg[303]  ( .D(ereg_next[303]), .CLK(clk), .RST(rst), .I(e[303]), 
        .Q(ein[303]) );
  DFF \ereg_reg[304]  ( .D(ereg_next[304]), .CLK(clk), .RST(rst), .I(e[304]), 
        .Q(ein[304]) );
  DFF \ereg_reg[305]  ( .D(ereg_next[305]), .CLK(clk), .RST(rst), .I(e[305]), 
        .Q(ein[305]) );
  DFF \ereg_reg[306]  ( .D(ereg_next[306]), .CLK(clk), .RST(rst), .I(e[306]), 
        .Q(ein[306]) );
  DFF \ereg_reg[307]  ( .D(ereg_next[307]), .CLK(clk), .RST(rst), .I(e[307]), 
        .Q(ein[307]) );
  DFF \ereg_reg[308]  ( .D(ereg_next[308]), .CLK(clk), .RST(rst), .I(e[308]), 
        .Q(ein[308]) );
  DFF \ereg_reg[309]  ( .D(ereg_next[309]), .CLK(clk), .RST(rst), .I(e[309]), 
        .Q(ein[309]) );
  DFF \ereg_reg[310]  ( .D(ereg_next[310]), .CLK(clk), .RST(rst), .I(e[310]), 
        .Q(ein[310]) );
  DFF \ereg_reg[311]  ( .D(ereg_next[311]), .CLK(clk), .RST(rst), .I(e[311]), 
        .Q(ein[311]) );
  DFF \ereg_reg[312]  ( .D(ereg_next[312]), .CLK(clk), .RST(rst), .I(e[312]), 
        .Q(ein[312]) );
  DFF \ereg_reg[313]  ( .D(ereg_next[313]), .CLK(clk), .RST(rst), .I(e[313]), 
        .Q(ein[313]) );
  DFF \ereg_reg[314]  ( .D(ereg_next[314]), .CLK(clk), .RST(rst), .I(e[314]), 
        .Q(ein[314]) );
  DFF \ereg_reg[315]  ( .D(ereg_next[315]), .CLK(clk), .RST(rst), .I(e[315]), 
        .Q(ein[315]) );
  DFF \ereg_reg[316]  ( .D(ereg_next[316]), .CLK(clk), .RST(rst), .I(e[316]), 
        .Q(ein[316]) );
  DFF \ereg_reg[317]  ( .D(ereg_next[317]), .CLK(clk), .RST(rst), .I(e[317]), 
        .Q(ein[317]) );
  DFF \ereg_reg[318]  ( .D(ereg_next[318]), .CLK(clk), .RST(rst), .I(e[318]), 
        .Q(ein[318]) );
  DFF \ereg_reg[319]  ( .D(ereg_next[319]), .CLK(clk), .RST(rst), .I(e[319]), 
        .Q(ein[319]) );
  DFF \ereg_reg[320]  ( .D(ereg_next[320]), .CLK(clk), .RST(rst), .I(e[320]), 
        .Q(ein[320]) );
  DFF \ereg_reg[321]  ( .D(ereg_next[321]), .CLK(clk), .RST(rst), .I(e[321]), 
        .Q(ein[321]) );
  DFF \ereg_reg[322]  ( .D(ereg_next[322]), .CLK(clk), .RST(rst), .I(e[322]), 
        .Q(ein[322]) );
  DFF \ereg_reg[323]  ( .D(ereg_next[323]), .CLK(clk), .RST(rst), .I(e[323]), 
        .Q(ein[323]) );
  DFF \ereg_reg[324]  ( .D(ereg_next[324]), .CLK(clk), .RST(rst), .I(e[324]), 
        .Q(ein[324]) );
  DFF \ereg_reg[325]  ( .D(ereg_next[325]), .CLK(clk), .RST(rst), .I(e[325]), 
        .Q(ein[325]) );
  DFF \ereg_reg[326]  ( .D(ereg_next[326]), .CLK(clk), .RST(rst), .I(e[326]), 
        .Q(ein[326]) );
  DFF \ereg_reg[327]  ( .D(ereg_next[327]), .CLK(clk), .RST(rst), .I(e[327]), 
        .Q(ein[327]) );
  DFF \ereg_reg[328]  ( .D(ereg_next[328]), .CLK(clk), .RST(rst), .I(e[328]), 
        .Q(ein[328]) );
  DFF \ereg_reg[329]  ( .D(ereg_next[329]), .CLK(clk), .RST(rst), .I(e[329]), 
        .Q(ein[329]) );
  DFF \ereg_reg[330]  ( .D(ereg_next[330]), .CLK(clk), .RST(rst), .I(e[330]), 
        .Q(ein[330]) );
  DFF \ereg_reg[331]  ( .D(ereg_next[331]), .CLK(clk), .RST(rst), .I(e[331]), 
        .Q(ein[331]) );
  DFF \ereg_reg[332]  ( .D(ereg_next[332]), .CLK(clk), .RST(rst), .I(e[332]), 
        .Q(ein[332]) );
  DFF \ereg_reg[333]  ( .D(ereg_next[333]), .CLK(clk), .RST(rst), .I(e[333]), 
        .Q(ein[333]) );
  DFF \ereg_reg[334]  ( .D(ereg_next[334]), .CLK(clk), .RST(rst), .I(e[334]), 
        .Q(ein[334]) );
  DFF \ereg_reg[335]  ( .D(ereg_next[335]), .CLK(clk), .RST(rst), .I(e[335]), 
        .Q(ein[335]) );
  DFF \ereg_reg[336]  ( .D(ereg_next[336]), .CLK(clk), .RST(rst), .I(e[336]), 
        .Q(ein[336]) );
  DFF \ereg_reg[337]  ( .D(ereg_next[337]), .CLK(clk), .RST(rst), .I(e[337]), 
        .Q(ein[337]) );
  DFF \ereg_reg[338]  ( .D(ereg_next[338]), .CLK(clk), .RST(rst), .I(e[338]), 
        .Q(ein[338]) );
  DFF \ereg_reg[339]  ( .D(ereg_next[339]), .CLK(clk), .RST(rst), .I(e[339]), 
        .Q(ein[339]) );
  DFF \ereg_reg[340]  ( .D(ereg_next[340]), .CLK(clk), .RST(rst), .I(e[340]), 
        .Q(ein[340]) );
  DFF \ereg_reg[341]  ( .D(ereg_next[341]), .CLK(clk), .RST(rst), .I(e[341]), 
        .Q(ein[341]) );
  DFF \ereg_reg[342]  ( .D(ereg_next[342]), .CLK(clk), .RST(rst), .I(e[342]), 
        .Q(ein[342]) );
  DFF \ereg_reg[343]  ( .D(ereg_next[343]), .CLK(clk), .RST(rst), .I(e[343]), 
        .Q(ein[343]) );
  DFF \ereg_reg[344]  ( .D(ereg_next[344]), .CLK(clk), .RST(rst), .I(e[344]), 
        .Q(ein[344]) );
  DFF \ereg_reg[345]  ( .D(ereg_next[345]), .CLK(clk), .RST(rst), .I(e[345]), 
        .Q(ein[345]) );
  DFF \ereg_reg[346]  ( .D(ereg_next[346]), .CLK(clk), .RST(rst), .I(e[346]), 
        .Q(ein[346]) );
  DFF \ereg_reg[347]  ( .D(ereg_next[347]), .CLK(clk), .RST(rst), .I(e[347]), 
        .Q(ein[347]) );
  DFF \ereg_reg[348]  ( .D(ereg_next[348]), .CLK(clk), .RST(rst), .I(e[348]), 
        .Q(ein[348]) );
  DFF \ereg_reg[349]  ( .D(ereg_next[349]), .CLK(clk), .RST(rst), .I(e[349]), 
        .Q(ein[349]) );
  DFF \ereg_reg[350]  ( .D(ereg_next[350]), .CLK(clk), .RST(rst), .I(e[350]), 
        .Q(ein[350]) );
  DFF \ereg_reg[351]  ( .D(ereg_next[351]), .CLK(clk), .RST(rst), .I(e[351]), 
        .Q(ein[351]) );
  DFF \ereg_reg[352]  ( .D(ereg_next[352]), .CLK(clk), .RST(rst), .I(e[352]), 
        .Q(ein[352]) );
  DFF \ereg_reg[353]  ( .D(ereg_next[353]), .CLK(clk), .RST(rst), .I(e[353]), 
        .Q(ein[353]) );
  DFF \ereg_reg[354]  ( .D(ereg_next[354]), .CLK(clk), .RST(rst), .I(e[354]), 
        .Q(ein[354]) );
  DFF \ereg_reg[355]  ( .D(ereg_next[355]), .CLK(clk), .RST(rst), .I(e[355]), 
        .Q(ein[355]) );
  DFF \ereg_reg[356]  ( .D(ereg_next[356]), .CLK(clk), .RST(rst), .I(e[356]), 
        .Q(ein[356]) );
  DFF \ereg_reg[357]  ( .D(ereg_next[357]), .CLK(clk), .RST(rst), .I(e[357]), 
        .Q(ein[357]) );
  DFF \ereg_reg[358]  ( .D(ereg_next[358]), .CLK(clk), .RST(rst), .I(e[358]), 
        .Q(ein[358]) );
  DFF \ereg_reg[359]  ( .D(ereg_next[359]), .CLK(clk), .RST(rst), .I(e[359]), 
        .Q(ein[359]) );
  DFF \ereg_reg[360]  ( .D(ereg_next[360]), .CLK(clk), .RST(rst), .I(e[360]), 
        .Q(ein[360]) );
  DFF \ereg_reg[361]  ( .D(ereg_next[361]), .CLK(clk), .RST(rst), .I(e[361]), 
        .Q(ein[361]) );
  DFF \ereg_reg[362]  ( .D(ereg_next[362]), .CLK(clk), .RST(rst), .I(e[362]), 
        .Q(ein[362]) );
  DFF \ereg_reg[363]  ( .D(ereg_next[363]), .CLK(clk), .RST(rst), .I(e[363]), 
        .Q(ein[363]) );
  DFF \ereg_reg[364]  ( .D(ereg_next[364]), .CLK(clk), .RST(rst), .I(e[364]), 
        .Q(ein[364]) );
  DFF \ereg_reg[365]  ( .D(ereg_next[365]), .CLK(clk), .RST(rst), .I(e[365]), 
        .Q(ein[365]) );
  DFF \ereg_reg[366]  ( .D(ereg_next[366]), .CLK(clk), .RST(rst), .I(e[366]), 
        .Q(ein[366]) );
  DFF \ereg_reg[367]  ( .D(ereg_next[367]), .CLK(clk), .RST(rst), .I(e[367]), 
        .Q(ein[367]) );
  DFF \ereg_reg[368]  ( .D(ereg_next[368]), .CLK(clk), .RST(rst), .I(e[368]), 
        .Q(ein[368]) );
  DFF \ereg_reg[369]  ( .D(ereg_next[369]), .CLK(clk), .RST(rst), .I(e[369]), 
        .Q(ein[369]) );
  DFF \ereg_reg[370]  ( .D(ereg_next[370]), .CLK(clk), .RST(rst), .I(e[370]), 
        .Q(ein[370]) );
  DFF \ereg_reg[371]  ( .D(ereg_next[371]), .CLK(clk), .RST(rst), .I(e[371]), 
        .Q(ein[371]) );
  DFF \ereg_reg[372]  ( .D(ereg_next[372]), .CLK(clk), .RST(rst), .I(e[372]), 
        .Q(ein[372]) );
  DFF \ereg_reg[373]  ( .D(ereg_next[373]), .CLK(clk), .RST(rst), .I(e[373]), 
        .Q(ein[373]) );
  DFF \ereg_reg[374]  ( .D(ereg_next[374]), .CLK(clk), .RST(rst), .I(e[374]), 
        .Q(ein[374]) );
  DFF \ereg_reg[375]  ( .D(ereg_next[375]), .CLK(clk), .RST(rst), .I(e[375]), 
        .Q(ein[375]) );
  DFF \ereg_reg[376]  ( .D(ereg_next[376]), .CLK(clk), .RST(rst), .I(e[376]), 
        .Q(ein[376]) );
  DFF \ereg_reg[377]  ( .D(ereg_next[377]), .CLK(clk), .RST(rst), .I(e[377]), 
        .Q(ein[377]) );
  DFF \ereg_reg[378]  ( .D(ereg_next[378]), .CLK(clk), .RST(rst), .I(e[378]), 
        .Q(ein[378]) );
  DFF \ereg_reg[379]  ( .D(ereg_next[379]), .CLK(clk), .RST(rst), .I(e[379]), 
        .Q(ein[379]) );
  DFF \ereg_reg[380]  ( .D(ereg_next[380]), .CLK(clk), .RST(rst), .I(e[380]), 
        .Q(ein[380]) );
  DFF \ereg_reg[381]  ( .D(ereg_next[381]), .CLK(clk), .RST(rst), .I(e[381]), 
        .Q(ein[381]) );
  DFF \ereg_reg[382]  ( .D(ereg_next[382]), .CLK(clk), .RST(rst), .I(e[382]), 
        .Q(ein[382]) );
  DFF \ereg_reg[383]  ( .D(ereg_next[383]), .CLK(clk), .RST(rst), .I(e[383]), 
        .Q(ein[383]) );
  DFF \ereg_reg[384]  ( .D(ereg_next[384]), .CLK(clk), .RST(rst), .I(e[384]), 
        .Q(ein[384]) );
  DFF \ereg_reg[385]  ( .D(ereg_next[385]), .CLK(clk), .RST(rst), .I(e[385]), 
        .Q(ein[385]) );
  DFF \ereg_reg[386]  ( .D(ereg_next[386]), .CLK(clk), .RST(rst), .I(e[386]), 
        .Q(ein[386]) );
  DFF \ereg_reg[387]  ( .D(ereg_next[387]), .CLK(clk), .RST(rst), .I(e[387]), 
        .Q(ein[387]) );
  DFF \ereg_reg[388]  ( .D(ereg_next[388]), .CLK(clk), .RST(rst), .I(e[388]), 
        .Q(ein[388]) );
  DFF \ereg_reg[389]  ( .D(ereg_next[389]), .CLK(clk), .RST(rst), .I(e[389]), 
        .Q(ein[389]) );
  DFF \ereg_reg[390]  ( .D(ereg_next[390]), .CLK(clk), .RST(rst), .I(e[390]), 
        .Q(ein[390]) );
  DFF \ereg_reg[391]  ( .D(ereg_next[391]), .CLK(clk), .RST(rst), .I(e[391]), 
        .Q(ein[391]) );
  DFF \ereg_reg[392]  ( .D(ereg_next[392]), .CLK(clk), .RST(rst), .I(e[392]), 
        .Q(ein[392]) );
  DFF \ereg_reg[393]  ( .D(ereg_next[393]), .CLK(clk), .RST(rst), .I(e[393]), 
        .Q(ein[393]) );
  DFF \ereg_reg[394]  ( .D(ereg_next[394]), .CLK(clk), .RST(rst), .I(e[394]), 
        .Q(ein[394]) );
  DFF \ereg_reg[395]  ( .D(ereg_next[395]), .CLK(clk), .RST(rst), .I(e[395]), 
        .Q(ein[395]) );
  DFF \ereg_reg[396]  ( .D(ereg_next[396]), .CLK(clk), .RST(rst), .I(e[396]), 
        .Q(ein[396]) );
  DFF \ereg_reg[397]  ( .D(ereg_next[397]), .CLK(clk), .RST(rst), .I(e[397]), 
        .Q(ein[397]) );
  DFF \ereg_reg[398]  ( .D(ereg_next[398]), .CLK(clk), .RST(rst), .I(e[398]), 
        .Q(ein[398]) );
  DFF \ereg_reg[399]  ( .D(ereg_next[399]), .CLK(clk), .RST(rst), .I(e[399]), 
        .Q(ein[399]) );
  DFF \ereg_reg[400]  ( .D(ereg_next[400]), .CLK(clk), .RST(rst), .I(e[400]), 
        .Q(ein[400]) );
  DFF \ereg_reg[401]  ( .D(ereg_next[401]), .CLK(clk), .RST(rst), .I(e[401]), 
        .Q(ein[401]) );
  DFF \ereg_reg[402]  ( .D(ereg_next[402]), .CLK(clk), .RST(rst), .I(e[402]), 
        .Q(ein[402]) );
  DFF \ereg_reg[403]  ( .D(ereg_next[403]), .CLK(clk), .RST(rst), .I(e[403]), 
        .Q(ein[403]) );
  DFF \ereg_reg[404]  ( .D(ereg_next[404]), .CLK(clk), .RST(rst), .I(e[404]), 
        .Q(ein[404]) );
  DFF \ereg_reg[405]  ( .D(ereg_next[405]), .CLK(clk), .RST(rst), .I(e[405]), 
        .Q(ein[405]) );
  DFF \ereg_reg[406]  ( .D(ereg_next[406]), .CLK(clk), .RST(rst), .I(e[406]), 
        .Q(ein[406]) );
  DFF \ereg_reg[407]  ( .D(ereg_next[407]), .CLK(clk), .RST(rst), .I(e[407]), 
        .Q(ein[407]) );
  DFF \ereg_reg[408]  ( .D(ereg_next[408]), .CLK(clk), .RST(rst), .I(e[408]), 
        .Q(ein[408]) );
  DFF \ereg_reg[409]  ( .D(ereg_next[409]), .CLK(clk), .RST(rst), .I(e[409]), 
        .Q(ein[409]) );
  DFF \ereg_reg[410]  ( .D(ereg_next[410]), .CLK(clk), .RST(rst), .I(e[410]), 
        .Q(ein[410]) );
  DFF \ereg_reg[411]  ( .D(ereg_next[411]), .CLK(clk), .RST(rst), .I(e[411]), 
        .Q(ein[411]) );
  DFF \ereg_reg[412]  ( .D(ereg_next[412]), .CLK(clk), .RST(rst), .I(e[412]), 
        .Q(ein[412]) );
  DFF \ereg_reg[413]  ( .D(ereg_next[413]), .CLK(clk), .RST(rst), .I(e[413]), 
        .Q(ein[413]) );
  DFF \ereg_reg[414]  ( .D(ereg_next[414]), .CLK(clk), .RST(rst), .I(e[414]), 
        .Q(ein[414]) );
  DFF \ereg_reg[415]  ( .D(ereg_next[415]), .CLK(clk), .RST(rst), .I(e[415]), 
        .Q(ein[415]) );
  DFF \ereg_reg[416]  ( .D(ereg_next[416]), .CLK(clk), .RST(rst), .I(e[416]), 
        .Q(ein[416]) );
  DFF \ereg_reg[417]  ( .D(ereg_next[417]), .CLK(clk), .RST(rst), .I(e[417]), 
        .Q(ein[417]) );
  DFF \ereg_reg[418]  ( .D(ereg_next[418]), .CLK(clk), .RST(rst), .I(e[418]), 
        .Q(ein[418]) );
  DFF \ereg_reg[419]  ( .D(ereg_next[419]), .CLK(clk), .RST(rst), .I(e[419]), 
        .Q(ein[419]) );
  DFF \ereg_reg[420]  ( .D(ereg_next[420]), .CLK(clk), .RST(rst), .I(e[420]), 
        .Q(ein[420]) );
  DFF \ereg_reg[421]  ( .D(ereg_next[421]), .CLK(clk), .RST(rst), .I(e[421]), 
        .Q(ein[421]) );
  DFF \ereg_reg[422]  ( .D(ereg_next[422]), .CLK(clk), .RST(rst), .I(e[422]), 
        .Q(ein[422]) );
  DFF \ereg_reg[423]  ( .D(ereg_next[423]), .CLK(clk), .RST(rst), .I(e[423]), 
        .Q(ein[423]) );
  DFF \ereg_reg[424]  ( .D(ereg_next[424]), .CLK(clk), .RST(rst), .I(e[424]), 
        .Q(ein[424]) );
  DFF \ereg_reg[425]  ( .D(ereg_next[425]), .CLK(clk), .RST(rst), .I(e[425]), 
        .Q(ein[425]) );
  DFF \ereg_reg[426]  ( .D(ereg_next[426]), .CLK(clk), .RST(rst), .I(e[426]), 
        .Q(ein[426]) );
  DFF \ereg_reg[427]  ( .D(ereg_next[427]), .CLK(clk), .RST(rst), .I(e[427]), 
        .Q(ein[427]) );
  DFF \ereg_reg[428]  ( .D(ereg_next[428]), .CLK(clk), .RST(rst), .I(e[428]), 
        .Q(ein[428]) );
  DFF \ereg_reg[429]  ( .D(ereg_next[429]), .CLK(clk), .RST(rst), .I(e[429]), 
        .Q(ein[429]) );
  DFF \ereg_reg[430]  ( .D(ereg_next[430]), .CLK(clk), .RST(rst), .I(e[430]), 
        .Q(ein[430]) );
  DFF \ereg_reg[431]  ( .D(ereg_next[431]), .CLK(clk), .RST(rst), .I(e[431]), 
        .Q(ein[431]) );
  DFF \ereg_reg[432]  ( .D(ereg_next[432]), .CLK(clk), .RST(rst), .I(e[432]), 
        .Q(ein[432]) );
  DFF \ereg_reg[433]  ( .D(ereg_next[433]), .CLK(clk), .RST(rst), .I(e[433]), 
        .Q(ein[433]) );
  DFF \ereg_reg[434]  ( .D(ereg_next[434]), .CLK(clk), .RST(rst), .I(e[434]), 
        .Q(ein[434]) );
  DFF \ereg_reg[435]  ( .D(ereg_next[435]), .CLK(clk), .RST(rst), .I(e[435]), 
        .Q(ein[435]) );
  DFF \ereg_reg[436]  ( .D(ereg_next[436]), .CLK(clk), .RST(rst), .I(e[436]), 
        .Q(ein[436]) );
  DFF \ereg_reg[437]  ( .D(ereg_next[437]), .CLK(clk), .RST(rst), .I(e[437]), 
        .Q(ein[437]) );
  DFF \ereg_reg[438]  ( .D(ereg_next[438]), .CLK(clk), .RST(rst), .I(e[438]), 
        .Q(ein[438]) );
  DFF \ereg_reg[439]  ( .D(ereg_next[439]), .CLK(clk), .RST(rst), .I(e[439]), 
        .Q(ein[439]) );
  DFF \ereg_reg[440]  ( .D(ereg_next[440]), .CLK(clk), .RST(rst), .I(e[440]), 
        .Q(ein[440]) );
  DFF \ereg_reg[441]  ( .D(ereg_next[441]), .CLK(clk), .RST(rst), .I(e[441]), 
        .Q(ein[441]) );
  DFF \ereg_reg[442]  ( .D(ereg_next[442]), .CLK(clk), .RST(rst), .I(e[442]), 
        .Q(ein[442]) );
  DFF \ereg_reg[443]  ( .D(ereg_next[443]), .CLK(clk), .RST(rst), .I(e[443]), 
        .Q(ein[443]) );
  DFF \ereg_reg[444]  ( .D(ereg_next[444]), .CLK(clk), .RST(rst), .I(e[444]), 
        .Q(ein[444]) );
  DFF \ereg_reg[445]  ( .D(ereg_next[445]), .CLK(clk), .RST(rst), .I(e[445]), 
        .Q(ein[445]) );
  DFF \ereg_reg[446]  ( .D(ereg_next[446]), .CLK(clk), .RST(rst), .I(e[446]), 
        .Q(ein[446]) );
  DFF \ereg_reg[447]  ( .D(ereg_next[447]), .CLK(clk), .RST(rst), .I(e[447]), 
        .Q(ein[447]) );
  DFF \ereg_reg[448]  ( .D(ereg_next[448]), .CLK(clk), .RST(rst), .I(e[448]), 
        .Q(ein[448]) );
  DFF \ereg_reg[449]  ( .D(ereg_next[449]), .CLK(clk), .RST(rst), .I(e[449]), 
        .Q(ein[449]) );
  DFF \ereg_reg[450]  ( .D(ereg_next[450]), .CLK(clk), .RST(rst), .I(e[450]), 
        .Q(ein[450]) );
  DFF \ereg_reg[451]  ( .D(ereg_next[451]), .CLK(clk), .RST(rst), .I(e[451]), 
        .Q(ein[451]) );
  DFF \ereg_reg[452]  ( .D(ereg_next[452]), .CLK(clk), .RST(rst), .I(e[452]), 
        .Q(ein[452]) );
  DFF \ereg_reg[453]  ( .D(ereg_next[453]), .CLK(clk), .RST(rst), .I(e[453]), 
        .Q(ein[453]) );
  DFF \ereg_reg[454]  ( .D(ereg_next[454]), .CLK(clk), .RST(rst), .I(e[454]), 
        .Q(ein[454]) );
  DFF \ereg_reg[455]  ( .D(ereg_next[455]), .CLK(clk), .RST(rst), .I(e[455]), 
        .Q(ein[455]) );
  DFF \ereg_reg[456]  ( .D(ereg_next[456]), .CLK(clk), .RST(rst), .I(e[456]), 
        .Q(ein[456]) );
  DFF \ereg_reg[457]  ( .D(ereg_next[457]), .CLK(clk), .RST(rst), .I(e[457]), 
        .Q(ein[457]) );
  DFF \ereg_reg[458]  ( .D(ereg_next[458]), .CLK(clk), .RST(rst), .I(e[458]), 
        .Q(ein[458]) );
  DFF \ereg_reg[459]  ( .D(ereg_next[459]), .CLK(clk), .RST(rst), .I(e[459]), 
        .Q(ein[459]) );
  DFF \ereg_reg[460]  ( .D(ereg_next[460]), .CLK(clk), .RST(rst), .I(e[460]), 
        .Q(ein[460]) );
  DFF \ereg_reg[461]  ( .D(ereg_next[461]), .CLK(clk), .RST(rst), .I(e[461]), 
        .Q(ein[461]) );
  DFF \ereg_reg[462]  ( .D(ereg_next[462]), .CLK(clk), .RST(rst), .I(e[462]), 
        .Q(ein[462]) );
  DFF \ereg_reg[463]  ( .D(ereg_next[463]), .CLK(clk), .RST(rst), .I(e[463]), 
        .Q(ein[463]) );
  DFF \ereg_reg[464]  ( .D(ereg_next[464]), .CLK(clk), .RST(rst), .I(e[464]), 
        .Q(ein[464]) );
  DFF \ereg_reg[465]  ( .D(ereg_next[465]), .CLK(clk), .RST(rst), .I(e[465]), 
        .Q(ein[465]) );
  DFF \ereg_reg[466]  ( .D(ereg_next[466]), .CLK(clk), .RST(rst), .I(e[466]), 
        .Q(ein[466]) );
  DFF \ereg_reg[467]  ( .D(ereg_next[467]), .CLK(clk), .RST(rst), .I(e[467]), 
        .Q(ein[467]) );
  DFF \ereg_reg[468]  ( .D(ereg_next[468]), .CLK(clk), .RST(rst), .I(e[468]), 
        .Q(ein[468]) );
  DFF \ereg_reg[469]  ( .D(ereg_next[469]), .CLK(clk), .RST(rst), .I(e[469]), 
        .Q(ein[469]) );
  DFF \ereg_reg[470]  ( .D(ereg_next[470]), .CLK(clk), .RST(rst), .I(e[470]), 
        .Q(ein[470]) );
  DFF \ereg_reg[471]  ( .D(ereg_next[471]), .CLK(clk), .RST(rst), .I(e[471]), 
        .Q(ein[471]) );
  DFF \ereg_reg[472]  ( .D(ereg_next[472]), .CLK(clk), .RST(rst), .I(e[472]), 
        .Q(ein[472]) );
  DFF \ereg_reg[473]  ( .D(ereg_next[473]), .CLK(clk), .RST(rst), .I(e[473]), 
        .Q(ein[473]) );
  DFF \ereg_reg[474]  ( .D(ereg_next[474]), .CLK(clk), .RST(rst), .I(e[474]), 
        .Q(ein[474]) );
  DFF \ereg_reg[475]  ( .D(ereg_next[475]), .CLK(clk), .RST(rst), .I(e[475]), 
        .Q(ein[475]) );
  DFF \ereg_reg[476]  ( .D(ereg_next[476]), .CLK(clk), .RST(rst), .I(e[476]), 
        .Q(ein[476]) );
  DFF \ereg_reg[477]  ( .D(ereg_next[477]), .CLK(clk), .RST(rst), .I(e[477]), 
        .Q(ein[477]) );
  DFF \ereg_reg[478]  ( .D(ereg_next[478]), .CLK(clk), .RST(rst), .I(e[478]), 
        .Q(ein[478]) );
  DFF \ereg_reg[479]  ( .D(ereg_next[479]), .CLK(clk), .RST(rst), .I(e[479]), 
        .Q(ein[479]) );
  DFF \ereg_reg[480]  ( .D(ereg_next[480]), .CLK(clk), .RST(rst), .I(e[480]), 
        .Q(ein[480]) );
  DFF \ereg_reg[481]  ( .D(ereg_next[481]), .CLK(clk), .RST(rst), .I(e[481]), 
        .Q(ein[481]) );
  DFF \ereg_reg[482]  ( .D(ereg_next[482]), .CLK(clk), .RST(rst), .I(e[482]), 
        .Q(ein[482]) );
  DFF \ereg_reg[483]  ( .D(ereg_next[483]), .CLK(clk), .RST(rst), .I(e[483]), 
        .Q(ein[483]) );
  DFF \ereg_reg[484]  ( .D(ereg_next[484]), .CLK(clk), .RST(rst), .I(e[484]), 
        .Q(ein[484]) );
  DFF \ereg_reg[485]  ( .D(ereg_next[485]), .CLK(clk), .RST(rst), .I(e[485]), 
        .Q(ein[485]) );
  DFF \ereg_reg[486]  ( .D(ereg_next[486]), .CLK(clk), .RST(rst), .I(e[486]), 
        .Q(ein[486]) );
  DFF \ereg_reg[487]  ( .D(ereg_next[487]), .CLK(clk), .RST(rst), .I(e[487]), 
        .Q(ein[487]) );
  DFF \ereg_reg[488]  ( .D(ereg_next[488]), .CLK(clk), .RST(rst), .I(e[488]), 
        .Q(ein[488]) );
  DFF \ereg_reg[489]  ( .D(ereg_next[489]), .CLK(clk), .RST(rst), .I(e[489]), 
        .Q(ein[489]) );
  DFF \ereg_reg[490]  ( .D(ereg_next[490]), .CLK(clk), .RST(rst), .I(e[490]), 
        .Q(ein[490]) );
  DFF \ereg_reg[491]  ( .D(ereg_next[491]), .CLK(clk), .RST(rst), .I(e[491]), 
        .Q(ein[491]) );
  DFF \ereg_reg[492]  ( .D(ereg_next[492]), .CLK(clk), .RST(rst), .I(e[492]), 
        .Q(ein[492]) );
  DFF \ereg_reg[493]  ( .D(ereg_next[493]), .CLK(clk), .RST(rst), .I(e[493]), 
        .Q(ein[493]) );
  DFF \ereg_reg[494]  ( .D(ereg_next[494]), .CLK(clk), .RST(rst), .I(e[494]), 
        .Q(ein[494]) );
  DFF \ereg_reg[495]  ( .D(ereg_next[495]), .CLK(clk), .RST(rst), .I(e[495]), 
        .Q(ein[495]) );
  DFF \ereg_reg[496]  ( .D(ereg_next[496]), .CLK(clk), .RST(rst), .I(e[496]), 
        .Q(ein[496]) );
  DFF \ereg_reg[497]  ( .D(ereg_next[497]), .CLK(clk), .RST(rst), .I(e[497]), 
        .Q(ein[497]) );
  DFF \ereg_reg[498]  ( .D(ereg_next[498]), .CLK(clk), .RST(rst), .I(e[498]), 
        .Q(ein[498]) );
  DFF \ereg_reg[499]  ( .D(ereg_next[499]), .CLK(clk), .RST(rst), .I(e[499]), 
        .Q(ein[499]) );
  DFF \ereg_reg[500]  ( .D(ereg_next[500]), .CLK(clk), .RST(rst), .I(e[500]), 
        .Q(ein[500]) );
  DFF \ereg_reg[501]  ( .D(ereg_next[501]), .CLK(clk), .RST(rst), .I(e[501]), 
        .Q(ein[501]) );
  DFF \ereg_reg[502]  ( .D(ereg_next[502]), .CLK(clk), .RST(rst), .I(e[502]), 
        .Q(ein[502]) );
  DFF \ereg_reg[503]  ( .D(ereg_next[503]), .CLK(clk), .RST(rst), .I(e[503]), 
        .Q(ein[503]) );
  DFF \ereg_reg[504]  ( .D(ereg_next[504]), .CLK(clk), .RST(rst), .I(e[504]), 
        .Q(ein[504]) );
  DFF \ereg_reg[505]  ( .D(ereg_next[505]), .CLK(clk), .RST(rst), .I(e[505]), 
        .Q(ein[505]) );
  DFF \ereg_reg[506]  ( .D(ereg_next[506]), .CLK(clk), .RST(rst), .I(e[506]), 
        .Q(ein[506]) );
  DFF \ereg_reg[507]  ( .D(ereg_next[507]), .CLK(clk), .RST(rst), .I(e[507]), 
        .Q(ein[507]) );
  DFF \ereg_reg[508]  ( .D(ereg_next[508]), .CLK(clk), .RST(rst), .I(e[508]), 
        .Q(ein[508]) );
  DFF \ereg_reg[509]  ( .D(ereg_next[509]), .CLK(clk), .RST(rst), .I(e[509]), 
        .Q(ein[509]) );
  DFF \ereg_reg[510]  ( .D(ereg_next[510]), .CLK(clk), .RST(rst), .I(e[510]), 
        .Q(ein[510]) );
  DFF \ereg_reg[511]  ( .D(ereg_next[511]), .CLK(clk), .RST(rst), .I(e[511]), 
        .Q(ein[511]) );
  DFF first_one_reg ( .D(n6), .CLK(clk), .RST(rst), .I(1'b0), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(creg_next[0]), .CLK(clk), .RST(rst), .I(m[0]), .Q(
        c[0]) );
  DFF \creg_reg[1]  ( .D(creg_next[1]), .CLK(clk), .RST(rst), .I(m[1]), .Q(
        c[1]) );
  DFF \creg_reg[2]  ( .D(creg_next[2]), .CLK(clk), .RST(rst), .I(m[2]), .Q(
        c[2]) );
  DFF \creg_reg[3]  ( .D(creg_next[3]), .CLK(clk), .RST(rst), .I(m[3]), .Q(
        c[3]) );
  DFF \creg_reg[4]  ( .D(creg_next[4]), .CLK(clk), .RST(rst), .I(m[4]), .Q(
        c[4]) );
  DFF \creg_reg[5]  ( .D(creg_next[5]), .CLK(clk), .RST(rst), .I(m[5]), .Q(
        c[5]) );
  DFF \creg_reg[6]  ( .D(creg_next[6]), .CLK(clk), .RST(rst), .I(m[6]), .Q(
        c[6]) );
  DFF \creg_reg[7]  ( .D(creg_next[7]), .CLK(clk), .RST(rst), .I(m[7]), .Q(
        c[7]) );
  DFF \creg_reg[8]  ( .D(creg_next[8]), .CLK(clk), .RST(rst), .I(m[8]), .Q(
        c[8]) );
  DFF \creg_reg[9]  ( .D(creg_next[9]), .CLK(clk), .RST(rst), .I(m[9]), .Q(
        c[9]) );
  DFF \creg_reg[10]  ( .D(creg_next[10]), .CLK(clk), .RST(rst), .I(m[10]), .Q(
        c[10]) );
  DFF \creg_reg[11]  ( .D(creg_next[11]), .CLK(clk), .RST(rst), .I(m[11]), .Q(
        c[11]) );
  DFF \creg_reg[12]  ( .D(creg_next[12]), .CLK(clk), .RST(rst), .I(m[12]), .Q(
        c[12]) );
  DFF \creg_reg[13]  ( .D(creg_next[13]), .CLK(clk), .RST(rst), .I(m[13]), .Q(
        c[13]) );
  DFF \creg_reg[14]  ( .D(creg_next[14]), .CLK(clk), .RST(rst), .I(m[14]), .Q(
        c[14]) );
  DFF \creg_reg[15]  ( .D(creg_next[15]), .CLK(clk), .RST(rst), .I(m[15]), .Q(
        c[15]) );
  DFF \creg_reg[16]  ( .D(creg_next[16]), .CLK(clk), .RST(rst), .I(m[16]), .Q(
        c[16]) );
  DFF \creg_reg[17]  ( .D(creg_next[17]), .CLK(clk), .RST(rst), .I(m[17]), .Q(
        c[17]) );
  DFF \creg_reg[18]  ( .D(creg_next[18]), .CLK(clk), .RST(rst), .I(m[18]), .Q(
        c[18]) );
  DFF \creg_reg[19]  ( .D(creg_next[19]), .CLK(clk), .RST(rst), .I(m[19]), .Q(
        c[19]) );
  DFF \creg_reg[20]  ( .D(creg_next[20]), .CLK(clk), .RST(rst), .I(m[20]), .Q(
        c[20]) );
  DFF \creg_reg[21]  ( .D(creg_next[21]), .CLK(clk), .RST(rst), .I(m[21]), .Q(
        c[21]) );
  DFF \creg_reg[22]  ( .D(creg_next[22]), .CLK(clk), .RST(rst), .I(m[22]), .Q(
        c[22]) );
  DFF \creg_reg[23]  ( .D(creg_next[23]), .CLK(clk), .RST(rst), .I(m[23]), .Q(
        c[23]) );
  DFF \creg_reg[24]  ( .D(creg_next[24]), .CLK(clk), .RST(rst), .I(m[24]), .Q(
        c[24]) );
  DFF \creg_reg[25]  ( .D(creg_next[25]), .CLK(clk), .RST(rst), .I(m[25]), .Q(
        c[25]) );
  DFF \creg_reg[26]  ( .D(creg_next[26]), .CLK(clk), .RST(rst), .I(m[26]), .Q(
        c[26]) );
  DFF \creg_reg[27]  ( .D(creg_next[27]), .CLK(clk), .RST(rst), .I(m[27]), .Q(
        c[27]) );
  DFF \creg_reg[28]  ( .D(creg_next[28]), .CLK(clk), .RST(rst), .I(m[28]), .Q(
        c[28]) );
  DFF \creg_reg[29]  ( .D(creg_next[29]), .CLK(clk), .RST(rst), .I(m[29]), .Q(
        c[29]) );
  DFF \creg_reg[30]  ( .D(creg_next[30]), .CLK(clk), .RST(rst), .I(m[30]), .Q(
        c[30]) );
  DFF \creg_reg[31]  ( .D(creg_next[31]), .CLK(clk), .RST(rst), .I(m[31]), .Q(
        c[31]) );
  DFF \creg_reg[32]  ( .D(creg_next[32]), .CLK(clk), .RST(rst), .I(m[32]), .Q(
        c[32]) );
  DFF \creg_reg[33]  ( .D(creg_next[33]), .CLK(clk), .RST(rst), .I(m[33]), .Q(
        c[33]) );
  DFF \creg_reg[34]  ( .D(creg_next[34]), .CLK(clk), .RST(rst), .I(m[34]), .Q(
        c[34]) );
  DFF \creg_reg[35]  ( .D(creg_next[35]), .CLK(clk), .RST(rst), .I(m[35]), .Q(
        c[35]) );
  DFF \creg_reg[36]  ( .D(creg_next[36]), .CLK(clk), .RST(rst), .I(m[36]), .Q(
        c[36]) );
  DFF \creg_reg[37]  ( .D(creg_next[37]), .CLK(clk), .RST(rst), .I(m[37]), .Q(
        c[37]) );
  DFF \creg_reg[38]  ( .D(creg_next[38]), .CLK(clk), .RST(rst), .I(m[38]), .Q(
        c[38]) );
  DFF \creg_reg[39]  ( .D(creg_next[39]), .CLK(clk), .RST(rst), .I(m[39]), .Q(
        c[39]) );
  DFF \creg_reg[40]  ( .D(creg_next[40]), .CLK(clk), .RST(rst), .I(m[40]), .Q(
        c[40]) );
  DFF \creg_reg[41]  ( .D(creg_next[41]), .CLK(clk), .RST(rst), .I(m[41]), .Q(
        c[41]) );
  DFF \creg_reg[42]  ( .D(creg_next[42]), .CLK(clk), .RST(rst), .I(m[42]), .Q(
        c[42]) );
  DFF \creg_reg[43]  ( .D(creg_next[43]), .CLK(clk), .RST(rst), .I(m[43]), .Q(
        c[43]) );
  DFF \creg_reg[44]  ( .D(creg_next[44]), .CLK(clk), .RST(rst), .I(m[44]), .Q(
        c[44]) );
  DFF \creg_reg[45]  ( .D(creg_next[45]), .CLK(clk), .RST(rst), .I(m[45]), .Q(
        c[45]) );
  DFF \creg_reg[46]  ( .D(creg_next[46]), .CLK(clk), .RST(rst), .I(m[46]), .Q(
        c[46]) );
  DFF \creg_reg[47]  ( .D(creg_next[47]), .CLK(clk), .RST(rst), .I(m[47]), .Q(
        c[47]) );
  DFF \creg_reg[48]  ( .D(creg_next[48]), .CLK(clk), .RST(rst), .I(m[48]), .Q(
        c[48]) );
  DFF \creg_reg[49]  ( .D(creg_next[49]), .CLK(clk), .RST(rst), .I(m[49]), .Q(
        c[49]) );
  DFF \creg_reg[50]  ( .D(creg_next[50]), .CLK(clk), .RST(rst), .I(m[50]), .Q(
        c[50]) );
  DFF \creg_reg[51]  ( .D(creg_next[51]), .CLK(clk), .RST(rst), .I(m[51]), .Q(
        c[51]) );
  DFF \creg_reg[52]  ( .D(creg_next[52]), .CLK(clk), .RST(rst), .I(m[52]), .Q(
        c[52]) );
  DFF \creg_reg[53]  ( .D(creg_next[53]), .CLK(clk), .RST(rst), .I(m[53]), .Q(
        c[53]) );
  DFF \creg_reg[54]  ( .D(creg_next[54]), .CLK(clk), .RST(rst), .I(m[54]), .Q(
        c[54]) );
  DFF \creg_reg[55]  ( .D(creg_next[55]), .CLK(clk), .RST(rst), .I(m[55]), .Q(
        c[55]) );
  DFF \creg_reg[56]  ( .D(creg_next[56]), .CLK(clk), .RST(rst), .I(m[56]), .Q(
        c[56]) );
  DFF \creg_reg[57]  ( .D(creg_next[57]), .CLK(clk), .RST(rst), .I(m[57]), .Q(
        c[57]) );
  DFF \creg_reg[58]  ( .D(creg_next[58]), .CLK(clk), .RST(rst), .I(m[58]), .Q(
        c[58]) );
  DFF \creg_reg[59]  ( .D(creg_next[59]), .CLK(clk), .RST(rst), .I(m[59]), .Q(
        c[59]) );
  DFF \creg_reg[60]  ( .D(creg_next[60]), .CLK(clk), .RST(rst), .I(m[60]), .Q(
        c[60]) );
  DFF \creg_reg[61]  ( .D(creg_next[61]), .CLK(clk), .RST(rst), .I(m[61]), .Q(
        c[61]) );
  DFF \creg_reg[62]  ( .D(creg_next[62]), .CLK(clk), .RST(rst), .I(m[62]), .Q(
        c[62]) );
  DFF \creg_reg[63]  ( .D(creg_next[63]), .CLK(clk), .RST(rst), .I(m[63]), .Q(
        c[63]) );
  DFF \creg_reg[64]  ( .D(creg_next[64]), .CLK(clk), .RST(rst), .I(m[64]), .Q(
        c[64]) );
  DFF \creg_reg[65]  ( .D(creg_next[65]), .CLK(clk), .RST(rst), .I(m[65]), .Q(
        c[65]) );
  DFF \creg_reg[66]  ( .D(creg_next[66]), .CLK(clk), .RST(rst), .I(m[66]), .Q(
        c[66]) );
  DFF \creg_reg[67]  ( .D(creg_next[67]), .CLK(clk), .RST(rst), .I(m[67]), .Q(
        c[67]) );
  DFF \creg_reg[68]  ( .D(creg_next[68]), .CLK(clk), .RST(rst), .I(m[68]), .Q(
        c[68]) );
  DFF \creg_reg[69]  ( .D(creg_next[69]), .CLK(clk), .RST(rst), .I(m[69]), .Q(
        c[69]) );
  DFF \creg_reg[70]  ( .D(creg_next[70]), .CLK(clk), .RST(rst), .I(m[70]), .Q(
        c[70]) );
  DFF \creg_reg[71]  ( .D(creg_next[71]), .CLK(clk), .RST(rst), .I(m[71]), .Q(
        c[71]) );
  DFF \creg_reg[72]  ( .D(creg_next[72]), .CLK(clk), .RST(rst), .I(m[72]), .Q(
        c[72]) );
  DFF \creg_reg[73]  ( .D(creg_next[73]), .CLK(clk), .RST(rst), .I(m[73]), .Q(
        c[73]) );
  DFF \creg_reg[74]  ( .D(creg_next[74]), .CLK(clk), .RST(rst), .I(m[74]), .Q(
        c[74]) );
  DFF \creg_reg[75]  ( .D(creg_next[75]), .CLK(clk), .RST(rst), .I(m[75]), .Q(
        c[75]) );
  DFF \creg_reg[76]  ( .D(creg_next[76]), .CLK(clk), .RST(rst), .I(m[76]), .Q(
        c[76]) );
  DFF \creg_reg[77]  ( .D(creg_next[77]), .CLK(clk), .RST(rst), .I(m[77]), .Q(
        c[77]) );
  DFF \creg_reg[78]  ( .D(creg_next[78]), .CLK(clk), .RST(rst), .I(m[78]), .Q(
        c[78]) );
  DFF \creg_reg[79]  ( .D(creg_next[79]), .CLK(clk), .RST(rst), .I(m[79]), .Q(
        c[79]) );
  DFF \creg_reg[80]  ( .D(creg_next[80]), .CLK(clk), .RST(rst), .I(m[80]), .Q(
        c[80]) );
  DFF \creg_reg[81]  ( .D(creg_next[81]), .CLK(clk), .RST(rst), .I(m[81]), .Q(
        c[81]) );
  DFF \creg_reg[82]  ( .D(creg_next[82]), .CLK(clk), .RST(rst), .I(m[82]), .Q(
        c[82]) );
  DFF \creg_reg[83]  ( .D(creg_next[83]), .CLK(clk), .RST(rst), .I(m[83]), .Q(
        c[83]) );
  DFF \creg_reg[84]  ( .D(creg_next[84]), .CLK(clk), .RST(rst), .I(m[84]), .Q(
        c[84]) );
  DFF \creg_reg[85]  ( .D(creg_next[85]), .CLK(clk), .RST(rst), .I(m[85]), .Q(
        c[85]) );
  DFF \creg_reg[86]  ( .D(creg_next[86]), .CLK(clk), .RST(rst), .I(m[86]), .Q(
        c[86]) );
  DFF \creg_reg[87]  ( .D(creg_next[87]), .CLK(clk), .RST(rst), .I(m[87]), .Q(
        c[87]) );
  DFF \creg_reg[88]  ( .D(creg_next[88]), .CLK(clk), .RST(rst), .I(m[88]), .Q(
        c[88]) );
  DFF \creg_reg[89]  ( .D(creg_next[89]), .CLK(clk), .RST(rst), .I(m[89]), .Q(
        c[89]) );
  DFF \creg_reg[90]  ( .D(creg_next[90]), .CLK(clk), .RST(rst), .I(m[90]), .Q(
        c[90]) );
  DFF \creg_reg[91]  ( .D(creg_next[91]), .CLK(clk), .RST(rst), .I(m[91]), .Q(
        c[91]) );
  DFF \creg_reg[92]  ( .D(creg_next[92]), .CLK(clk), .RST(rst), .I(m[92]), .Q(
        c[92]) );
  DFF \creg_reg[93]  ( .D(creg_next[93]), .CLK(clk), .RST(rst), .I(m[93]), .Q(
        c[93]) );
  DFF \creg_reg[94]  ( .D(creg_next[94]), .CLK(clk), .RST(rst), .I(m[94]), .Q(
        c[94]) );
  DFF \creg_reg[95]  ( .D(creg_next[95]), .CLK(clk), .RST(rst), .I(m[95]), .Q(
        c[95]) );
  DFF \creg_reg[96]  ( .D(creg_next[96]), .CLK(clk), .RST(rst), .I(m[96]), .Q(
        c[96]) );
  DFF \creg_reg[97]  ( .D(creg_next[97]), .CLK(clk), .RST(rst), .I(m[97]), .Q(
        c[97]) );
  DFF \creg_reg[98]  ( .D(creg_next[98]), .CLK(clk), .RST(rst), .I(m[98]), .Q(
        c[98]) );
  DFF \creg_reg[99]  ( .D(creg_next[99]), .CLK(clk), .RST(rst), .I(m[99]), .Q(
        c[99]) );
  DFF \creg_reg[100]  ( .D(creg_next[100]), .CLK(clk), .RST(rst), .I(m[100]), 
        .Q(c[100]) );
  DFF \creg_reg[101]  ( .D(creg_next[101]), .CLK(clk), .RST(rst), .I(m[101]), 
        .Q(c[101]) );
  DFF \creg_reg[102]  ( .D(creg_next[102]), .CLK(clk), .RST(rst), .I(m[102]), 
        .Q(c[102]) );
  DFF \creg_reg[103]  ( .D(creg_next[103]), .CLK(clk), .RST(rst), .I(m[103]), 
        .Q(c[103]) );
  DFF \creg_reg[104]  ( .D(creg_next[104]), .CLK(clk), .RST(rst), .I(m[104]), 
        .Q(c[104]) );
  DFF \creg_reg[105]  ( .D(creg_next[105]), .CLK(clk), .RST(rst), .I(m[105]), 
        .Q(c[105]) );
  DFF \creg_reg[106]  ( .D(creg_next[106]), .CLK(clk), .RST(rst), .I(m[106]), 
        .Q(c[106]) );
  DFF \creg_reg[107]  ( .D(creg_next[107]), .CLK(clk), .RST(rst), .I(m[107]), 
        .Q(c[107]) );
  DFF \creg_reg[108]  ( .D(creg_next[108]), .CLK(clk), .RST(rst), .I(m[108]), 
        .Q(c[108]) );
  DFF \creg_reg[109]  ( .D(creg_next[109]), .CLK(clk), .RST(rst), .I(m[109]), 
        .Q(c[109]) );
  DFF \creg_reg[110]  ( .D(creg_next[110]), .CLK(clk), .RST(rst), .I(m[110]), 
        .Q(c[110]) );
  DFF \creg_reg[111]  ( .D(creg_next[111]), .CLK(clk), .RST(rst), .I(m[111]), 
        .Q(c[111]) );
  DFF \creg_reg[112]  ( .D(creg_next[112]), .CLK(clk), .RST(rst), .I(m[112]), 
        .Q(c[112]) );
  DFF \creg_reg[113]  ( .D(creg_next[113]), .CLK(clk), .RST(rst), .I(m[113]), 
        .Q(c[113]) );
  DFF \creg_reg[114]  ( .D(creg_next[114]), .CLK(clk), .RST(rst), .I(m[114]), 
        .Q(c[114]) );
  DFF \creg_reg[115]  ( .D(creg_next[115]), .CLK(clk), .RST(rst), .I(m[115]), 
        .Q(c[115]) );
  DFF \creg_reg[116]  ( .D(creg_next[116]), .CLK(clk), .RST(rst), .I(m[116]), 
        .Q(c[116]) );
  DFF \creg_reg[117]  ( .D(creg_next[117]), .CLK(clk), .RST(rst), .I(m[117]), 
        .Q(c[117]) );
  DFF \creg_reg[118]  ( .D(creg_next[118]), .CLK(clk), .RST(rst), .I(m[118]), 
        .Q(c[118]) );
  DFF \creg_reg[119]  ( .D(creg_next[119]), .CLK(clk), .RST(rst), .I(m[119]), 
        .Q(c[119]) );
  DFF \creg_reg[120]  ( .D(creg_next[120]), .CLK(clk), .RST(rst), .I(m[120]), 
        .Q(c[120]) );
  DFF \creg_reg[121]  ( .D(creg_next[121]), .CLK(clk), .RST(rst), .I(m[121]), 
        .Q(c[121]) );
  DFF \creg_reg[122]  ( .D(creg_next[122]), .CLK(clk), .RST(rst), .I(m[122]), 
        .Q(c[122]) );
  DFF \creg_reg[123]  ( .D(creg_next[123]), .CLK(clk), .RST(rst), .I(m[123]), 
        .Q(c[123]) );
  DFF \creg_reg[124]  ( .D(creg_next[124]), .CLK(clk), .RST(rst), .I(m[124]), 
        .Q(c[124]) );
  DFF \creg_reg[125]  ( .D(creg_next[125]), .CLK(clk), .RST(rst), .I(m[125]), 
        .Q(c[125]) );
  DFF \creg_reg[126]  ( .D(creg_next[126]), .CLK(clk), .RST(rst), .I(m[126]), 
        .Q(c[126]) );
  DFF \creg_reg[127]  ( .D(creg_next[127]), .CLK(clk), .RST(rst), .I(m[127]), 
        .Q(c[127]) );
  DFF \creg_reg[128]  ( .D(creg_next[128]), .CLK(clk), .RST(rst), .I(m[128]), 
        .Q(c[128]) );
  DFF \creg_reg[129]  ( .D(creg_next[129]), .CLK(clk), .RST(rst), .I(m[129]), 
        .Q(c[129]) );
  DFF \creg_reg[130]  ( .D(creg_next[130]), .CLK(clk), .RST(rst), .I(m[130]), 
        .Q(c[130]) );
  DFF \creg_reg[131]  ( .D(creg_next[131]), .CLK(clk), .RST(rst), .I(m[131]), 
        .Q(c[131]) );
  DFF \creg_reg[132]  ( .D(creg_next[132]), .CLK(clk), .RST(rst), .I(m[132]), 
        .Q(c[132]) );
  DFF \creg_reg[133]  ( .D(creg_next[133]), .CLK(clk), .RST(rst), .I(m[133]), 
        .Q(c[133]) );
  DFF \creg_reg[134]  ( .D(creg_next[134]), .CLK(clk), .RST(rst), .I(m[134]), 
        .Q(c[134]) );
  DFF \creg_reg[135]  ( .D(creg_next[135]), .CLK(clk), .RST(rst), .I(m[135]), 
        .Q(c[135]) );
  DFF \creg_reg[136]  ( .D(creg_next[136]), .CLK(clk), .RST(rst), .I(m[136]), 
        .Q(c[136]) );
  DFF \creg_reg[137]  ( .D(creg_next[137]), .CLK(clk), .RST(rst), .I(m[137]), 
        .Q(c[137]) );
  DFF \creg_reg[138]  ( .D(creg_next[138]), .CLK(clk), .RST(rst), .I(m[138]), 
        .Q(c[138]) );
  DFF \creg_reg[139]  ( .D(creg_next[139]), .CLK(clk), .RST(rst), .I(m[139]), 
        .Q(c[139]) );
  DFF \creg_reg[140]  ( .D(creg_next[140]), .CLK(clk), .RST(rst), .I(m[140]), 
        .Q(c[140]) );
  DFF \creg_reg[141]  ( .D(creg_next[141]), .CLK(clk), .RST(rst), .I(m[141]), 
        .Q(c[141]) );
  DFF \creg_reg[142]  ( .D(creg_next[142]), .CLK(clk), .RST(rst), .I(m[142]), 
        .Q(c[142]) );
  DFF \creg_reg[143]  ( .D(creg_next[143]), .CLK(clk), .RST(rst), .I(m[143]), 
        .Q(c[143]) );
  DFF \creg_reg[144]  ( .D(creg_next[144]), .CLK(clk), .RST(rst), .I(m[144]), 
        .Q(c[144]) );
  DFF \creg_reg[145]  ( .D(creg_next[145]), .CLK(clk), .RST(rst), .I(m[145]), 
        .Q(c[145]) );
  DFF \creg_reg[146]  ( .D(creg_next[146]), .CLK(clk), .RST(rst), .I(m[146]), 
        .Q(c[146]) );
  DFF \creg_reg[147]  ( .D(creg_next[147]), .CLK(clk), .RST(rst), .I(m[147]), 
        .Q(c[147]) );
  DFF \creg_reg[148]  ( .D(creg_next[148]), .CLK(clk), .RST(rst), .I(m[148]), 
        .Q(c[148]) );
  DFF \creg_reg[149]  ( .D(creg_next[149]), .CLK(clk), .RST(rst), .I(m[149]), 
        .Q(c[149]) );
  DFF \creg_reg[150]  ( .D(creg_next[150]), .CLK(clk), .RST(rst), .I(m[150]), 
        .Q(c[150]) );
  DFF \creg_reg[151]  ( .D(creg_next[151]), .CLK(clk), .RST(rst), .I(m[151]), 
        .Q(c[151]) );
  DFF \creg_reg[152]  ( .D(creg_next[152]), .CLK(clk), .RST(rst), .I(m[152]), 
        .Q(c[152]) );
  DFF \creg_reg[153]  ( .D(creg_next[153]), .CLK(clk), .RST(rst), .I(m[153]), 
        .Q(c[153]) );
  DFF \creg_reg[154]  ( .D(creg_next[154]), .CLK(clk), .RST(rst), .I(m[154]), 
        .Q(c[154]) );
  DFF \creg_reg[155]  ( .D(creg_next[155]), .CLK(clk), .RST(rst), .I(m[155]), 
        .Q(c[155]) );
  DFF \creg_reg[156]  ( .D(creg_next[156]), .CLK(clk), .RST(rst), .I(m[156]), 
        .Q(c[156]) );
  DFF \creg_reg[157]  ( .D(creg_next[157]), .CLK(clk), .RST(rst), .I(m[157]), 
        .Q(c[157]) );
  DFF \creg_reg[158]  ( .D(creg_next[158]), .CLK(clk), .RST(rst), .I(m[158]), 
        .Q(c[158]) );
  DFF \creg_reg[159]  ( .D(creg_next[159]), .CLK(clk), .RST(rst), .I(m[159]), 
        .Q(c[159]) );
  DFF \creg_reg[160]  ( .D(creg_next[160]), .CLK(clk), .RST(rst), .I(m[160]), 
        .Q(c[160]) );
  DFF \creg_reg[161]  ( .D(creg_next[161]), .CLK(clk), .RST(rst), .I(m[161]), 
        .Q(c[161]) );
  DFF \creg_reg[162]  ( .D(creg_next[162]), .CLK(clk), .RST(rst), .I(m[162]), 
        .Q(c[162]) );
  DFF \creg_reg[163]  ( .D(creg_next[163]), .CLK(clk), .RST(rst), .I(m[163]), 
        .Q(c[163]) );
  DFF \creg_reg[164]  ( .D(creg_next[164]), .CLK(clk), .RST(rst), .I(m[164]), 
        .Q(c[164]) );
  DFF \creg_reg[165]  ( .D(creg_next[165]), .CLK(clk), .RST(rst), .I(m[165]), 
        .Q(c[165]) );
  DFF \creg_reg[166]  ( .D(creg_next[166]), .CLK(clk), .RST(rst), .I(m[166]), 
        .Q(c[166]) );
  DFF \creg_reg[167]  ( .D(creg_next[167]), .CLK(clk), .RST(rst), .I(m[167]), 
        .Q(c[167]) );
  DFF \creg_reg[168]  ( .D(creg_next[168]), .CLK(clk), .RST(rst), .I(m[168]), 
        .Q(c[168]) );
  DFF \creg_reg[169]  ( .D(creg_next[169]), .CLK(clk), .RST(rst), .I(m[169]), 
        .Q(c[169]) );
  DFF \creg_reg[170]  ( .D(creg_next[170]), .CLK(clk), .RST(rst), .I(m[170]), 
        .Q(c[170]) );
  DFF \creg_reg[171]  ( .D(creg_next[171]), .CLK(clk), .RST(rst), .I(m[171]), 
        .Q(c[171]) );
  DFF \creg_reg[172]  ( .D(creg_next[172]), .CLK(clk), .RST(rst), .I(m[172]), 
        .Q(c[172]) );
  DFF \creg_reg[173]  ( .D(creg_next[173]), .CLK(clk), .RST(rst), .I(m[173]), 
        .Q(c[173]) );
  DFF \creg_reg[174]  ( .D(creg_next[174]), .CLK(clk), .RST(rst), .I(m[174]), 
        .Q(c[174]) );
  DFF \creg_reg[175]  ( .D(creg_next[175]), .CLK(clk), .RST(rst), .I(m[175]), 
        .Q(c[175]) );
  DFF \creg_reg[176]  ( .D(creg_next[176]), .CLK(clk), .RST(rst), .I(m[176]), 
        .Q(c[176]) );
  DFF \creg_reg[177]  ( .D(creg_next[177]), .CLK(clk), .RST(rst), .I(m[177]), 
        .Q(c[177]) );
  DFF \creg_reg[178]  ( .D(creg_next[178]), .CLK(clk), .RST(rst), .I(m[178]), 
        .Q(c[178]) );
  DFF \creg_reg[179]  ( .D(creg_next[179]), .CLK(clk), .RST(rst), .I(m[179]), 
        .Q(c[179]) );
  DFF \creg_reg[180]  ( .D(creg_next[180]), .CLK(clk), .RST(rst), .I(m[180]), 
        .Q(c[180]) );
  DFF \creg_reg[181]  ( .D(creg_next[181]), .CLK(clk), .RST(rst), .I(m[181]), 
        .Q(c[181]) );
  DFF \creg_reg[182]  ( .D(creg_next[182]), .CLK(clk), .RST(rst), .I(m[182]), 
        .Q(c[182]) );
  DFF \creg_reg[183]  ( .D(creg_next[183]), .CLK(clk), .RST(rst), .I(m[183]), 
        .Q(c[183]) );
  DFF \creg_reg[184]  ( .D(creg_next[184]), .CLK(clk), .RST(rst), .I(m[184]), 
        .Q(c[184]) );
  DFF \creg_reg[185]  ( .D(creg_next[185]), .CLK(clk), .RST(rst), .I(m[185]), 
        .Q(c[185]) );
  DFF \creg_reg[186]  ( .D(creg_next[186]), .CLK(clk), .RST(rst), .I(m[186]), 
        .Q(c[186]) );
  DFF \creg_reg[187]  ( .D(creg_next[187]), .CLK(clk), .RST(rst), .I(m[187]), 
        .Q(c[187]) );
  DFF \creg_reg[188]  ( .D(creg_next[188]), .CLK(clk), .RST(rst), .I(m[188]), 
        .Q(c[188]) );
  DFF \creg_reg[189]  ( .D(creg_next[189]), .CLK(clk), .RST(rst), .I(m[189]), 
        .Q(c[189]) );
  DFF \creg_reg[190]  ( .D(creg_next[190]), .CLK(clk), .RST(rst), .I(m[190]), 
        .Q(c[190]) );
  DFF \creg_reg[191]  ( .D(creg_next[191]), .CLK(clk), .RST(rst), .I(m[191]), 
        .Q(c[191]) );
  DFF \creg_reg[192]  ( .D(creg_next[192]), .CLK(clk), .RST(rst), .I(m[192]), 
        .Q(c[192]) );
  DFF \creg_reg[193]  ( .D(creg_next[193]), .CLK(clk), .RST(rst), .I(m[193]), 
        .Q(c[193]) );
  DFF \creg_reg[194]  ( .D(creg_next[194]), .CLK(clk), .RST(rst), .I(m[194]), 
        .Q(c[194]) );
  DFF \creg_reg[195]  ( .D(creg_next[195]), .CLK(clk), .RST(rst), .I(m[195]), 
        .Q(c[195]) );
  DFF \creg_reg[196]  ( .D(creg_next[196]), .CLK(clk), .RST(rst), .I(m[196]), 
        .Q(c[196]) );
  DFF \creg_reg[197]  ( .D(creg_next[197]), .CLK(clk), .RST(rst), .I(m[197]), 
        .Q(c[197]) );
  DFF \creg_reg[198]  ( .D(creg_next[198]), .CLK(clk), .RST(rst), .I(m[198]), 
        .Q(c[198]) );
  DFF \creg_reg[199]  ( .D(creg_next[199]), .CLK(clk), .RST(rst), .I(m[199]), 
        .Q(c[199]) );
  DFF \creg_reg[200]  ( .D(creg_next[200]), .CLK(clk), .RST(rst), .I(m[200]), 
        .Q(c[200]) );
  DFF \creg_reg[201]  ( .D(creg_next[201]), .CLK(clk), .RST(rst), .I(m[201]), 
        .Q(c[201]) );
  DFF \creg_reg[202]  ( .D(creg_next[202]), .CLK(clk), .RST(rst), .I(m[202]), 
        .Q(c[202]) );
  DFF \creg_reg[203]  ( .D(creg_next[203]), .CLK(clk), .RST(rst), .I(m[203]), 
        .Q(c[203]) );
  DFF \creg_reg[204]  ( .D(creg_next[204]), .CLK(clk), .RST(rst), .I(m[204]), 
        .Q(c[204]) );
  DFF \creg_reg[205]  ( .D(creg_next[205]), .CLK(clk), .RST(rst), .I(m[205]), 
        .Q(c[205]) );
  DFF \creg_reg[206]  ( .D(creg_next[206]), .CLK(clk), .RST(rst), .I(m[206]), 
        .Q(c[206]) );
  DFF \creg_reg[207]  ( .D(creg_next[207]), .CLK(clk), .RST(rst), .I(m[207]), 
        .Q(c[207]) );
  DFF \creg_reg[208]  ( .D(creg_next[208]), .CLK(clk), .RST(rst), .I(m[208]), 
        .Q(c[208]) );
  DFF \creg_reg[209]  ( .D(creg_next[209]), .CLK(clk), .RST(rst), .I(m[209]), 
        .Q(c[209]) );
  DFF \creg_reg[210]  ( .D(creg_next[210]), .CLK(clk), .RST(rst), .I(m[210]), 
        .Q(c[210]) );
  DFF \creg_reg[211]  ( .D(creg_next[211]), .CLK(clk), .RST(rst), .I(m[211]), 
        .Q(c[211]) );
  DFF \creg_reg[212]  ( .D(creg_next[212]), .CLK(clk), .RST(rst), .I(m[212]), 
        .Q(c[212]) );
  DFF \creg_reg[213]  ( .D(creg_next[213]), .CLK(clk), .RST(rst), .I(m[213]), 
        .Q(c[213]) );
  DFF \creg_reg[214]  ( .D(creg_next[214]), .CLK(clk), .RST(rst), .I(m[214]), 
        .Q(c[214]) );
  DFF \creg_reg[215]  ( .D(creg_next[215]), .CLK(clk), .RST(rst), .I(m[215]), 
        .Q(c[215]) );
  DFF \creg_reg[216]  ( .D(creg_next[216]), .CLK(clk), .RST(rst), .I(m[216]), 
        .Q(c[216]) );
  DFF \creg_reg[217]  ( .D(creg_next[217]), .CLK(clk), .RST(rst), .I(m[217]), 
        .Q(c[217]) );
  DFF \creg_reg[218]  ( .D(creg_next[218]), .CLK(clk), .RST(rst), .I(m[218]), 
        .Q(c[218]) );
  DFF \creg_reg[219]  ( .D(creg_next[219]), .CLK(clk), .RST(rst), .I(m[219]), 
        .Q(c[219]) );
  DFF \creg_reg[220]  ( .D(creg_next[220]), .CLK(clk), .RST(rst), .I(m[220]), 
        .Q(c[220]) );
  DFF \creg_reg[221]  ( .D(creg_next[221]), .CLK(clk), .RST(rst), .I(m[221]), 
        .Q(c[221]) );
  DFF \creg_reg[222]  ( .D(creg_next[222]), .CLK(clk), .RST(rst), .I(m[222]), 
        .Q(c[222]) );
  DFF \creg_reg[223]  ( .D(creg_next[223]), .CLK(clk), .RST(rst), .I(m[223]), 
        .Q(c[223]) );
  DFF \creg_reg[224]  ( .D(creg_next[224]), .CLK(clk), .RST(rst), .I(m[224]), 
        .Q(c[224]) );
  DFF \creg_reg[225]  ( .D(creg_next[225]), .CLK(clk), .RST(rst), .I(m[225]), 
        .Q(c[225]) );
  DFF \creg_reg[226]  ( .D(creg_next[226]), .CLK(clk), .RST(rst), .I(m[226]), 
        .Q(c[226]) );
  DFF \creg_reg[227]  ( .D(creg_next[227]), .CLK(clk), .RST(rst), .I(m[227]), 
        .Q(c[227]) );
  DFF \creg_reg[228]  ( .D(creg_next[228]), .CLK(clk), .RST(rst), .I(m[228]), 
        .Q(c[228]) );
  DFF \creg_reg[229]  ( .D(creg_next[229]), .CLK(clk), .RST(rst), .I(m[229]), 
        .Q(c[229]) );
  DFF \creg_reg[230]  ( .D(creg_next[230]), .CLK(clk), .RST(rst), .I(m[230]), 
        .Q(c[230]) );
  DFF \creg_reg[231]  ( .D(creg_next[231]), .CLK(clk), .RST(rst), .I(m[231]), 
        .Q(c[231]) );
  DFF \creg_reg[232]  ( .D(creg_next[232]), .CLK(clk), .RST(rst), .I(m[232]), 
        .Q(c[232]) );
  DFF \creg_reg[233]  ( .D(creg_next[233]), .CLK(clk), .RST(rst), .I(m[233]), 
        .Q(c[233]) );
  DFF \creg_reg[234]  ( .D(creg_next[234]), .CLK(clk), .RST(rst), .I(m[234]), 
        .Q(c[234]) );
  DFF \creg_reg[235]  ( .D(creg_next[235]), .CLK(clk), .RST(rst), .I(m[235]), 
        .Q(c[235]) );
  DFF \creg_reg[236]  ( .D(creg_next[236]), .CLK(clk), .RST(rst), .I(m[236]), 
        .Q(c[236]) );
  DFF \creg_reg[237]  ( .D(creg_next[237]), .CLK(clk), .RST(rst), .I(m[237]), 
        .Q(c[237]) );
  DFF \creg_reg[238]  ( .D(creg_next[238]), .CLK(clk), .RST(rst), .I(m[238]), 
        .Q(c[238]) );
  DFF \creg_reg[239]  ( .D(creg_next[239]), .CLK(clk), .RST(rst), .I(m[239]), 
        .Q(c[239]) );
  DFF \creg_reg[240]  ( .D(creg_next[240]), .CLK(clk), .RST(rst), .I(m[240]), 
        .Q(c[240]) );
  DFF \creg_reg[241]  ( .D(creg_next[241]), .CLK(clk), .RST(rst), .I(m[241]), 
        .Q(c[241]) );
  DFF \creg_reg[242]  ( .D(creg_next[242]), .CLK(clk), .RST(rst), .I(m[242]), 
        .Q(c[242]) );
  DFF \creg_reg[243]  ( .D(creg_next[243]), .CLK(clk), .RST(rst), .I(m[243]), 
        .Q(c[243]) );
  DFF \creg_reg[244]  ( .D(creg_next[244]), .CLK(clk), .RST(rst), .I(m[244]), 
        .Q(c[244]) );
  DFF \creg_reg[245]  ( .D(creg_next[245]), .CLK(clk), .RST(rst), .I(m[245]), 
        .Q(c[245]) );
  DFF \creg_reg[246]  ( .D(creg_next[246]), .CLK(clk), .RST(rst), .I(m[246]), 
        .Q(c[246]) );
  DFF \creg_reg[247]  ( .D(creg_next[247]), .CLK(clk), .RST(rst), .I(m[247]), 
        .Q(c[247]) );
  DFF \creg_reg[248]  ( .D(creg_next[248]), .CLK(clk), .RST(rst), .I(m[248]), 
        .Q(c[248]) );
  DFF \creg_reg[249]  ( .D(creg_next[249]), .CLK(clk), .RST(rst), .I(m[249]), 
        .Q(c[249]) );
  DFF \creg_reg[250]  ( .D(creg_next[250]), .CLK(clk), .RST(rst), .I(m[250]), 
        .Q(c[250]) );
  DFF \creg_reg[251]  ( .D(creg_next[251]), .CLK(clk), .RST(rst), .I(m[251]), 
        .Q(c[251]) );
  DFF \creg_reg[252]  ( .D(creg_next[252]), .CLK(clk), .RST(rst), .I(m[252]), 
        .Q(c[252]) );
  DFF \creg_reg[253]  ( .D(creg_next[253]), .CLK(clk), .RST(rst), .I(m[253]), 
        .Q(c[253]) );
  DFF \creg_reg[254]  ( .D(creg_next[254]), .CLK(clk), .RST(rst), .I(m[254]), 
        .Q(c[254]) );
  DFF \creg_reg[255]  ( .D(creg_next[255]), .CLK(clk), .RST(rst), .I(m[255]), 
        .Q(c[255]) );
  DFF \creg_reg[256]  ( .D(creg_next[256]), .CLK(clk), .RST(rst), .I(m[256]), 
        .Q(c[256]) );
  DFF \creg_reg[257]  ( .D(creg_next[257]), .CLK(clk), .RST(rst), .I(m[257]), 
        .Q(c[257]) );
  DFF \creg_reg[258]  ( .D(creg_next[258]), .CLK(clk), .RST(rst), .I(m[258]), 
        .Q(c[258]) );
  DFF \creg_reg[259]  ( .D(creg_next[259]), .CLK(clk), .RST(rst), .I(m[259]), 
        .Q(c[259]) );
  DFF \creg_reg[260]  ( .D(creg_next[260]), .CLK(clk), .RST(rst), .I(m[260]), 
        .Q(c[260]) );
  DFF \creg_reg[261]  ( .D(creg_next[261]), .CLK(clk), .RST(rst), .I(m[261]), 
        .Q(c[261]) );
  DFF \creg_reg[262]  ( .D(creg_next[262]), .CLK(clk), .RST(rst), .I(m[262]), 
        .Q(c[262]) );
  DFF \creg_reg[263]  ( .D(creg_next[263]), .CLK(clk), .RST(rst), .I(m[263]), 
        .Q(c[263]) );
  DFF \creg_reg[264]  ( .D(creg_next[264]), .CLK(clk), .RST(rst), .I(m[264]), 
        .Q(c[264]) );
  DFF \creg_reg[265]  ( .D(creg_next[265]), .CLK(clk), .RST(rst), .I(m[265]), 
        .Q(c[265]) );
  DFF \creg_reg[266]  ( .D(creg_next[266]), .CLK(clk), .RST(rst), .I(m[266]), 
        .Q(c[266]) );
  DFF \creg_reg[267]  ( .D(creg_next[267]), .CLK(clk), .RST(rst), .I(m[267]), 
        .Q(c[267]) );
  DFF \creg_reg[268]  ( .D(creg_next[268]), .CLK(clk), .RST(rst), .I(m[268]), 
        .Q(c[268]) );
  DFF \creg_reg[269]  ( .D(creg_next[269]), .CLK(clk), .RST(rst), .I(m[269]), 
        .Q(c[269]) );
  DFF \creg_reg[270]  ( .D(creg_next[270]), .CLK(clk), .RST(rst), .I(m[270]), 
        .Q(c[270]) );
  DFF \creg_reg[271]  ( .D(creg_next[271]), .CLK(clk), .RST(rst), .I(m[271]), 
        .Q(c[271]) );
  DFF \creg_reg[272]  ( .D(creg_next[272]), .CLK(clk), .RST(rst), .I(m[272]), 
        .Q(c[272]) );
  DFF \creg_reg[273]  ( .D(creg_next[273]), .CLK(clk), .RST(rst), .I(m[273]), 
        .Q(c[273]) );
  DFF \creg_reg[274]  ( .D(creg_next[274]), .CLK(clk), .RST(rst), .I(m[274]), 
        .Q(c[274]) );
  DFF \creg_reg[275]  ( .D(creg_next[275]), .CLK(clk), .RST(rst), .I(m[275]), 
        .Q(c[275]) );
  DFF \creg_reg[276]  ( .D(creg_next[276]), .CLK(clk), .RST(rst), .I(m[276]), 
        .Q(c[276]) );
  DFF \creg_reg[277]  ( .D(creg_next[277]), .CLK(clk), .RST(rst), .I(m[277]), 
        .Q(c[277]) );
  DFF \creg_reg[278]  ( .D(creg_next[278]), .CLK(clk), .RST(rst), .I(m[278]), 
        .Q(c[278]) );
  DFF \creg_reg[279]  ( .D(creg_next[279]), .CLK(clk), .RST(rst), .I(m[279]), 
        .Q(c[279]) );
  DFF \creg_reg[280]  ( .D(creg_next[280]), .CLK(clk), .RST(rst), .I(m[280]), 
        .Q(c[280]) );
  DFF \creg_reg[281]  ( .D(creg_next[281]), .CLK(clk), .RST(rst), .I(m[281]), 
        .Q(c[281]) );
  DFF \creg_reg[282]  ( .D(creg_next[282]), .CLK(clk), .RST(rst), .I(m[282]), 
        .Q(c[282]) );
  DFF \creg_reg[283]  ( .D(creg_next[283]), .CLK(clk), .RST(rst), .I(m[283]), 
        .Q(c[283]) );
  DFF \creg_reg[284]  ( .D(creg_next[284]), .CLK(clk), .RST(rst), .I(m[284]), 
        .Q(c[284]) );
  DFF \creg_reg[285]  ( .D(creg_next[285]), .CLK(clk), .RST(rst), .I(m[285]), 
        .Q(c[285]) );
  DFF \creg_reg[286]  ( .D(creg_next[286]), .CLK(clk), .RST(rst), .I(m[286]), 
        .Q(c[286]) );
  DFF \creg_reg[287]  ( .D(creg_next[287]), .CLK(clk), .RST(rst), .I(m[287]), 
        .Q(c[287]) );
  DFF \creg_reg[288]  ( .D(creg_next[288]), .CLK(clk), .RST(rst), .I(m[288]), 
        .Q(c[288]) );
  DFF \creg_reg[289]  ( .D(creg_next[289]), .CLK(clk), .RST(rst), .I(m[289]), 
        .Q(c[289]) );
  DFF \creg_reg[290]  ( .D(creg_next[290]), .CLK(clk), .RST(rst), .I(m[290]), 
        .Q(c[290]) );
  DFF \creg_reg[291]  ( .D(creg_next[291]), .CLK(clk), .RST(rst), .I(m[291]), 
        .Q(c[291]) );
  DFF \creg_reg[292]  ( .D(creg_next[292]), .CLK(clk), .RST(rst), .I(m[292]), 
        .Q(c[292]) );
  DFF \creg_reg[293]  ( .D(creg_next[293]), .CLK(clk), .RST(rst), .I(m[293]), 
        .Q(c[293]) );
  DFF \creg_reg[294]  ( .D(creg_next[294]), .CLK(clk), .RST(rst), .I(m[294]), 
        .Q(c[294]) );
  DFF \creg_reg[295]  ( .D(creg_next[295]), .CLK(clk), .RST(rst), .I(m[295]), 
        .Q(c[295]) );
  DFF \creg_reg[296]  ( .D(creg_next[296]), .CLK(clk), .RST(rst), .I(m[296]), 
        .Q(c[296]) );
  DFF \creg_reg[297]  ( .D(creg_next[297]), .CLK(clk), .RST(rst), .I(m[297]), 
        .Q(c[297]) );
  DFF \creg_reg[298]  ( .D(creg_next[298]), .CLK(clk), .RST(rst), .I(m[298]), 
        .Q(c[298]) );
  DFF \creg_reg[299]  ( .D(creg_next[299]), .CLK(clk), .RST(rst), .I(m[299]), 
        .Q(c[299]) );
  DFF \creg_reg[300]  ( .D(creg_next[300]), .CLK(clk), .RST(rst), .I(m[300]), 
        .Q(c[300]) );
  DFF \creg_reg[301]  ( .D(creg_next[301]), .CLK(clk), .RST(rst), .I(m[301]), 
        .Q(c[301]) );
  DFF \creg_reg[302]  ( .D(creg_next[302]), .CLK(clk), .RST(rst), .I(m[302]), 
        .Q(c[302]) );
  DFF \creg_reg[303]  ( .D(creg_next[303]), .CLK(clk), .RST(rst), .I(m[303]), 
        .Q(c[303]) );
  DFF \creg_reg[304]  ( .D(creg_next[304]), .CLK(clk), .RST(rst), .I(m[304]), 
        .Q(c[304]) );
  DFF \creg_reg[305]  ( .D(creg_next[305]), .CLK(clk), .RST(rst), .I(m[305]), 
        .Q(c[305]) );
  DFF \creg_reg[306]  ( .D(creg_next[306]), .CLK(clk), .RST(rst), .I(m[306]), 
        .Q(c[306]) );
  DFF \creg_reg[307]  ( .D(creg_next[307]), .CLK(clk), .RST(rst), .I(m[307]), 
        .Q(c[307]) );
  DFF \creg_reg[308]  ( .D(creg_next[308]), .CLK(clk), .RST(rst), .I(m[308]), 
        .Q(c[308]) );
  DFF \creg_reg[309]  ( .D(creg_next[309]), .CLK(clk), .RST(rst), .I(m[309]), 
        .Q(c[309]) );
  DFF \creg_reg[310]  ( .D(creg_next[310]), .CLK(clk), .RST(rst), .I(m[310]), 
        .Q(c[310]) );
  DFF \creg_reg[311]  ( .D(creg_next[311]), .CLK(clk), .RST(rst), .I(m[311]), 
        .Q(c[311]) );
  DFF \creg_reg[312]  ( .D(creg_next[312]), .CLK(clk), .RST(rst), .I(m[312]), 
        .Q(c[312]) );
  DFF \creg_reg[313]  ( .D(creg_next[313]), .CLK(clk), .RST(rst), .I(m[313]), 
        .Q(c[313]) );
  DFF \creg_reg[314]  ( .D(creg_next[314]), .CLK(clk), .RST(rst), .I(m[314]), 
        .Q(c[314]) );
  DFF \creg_reg[315]  ( .D(creg_next[315]), .CLK(clk), .RST(rst), .I(m[315]), 
        .Q(c[315]) );
  DFF \creg_reg[316]  ( .D(creg_next[316]), .CLK(clk), .RST(rst), .I(m[316]), 
        .Q(c[316]) );
  DFF \creg_reg[317]  ( .D(creg_next[317]), .CLK(clk), .RST(rst), .I(m[317]), 
        .Q(c[317]) );
  DFF \creg_reg[318]  ( .D(creg_next[318]), .CLK(clk), .RST(rst), .I(m[318]), 
        .Q(c[318]) );
  DFF \creg_reg[319]  ( .D(creg_next[319]), .CLK(clk), .RST(rst), .I(m[319]), 
        .Q(c[319]) );
  DFF \creg_reg[320]  ( .D(creg_next[320]), .CLK(clk), .RST(rst), .I(m[320]), 
        .Q(c[320]) );
  DFF \creg_reg[321]  ( .D(creg_next[321]), .CLK(clk), .RST(rst), .I(m[321]), 
        .Q(c[321]) );
  DFF \creg_reg[322]  ( .D(creg_next[322]), .CLK(clk), .RST(rst), .I(m[322]), 
        .Q(c[322]) );
  DFF \creg_reg[323]  ( .D(creg_next[323]), .CLK(clk), .RST(rst), .I(m[323]), 
        .Q(c[323]) );
  DFF \creg_reg[324]  ( .D(creg_next[324]), .CLK(clk), .RST(rst), .I(m[324]), 
        .Q(c[324]) );
  DFF \creg_reg[325]  ( .D(creg_next[325]), .CLK(clk), .RST(rst), .I(m[325]), 
        .Q(c[325]) );
  DFF \creg_reg[326]  ( .D(creg_next[326]), .CLK(clk), .RST(rst), .I(m[326]), 
        .Q(c[326]) );
  DFF \creg_reg[327]  ( .D(creg_next[327]), .CLK(clk), .RST(rst), .I(m[327]), 
        .Q(c[327]) );
  DFF \creg_reg[328]  ( .D(creg_next[328]), .CLK(clk), .RST(rst), .I(m[328]), 
        .Q(c[328]) );
  DFF \creg_reg[329]  ( .D(creg_next[329]), .CLK(clk), .RST(rst), .I(m[329]), 
        .Q(c[329]) );
  DFF \creg_reg[330]  ( .D(creg_next[330]), .CLK(clk), .RST(rst), .I(m[330]), 
        .Q(c[330]) );
  DFF \creg_reg[331]  ( .D(creg_next[331]), .CLK(clk), .RST(rst), .I(m[331]), 
        .Q(c[331]) );
  DFF \creg_reg[332]  ( .D(creg_next[332]), .CLK(clk), .RST(rst), .I(m[332]), 
        .Q(c[332]) );
  DFF \creg_reg[333]  ( .D(creg_next[333]), .CLK(clk), .RST(rst), .I(m[333]), 
        .Q(c[333]) );
  DFF \creg_reg[334]  ( .D(creg_next[334]), .CLK(clk), .RST(rst), .I(m[334]), 
        .Q(c[334]) );
  DFF \creg_reg[335]  ( .D(creg_next[335]), .CLK(clk), .RST(rst), .I(m[335]), 
        .Q(c[335]) );
  DFF \creg_reg[336]  ( .D(creg_next[336]), .CLK(clk), .RST(rst), .I(m[336]), 
        .Q(c[336]) );
  DFF \creg_reg[337]  ( .D(creg_next[337]), .CLK(clk), .RST(rst), .I(m[337]), 
        .Q(c[337]) );
  DFF \creg_reg[338]  ( .D(creg_next[338]), .CLK(clk), .RST(rst), .I(m[338]), 
        .Q(c[338]) );
  DFF \creg_reg[339]  ( .D(creg_next[339]), .CLK(clk), .RST(rst), .I(m[339]), 
        .Q(c[339]) );
  DFF \creg_reg[340]  ( .D(creg_next[340]), .CLK(clk), .RST(rst), .I(m[340]), 
        .Q(c[340]) );
  DFF \creg_reg[341]  ( .D(creg_next[341]), .CLK(clk), .RST(rst), .I(m[341]), 
        .Q(c[341]) );
  DFF \creg_reg[342]  ( .D(creg_next[342]), .CLK(clk), .RST(rst), .I(m[342]), 
        .Q(c[342]) );
  DFF \creg_reg[343]  ( .D(creg_next[343]), .CLK(clk), .RST(rst), .I(m[343]), 
        .Q(c[343]) );
  DFF \creg_reg[344]  ( .D(creg_next[344]), .CLK(clk), .RST(rst), .I(m[344]), 
        .Q(c[344]) );
  DFF \creg_reg[345]  ( .D(creg_next[345]), .CLK(clk), .RST(rst), .I(m[345]), 
        .Q(c[345]) );
  DFF \creg_reg[346]  ( .D(creg_next[346]), .CLK(clk), .RST(rst), .I(m[346]), 
        .Q(c[346]) );
  DFF \creg_reg[347]  ( .D(creg_next[347]), .CLK(clk), .RST(rst), .I(m[347]), 
        .Q(c[347]) );
  DFF \creg_reg[348]  ( .D(creg_next[348]), .CLK(clk), .RST(rst), .I(m[348]), 
        .Q(c[348]) );
  DFF \creg_reg[349]  ( .D(creg_next[349]), .CLK(clk), .RST(rst), .I(m[349]), 
        .Q(c[349]) );
  DFF \creg_reg[350]  ( .D(creg_next[350]), .CLK(clk), .RST(rst), .I(m[350]), 
        .Q(c[350]) );
  DFF \creg_reg[351]  ( .D(creg_next[351]), .CLK(clk), .RST(rst), .I(m[351]), 
        .Q(c[351]) );
  DFF \creg_reg[352]  ( .D(creg_next[352]), .CLK(clk), .RST(rst), .I(m[352]), 
        .Q(c[352]) );
  DFF \creg_reg[353]  ( .D(creg_next[353]), .CLK(clk), .RST(rst), .I(m[353]), 
        .Q(c[353]) );
  DFF \creg_reg[354]  ( .D(creg_next[354]), .CLK(clk), .RST(rst), .I(m[354]), 
        .Q(c[354]) );
  DFF \creg_reg[355]  ( .D(creg_next[355]), .CLK(clk), .RST(rst), .I(m[355]), 
        .Q(c[355]) );
  DFF \creg_reg[356]  ( .D(creg_next[356]), .CLK(clk), .RST(rst), .I(m[356]), 
        .Q(c[356]) );
  DFF \creg_reg[357]  ( .D(creg_next[357]), .CLK(clk), .RST(rst), .I(m[357]), 
        .Q(c[357]) );
  DFF \creg_reg[358]  ( .D(creg_next[358]), .CLK(clk), .RST(rst), .I(m[358]), 
        .Q(c[358]) );
  DFF \creg_reg[359]  ( .D(creg_next[359]), .CLK(clk), .RST(rst), .I(m[359]), 
        .Q(c[359]) );
  DFF \creg_reg[360]  ( .D(creg_next[360]), .CLK(clk), .RST(rst), .I(m[360]), 
        .Q(c[360]) );
  DFF \creg_reg[361]  ( .D(creg_next[361]), .CLK(clk), .RST(rst), .I(m[361]), 
        .Q(c[361]) );
  DFF \creg_reg[362]  ( .D(creg_next[362]), .CLK(clk), .RST(rst), .I(m[362]), 
        .Q(c[362]) );
  DFF \creg_reg[363]  ( .D(creg_next[363]), .CLK(clk), .RST(rst), .I(m[363]), 
        .Q(c[363]) );
  DFF \creg_reg[364]  ( .D(creg_next[364]), .CLK(clk), .RST(rst), .I(m[364]), 
        .Q(c[364]) );
  DFF \creg_reg[365]  ( .D(creg_next[365]), .CLK(clk), .RST(rst), .I(m[365]), 
        .Q(c[365]) );
  DFF \creg_reg[366]  ( .D(creg_next[366]), .CLK(clk), .RST(rst), .I(m[366]), 
        .Q(c[366]) );
  DFF \creg_reg[367]  ( .D(creg_next[367]), .CLK(clk), .RST(rst), .I(m[367]), 
        .Q(c[367]) );
  DFF \creg_reg[368]  ( .D(creg_next[368]), .CLK(clk), .RST(rst), .I(m[368]), 
        .Q(c[368]) );
  DFF \creg_reg[369]  ( .D(creg_next[369]), .CLK(clk), .RST(rst), .I(m[369]), 
        .Q(c[369]) );
  DFF \creg_reg[370]  ( .D(creg_next[370]), .CLK(clk), .RST(rst), .I(m[370]), 
        .Q(c[370]) );
  DFF \creg_reg[371]  ( .D(creg_next[371]), .CLK(clk), .RST(rst), .I(m[371]), 
        .Q(c[371]) );
  DFF \creg_reg[372]  ( .D(creg_next[372]), .CLK(clk), .RST(rst), .I(m[372]), 
        .Q(c[372]) );
  DFF \creg_reg[373]  ( .D(creg_next[373]), .CLK(clk), .RST(rst), .I(m[373]), 
        .Q(c[373]) );
  DFF \creg_reg[374]  ( .D(creg_next[374]), .CLK(clk), .RST(rst), .I(m[374]), 
        .Q(c[374]) );
  DFF \creg_reg[375]  ( .D(creg_next[375]), .CLK(clk), .RST(rst), .I(m[375]), 
        .Q(c[375]) );
  DFF \creg_reg[376]  ( .D(creg_next[376]), .CLK(clk), .RST(rst), .I(m[376]), 
        .Q(c[376]) );
  DFF \creg_reg[377]  ( .D(creg_next[377]), .CLK(clk), .RST(rst), .I(m[377]), 
        .Q(c[377]) );
  DFF \creg_reg[378]  ( .D(creg_next[378]), .CLK(clk), .RST(rst), .I(m[378]), 
        .Q(c[378]) );
  DFF \creg_reg[379]  ( .D(creg_next[379]), .CLK(clk), .RST(rst), .I(m[379]), 
        .Q(c[379]) );
  DFF \creg_reg[380]  ( .D(creg_next[380]), .CLK(clk), .RST(rst), .I(m[380]), 
        .Q(c[380]) );
  DFF \creg_reg[381]  ( .D(creg_next[381]), .CLK(clk), .RST(rst), .I(m[381]), 
        .Q(c[381]) );
  DFF \creg_reg[382]  ( .D(creg_next[382]), .CLK(clk), .RST(rst), .I(m[382]), 
        .Q(c[382]) );
  DFF \creg_reg[383]  ( .D(creg_next[383]), .CLK(clk), .RST(rst), .I(m[383]), 
        .Q(c[383]) );
  DFF \creg_reg[384]  ( .D(creg_next[384]), .CLK(clk), .RST(rst), .I(m[384]), 
        .Q(c[384]) );
  DFF \creg_reg[385]  ( .D(creg_next[385]), .CLK(clk), .RST(rst), .I(m[385]), 
        .Q(c[385]) );
  DFF \creg_reg[386]  ( .D(creg_next[386]), .CLK(clk), .RST(rst), .I(m[386]), 
        .Q(c[386]) );
  DFF \creg_reg[387]  ( .D(creg_next[387]), .CLK(clk), .RST(rst), .I(m[387]), 
        .Q(c[387]) );
  DFF \creg_reg[388]  ( .D(creg_next[388]), .CLK(clk), .RST(rst), .I(m[388]), 
        .Q(c[388]) );
  DFF \creg_reg[389]  ( .D(creg_next[389]), .CLK(clk), .RST(rst), .I(m[389]), 
        .Q(c[389]) );
  DFF \creg_reg[390]  ( .D(creg_next[390]), .CLK(clk), .RST(rst), .I(m[390]), 
        .Q(c[390]) );
  DFF \creg_reg[391]  ( .D(creg_next[391]), .CLK(clk), .RST(rst), .I(m[391]), 
        .Q(c[391]) );
  DFF \creg_reg[392]  ( .D(creg_next[392]), .CLK(clk), .RST(rst), .I(m[392]), 
        .Q(c[392]) );
  DFF \creg_reg[393]  ( .D(creg_next[393]), .CLK(clk), .RST(rst), .I(m[393]), 
        .Q(c[393]) );
  DFF \creg_reg[394]  ( .D(creg_next[394]), .CLK(clk), .RST(rst), .I(m[394]), 
        .Q(c[394]) );
  DFF \creg_reg[395]  ( .D(creg_next[395]), .CLK(clk), .RST(rst), .I(m[395]), 
        .Q(c[395]) );
  DFF \creg_reg[396]  ( .D(creg_next[396]), .CLK(clk), .RST(rst), .I(m[396]), 
        .Q(c[396]) );
  DFF \creg_reg[397]  ( .D(creg_next[397]), .CLK(clk), .RST(rst), .I(m[397]), 
        .Q(c[397]) );
  DFF \creg_reg[398]  ( .D(creg_next[398]), .CLK(clk), .RST(rst), .I(m[398]), 
        .Q(c[398]) );
  DFF \creg_reg[399]  ( .D(creg_next[399]), .CLK(clk), .RST(rst), .I(m[399]), 
        .Q(c[399]) );
  DFF \creg_reg[400]  ( .D(creg_next[400]), .CLK(clk), .RST(rst), .I(m[400]), 
        .Q(c[400]) );
  DFF \creg_reg[401]  ( .D(creg_next[401]), .CLK(clk), .RST(rst), .I(m[401]), 
        .Q(c[401]) );
  DFF \creg_reg[402]  ( .D(creg_next[402]), .CLK(clk), .RST(rst), .I(m[402]), 
        .Q(c[402]) );
  DFF \creg_reg[403]  ( .D(creg_next[403]), .CLK(clk), .RST(rst), .I(m[403]), 
        .Q(c[403]) );
  DFF \creg_reg[404]  ( .D(creg_next[404]), .CLK(clk), .RST(rst), .I(m[404]), 
        .Q(c[404]) );
  DFF \creg_reg[405]  ( .D(creg_next[405]), .CLK(clk), .RST(rst), .I(m[405]), 
        .Q(c[405]) );
  DFF \creg_reg[406]  ( .D(creg_next[406]), .CLK(clk), .RST(rst), .I(m[406]), 
        .Q(c[406]) );
  DFF \creg_reg[407]  ( .D(creg_next[407]), .CLK(clk), .RST(rst), .I(m[407]), 
        .Q(c[407]) );
  DFF \creg_reg[408]  ( .D(creg_next[408]), .CLK(clk), .RST(rst), .I(m[408]), 
        .Q(c[408]) );
  DFF \creg_reg[409]  ( .D(creg_next[409]), .CLK(clk), .RST(rst), .I(m[409]), 
        .Q(c[409]) );
  DFF \creg_reg[410]  ( .D(creg_next[410]), .CLK(clk), .RST(rst), .I(m[410]), 
        .Q(c[410]) );
  DFF \creg_reg[411]  ( .D(creg_next[411]), .CLK(clk), .RST(rst), .I(m[411]), 
        .Q(c[411]) );
  DFF \creg_reg[412]  ( .D(creg_next[412]), .CLK(clk), .RST(rst), .I(m[412]), 
        .Q(c[412]) );
  DFF \creg_reg[413]  ( .D(creg_next[413]), .CLK(clk), .RST(rst), .I(m[413]), 
        .Q(c[413]) );
  DFF \creg_reg[414]  ( .D(creg_next[414]), .CLK(clk), .RST(rst), .I(m[414]), 
        .Q(c[414]) );
  DFF \creg_reg[415]  ( .D(creg_next[415]), .CLK(clk), .RST(rst), .I(m[415]), 
        .Q(c[415]) );
  DFF \creg_reg[416]  ( .D(creg_next[416]), .CLK(clk), .RST(rst), .I(m[416]), 
        .Q(c[416]) );
  DFF \creg_reg[417]  ( .D(creg_next[417]), .CLK(clk), .RST(rst), .I(m[417]), 
        .Q(c[417]) );
  DFF \creg_reg[418]  ( .D(creg_next[418]), .CLK(clk), .RST(rst), .I(m[418]), 
        .Q(c[418]) );
  DFF \creg_reg[419]  ( .D(creg_next[419]), .CLK(clk), .RST(rst), .I(m[419]), 
        .Q(c[419]) );
  DFF \creg_reg[420]  ( .D(creg_next[420]), .CLK(clk), .RST(rst), .I(m[420]), 
        .Q(c[420]) );
  DFF \creg_reg[421]  ( .D(creg_next[421]), .CLK(clk), .RST(rst), .I(m[421]), 
        .Q(c[421]) );
  DFF \creg_reg[422]  ( .D(creg_next[422]), .CLK(clk), .RST(rst), .I(m[422]), 
        .Q(c[422]) );
  DFF \creg_reg[423]  ( .D(creg_next[423]), .CLK(clk), .RST(rst), .I(m[423]), 
        .Q(c[423]) );
  DFF \creg_reg[424]  ( .D(creg_next[424]), .CLK(clk), .RST(rst), .I(m[424]), 
        .Q(c[424]) );
  DFF \creg_reg[425]  ( .D(creg_next[425]), .CLK(clk), .RST(rst), .I(m[425]), 
        .Q(c[425]) );
  DFF \creg_reg[426]  ( .D(creg_next[426]), .CLK(clk), .RST(rst), .I(m[426]), 
        .Q(c[426]) );
  DFF \creg_reg[427]  ( .D(creg_next[427]), .CLK(clk), .RST(rst), .I(m[427]), 
        .Q(c[427]) );
  DFF \creg_reg[428]  ( .D(creg_next[428]), .CLK(clk), .RST(rst), .I(m[428]), 
        .Q(c[428]) );
  DFF \creg_reg[429]  ( .D(creg_next[429]), .CLK(clk), .RST(rst), .I(m[429]), 
        .Q(c[429]) );
  DFF \creg_reg[430]  ( .D(creg_next[430]), .CLK(clk), .RST(rst), .I(m[430]), 
        .Q(c[430]) );
  DFF \creg_reg[431]  ( .D(creg_next[431]), .CLK(clk), .RST(rst), .I(m[431]), 
        .Q(c[431]) );
  DFF \creg_reg[432]  ( .D(creg_next[432]), .CLK(clk), .RST(rst), .I(m[432]), 
        .Q(c[432]) );
  DFF \creg_reg[433]  ( .D(creg_next[433]), .CLK(clk), .RST(rst), .I(m[433]), 
        .Q(c[433]) );
  DFF \creg_reg[434]  ( .D(creg_next[434]), .CLK(clk), .RST(rst), .I(m[434]), 
        .Q(c[434]) );
  DFF \creg_reg[435]  ( .D(creg_next[435]), .CLK(clk), .RST(rst), .I(m[435]), 
        .Q(c[435]) );
  DFF \creg_reg[436]  ( .D(creg_next[436]), .CLK(clk), .RST(rst), .I(m[436]), 
        .Q(c[436]) );
  DFF \creg_reg[437]  ( .D(creg_next[437]), .CLK(clk), .RST(rst), .I(m[437]), 
        .Q(c[437]) );
  DFF \creg_reg[438]  ( .D(creg_next[438]), .CLK(clk), .RST(rst), .I(m[438]), 
        .Q(c[438]) );
  DFF \creg_reg[439]  ( .D(creg_next[439]), .CLK(clk), .RST(rst), .I(m[439]), 
        .Q(c[439]) );
  DFF \creg_reg[440]  ( .D(creg_next[440]), .CLK(clk), .RST(rst), .I(m[440]), 
        .Q(c[440]) );
  DFF \creg_reg[441]  ( .D(creg_next[441]), .CLK(clk), .RST(rst), .I(m[441]), 
        .Q(c[441]) );
  DFF \creg_reg[442]  ( .D(creg_next[442]), .CLK(clk), .RST(rst), .I(m[442]), 
        .Q(c[442]) );
  DFF \creg_reg[443]  ( .D(creg_next[443]), .CLK(clk), .RST(rst), .I(m[443]), 
        .Q(c[443]) );
  DFF \creg_reg[444]  ( .D(creg_next[444]), .CLK(clk), .RST(rst), .I(m[444]), 
        .Q(c[444]) );
  DFF \creg_reg[445]  ( .D(creg_next[445]), .CLK(clk), .RST(rst), .I(m[445]), 
        .Q(c[445]) );
  DFF \creg_reg[446]  ( .D(creg_next[446]), .CLK(clk), .RST(rst), .I(m[446]), 
        .Q(c[446]) );
  DFF \creg_reg[447]  ( .D(creg_next[447]), .CLK(clk), .RST(rst), .I(m[447]), 
        .Q(c[447]) );
  DFF \creg_reg[448]  ( .D(creg_next[448]), .CLK(clk), .RST(rst), .I(m[448]), 
        .Q(c[448]) );
  DFF \creg_reg[449]  ( .D(creg_next[449]), .CLK(clk), .RST(rst), .I(m[449]), 
        .Q(c[449]) );
  DFF \creg_reg[450]  ( .D(creg_next[450]), .CLK(clk), .RST(rst), .I(m[450]), 
        .Q(c[450]) );
  DFF \creg_reg[451]  ( .D(creg_next[451]), .CLK(clk), .RST(rst), .I(m[451]), 
        .Q(c[451]) );
  DFF \creg_reg[452]  ( .D(creg_next[452]), .CLK(clk), .RST(rst), .I(m[452]), 
        .Q(c[452]) );
  DFF \creg_reg[453]  ( .D(creg_next[453]), .CLK(clk), .RST(rst), .I(m[453]), 
        .Q(c[453]) );
  DFF \creg_reg[454]  ( .D(creg_next[454]), .CLK(clk), .RST(rst), .I(m[454]), 
        .Q(c[454]) );
  DFF \creg_reg[455]  ( .D(creg_next[455]), .CLK(clk), .RST(rst), .I(m[455]), 
        .Q(c[455]) );
  DFF \creg_reg[456]  ( .D(creg_next[456]), .CLK(clk), .RST(rst), .I(m[456]), 
        .Q(c[456]) );
  DFF \creg_reg[457]  ( .D(creg_next[457]), .CLK(clk), .RST(rst), .I(m[457]), 
        .Q(c[457]) );
  DFF \creg_reg[458]  ( .D(creg_next[458]), .CLK(clk), .RST(rst), .I(m[458]), 
        .Q(c[458]) );
  DFF \creg_reg[459]  ( .D(creg_next[459]), .CLK(clk), .RST(rst), .I(m[459]), 
        .Q(c[459]) );
  DFF \creg_reg[460]  ( .D(creg_next[460]), .CLK(clk), .RST(rst), .I(m[460]), 
        .Q(c[460]) );
  DFF \creg_reg[461]  ( .D(creg_next[461]), .CLK(clk), .RST(rst), .I(m[461]), 
        .Q(c[461]) );
  DFF \creg_reg[462]  ( .D(creg_next[462]), .CLK(clk), .RST(rst), .I(m[462]), 
        .Q(c[462]) );
  DFF \creg_reg[463]  ( .D(creg_next[463]), .CLK(clk), .RST(rst), .I(m[463]), 
        .Q(c[463]) );
  DFF \creg_reg[464]  ( .D(creg_next[464]), .CLK(clk), .RST(rst), .I(m[464]), 
        .Q(c[464]) );
  DFF \creg_reg[465]  ( .D(creg_next[465]), .CLK(clk), .RST(rst), .I(m[465]), 
        .Q(c[465]) );
  DFF \creg_reg[466]  ( .D(creg_next[466]), .CLK(clk), .RST(rst), .I(m[466]), 
        .Q(c[466]) );
  DFF \creg_reg[467]  ( .D(creg_next[467]), .CLK(clk), .RST(rst), .I(m[467]), 
        .Q(c[467]) );
  DFF \creg_reg[468]  ( .D(creg_next[468]), .CLK(clk), .RST(rst), .I(m[468]), 
        .Q(c[468]) );
  DFF \creg_reg[469]  ( .D(creg_next[469]), .CLK(clk), .RST(rst), .I(m[469]), 
        .Q(c[469]) );
  DFF \creg_reg[470]  ( .D(creg_next[470]), .CLK(clk), .RST(rst), .I(m[470]), 
        .Q(c[470]) );
  DFF \creg_reg[471]  ( .D(creg_next[471]), .CLK(clk), .RST(rst), .I(m[471]), 
        .Q(c[471]) );
  DFF \creg_reg[472]  ( .D(creg_next[472]), .CLK(clk), .RST(rst), .I(m[472]), 
        .Q(c[472]) );
  DFF \creg_reg[473]  ( .D(creg_next[473]), .CLK(clk), .RST(rst), .I(m[473]), 
        .Q(c[473]) );
  DFF \creg_reg[474]  ( .D(creg_next[474]), .CLK(clk), .RST(rst), .I(m[474]), 
        .Q(c[474]) );
  DFF \creg_reg[475]  ( .D(creg_next[475]), .CLK(clk), .RST(rst), .I(m[475]), 
        .Q(c[475]) );
  DFF \creg_reg[476]  ( .D(creg_next[476]), .CLK(clk), .RST(rst), .I(m[476]), 
        .Q(c[476]) );
  DFF \creg_reg[477]  ( .D(creg_next[477]), .CLK(clk), .RST(rst), .I(m[477]), 
        .Q(c[477]) );
  DFF \creg_reg[478]  ( .D(creg_next[478]), .CLK(clk), .RST(rst), .I(m[478]), 
        .Q(c[478]) );
  DFF \creg_reg[479]  ( .D(creg_next[479]), .CLK(clk), .RST(rst), .I(m[479]), 
        .Q(c[479]) );
  DFF \creg_reg[480]  ( .D(creg_next[480]), .CLK(clk), .RST(rst), .I(m[480]), 
        .Q(c[480]) );
  DFF \creg_reg[481]  ( .D(creg_next[481]), .CLK(clk), .RST(rst), .I(m[481]), 
        .Q(c[481]) );
  DFF \creg_reg[482]  ( .D(creg_next[482]), .CLK(clk), .RST(rst), .I(m[482]), 
        .Q(c[482]) );
  DFF \creg_reg[483]  ( .D(creg_next[483]), .CLK(clk), .RST(rst), .I(m[483]), 
        .Q(c[483]) );
  DFF \creg_reg[484]  ( .D(creg_next[484]), .CLK(clk), .RST(rst), .I(m[484]), 
        .Q(c[484]) );
  DFF \creg_reg[485]  ( .D(creg_next[485]), .CLK(clk), .RST(rst), .I(m[485]), 
        .Q(c[485]) );
  DFF \creg_reg[486]  ( .D(creg_next[486]), .CLK(clk), .RST(rst), .I(m[486]), 
        .Q(c[486]) );
  DFF \creg_reg[487]  ( .D(creg_next[487]), .CLK(clk), .RST(rst), .I(m[487]), 
        .Q(c[487]) );
  DFF \creg_reg[488]  ( .D(creg_next[488]), .CLK(clk), .RST(rst), .I(m[488]), 
        .Q(c[488]) );
  DFF \creg_reg[489]  ( .D(creg_next[489]), .CLK(clk), .RST(rst), .I(m[489]), 
        .Q(c[489]) );
  DFF \creg_reg[490]  ( .D(creg_next[490]), .CLK(clk), .RST(rst), .I(m[490]), 
        .Q(c[490]) );
  DFF \creg_reg[491]  ( .D(creg_next[491]), .CLK(clk), .RST(rst), .I(m[491]), 
        .Q(c[491]) );
  DFF \creg_reg[492]  ( .D(creg_next[492]), .CLK(clk), .RST(rst), .I(m[492]), 
        .Q(c[492]) );
  DFF \creg_reg[493]  ( .D(creg_next[493]), .CLK(clk), .RST(rst), .I(m[493]), 
        .Q(c[493]) );
  DFF \creg_reg[494]  ( .D(creg_next[494]), .CLK(clk), .RST(rst), .I(m[494]), 
        .Q(c[494]) );
  DFF \creg_reg[495]  ( .D(creg_next[495]), .CLK(clk), .RST(rst), .I(m[495]), 
        .Q(c[495]) );
  DFF \creg_reg[496]  ( .D(creg_next[496]), .CLK(clk), .RST(rst), .I(m[496]), 
        .Q(c[496]) );
  DFF \creg_reg[497]  ( .D(creg_next[497]), .CLK(clk), .RST(rst), .I(m[497]), 
        .Q(c[497]) );
  DFF \creg_reg[498]  ( .D(creg_next[498]), .CLK(clk), .RST(rst), .I(m[498]), 
        .Q(c[498]) );
  DFF \creg_reg[499]  ( .D(creg_next[499]), .CLK(clk), .RST(rst), .I(m[499]), 
        .Q(c[499]) );
  DFF \creg_reg[500]  ( .D(creg_next[500]), .CLK(clk), .RST(rst), .I(m[500]), 
        .Q(c[500]) );
  DFF \creg_reg[501]  ( .D(creg_next[501]), .CLK(clk), .RST(rst), .I(m[501]), 
        .Q(c[501]) );
  DFF \creg_reg[502]  ( .D(creg_next[502]), .CLK(clk), .RST(rst), .I(m[502]), 
        .Q(c[502]) );
  DFF \creg_reg[503]  ( .D(creg_next[503]), .CLK(clk), .RST(rst), .I(m[503]), 
        .Q(c[503]) );
  DFF \creg_reg[504]  ( .D(creg_next[504]), .CLK(clk), .RST(rst), .I(m[504]), 
        .Q(c[504]) );
  DFF \creg_reg[505]  ( .D(creg_next[505]), .CLK(clk), .RST(rst), .I(m[505]), 
        .Q(c[505]) );
  DFF \creg_reg[506]  ( .D(creg_next[506]), .CLK(clk), .RST(rst), .I(m[506]), 
        .Q(c[506]) );
  DFF \creg_reg[507]  ( .D(creg_next[507]), .CLK(clk), .RST(rst), .I(m[507]), 
        .Q(c[507]) );
  DFF \creg_reg[508]  ( .D(creg_next[508]), .CLK(clk), .RST(rst), .I(m[508]), 
        .Q(c[508]) );
  DFF \creg_reg[509]  ( .D(creg_next[509]), .CLK(clk), .RST(rst), .I(m[509]), 
        .Q(c[509]) );
  DFF \creg_reg[510]  ( .D(creg_next[510]), .CLK(clk), .RST(rst), .I(m[510]), 
        .Q(c[510]) );
  DFF \creg_reg[511]  ( .D(creg_next[511]), .CLK(clk), .RST(rst), .I(m[511]), 
        .Q(c[511]) );
  XOR U524 ( .A(start_in[511]), .B(mul_pow), .Z(n8) );
  NANDN U525 ( .A(first_one), .B(n521), .Z(n6) );
  NAND U526 ( .A(n522), .B(ein[511]), .Z(n521) );
  AND U527 ( .A(mul_pow), .B(start_in[511]), .Z(n522) );
  NAND U528 ( .A(n523), .B(n524), .Z(_0_net_) );
  NANDN U529 ( .A(mul_pow), .B(first_one), .Z(n524) );
  NAND U530 ( .A(first_one), .B(ein[511]), .Z(n523) );
endmodule

