
module sum_N16384_CC8 ( clk, rst, a, b, c );
  input [2047:0] a;
  input [2047:0] b;
  output [2047:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        carry_on) );
  XOR U4 ( .A(n2), .B(n3), .Z(carry_on_d) );
  ANDN U5 ( .B(n4), .A(n5), .Z(n2) );
  XOR U6 ( .A(b[2047]), .B(n3), .Z(n4) );
  XNOR U7 ( .A(b[9]), .B(n6), .Z(c[9]) );
  XNOR U8 ( .A(b[99]), .B(n7), .Z(c[99]) );
  XNOR U9 ( .A(b[999]), .B(n8), .Z(c[999]) );
  XNOR U10 ( .A(b[998]), .B(n9), .Z(c[998]) );
  XNOR U11 ( .A(b[997]), .B(n10), .Z(c[997]) );
  XNOR U12 ( .A(b[996]), .B(n11), .Z(c[996]) );
  XNOR U13 ( .A(b[995]), .B(n12), .Z(c[995]) );
  XNOR U14 ( .A(b[994]), .B(n13), .Z(c[994]) );
  XNOR U15 ( .A(b[993]), .B(n14), .Z(c[993]) );
  XNOR U16 ( .A(b[992]), .B(n15), .Z(c[992]) );
  XNOR U17 ( .A(b[991]), .B(n16), .Z(c[991]) );
  XNOR U18 ( .A(b[990]), .B(n17), .Z(c[990]) );
  XNOR U19 ( .A(b[98]), .B(n18), .Z(c[98]) );
  XNOR U20 ( .A(b[989]), .B(n19), .Z(c[989]) );
  XNOR U21 ( .A(b[988]), .B(n20), .Z(c[988]) );
  XNOR U22 ( .A(b[987]), .B(n21), .Z(c[987]) );
  XNOR U23 ( .A(b[986]), .B(n22), .Z(c[986]) );
  XNOR U24 ( .A(b[985]), .B(n23), .Z(c[985]) );
  XNOR U25 ( .A(b[984]), .B(n24), .Z(c[984]) );
  XNOR U26 ( .A(b[983]), .B(n25), .Z(c[983]) );
  XNOR U27 ( .A(b[982]), .B(n26), .Z(c[982]) );
  XNOR U28 ( .A(b[981]), .B(n27), .Z(c[981]) );
  XNOR U29 ( .A(b[980]), .B(n28), .Z(c[980]) );
  XNOR U30 ( .A(b[97]), .B(n29), .Z(c[97]) );
  XNOR U31 ( .A(b[979]), .B(n30), .Z(c[979]) );
  XNOR U32 ( .A(b[978]), .B(n31), .Z(c[978]) );
  XNOR U33 ( .A(b[977]), .B(n32), .Z(c[977]) );
  XNOR U34 ( .A(b[976]), .B(n33), .Z(c[976]) );
  XNOR U35 ( .A(b[975]), .B(n34), .Z(c[975]) );
  XNOR U36 ( .A(b[974]), .B(n35), .Z(c[974]) );
  XNOR U37 ( .A(b[973]), .B(n36), .Z(c[973]) );
  XNOR U38 ( .A(b[972]), .B(n37), .Z(c[972]) );
  XNOR U39 ( .A(b[971]), .B(n38), .Z(c[971]) );
  XNOR U40 ( .A(b[970]), .B(n39), .Z(c[970]) );
  XNOR U41 ( .A(b[96]), .B(n40), .Z(c[96]) );
  XNOR U42 ( .A(b[969]), .B(n41), .Z(c[969]) );
  XNOR U43 ( .A(b[968]), .B(n42), .Z(c[968]) );
  XNOR U44 ( .A(b[967]), .B(n43), .Z(c[967]) );
  XNOR U45 ( .A(b[966]), .B(n44), .Z(c[966]) );
  XNOR U46 ( .A(b[965]), .B(n45), .Z(c[965]) );
  XNOR U47 ( .A(b[964]), .B(n46), .Z(c[964]) );
  XNOR U48 ( .A(b[963]), .B(n47), .Z(c[963]) );
  XNOR U49 ( .A(b[962]), .B(n48), .Z(c[962]) );
  XNOR U50 ( .A(b[961]), .B(n49), .Z(c[961]) );
  XNOR U51 ( .A(b[960]), .B(n50), .Z(c[960]) );
  XNOR U52 ( .A(b[95]), .B(n51), .Z(c[95]) );
  XNOR U53 ( .A(b[959]), .B(n52), .Z(c[959]) );
  XNOR U54 ( .A(b[958]), .B(n53), .Z(c[958]) );
  XNOR U55 ( .A(b[957]), .B(n54), .Z(c[957]) );
  XNOR U56 ( .A(b[956]), .B(n55), .Z(c[956]) );
  XNOR U57 ( .A(b[955]), .B(n56), .Z(c[955]) );
  XNOR U58 ( .A(b[954]), .B(n57), .Z(c[954]) );
  XNOR U59 ( .A(b[953]), .B(n58), .Z(c[953]) );
  XNOR U60 ( .A(b[952]), .B(n59), .Z(c[952]) );
  XNOR U61 ( .A(b[951]), .B(n60), .Z(c[951]) );
  XNOR U62 ( .A(b[950]), .B(n61), .Z(c[950]) );
  XNOR U63 ( .A(b[94]), .B(n62), .Z(c[94]) );
  XNOR U64 ( .A(b[949]), .B(n63), .Z(c[949]) );
  XNOR U65 ( .A(b[948]), .B(n64), .Z(c[948]) );
  XNOR U66 ( .A(b[947]), .B(n65), .Z(c[947]) );
  XNOR U67 ( .A(b[946]), .B(n66), .Z(c[946]) );
  XNOR U68 ( .A(b[945]), .B(n67), .Z(c[945]) );
  XNOR U69 ( .A(b[944]), .B(n68), .Z(c[944]) );
  XNOR U70 ( .A(b[943]), .B(n69), .Z(c[943]) );
  XNOR U71 ( .A(b[942]), .B(n70), .Z(c[942]) );
  XNOR U72 ( .A(b[941]), .B(n71), .Z(c[941]) );
  XNOR U73 ( .A(b[940]), .B(n72), .Z(c[940]) );
  XNOR U74 ( .A(b[93]), .B(n73), .Z(c[93]) );
  XNOR U75 ( .A(b[939]), .B(n74), .Z(c[939]) );
  XNOR U76 ( .A(b[938]), .B(n75), .Z(c[938]) );
  XNOR U77 ( .A(b[937]), .B(n76), .Z(c[937]) );
  XNOR U78 ( .A(b[936]), .B(n77), .Z(c[936]) );
  XNOR U79 ( .A(b[935]), .B(n78), .Z(c[935]) );
  XNOR U80 ( .A(b[934]), .B(n79), .Z(c[934]) );
  XNOR U81 ( .A(b[933]), .B(n80), .Z(c[933]) );
  XNOR U82 ( .A(b[932]), .B(n81), .Z(c[932]) );
  XNOR U83 ( .A(b[931]), .B(n82), .Z(c[931]) );
  XNOR U84 ( .A(b[930]), .B(n83), .Z(c[930]) );
  XNOR U85 ( .A(b[92]), .B(n84), .Z(c[92]) );
  XNOR U86 ( .A(b[929]), .B(n85), .Z(c[929]) );
  XNOR U87 ( .A(b[928]), .B(n86), .Z(c[928]) );
  XNOR U88 ( .A(b[927]), .B(n87), .Z(c[927]) );
  XNOR U89 ( .A(b[926]), .B(n88), .Z(c[926]) );
  XNOR U90 ( .A(b[925]), .B(n89), .Z(c[925]) );
  XNOR U91 ( .A(b[924]), .B(n90), .Z(c[924]) );
  XNOR U92 ( .A(b[923]), .B(n91), .Z(c[923]) );
  XNOR U93 ( .A(b[922]), .B(n92), .Z(c[922]) );
  XNOR U94 ( .A(b[921]), .B(n93), .Z(c[921]) );
  XNOR U95 ( .A(b[920]), .B(n94), .Z(c[920]) );
  XNOR U96 ( .A(b[91]), .B(n95), .Z(c[91]) );
  XNOR U97 ( .A(b[919]), .B(n96), .Z(c[919]) );
  XNOR U98 ( .A(b[918]), .B(n97), .Z(c[918]) );
  XNOR U99 ( .A(b[917]), .B(n98), .Z(c[917]) );
  XNOR U100 ( .A(b[916]), .B(n99), .Z(c[916]) );
  XNOR U101 ( .A(b[915]), .B(n100), .Z(c[915]) );
  XNOR U102 ( .A(b[914]), .B(n101), .Z(c[914]) );
  XNOR U103 ( .A(b[913]), .B(n102), .Z(c[913]) );
  XNOR U104 ( .A(b[912]), .B(n103), .Z(c[912]) );
  XNOR U105 ( .A(b[911]), .B(n104), .Z(c[911]) );
  XNOR U106 ( .A(b[910]), .B(n105), .Z(c[910]) );
  XNOR U107 ( .A(b[90]), .B(n106), .Z(c[90]) );
  XNOR U108 ( .A(b[909]), .B(n107), .Z(c[909]) );
  XNOR U109 ( .A(b[908]), .B(n108), .Z(c[908]) );
  XNOR U110 ( .A(b[907]), .B(n109), .Z(c[907]) );
  XNOR U111 ( .A(b[906]), .B(n110), .Z(c[906]) );
  XNOR U112 ( .A(b[905]), .B(n111), .Z(c[905]) );
  XNOR U113 ( .A(b[904]), .B(n112), .Z(c[904]) );
  XNOR U114 ( .A(b[903]), .B(n113), .Z(c[903]) );
  XNOR U115 ( .A(b[902]), .B(n114), .Z(c[902]) );
  XNOR U116 ( .A(b[901]), .B(n115), .Z(c[901]) );
  XNOR U117 ( .A(b[900]), .B(n116), .Z(c[900]) );
  XNOR U118 ( .A(b[8]), .B(n117), .Z(c[8]) );
  XNOR U119 ( .A(b[89]), .B(n118), .Z(c[89]) );
  XNOR U120 ( .A(b[899]), .B(n119), .Z(c[899]) );
  XNOR U121 ( .A(b[898]), .B(n120), .Z(c[898]) );
  XNOR U122 ( .A(b[897]), .B(n121), .Z(c[897]) );
  XNOR U123 ( .A(b[896]), .B(n122), .Z(c[896]) );
  XNOR U124 ( .A(b[895]), .B(n123), .Z(c[895]) );
  XNOR U125 ( .A(b[894]), .B(n124), .Z(c[894]) );
  XNOR U126 ( .A(b[893]), .B(n125), .Z(c[893]) );
  XNOR U127 ( .A(b[892]), .B(n126), .Z(c[892]) );
  XNOR U128 ( .A(b[891]), .B(n127), .Z(c[891]) );
  XNOR U129 ( .A(b[890]), .B(n128), .Z(c[890]) );
  XNOR U130 ( .A(b[88]), .B(n129), .Z(c[88]) );
  XNOR U131 ( .A(b[889]), .B(n130), .Z(c[889]) );
  XNOR U132 ( .A(b[888]), .B(n131), .Z(c[888]) );
  XNOR U133 ( .A(b[887]), .B(n132), .Z(c[887]) );
  XNOR U134 ( .A(b[886]), .B(n133), .Z(c[886]) );
  XNOR U135 ( .A(b[885]), .B(n134), .Z(c[885]) );
  XNOR U136 ( .A(b[884]), .B(n135), .Z(c[884]) );
  XNOR U137 ( .A(b[883]), .B(n136), .Z(c[883]) );
  XNOR U138 ( .A(b[882]), .B(n137), .Z(c[882]) );
  XNOR U139 ( .A(b[881]), .B(n138), .Z(c[881]) );
  XNOR U140 ( .A(b[880]), .B(n139), .Z(c[880]) );
  XNOR U141 ( .A(b[87]), .B(n140), .Z(c[87]) );
  XNOR U142 ( .A(b[879]), .B(n141), .Z(c[879]) );
  XNOR U143 ( .A(b[878]), .B(n142), .Z(c[878]) );
  XNOR U144 ( .A(b[877]), .B(n143), .Z(c[877]) );
  XNOR U145 ( .A(b[876]), .B(n144), .Z(c[876]) );
  XNOR U146 ( .A(b[875]), .B(n145), .Z(c[875]) );
  XNOR U147 ( .A(b[874]), .B(n146), .Z(c[874]) );
  XNOR U148 ( .A(b[873]), .B(n147), .Z(c[873]) );
  XNOR U149 ( .A(b[872]), .B(n148), .Z(c[872]) );
  XNOR U150 ( .A(b[871]), .B(n149), .Z(c[871]) );
  XNOR U151 ( .A(b[870]), .B(n150), .Z(c[870]) );
  XNOR U152 ( .A(b[86]), .B(n151), .Z(c[86]) );
  XNOR U153 ( .A(b[869]), .B(n152), .Z(c[869]) );
  XNOR U154 ( .A(b[868]), .B(n153), .Z(c[868]) );
  XNOR U155 ( .A(b[867]), .B(n154), .Z(c[867]) );
  XNOR U156 ( .A(b[866]), .B(n155), .Z(c[866]) );
  XNOR U157 ( .A(b[865]), .B(n156), .Z(c[865]) );
  XNOR U158 ( .A(b[864]), .B(n157), .Z(c[864]) );
  XNOR U159 ( .A(b[863]), .B(n158), .Z(c[863]) );
  XNOR U160 ( .A(b[862]), .B(n159), .Z(c[862]) );
  XNOR U161 ( .A(b[861]), .B(n160), .Z(c[861]) );
  XNOR U162 ( .A(b[860]), .B(n161), .Z(c[860]) );
  XNOR U163 ( .A(b[85]), .B(n162), .Z(c[85]) );
  XNOR U164 ( .A(b[859]), .B(n163), .Z(c[859]) );
  XNOR U165 ( .A(b[858]), .B(n164), .Z(c[858]) );
  XNOR U166 ( .A(b[857]), .B(n165), .Z(c[857]) );
  XNOR U167 ( .A(b[856]), .B(n166), .Z(c[856]) );
  XNOR U168 ( .A(b[855]), .B(n167), .Z(c[855]) );
  XNOR U169 ( .A(b[854]), .B(n168), .Z(c[854]) );
  XNOR U170 ( .A(b[853]), .B(n169), .Z(c[853]) );
  XNOR U171 ( .A(b[852]), .B(n170), .Z(c[852]) );
  XNOR U172 ( .A(b[851]), .B(n171), .Z(c[851]) );
  XNOR U173 ( .A(b[850]), .B(n172), .Z(c[850]) );
  XNOR U174 ( .A(b[84]), .B(n173), .Z(c[84]) );
  XNOR U175 ( .A(b[849]), .B(n174), .Z(c[849]) );
  XNOR U176 ( .A(b[848]), .B(n175), .Z(c[848]) );
  XNOR U177 ( .A(b[847]), .B(n176), .Z(c[847]) );
  XNOR U178 ( .A(b[846]), .B(n177), .Z(c[846]) );
  XNOR U179 ( .A(b[845]), .B(n178), .Z(c[845]) );
  XNOR U180 ( .A(b[844]), .B(n179), .Z(c[844]) );
  XNOR U181 ( .A(b[843]), .B(n180), .Z(c[843]) );
  XNOR U182 ( .A(b[842]), .B(n181), .Z(c[842]) );
  XNOR U183 ( .A(b[841]), .B(n182), .Z(c[841]) );
  XNOR U184 ( .A(b[840]), .B(n183), .Z(c[840]) );
  XNOR U185 ( .A(b[83]), .B(n184), .Z(c[83]) );
  XNOR U186 ( .A(b[839]), .B(n185), .Z(c[839]) );
  XNOR U187 ( .A(b[838]), .B(n186), .Z(c[838]) );
  XNOR U188 ( .A(b[837]), .B(n187), .Z(c[837]) );
  XNOR U189 ( .A(b[836]), .B(n188), .Z(c[836]) );
  XNOR U190 ( .A(b[835]), .B(n189), .Z(c[835]) );
  XNOR U191 ( .A(b[834]), .B(n190), .Z(c[834]) );
  XNOR U192 ( .A(b[833]), .B(n191), .Z(c[833]) );
  XNOR U193 ( .A(b[832]), .B(n192), .Z(c[832]) );
  XNOR U194 ( .A(b[831]), .B(n193), .Z(c[831]) );
  XNOR U195 ( .A(b[830]), .B(n194), .Z(c[830]) );
  XNOR U196 ( .A(b[82]), .B(n195), .Z(c[82]) );
  XNOR U197 ( .A(b[829]), .B(n196), .Z(c[829]) );
  XNOR U198 ( .A(b[828]), .B(n197), .Z(c[828]) );
  XNOR U199 ( .A(b[827]), .B(n198), .Z(c[827]) );
  XNOR U200 ( .A(b[826]), .B(n199), .Z(c[826]) );
  XNOR U201 ( .A(b[825]), .B(n200), .Z(c[825]) );
  XNOR U202 ( .A(b[824]), .B(n201), .Z(c[824]) );
  XNOR U203 ( .A(b[823]), .B(n202), .Z(c[823]) );
  XNOR U204 ( .A(b[822]), .B(n203), .Z(c[822]) );
  XNOR U205 ( .A(b[821]), .B(n204), .Z(c[821]) );
  XNOR U206 ( .A(b[820]), .B(n205), .Z(c[820]) );
  XNOR U207 ( .A(b[81]), .B(n206), .Z(c[81]) );
  XNOR U208 ( .A(b[819]), .B(n207), .Z(c[819]) );
  XNOR U209 ( .A(b[818]), .B(n208), .Z(c[818]) );
  XNOR U210 ( .A(b[817]), .B(n209), .Z(c[817]) );
  XNOR U211 ( .A(b[816]), .B(n210), .Z(c[816]) );
  XNOR U212 ( .A(b[815]), .B(n211), .Z(c[815]) );
  XNOR U213 ( .A(b[814]), .B(n212), .Z(c[814]) );
  XNOR U214 ( .A(b[813]), .B(n213), .Z(c[813]) );
  XNOR U215 ( .A(b[812]), .B(n214), .Z(c[812]) );
  XNOR U216 ( .A(b[811]), .B(n215), .Z(c[811]) );
  XNOR U217 ( .A(b[810]), .B(n216), .Z(c[810]) );
  XNOR U218 ( .A(b[80]), .B(n217), .Z(c[80]) );
  XNOR U219 ( .A(b[809]), .B(n218), .Z(c[809]) );
  XNOR U220 ( .A(b[808]), .B(n219), .Z(c[808]) );
  XNOR U221 ( .A(b[807]), .B(n220), .Z(c[807]) );
  XNOR U222 ( .A(b[806]), .B(n221), .Z(c[806]) );
  XNOR U223 ( .A(b[805]), .B(n222), .Z(c[805]) );
  XNOR U224 ( .A(b[804]), .B(n223), .Z(c[804]) );
  XNOR U225 ( .A(b[803]), .B(n224), .Z(c[803]) );
  XNOR U226 ( .A(b[802]), .B(n225), .Z(c[802]) );
  XNOR U227 ( .A(b[801]), .B(n226), .Z(c[801]) );
  XNOR U228 ( .A(b[800]), .B(n227), .Z(c[800]) );
  XNOR U229 ( .A(b[7]), .B(n228), .Z(c[7]) );
  XNOR U230 ( .A(b[79]), .B(n229), .Z(c[79]) );
  XNOR U231 ( .A(b[799]), .B(n230), .Z(c[799]) );
  XNOR U232 ( .A(b[798]), .B(n231), .Z(c[798]) );
  XNOR U233 ( .A(b[797]), .B(n232), .Z(c[797]) );
  XNOR U234 ( .A(b[796]), .B(n233), .Z(c[796]) );
  XNOR U235 ( .A(b[795]), .B(n234), .Z(c[795]) );
  XNOR U236 ( .A(b[794]), .B(n235), .Z(c[794]) );
  XNOR U237 ( .A(b[793]), .B(n236), .Z(c[793]) );
  XNOR U238 ( .A(b[792]), .B(n237), .Z(c[792]) );
  XNOR U239 ( .A(b[791]), .B(n238), .Z(c[791]) );
  XNOR U240 ( .A(b[790]), .B(n239), .Z(c[790]) );
  XNOR U241 ( .A(b[78]), .B(n240), .Z(c[78]) );
  XNOR U242 ( .A(b[789]), .B(n241), .Z(c[789]) );
  XNOR U243 ( .A(b[788]), .B(n242), .Z(c[788]) );
  XNOR U244 ( .A(b[787]), .B(n243), .Z(c[787]) );
  XNOR U245 ( .A(b[786]), .B(n244), .Z(c[786]) );
  XNOR U246 ( .A(b[785]), .B(n245), .Z(c[785]) );
  XNOR U247 ( .A(b[784]), .B(n246), .Z(c[784]) );
  XNOR U248 ( .A(b[783]), .B(n247), .Z(c[783]) );
  XNOR U249 ( .A(b[782]), .B(n248), .Z(c[782]) );
  XNOR U250 ( .A(b[781]), .B(n249), .Z(c[781]) );
  XNOR U251 ( .A(b[780]), .B(n250), .Z(c[780]) );
  XNOR U252 ( .A(b[77]), .B(n251), .Z(c[77]) );
  XNOR U253 ( .A(b[779]), .B(n252), .Z(c[779]) );
  XNOR U254 ( .A(b[778]), .B(n253), .Z(c[778]) );
  XNOR U255 ( .A(b[777]), .B(n254), .Z(c[777]) );
  XNOR U256 ( .A(b[776]), .B(n255), .Z(c[776]) );
  XNOR U257 ( .A(b[775]), .B(n256), .Z(c[775]) );
  XNOR U258 ( .A(b[774]), .B(n257), .Z(c[774]) );
  XNOR U259 ( .A(b[773]), .B(n258), .Z(c[773]) );
  XNOR U260 ( .A(b[772]), .B(n259), .Z(c[772]) );
  XNOR U261 ( .A(b[771]), .B(n260), .Z(c[771]) );
  XNOR U262 ( .A(b[770]), .B(n261), .Z(c[770]) );
  XNOR U263 ( .A(b[76]), .B(n262), .Z(c[76]) );
  XNOR U264 ( .A(b[769]), .B(n263), .Z(c[769]) );
  XNOR U265 ( .A(b[768]), .B(n264), .Z(c[768]) );
  XNOR U266 ( .A(b[767]), .B(n265), .Z(c[767]) );
  XNOR U267 ( .A(b[766]), .B(n266), .Z(c[766]) );
  XNOR U268 ( .A(b[765]), .B(n267), .Z(c[765]) );
  XNOR U269 ( .A(b[764]), .B(n268), .Z(c[764]) );
  XNOR U270 ( .A(b[763]), .B(n269), .Z(c[763]) );
  XNOR U271 ( .A(b[762]), .B(n270), .Z(c[762]) );
  XNOR U272 ( .A(b[761]), .B(n271), .Z(c[761]) );
  XNOR U273 ( .A(b[760]), .B(n272), .Z(c[760]) );
  XNOR U274 ( .A(b[75]), .B(n273), .Z(c[75]) );
  XNOR U275 ( .A(b[759]), .B(n274), .Z(c[759]) );
  XNOR U276 ( .A(b[758]), .B(n275), .Z(c[758]) );
  XNOR U277 ( .A(b[757]), .B(n276), .Z(c[757]) );
  XNOR U278 ( .A(b[756]), .B(n277), .Z(c[756]) );
  XNOR U279 ( .A(b[755]), .B(n278), .Z(c[755]) );
  XNOR U280 ( .A(b[754]), .B(n279), .Z(c[754]) );
  XNOR U281 ( .A(b[753]), .B(n280), .Z(c[753]) );
  XNOR U282 ( .A(b[752]), .B(n281), .Z(c[752]) );
  XNOR U283 ( .A(b[751]), .B(n282), .Z(c[751]) );
  XNOR U284 ( .A(b[750]), .B(n283), .Z(c[750]) );
  XNOR U285 ( .A(b[74]), .B(n284), .Z(c[74]) );
  XNOR U286 ( .A(b[749]), .B(n285), .Z(c[749]) );
  XNOR U287 ( .A(b[748]), .B(n286), .Z(c[748]) );
  XNOR U288 ( .A(b[747]), .B(n287), .Z(c[747]) );
  XNOR U289 ( .A(b[746]), .B(n288), .Z(c[746]) );
  XNOR U290 ( .A(b[745]), .B(n289), .Z(c[745]) );
  XNOR U291 ( .A(b[744]), .B(n290), .Z(c[744]) );
  XNOR U292 ( .A(b[743]), .B(n291), .Z(c[743]) );
  XNOR U293 ( .A(b[742]), .B(n292), .Z(c[742]) );
  XNOR U294 ( .A(b[741]), .B(n293), .Z(c[741]) );
  XNOR U295 ( .A(b[740]), .B(n294), .Z(c[740]) );
  XNOR U296 ( .A(b[73]), .B(n295), .Z(c[73]) );
  XNOR U297 ( .A(b[739]), .B(n296), .Z(c[739]) );
  XNOR U298 ( .A(b[738]), .B(n297), .Z(c[738]) );
  XNOR U299 ( .A(b[737]), .B(n298), .Z(c[737]) );
  XNOR U300 ( .A(b[736]), .B(n299), .Z(c[736]) );
  XNOR U301 ( .A(b[735]), .B(n300), .Z(c[735]) );
  XNOR U302 ( .A(b[734]), .B(n301), .Z(c[734]) );
  XNOR U303 ( .A(b[733]), .B(n302), .Z(c[733]) );
  XNOR U304 ( .A(b[732]), .B(n303), .Z(c[732]) );
  XNOR U305 ( .A(b[731]), .B(n304), .Z(c[731]) );
  XNOR U306 ( .A(b[730]), .B(n305), .Z(c[730]) );
  XNOR U307 ( .A(b[72]), .B(n306), .Z(c[72]) );
  XNOR U308 ( .A(b[729]), .B(n307), .Z(c[729]) );
  XNOR U309 ( .A(b[728]), .B(n308), .Z(c[728]) );
  XNOR U310 ( .A(b[727]), .B(n309), .Z(c[727]) );
  XNOR U311 ( .A(b[726]), .B(n310), .Z(c[726]) );
  XNOR U312 ( .A(b[725]), .B(n311), .Z(c[725]) );
  XNOR U313 ( .A(b[724]), .B(n312), .Z(c[724]) );
  XNOR U314 ( .A(b[723]), .B(n313), .Z(c[723]) );
  XNOR U315 ( .A(b[722]), .B(n314), .Z(c[722]) );
  XNOR U316 ( .A(b[721]), .B(n315), .Z(c[721]) );
  XNOR U317 ( .A(b[720]), .B(n316), .Z(c[720]) );
  XNOR U318 ( .A(b[71]), .B(n317), .Z(c[71]) );
  XNOR U319 ( .A(b[719]), .B(n318), .Z(c[719]) );
  XNOR U320 ( .A(b[718]), .B(n319), .Z(c[718]) );
  XNOR U321 ( .A(b[717]), .B(n320), .Z(c[717]) );
  XNOR U322 ( .A(b[716]), .B(n321), .Z(c[716]) );
  XNOR U323 ( .A(b[715]), .B(n322), .Z(c[715]) );
  XNOR U324 ( .A(b[714]), .B(n323), .Z(c[714]) );
  XNOR U325 ( .A(b[713]), .B(n324), .Z(c[713]) );
  XNOR U326 ( .A(b[712]), .B(n325), .Z(c[712]) );
  XNOR U327 ( .A(b[711]), .B(n326), .Z(c[711]) );
  XNOR U328 ( .A(b[710]), .B(n327), .Z(c[710]) );
  XNOR U329 ( .A(b[70]), .B(n328), .Z(c[70]) );
  XNOR U330 ( .A(b[709]), .B(n329), .Z(c[709]) );
  XNOR U331 ( .A(b[708]), .B(n330), .Z(c[708]) );
  XNOR U332 ( .A(b[707]), .B(n331), .Z(c[707]) );
  XNOR U333 ( .A(b[706]), .B(n332), .Z(c[706]) );
  XNOR U334 ( .A(b[705]), .B(n333), .Z(c[705]) );
  XNOR U335 ( .A(b[704]), .B(n334), .Z(c[704]) );
  XNOR U336 ( .A(b[703]), .B(n335), .Z(c[703]) );
  XNOR U337 ( .A(b[702]), .B(n336), .Z(c[702]) );
  XNOR U338 ( .A(b[701]), .B(n337), .Z(c[701]) );
  XNOR U339 ( .A(b[700]), .B(n338), .Z(c[700]) );
  XNOR U340 ( .A(b[6]), .B(n339), .Z(c[6]) );
  XNOR U341 ( .A(b[69]), .B(n340), .Z(c[69]) );
  XNOR U342 ( .A(b[699]), .B(n341), .Z(c[699]) );
  XNOR U343 ( .A(b[698]), .B(n342), .Z(c[698]) );
  XNOR U344 ( .A(b[697]), .B(n343), .Z(c[697]) );
  XNOR U345 ( .A(b[696]), .B(n344), .Z(c[696]) );
  XNOR U346 ( .A(b[695]), .B(n345), .Z(c[695]) );
  XNOR U347 ( .A(b[694]), .B(n346), .Z(c[694]) );
  XNOR U348 ( .A(b[693]), .B(n347), .Z(c[693]) );
  XNOR U349 ( .A(b[692]), .B(n348), .Z(c[692]) );
  XNOR U350 ( .A(b[691]), .B(n349), .Z(c[691]) );
  XNOR U351 ( .A(b[690]), .B(n350), .Z(c[690]) );
  XNOR U352 ( .A(b[68]), .B(n351), .Z(c[68]) );
  XNOR U353 ( .A(b[689]), .B(n352), .Z(c[689]) );
  XNOR U354 ( .A(b[688]), .B(n353), .Z(c[688]) );
  XNOR U355 ( .A(b[687]), .B(n354), .Z(c[687]) );
  XNOR U356 ( .A(b[686]), .B(n355), .Z(c[686]) );
  XNOR U357 ( .A(b[685]), .B(n356), .Z(c[685]) );
  XNOR U358 ( .A(b[684]), .B(n357), .Z(c[684]) );
  XNOR U359 ( .A(b[683]), .B(n358), .Z(c[683]) );
  XNOR U360 ( .A(b[682]), .B(n359), .Z(c[682]) );
  XNOR U361 ( .A(b[681]), .B(n360), .Z(c[681]) );
  XNOR U362 ( .A(b[680]), .B(n361), .Z(c[680]) );
  XNOR U363 ( .A(b[67]), .B(n362), .Z(c[67]) );
  XNOR U364 ( .A(b[679]), .B(n363), .Z(c[679]) );
  XNOR U365 ( .A(b[678]), .B(n364), .Z(c[678]) );
  XNOR U366 ( .A(b[677]), .B(n365), .Z(c[677]) );
  XNOR U367 ( .A(b[676]), .B(n366), .Z(c[676]) );
  XNOR U368 ( .A(b[675]), .B(n367), .Z(c[675]) );
  XNOR U369 ( .A(b[674]), .B(n368), .Z(c[674]) );
  XNOR U370 ( .A(b[673]), .B(n369), .Z(c[673]) );
  XNOR U371 ( .A(b[672]), .B(n370), .Z(c[672]) );
  XNOR U372 ( .A(b[671]), .B(n371), .Z(c[671]) );
  XNOR U373 ( .A(b[670]), .B(n372), .Z(c[670]) );
  XNOR U374 ( .A(b[66]), .B(n373), .Z(c[66]) );
  XNOR U375 ( .A(b[669]), .B(n374), .Z(c[669]) );
  XNOR U376 ( .A(b[668]), .B(n375), .Z(c[668]) );
  XNOR U377 ( .A(b[667]), .B(n376), .Z(c[667]) );
  XNOR U378 ( .A(b[666]), .B(n377), .Z(c[666]) );
  XNOR U379 ( .A(b[665]), .B(n378), .Z(c[665]) );
  XNOR U380 ( .A(b[664]), .B(n379), .Z(c[664]) );
  XNOR U381 ( .A(b[663]), .B(n380), .Z(c[663]) );
  XNOR U382 ( .A(b[662]), .B(n381), .Z(c[662]) );
  XNOR U383 ( .A(b[661]), .B(n382), .Z(c[661]) );
  XNOR U384 ( .A(b[660]), .B(n383), .Z(c[660]) );
  XNOR U385 ( .A(b[65]), .B(n384), .Z(c[65]) );
  XNOR U386 ( .A(b[659]), .B(n385), .Z(c[659]) );
  XNOR U387 ( .A(b[658]), .B(n386), .Z(c[658]) );
  XNOR U388 ( .A(b[657]), .B(n387), .Z(c[657]) );
  XNOR U389 ( .A(b[656]), .B(n388), .Z(c[656]) );
  XNOR U390 ( .A(b[655]), .B(n389), .Z(c[655]) );
  XNOR U391 ( .A(b[654]), .B(n390), .Z(c[654]) );
  XNOR U392 ( .A(b[653]), .B(n391), .Z(c[653]) );
  XNOR U393 ( .A(b[652]), .B(n392), .Z(c[652]) );
  XNOR U394 ( .A(b[651]), .B(n393), .Z(c[651]) );
  XNOR U395 ( .A(b[650]), .B(n394), .Z(c[650]) );
  XNOR U396 ( .A(b[64]), .B(n395), .Z(c[64]) );
  XNOR U397 ( .A(b[649]), .B(n396), .Z(c[649]) );
  XNOR U398 ( .A(b[648]), .B(n397), .Z(c[648]) );
  XNOR U399 ( .A(b[647]), .B(n398), .Z(c[647]) );
  XNOR U400 ( .A(b[646]), .B(n399), .Z(c[646]) );
  XNOR U401 ( .A(b[645]), .B(n400), .Z(c[645]) );
  XNOR U402 ( .A(b[644]), .B(n401), .Z(c[644]) );
  XNOR U403 ( .A(b[643]), .B(n402), .Z(c[643]) );
  XNOR U404 ( .A(b[642]), .B(n403), .Z(c[642]) );
  XNOR U405 ( .A(b[641]), .B(n404), .Z(c[641]) );
  XNOR U406 ( .A(b[640]), .B(n405), .Z(c[640]) );
  XNOR U407 ( .A(b[63]), .B(n406), .Z(c[63]) );
  XNOR U408 ( .A(b[639]), .B(n407), .Z(c[639]) );
  XNOR U409 ( .A(b[638]), .B(n408), .Z(c[638]) );
  XNOR U410 ( .A(b[637]), .B(n409), .Z(c[637]) );
  XNOR U411 ( .A(b[636]), .B(n410), .Z(c[636]) );
  XNOR U412 ( .A(b[635]), .B(n411), .Z(c[635]) );
  XNOR U413 ( .A(b[634]), .B(n412), .Z(c[634]) );
  XNOR U414 ( .A(b[633]), .B(n413), .Z(c[633]) );
  XNOR U415 ( .A(b[632]), .B(n414), .Z(c[632]) );
  XNOR U416 ( .A(b[631]), .B(n415), .Z(c[631]) );
  XNOR U417 ( .A(b[630]), .B(n416), .Z(c[630]) );
  XNOR U418 ( .A(b[62]), .B(n417), .Z(c[62]) );
  XNOR U419 ( .A(b[629]), .B(n418), .Z(c[629]) );
  XNOR U420 ( .A(b[628]), .B(n419), .Z(c[628]) );
  XNOR U421 ( .A(b[627]), .B(n420), .Z(c[627]) );
  XNOR U422 ( .A(b[626]), .B(n421), .Z(c[626]) );
  XNOR U423 ( .A(b[625]), .B(n422), .Z(c[625]) );
  XNOR U424 ( .A(b[624]), .B(n423), .Z(c[624]) );
  XNOR U425 ( .A(b[623]), .B(n424), .Z(c[623]) );
  XNOR U426 ( .A(b[622]), .B(n425), .Z(c[622]) );
  XNOR U427 ( .A(b[621]), .B(n426), .Z(c[621]) );
  XNOR U428 ( .A(b[620]), .B(n427), .Z(c[620]) );
  XNOR U429 ( .A(b[61]), .B(n428), .Z(c[61]) );
  XNOR U430 ( .A(b[619]), .B(n429), .Z(c[619]) );
  XNOR U431 ( .A(b[618]), .B(n430), .Z(c[618]) );
  XNOR U432 ( .A(b[617]), .B(n431), .Z(c[617]) );
  XNOR U433 ( .A(b[616]), .B(n432), .Z(c[616]) );
  XNOR U434 ( .A(b[615]), .B(n433), .Z(c[615]) );
  XNOR U435 ( .A(b[614]), .B(n434), .Z(c[614]) );
  XNOR U436 ( .A(b[613]), .B(n435), .Z(c[613]) );
  XNOR U437 ( .A(b[612]), .B(n436), .Z(c[612]) );
  XNOR U438 ( .A(b[611]), .B(n437), .Z(c[611]) );
  XNOR U439 ( .A(b[610]), .B(n438), .Z(c[610]) );
  XNOR U440 ( .A(b[60]), .B(n439), .Z(c[60]) );
  XNOR U441 ( .A(b[609]), .B(n440), .Z(c[609]) );
  XNOR U442 ( .A(b[608]), .B(n441), .Z(c[608]) );
  XNOR U443 ( .A(b[607]), .B(n442), .Z(c[607]) );
  XNOR U444 ( .A(b[606]), .B(n443), .Z(c[606]) );
  XNOR U445 ( .A(b[605]), .B(n444), .Z(c[605]) );
  XNOR U446 ( .A(b[604]), .B(n445), .Z(c[604]) );
  XNOR U447 ( .A(b[603]), .B(n446), .Z(c[603]) );
  XNOR U448 ( .A(b[602]), .B(n447), .Z(c[602]) );
  XNOR U449 ( .A(b[601]), .B(n448), .Z(c[601]) );
  XNOR U450 ( .A(b[600]), .B(n449), .Z(c[600]) );
  XNOR U451 ( .A(b[5]), .B(n450), .Z(c[5]) );
  XNOR U452 ( .A(b[59]), .B(n451), .Z(c[59]) );
  XNOR U453 ( .A(b[599]), .B(n452), .Z(c[599]) );
  XNOR U454 ( .A(b[598]), .B(n453), .Z(c[598]) );
  XNOR U455 ( .A(b[597]), .B(n454), .Z(c[597]) );
  XNOR U456 ( .A(b[596]), .B(n455), .Z(c[596]) );
  XNOR U457 ( .A(b[595]), .B(n456), .Z(c[595]) );
  XNOR U458 ( .A(b[594]), .B(n457), .Z(c[594]) );
  XNOR U459 ( .A(b[593]), .B(n458), .Z(c[593]) );
  XNOR U460 ( .A(b[592]), .B(n459), .Z(c[592]) );
  XNOR U461 ( .A(b[591]), .B(n460), .Z(c[591]) );
  XNOR U462 ( .A(b[590]), .B(n461), .Z(c[590]) );
  XNOR U463 ( .A(b[58]), .B(n462), .Z(c[58]) );
  XNOR U464 ( .A(b[589]), .B(n463), .Z(c[589]) );
  XNOR U465 ( .A(b[588]), .B(n464), .Z(c[588]) );
  XNOR U466 ( .A(b[587]), .B(n465), .Z(c[587]) );
  XNOR U467 ( .A(b[586]), .B(n466), .Z(c[586]) );
  XNOR U468 ( .A(b[585]), .B(n467), .Z(c[585]) );
  XNOR U469 ( .A(b[584]), .B(n468), .Z(c[584]) );
  XNOR U470 ( .A(b[583]), .B(n469), .Z(c[583]) );
  XNOR U471 ( .A(b[582]), .B(n470), .Z(c[582]) );
  XNOR U472 ( .A(b[581]), .B(n471), .Z(c[581]) );
  XNOR U473 ( .A(b[580]), .B(n472), .Z(c[580]) );
  XNOR U474 ( .A(b[57]), .B(n473), .Z(c[57]) );
  XNOR U475 ( .A(b[579]), .B(n474), .Z(c[579]) );
  XNOR U476 ( .A(b[578]), .B(n475), .Z(c[578]) );
  XNOR U477 ( .A(b[577]), .B(n476), .Z(c[577]) );
  XNOR U478 ( .A(b[576]), .B(n477), .Z(c[576]) );
  XNOR U479 ( .A(b[575]), .B(n478), .Z(c[575]) );
  XNOR U480 ( .A(b[574]), .B(n479), .Z(c[574]) );
  XNOR U481 ( .A(b[573]), .B(n480), .Z(c[573]) );
  XNOR U482 ( .A(b[572]), .B(n481), .Z(c[572]) );
  XNOR U483 ( .A(b[571]), .B(n482), .Z(c[571]) );
  XNOR U484 ( .A(b[570]), .B(n483), .Z(c[570]) );
  XNOR U485 ( .A(b[56]), .B(n484), .Z(c[56]) );
  XNOR U486 ( .A(b[569]), .B(n485), .Z(c[569]) );
  XNOR U487 ( .A(b[568]), .B(n486), .Z(c[568]) );
  XNOR U488 ( .A(b[567]), .B(n487), .Z(c[567]) );
  XNOR U489 ( .A(b[566]), .B(n488), .Z(c[566]) );
  XNOR U490 ( .A(b[565]), .B(n489), .Z(c[565]) );
  XNOR U491 ( .A(b[564]), .B(n490), .Z(c[564]) );
  XNOR U492 ( .A(b[563]), .B(n491), .Z(c[563]) );
  XNOR U493 ( .A(b[562]), .B(n492), .Z(c[562]) );
  XNOR U494 ( .A(b[561]), .B(n493), .Z(c[561]) );
  XNOR U495 ( .A(b[560]), .B(n494), .Z(c[560]) );
  XNOR U496 ( .A(b[55]), .B(n495), .Z(c[55]) );
  XNOR U497 ( .A(b[559]), .B(n496), .Z(c[559]) );
  XNOR U498 ( .A(b[558]), .B(n497), .Z(c[558]) );
  XNOR U499 ( .A(b[557]), .B(n498), .Z(c[557]) );
  XNOR U500 ( .A(b[556]), .B(n499), .Z(c[556]) );
  XNOR U501 ( .A(b[555]), .B(n500), .Z(c[555]) );
  XNOR U502 ( .A(b[554]), .B(n501), .Z(c[554]) );
  XNOR U503 ( .A(b[553]), .B(n502), .Z(c[553]) );
  XNOR U504 ( .A(b[552]), .B(n503), .Z(c[552]) );
  XNOR U505 ( .A(b[551]), .B(n504), .Z(c[551]) );
  XNOR U506 ( .A(b[550]), .B(n505), .Z(c[550]) );
  XNOR U507 ( .A(b[54]), .B(n506), .Z(c[54]) );
  XNOR U508 ( .A(b[549]), .B(n507), .Z(c[549]) );
  XNOR U509 ( .A(b[548]), .B(n508), .Z(c[548]) );
  XNOR U510 ( .A(b[547]), .B(n509), .Z(c[547]) );
  XNOR U511 ( .A(b[546]), .B(n510), .Z(c[546]) );
  XNOR U512 ( .A(b[545]), .B(n511), .Z(c[545]) );
  XNOR U513 ( .A(b[544]), .B(n512), .Z(c[544]) );
  XNOR U514 ( .A(b[543]), .B(n513), .Z(c[543]) );
  XNOR U515 ( .A(b[542]), .B(n514), .Z(c[542]) );
  XNOR U516 ( .A(b[541]), .B(n515), .Z(c[541]) );
  XNOR U517 ( .A(b[540]), .B(n516), .Z(c[540]) );
  XNOR U518 ( .A(b[53]), .B(n517), .Z(c[53]) );
  XNOR U519 ( .A(b[539]), .B(n518), .Z(c[539]) );
  XNOR U520 ( .A(b[538]), .B(n519), .Z(c[538]) );
  XNOR U521 ( .A(b[537]), .B(n520), .Z(c[537]) );
  XNOR U522 ( .A(b[536]), .B(n521), .Z(c[536]) );
  XNOR U523 ( .A(b[535]), .B(n522), .Z(c[535]) );
  XNOR U524 ( .A(b[534]), .B(n523), .Z(c[534]) );
  XNOR U525 ( .A(b[533]), .B(n524), .Z(c[533]) );
  XNOR U526 ( .A(b[532]), .B(n525), .Z(c[532]) );
  XNOR U527 ( .A(b[531]), .B(n526), .Z(c[531]) );
  XNOR U528 ( .A(b[530]), .B(n527), .Z(c[530]) );
  XNOR U529 ( .A(b[52]), .B(n528), .Z(c[52]) );
  XNOR U530 ( .A(b[529]), .B(n529), .Z(c[529]) );
  XNOR U531 ( .A(b[528]), .B(n530), .Z(c[528]) );
  XNOR U532 ( .A(b[527]), .B(n531), .Z(c[527]) );
  XNOR U533 ( .A(b[526]), .B(n532), .Z(c[526]) );
  XNOR U534 ( .A(b[525]), .B(n533), .Z(c[525]) );
  XNOR U535 ( .A(b[524]), .B(n534), .Z(c[524]) );
  XNOR U536 ( .A(b[523]), .B(n535), .Z(c[523]) );
  XNOR U537 ( .A(b[522]), .B(n536), .Z(c[522]) );
  XNOR U538 ( .A(b[521]), .B(n537), .Z(c[521]) );
  XNOR U539 ( .A(b[520]), .B(n538), .Z(c[520]) );
  XNOR U540 ( .A(b[51]), .B(n539), .Z(c[51]) );
  XNOR U541 ( .A(b[519]), .B(n540), .Z(c[519]) );
  XNOR U542 ( .A(b[518]), .B(n541), .Z(c[518]) );
  XNOR U543 ( .A(b[517]), .B(n542), .Z(c[517]) );
  XNOR U544 ( .A(b[516]), .B(n543), .Z(c[516]) );
  XNOR U545 ( .A(b[515]), .B(n544), .Z(c[515]) );
  XNOR U546 ( .A(b[514]), .B(n545), .Z(c[514]) );
  XNOR U547 ( .A(b[513]), .B(n546), .Z(c[513]) );
  XNOR U548 ( .A(b[512]), .B(n547), .Z(c[512]) );
  XNOR U549 ( .A(b[511]), .B(n548), .Z(c[511]) );
  XNOR U550 ( .A(b[510]), .B(n549), .Z(c[510]) );
  XNOR U551 ( .A(b[50]), .B(n550), .Z(c[50]) );
  XNOR U552 ( .A(b[509]), .B(n551), .Z(c[509]) );
  XNOR U553 ( .A(b[508]), .B(n552), .Z(c[508]) );
  XNOR U554 ( .A(b[507]), .B(n553), .Z(c[507]) );
  XNOR U555 ( .A(b[506]), .B(n554), .Z(c[506]) );
  XNOR U556 ( .A(b[505]), .B(n555), .Z(c[505]) );
  XNOR U557 ( .A(b[504]), .B(n556), .Z(c[504]) );
  XNOR U558 ( .A(b[503]), .B(n557), .Z(c[503]) );
  XNOR U559 ( .A(b[502]), .B(n558), .Z(c[502]) );
  XNOR U560 ( .A(b[501]), .B(n559), .Z(c[501]) );
  XNOR U561 ( .A(b[500]), .B(n560), .Z(c[500]) );
  XNOR U562 ( .A(b[4]), .B(n561), .Z(c[4]) );
  XNOR U563 ( .A(b[49]), .B(n562), .Z(c[49]) );
  XNOR U564 ( .A(b[499]), .B(n563), .Z(c[499]) );
  XNOR U565 ( .A(b[498]), .B(n564), .Z(c[498]) );
  XNOR U566 ( .A(b[497]), .B(n565), .Z(c[497]) );
  XNOR U567 ( .A(b[496]), .B(n566), .Z(c[496]) );
  XNOR U568 ( .A(b[495]), .B(n567), .Z(c[495]) );
  XNOR U569 ( .A(b[494]), .B(n568), .Z(c[494]) );
  XNOR U570 ( .A(b[493]), .B(n569), .Z(c[493]) );
  XNOR U571 ( .A(b[492]), .B(n570), .Z(c[492]) );
  XNOR U572 ( .A(b[491]), .B(n571), .Z(c[491]) );
  XNOR U573 ( .A(b[490]), .B(n572), .Z(c[490]) );
  XNOR U574 ( .A(b[48]), .B(n573), .Z(c[48]) );
  XNOR U575 ( .A(b[489]), .B(n574), .Z(c[489]) );
  XNOR U576 ( .A(b[488]), .B(n575), .Z(c[488]) );
  XNOR U577 ( .A(b[487]), .B(n576), .Z(c[487]) );
  XNOR U578 ( .A(b[486]), .B(n577), .Z(c[486]) );
  XNOR U579 ( .A(b[485]), .B(n578), .Z(c[485]) );
  XNOR U580 ( .A(b[484]), .B(n579), .Z(c[484]) );
  XNOR U581 ( .A(b[483]), .B(n580), .Z(c[483]) );
  XNOR U582 ( .A(b[482]), .B(n581), .Z(c[482]) );
  XNOR U583 ( .A(b[481]), .B(n582), .Z(c[481]) );
  XNOR U584 ( .A(b[480]), .B(n583), .Z(c[480]) );
  XNOR U585 ( .A(b[47]), .B(n584), .Z(c[47]) );
  XNOR U586 ( .A(b[479]), .B(n585), .Z(c[479]) );
  XNOR U587 ( .A(b[478]), .B(n586), .Z(c[478]) );
  XNOR U588 ( .A(b[477]), .B(n587), .Z(c[477]) );
  XNOR U589 ( .A(b[476]), .B(n588), .Z(c[476]) );
  XNOR U590 ( .A(b[475]), .B(n589), .Z(c[475]) );
  XNOR U591 ( .A(b[474]), .B(n590), .Z(c[474]) );
  XNOR U592 ( .A(b[473]), .B(n591), .Z(c[473]) );
  XNOR U593 ( .A(b[472]), .B(n592), .Z(c[472]) );
  XNOR U594 ( .A(b[471]), .B(n593), .Z(c[471]) );
  XNOR U595 ( .A(b[470]), .B(n594), .Z(c[470]) );
  XNOR U596 ( .A(b[46]), .B(n595), .Z(c[46]) );
  XNOR U597 ( .A(b[469]), .B(n596), .Z(c[469]) );
  XNOR U598 ( .A(b[468]), .B(n597), .Z(c[468]) );
  XNOR U599 ( .A(b[467]), .B(n598), .Z(c[467]) );
  XNOR U600 ( .A(b[466]), .B(n599), .Z(c[466]) );
  XNOR U601 ( .A(b[465]), .B(n600), .Z(c[465]) );
  XNOR U602 ( .A(b[464]), .B(n601), .Z(c[464]) );
  XNOR U603 ( .A(b[463]), .B(n602), .Z(c[463]) );
  XNOR U604 ( .A(b[462]), .B(n603), .Z(c[462]) );
  XNOR U605 ( .A(b[461]), .B(n604), .Z(c[461]) );
  XNOR U606 ( .A(b[460]), .B(n605), .Z(c[460]) );
  XNOR U607 ( .A(b[45]), .B(n606), .Z(c[45]) );
  XNOR U608 ( .A(b[459]), .B(n607), .Z(c[459]) );
  XNOR U609 ( .A(b[458]), .B(n608), .Z(c[458]) );
  XNOR U610 ( .A(b[457]), .B(n609), .Z(c[457]) );
  XNOR U611 ( .A(b[456]), .B(n610), .Z(c[456]) );
  XNOR U612 ( .A(b[455]), .B(n611), .Z(c[455]) );
  XNOR U613 ( .A(b[454]), .B(n612), .Z(c[454]) );
  XNOR U614 ( .A(b[453]), .B(n613), .Z(c[453]) );
  XNOR U615 ( .A(b[452]), .B(n614), .Z(c[452]) );
  XNOR U616 ( .A(b[451]), .B(n615), .Z(c[451]) );
  XNOR U617 ( .A(b[450]), .B(n616), .Z(c[450]) );
  XNOR U618 ( .A(b[44]), .B(n617), .Z(c[44]) );
  XNOR U619 ( .A(b[449]), .B(n618), .Z(c[449]) );
  XNOR U620 ( .A(b[448]), .B(n619), .Z(c[448]) );
  XNOR U621 ( .A(b[447]), .B(n620), .Z(c[447]) );
  XNOR U622 ( .A(b[446]), .B(n621), .Z(c[446]) );
  XNOR U623 ( .A(b[445]), .B(n622), .Z(c[445]) );
  XNOR U624 ( .A(b[444]), .B(n623), .Z(c[444]) );
  XNOR U625 ( .A(b[443]), .B(n624), .Z(c[443]) );
  XNOR U626 ( .A(b[442]), .B(n625), .Z(c[442]) );
  XNOR U627 ( .A(b[441]), .B(n626), .Z(c[441]) );
  XNOR U628 ( .A(b[440]), .B(n627), .Z(c[440]) );
  XNOR U629 ( .A(b[43]), .B(n628), .Z(c[43]) );
  XNOR U630 ( .A(b[439]), .B(n629), .Z(c[439]) );
  XNOR U631 ( .A(b[438]), .B(n630), .Z(c[438]) );
  XNOR U632 ( .A(b[437]), .B(n631), .Z(c[437]) );
  XNOR U633 ( .A(b[436]), .B(n632), .Z(c[436]) );
  XNOR U634 ( .A(b[435]), .B(n633), .Z(c[435]) );
  XNOR U635 ( .A(b[434]), .B(n634), .Z(c[434]) );
  XNOR U636 ( .A(b[433]), .B(n635), .Z(c[433]) );
  XNOR U637 ( .A(b[432]), .B(n636), .Z(c[432]) );
  XNOR U638 ( .A(b[431]), .B(n637), .Z(c[431]) );
  XNOR U639 ( .A(b[430]), .B(n638), .Z(c[430]) );
  XNOR U640 ( .A(b[42]), .B(n639), .Z(c[42]) );
  XNOR U641 ( .A(b[429]), .B(n640), .Z(c[429]) );
  XNOR U642 ( .A(b[428]), .B(n641), .Z(c[428]) );
  XNOR U643 ( .A(b[427]), .B(n642), .Z(c[427]) );
  XNOR U644 ( .A(b[426]), .B(n643), .Z(c[426]) );
  XNOR U645 ( .A(b[425]), .B(n644), .Z(c[425]) );
  XNOR U646 ( .A(b[424]), .B(n645), .Z(c[424]) );
  XNOR U647 ( .A(b[423]), .B(n646), .Z(c[423]) );
  XNOR U648 ( .A(b[422]), .B(n647), .Z(c[422]) );
  XNOR U649 ( .A(b[421]), .B(n648), .Z(c[421]) );
  XNOR U650 ( .A(b[420]), .B(n649), .Z(c[420]) );
  XNOR U651 ( .A(b[41]), .B(n650), .Z(c[41]) );
  XNOR U652 ( .A(b[419]), .B(n651), .Z(c[419]) );
  XNOR U653 ( .A(b[418]), .B(n652), .Z(c[418]) );
  XNOR U654 ( .A(b[417]), .B(n653), .Z(c[417]) );
  XNOR U655 ( .A(b[416]), .B(n654), .Z(c[416]) );
  XNOR U656 ( .A(b[415]), .B(n655), .Z(c[415]) );
  XNOR U657 ( .A(b[414]), .B(n656), .Z(c[414]) );
  XNOR U658 ( .A(b[413]), .B(n657), .Z(c[413]) );
  XNOR U659 ( .A(b[412]), .B(n658), .Z(c[412]) );
  XNOR U660 ( .A(b[411]), .B(n659), .Z(c[411]) );
  XNOR U661 ( .A(b[410]), .B(n660), .Z(c[410]) );
  XNOR U662 ( .A(b[40]), .B(n661), .Z(c[40]) );
  XNOR U663 ( .A(b[409]), .B(n662), .Z(c[409]) );
  XNOR U664 ( .A(b[408]), .B(n663), .Z(c[408]) );
  XNOR U665 ( .A(b[407]), .B(n664), .Z(c[407]) );
  XNOR U666 ( .A(b[406]), .B(n665), .Z(c[406]) );
  XNOR U667 ( .A(b[405]), .B(n666), .Z(c[405]) );
  XNOR U668 ( .A(b[404]), .B(n667), .Z(c[404]) );
  XNOR U669 ( .A(b[403]), .B(n668), .Z(c[403]) );
  XNOR U670 ( .A(b[402]), .B(n669), .Z(c[402]) );
  XNOR U671 ( .A(b[401]), .B(n670), .Z(c[401]) );
  XNOR U672 ( .A(b[400]), .B(n671), .Z(c[400]) );
  XNOR U673 ( .A(b[3]), .B(n672), .Z(c[3]) );
  XNOR U674 ( .A(b[39]), .B(n673), .Z(c[39]) );
  XNOR U675 ( .A(b[399]), .B(n674), .Z(c[399]) );
  XNOR U676 ( .A(b[398]), .B(n675), .Z(c[398]) );
  XNOR U677 ( .A(b[397]), .B(n676), .Z(c[397]) );
  XNOR U678 ( .A(b[396]), .B(n677), .Z(c[396]) );
  XNOR U679 ( .A(b[395]), .B(n678), .Z(c[395]) );
  XNOR U680 ( .A(b[394]), .B(n679), .Z(c[394]) );
  XNOR U681 ( .A(b[393]), .B(n680), .Z(c[393]) );
  XNOR U682 ( .A(b[392]), .B(n681), .Z(c[392]) );
  XNOR U683 ( .A(b[391]), .B(n682), .Z(c[391]) );
  XNOR U684 ( .A(b[390]), .B(n683), .Z(c[390]) );
  XNOR U685 ( .A(b[38]), .B(n684), .Z(c[38]) );
  XNOR U686 ( .A(b[389]), .B(n685), .Z(c[389]) );
  XNOR U687 ( .A(b[388]), .B(n686), .Z(c[388]) );
  XNOR U688 ( .A(b[387]), .B(n687), .Z(c[387]) );
  XNOR U689 ( .A(b[386]), .B(n688), .Z(c[386]) );
  XNOR U690 ( .A(b[385]), .B(n689), .Z(c[385]) );
  XNOR U691 ( .A(b[384]), .B(n690), .Z(c[384]) );
  XNOR U692 ( .A(b[383]), .B(n691), .Z(c[383]) );
  XNOR U693 ( .A(b[382]), .B(n692), .Z(c[382]) );
  XNOR U694 ( .A(b[381]), .B(n693), .Z(c[381]) );
  XNOR U695 ( .A(b[380]), .B(n694), .Z(c[380]) );
  XNOR U696 ( .A(b[37]), .B(n695), .Z(c[37]) );
  XNOR U697 ( .A(b[379]), .B(n696), .Z(c[379]) );
  XNOR U698 ( .A(b[378]), .B(n697), .Z(c[378]) );
  XNOR U699 ( .A(b[377]), .B(n698), .Z(c[377]) );
  XNOR U700 ( .A(b[376]), .B(n699), .Z(c[376]) );
  XNOR U701 ( .A(b[375]), .B(n700), .Z(c[375]) );
  XNOR U702 ( .A(b[374]), .B(n701), .Z(c[374]) );
  XNOR U703 ( .A(b[373]), .B(n702), .Z(c[373]) );
  XNOR U704 ( .A(b[372]), .B(n703), .Z(c[372]) );
  XNOR U705 ( .A(b[371]), .B(n704), .Z(c[371]) );
  XNOR U706 ( .A(b[370]), .B(n705), .Z(c[370]) );
  XNOR U707 ( .A(b[36]), .B(n706), .Z(c[36]) );
  XNOR U708 ( .A(b[369]), .B(n707), .Z(c[369]) );
  XNOR U709 ( .A(b[368]), .B(n708), .Z(c[368]) );
  XNOR U710 ( .A(b[367]), .B(n709), .Z(c[367]) );
  XNOR U711 ( .A(b[366]), .B(n710), .Z(c[366]) );
  XNOR U712 ( .A(b[365]), .B(n711), .Z(c[365]) );
  XNOR U713 ( .A(b[364]), .B(n712), .Z(c[364]) );
  XNOR U714 ( .A(b[363]), .B(n713), .Z(c[363]) );
  XNOR U715 ( .A(b[362]), .B(n714), .Z(c[362]) );
  XNOR U716 ( .A(b[361]), .B(n715), .Z(c[361]) );
  XNOR U717 ( .A(b[360]), .B(n716), .Z(c[360]) );
  XNOR U718 ( .A(b[35]), .B(n717), .Z(c[35]) );
  XNOR U719 ( .A(b[359]), .B(n718), .Z(c[359]) );
  XNOR U720 ( .A(b[358]), .B(n719), .Z(c[358]) );
  XNOR U721 ( .A(b[357]), .B(n720), .Z(c[357]) );
  XNOR U722 ( .A(b[356]), .B(n721), .Z(c[356]) );
  XNOR U723 ( .A(b[355]), .B(n722), .Z(c[355]) );
  XNOR U724 ( .A(b[354]), .B(n723), .Z(c[354]) );
  XNOR U725 ( .A(b[353]), .B(n724), .Z(c[353]) );
  XNOR U726 ( .A(b[352]), .B(n725), .Z(c[352]) );
  XNOR U727 ( .A(b[351]), .B(n726), .Z(c[351]) );
  XNOR U728 ( .A(b[350]), .B(n727), .Z(c[350]) );
  XNOR U729 ( .A(b[34]), .B(n728), .Z(c[34]) );
  XNOR U730 ( .A(b[349]), .B(n729), .Z(c[349]) );
  XNOR U731 ( .A(b[348]), .B(n730), .Z(c[348]) );
  XNOR U732 ( .A(b[347]), .B(n731), .Z(c[347]) );
  XNOR U733 ( .A(b[346]), .B(n732), .Z(c[346]) );
  XNOR U734 ( .A(b[345]), .B(n733), .Z(c[345]) );
  XNOR U735 ( .A(b[344]), .B(n734), .Z(c[344]) );
  XNOR U736 ( .A(b[343]), .B(n735), .Z(c[343]) );
  XNOR U737 ( .A(b[342]), .B(n736), .Z(c[342]) );
  XNOR U738 ( .A(b[341]), .B(n737), .Z(c[341]) );
  XNOR U739 ( .A(b[340]), .B(n738), .Z(c[340]) );
  XNOR U740 ( .A(b[33]), .B(n739), .Z(c[33]) );
  XNOR U741 ( .A(b[339]), .B(n740), .Z(c[339]) );
  XNOR U742 ( .A(b[338]), .B(n741), .Z(c[338]) );
  XNOR U743 ( .A(b[337]), .B(n742), .Z(c[337]) );
  XNOR U744 ( .A(b[336]), .B(n743), .Z(c[336]) );
  XNOR U745 ( .A(b[335]), .B(n744), .Z(c[335]) );
  XNOR U746 ( .A(b[334]), .B(n745), .Z(c[334]) );
  XNOR U747 ( .A(b[333]), .B(n746), .Z(c[333]) );
  XNOR U748 ( .A(b[332]), .B(n747), .Z(c[332]) );
  XNOR U749 ( .A(b[331]), .B(n748), .Z(c[331]) );
  XNOR U750 ( .A(b[330]), .B(n749), .Z(c[330]) );
  XNOR U751 ( .A(b[32]), .B(n750), .Z(c[32]) );
  XNOR U752 ( .A(b[329]), .B(n751), .Z(c[329]) );
  XNOR U753 ( .A(b[328]), .B(n752), .Z(c[328]) );
  XNOR U754 ( .A(b[327]), .B(n753), .Z(c[327]) );
  XNOR U755 ( .A(b[326]), .B(n754), .Z(c[326]) );
  XNOR U756 ( .A(b[325]), .B(n755), .Z(c[325]) );
  XNOR U757 ( .A(b[324]), .B(n756), .Z(c[324]) );
  XNOR U758 ( .A(b[323]), .B(n757), .Z(c[323]) );
  XNOR U759 ( .A(b[322]), .B(n758), .Z(c[322]) );
  XNOR U760 ( .A(b[321]), .B(n759), .Z(c[321]) );
  XNOR U761 ( .A(b[320]), .B(n760), .Z(c[320]) );
  XNOR U762 ( .A(b[31]), .B(n761), .Z(c[31]) );
  XNOR U763 ( .A(b[319]), .B(n762), .Z(c[319]) );
  XNOR U764 ( .A(b[318]), .B(n763), .Z(c[318]) );
  XNOR U765 ( .A(b[317]), .B(n764), .Z(c[317]) );
  XNOR U766 ( .A(b[316]), .B(n765), .Z(c[316]) );
  XNOR U767 ( .A(b[315]), .B(n766), .Z(c[315]) );
  XNOR U768 ( .A(b[314]), .B(n767), .Z(c[314]) );
  XNOR U769 ( .A(b[313]), .B(n768), .Z(c[313]) );
  XNOR U770 ( .A(b[312]), .B(n769), .Z(c[312]) );
  XNOR U771 ( .A(b[311]), .B(n770), .Z(c[311]) );
  XNOR U772 ( .A(b[310]), .B(n771), .Z(c[310]) );
  XNOR U773 ( .A(b[30]), .B(n772), .Z(c[30]) );
  XNOR U774 ( .A(b[309]), .B(n773), .Z(c[309]) );
  XNOR U775 ( .A(b[308]), .B(n774), .Z(c[308]) );
  XNOR U776 ( .A(b[307]), .B(n775), .Z(c[307]) );
  XNOR U777 ( .A(b[306]), .B(n776), .Z(c[306]) );
  XNOR U778 ( .A(b[305]), .B(n777), .Z(c[305]) );
  XNOR U779 ( .A(b[304]), .B(n778), .Z(c[304]) );
  XNOR U780 ( .A(b[303]), .B(n779), .Z(c[303]) );
  XNOR U781 ( .A(b[302]), .B(n780), .Z(c[302]) );
  XNOR U782 ( .A(b[301]), .B(n781), .Z(c[301]) );
  XNOR U783 ( .A(b[300]), .B(n782), .Z(c[300]) );
  XNOR U784 ( .A(b[2]), .B(n783), .Z(c[2]) );
  XNOR U785 ( .A(b[29]), .B(n784), .Z(c[29]) );
  XNOR U786 ( .A(b[299]), .B(n785), .Z(c[299]) );
  XNOR U787 ( .A(b[298]), .B(n786), .Z(c[298]) );
  XNOR U788 ( .A(b[297]), .B(n787), .Z(c[297]) );
  XNOR U789 ( .A(b[296]), .B(n788), .Z(c[296]) );
  XNOR U790 ( .A(b[295]), .B(n789), .Z(c[295]) );
  XNOR U791 ( .A(b[294]), .B(n790), .Z(c[294]) );
  XNOR U792 ( .A(b[293]), .B(n791), .Z(c[293]) );
  XNOR U793 ( .A(b[292]), .B(n792), .Z(c[292]) );
  XNOR U794 ( .A(b[291]), .B(n793), .Z(c[291]) );
  XNOR U795 ( .A(b[290]), .B(n794), .Z(c[290]) );
  XNOR U796 ( .A(b[28]), .B(n795), .Z(c[28]) );
  XNOR U797 ( .A(b[289]), .B(n796), .Z(c[289]) );
  XNOR U798 ( .A(b[288]), .B(n797), .Z(c[288]) );
  XNOR U799 ( .A(b[287]), .B(n798), .Z(c[287]) );
  XNOR U800 ( .A(b[286]), .B(n799), .Z(c[286]) );
  XNOR U801 ( .A(b[285]), .B(n800), .Z(c[285]) );
  XNOR U802 ( .A(b[284]), .B(n801), .Z(c[284]) );
  XNOR U803 ( .A(b[283]), .B(n802), .Z(c[283]) );
  XNOR U804 ( .A(b[282]), .B(n803), .Z(c[282]) );
  XNOR U805 ( .A(b[281]), .B(n804), .Z(c[281]) );
  XNOR U806 ( .A(b[280]), .B(n805), .Z(c[280]) );
  XNOR U807 ( .A(b[27]), .B(n806), .Z(c[27]) );
  XNOR U808 ( .A(b[279]), .B(n807), .Z(c[279]) );
  XNOR U809 ( .A(b[278]), .B(n808), .Z(c[278]) );
  XNOR U810 ( .A(b[277]), .B(n809), .Z(c[277]) );
  XNOR U811 ( .A(b[276]), .B(n810), .Z(c[276]) );
  XNOR U812 ( .A(b[275]), .B(n811), .Z(c[275]) );
  XNOR U813 ( .A(b[274]), .B(n812), .Z(c[274]) );
  XNOR U814 ( .A(b[273]), .B(n813), .Z(c[273]) );
  XNOR U815 ( .A(b[272]), .B(n814), .Z(c[272]) );
  XNOR U816 ( .A(b[271]), .B(n815), .Z(c[271]) );
  XNOR U817 ( .A(b[270]), .B(n816), .Z(c[270]) );
  XNOR U818 ( .A(b[26]), .B(n817), .Z(c[26]) );
  XNOR U819 ( .A(b[269]), .B(n818), .Z(c[269]) );
  XNOR U820 ( .A(b[268]), .B(n819), .Z(c[268]) );
  XNOR U821 ( .A(b[267]), .B(n820), .Z(c[267]) );
  XNOR U822 ( .A(b[266]), .B(n821), .Z(c[266]) );
  XNOR U823 ( .A(b[265]), .B(n822), .Z(c[265]) );
  XNOR U824 ( .A(b[264]), .B(n823), .Z(c[264]) );
  XNOR U825 ( .A(b[263]), .B(n824), .Z(c[263]) );
  XNOR U826 ( .A(b[262]), .B(n825), .Z(c[262]) );
  XNOR U827 ( .A(b[261]), .B(n826), .Z(c[261]) );
  XNOR U828 ( .A(b[260]), .B(n827), .Z(c[260]) );
  XNOR U829 ( .A(b[25]), .B(n828), .Z(c[25]) );
  XNOR U830 ( .A(b[259]), .B(n829), .Z(c[259]) );
  XNOR U831 ( .A(b[258]), .B(n830), .Z(c[258]) );
  XNOR U832 ( .A(b[257]), .B(n831), .Z(c[257]) );
  XNOR U833 ( .A(b[256]), .B(n832), .Z(c[256]) );
  XNOR U834 ( .A(b[255]), .B(n833), .Z(c[255]) );
  XNOR U835 ( .A(b[254]), .B(n834), .Z(c[254]) );
  XNOR U836 ( .A(b[253]), .B(n835), .Z(c[253]) );
  XNOR U837 ( .A(b[252]), .B(n836), .Z(c[252]) );
  XNOR U838 ( .A(b[251]), .B(n837), .Z(c[251]) );
  XNOR U839 ( .A(b[250]), .B(n838), .Z(c[250]) );
  XNOR U840 ( .A(b[24]), .B(n839), .Z(c[24]) );
  XNOR U841 ( .A(b[249]), .B(n840), .Z(c[249]) );
  XNOR U842 ( .A(b[248]), .B(n841), .Z(c[248]) );
  XNOR U843 ( .A(b[247]), .B(n842), .Z(c[247]) );
  XNOR U844 ( .A(b[246]), .B(n843), .Z(c[246]) );
  XNOR U845 ( .A(b[245]), .B(n844), .Z(c[245]) );
  XNOR U846 ( .A(b[244]), .B(n845), .Z(c[244]) );
  XNOR U847 ( .A(b[243]), .B(n846), .Z(c[243]) );
  XNOR U848 ( .A(b[242]), .B(n847), .Z(c[242]) );
  XNOR U849 ( .A(b[241]), .B(n848), .Z(c[241]) );
  XNOR U850 ( .A(b[240]), .B(n849), .Z(c[240]) );
  XNOR U851 ( .A(b[23]), .B(n850), .Z(c[23]) );
  XNOR U852 ( .A(b[239]), .B(n851), .Z(c[239]) );
  XNOR U853 ( .A(b[238]), .B(n852), .Z(c[238]) );
  XNOR U854 ( .A(b[237]), .B(n853), .Z(c[237]) );
  XNOR U855 ( .A(b[236]), .B(n854), .Z(c[236]) );
  XNOR U856 ( .A(b[235]), .B(n855), .Z(c[235]) );
  XNOR U857 ( .A(b[234]), .B(n856), .Z(c[234]) );
  XNOR U858 ( .A(b[233]), .B(n857), .Z(c[233]) );
  XNOR U859 ( .A(b[232]), .B(n858), .Z(c[232]) );
  XNOR U860 ( .A(b[231]), .B(n859), .Z(c[231]) );
  XNOR U861 ( .A(b[230]), .B(n860), .Z(c[230]) );
  XNOR U862 ( .A(b[22]), .B(n861), .Z(c[22]) );
  XNOR U863 ( .A(b[229]), .B(n862), .Z(c[229]) );
  XNOR U864 ( .A(b[228]), .B(n863), .Z(c[228]) );
  XNOR U865 ( .A(b[227]), .B(n864), .Z(c[227]) );
  XNOR U866 ( .A(b[226]), .B(n865), .Z(c[226]) );
  XNOR U867 ( .A(b[225]), .B(n866), .Z(c[225]) );
  XNOR U868 ( .A(b[224]), .B(n867), .Z(c[224]) );
  XNOR U869 ( .A(b[223]), .B(n868), .Z(c[223]) );
  XNOR U870 ( .A(b[222]), .B(n869), .Z(c[222]) );
  XNOR U871 ( .A(b[221]), .B(n870), .Z(c[221]) );
  XNOR U872 ( .A(b[220]), .B(n871), .Z(c[220]) );
  XNOR U873 ( .A(b[21]), .B(n872), .Z(c[21]) );
  XNOR U874 ( .A(b[219]), .B(n873), .Z(c[219]) );
  XNOR U875 ( .A(b[218]), .B(n874), .Z(c[218]) );
  XNOR U876 ( .A(b[217]), .B(n875), .Z(c[217]) );
  XNOR U877 ( .A(b[216]), .B(n876), .Z(c[216]) );
  XNOR U878 ( .A(b[215]), .B(n877), .Z(c[215]) );
  XNOR U879 ( .A(b[214]), .B(n878), .Z(c[214]) );
  XNOR U880 ( .A(b[213]), .B(n879), .Z(c[213]) );
  XNOR U881 ( .A(b[212]), .B(n880), .Z(c[212]) );
  XNOR U882 ( .A(b[211]), .B(n881), .Z(c[211]) );
  XNOR U883 ( .A(b[210]), .B(n882), .Z(c[210]) );
  XNOR U884 ( .A(b[20]), .B(n883), .Z(c[20]) );
  XNOR U885 ( .A(b[209]), .B(n884), .Z(c[209]) );
  XNOR U886 ( .A(b[208]), .B(n885), .Z(c[208]) );
  XNOR U887 ( .A(b[207]), .B(n886), .Z(c[207]) );
  XNOR U888 ( .A(b[206]), .B(n887), .Z(c[206]) );
  XNOR U889 ( .A(b[205]), .B(n888), .Z(c[205]) );
  XNOR U890 ( .A(b[204]), .B(n889), .Z(c[204]) );
  XNOR U891 ( .A(b[2047]), .B(n5), .Z(c[2047]) );
  XNOR U892 ( .A(a[2047]), .B(n3), .Z(n5) );
  XNOR U893 ( .A(n890), .B(n891), .Z(n3) );
  ANDN U894 ( .B(n892), .A(n893), .Z(n890) );
  XNOR U895 ( .A(b[2046]), .B(n891), .Z(n892) );
  XNOR U896 ( .A(b[2046]), .B(n893), .Z(c[2046]) );
  XNOR U897 ( .A(a[2046]), .B(n894), .Z(n893) );
  IV U898 ( .A(n891), .Z(n894) );
  XOR U899 ( .A(n895), .B(n896), .Z(n891) );
  ANDN U900 ( .B(n897), .A(n898), .Z(n895) );
  XNOR U901 ( .A(b[2045]), .B(n896), .Z(n897) );
  XNOR U902 ( .A(b[2045]), .B(n898), .Z(c[2045]) );
  XNOR U903 ( .A(a[2045]), .B(n899), .Z(n898) );
  IV U904 ( .A(n896), .Z(n899) );
  XOR U905 ( .A(n900), .B(n901), .Z(n896) );
  ANDN U906 ( .B(n902), .A(n903), .Z(n900) );
  XNOR U907 ( .A(b[2044]), .B(n901), .Z(n902) );
  XNOR U908 ( .A(b[2044]), .B(n903), .Z(c[2044]) );
  XNOR U909 ( .A(a[2044]), .B(n904), .Z(n903) );
  IV U910 ( .A(n901), .Z(n904) );
  XOR U911 ( .A(n905), .B(n906), .Z(n901) );
  ANDN U912 ( .B(n907), .A(n908), .Z(n905) );
  XNOR U913 ( .A(b[2043]), .B(n906), .Z(n907) );
  XNOR U914 ( .A(b[2043]), .B(n908), .Z(c[2043]) );
  XNOR U915 ( .A(a[2043]), .B(n909), .Z(n908) );
  IV U916 ( .A(n906), .Z(n909) );
  XOR U917 ( .A(n910), .B(n911), .Z(n906) );
  ANDN U918 ( .B(n912), .A(n913), .Z(n910) );
  XNOR U919 ( .A(b[2042]), .B(n911), .Z(n912) );
  XNOR U920 ( .A(b[2042]), .B(n913), .Z(c[2042]) );
  XNOR U921 ( .A(a[2042]), .B(n914), .Z(n913) );
  IV U922 ( .A(n911), .Z(n914) );
  XOR U923 ( .A(n915), .B(n916), .Z(n911) );
  ANDN U924 ( .B(n917), .A(n918), .Z(n915) );
  XNOR U925 ( .A(b[2041]), .B(n916), .Z(n917) );
  XNOR U926 ( .A(b[2041]), .B(n918), .Z(c[2041]) );
  XNOR U927 ( .A(a[2041]), .B(n919), .Z(n918) );
  IV U928 ( .A(n916), .Z(n919) );
  XOR U929 ( .A(n920), .B(n921), .Z(n916) );
  ANDN U930 ( .B(n922), .A(n923), .Z(n920) );
  XNOR U931 ( .A(b[2040]), .B(n921), .Z(n922) );
  XNOR U932 ( .A(b[2040]), .B(n923), .Z(c[2040]) );
  XNOR U933 ( .A(a[2040]), .B(n924), .Z(n923) );
  IV U934 ( .A(n921), .Z(n924) );
  XOR U935 ( .A(n925), .B(n926), .Z(n921) );
  ANDN U936 ( .B(n927), .A(n928), .Z(n925) );
  XNOR U937 ( .A(b[2039]), .B(n926), .Z(n927) );
  XNOR U938 ( .A(b[203]), .B(n929), .Z(c[203]) );
  XNOR U939 ( .A(b[2039]), .B(n928), .Z(c[2039]) );
  XNOR U940 ( .A(a[2039]), .B(n930), .Z(n928) );
  IV U941 ( .A(n926), .Z(n930) );
  XOR U942 ( .A(n931), .B(n932), .Z(n926) );
  ANDN U943 ( .B(n933), .A(n934), .Z(n931) );
  XNOR U944 ( .A(b[2038]), .B(n932), .Z(n933) );
  XNOR U945 ( .A(b[2038]), .B(n934), .Z(c[2038]) );
  XNOR U946 ( .A(a[2038]), .B(n935), .Z(n934) );
  IV U947 ( .A(n932), .Z(n935) );
  XOR U948 ( .A(n936), .B(n937), .Z(n932) );
  ANDN U949 ( .B(n938), .A(n939), .Z(n936) );
  XNOR U950 ( .A(b[2037]), .B(n937), .Z(n938) );
  XNOR U951 ( .A(b[2037]), .B(n939), .Z(c[2037]) );
  XNOR U952 ( .A(a[2037]), .B(n940), .Z(n939) );
  IV U953 ( .A(n937), .Z(n940) );
  XOR U954 ( .A(n941), .B(n942), .Z(n937) );
  ANDN U955 ( .B(n943), .A(n944), .Z(n941) );
  XNOR U956 ( .A(b[2036]), .B(n942), .Z(n943) );
  XNOR U957 ( .A(b[2036]), .B(n944), .Z(c[2036]) );
  XNOR U958 ( .A(a[2036]), .B(n945), .Z(n944) );
  IV U959 ( .A(n942), .Z(n945) );
  XOR U960 ( .A(n946), .B(n947), .Z(n942) );
  ANDN U961 ( .B(n948), .A(n949), .Z(n946) );
  XNOR U962 ( .A(b[2035]), .B(n947), .Z(n948) );
  XNOR U963 ( .A(b[2035]), .B(n949), .Z(c[2035]) );
  XNOR U964 ( .A(a[2035]), .B(n950), .Z(n949) );
  IV U965 ( .A(n947), .Z(n950) );
  XOR U966 ( .A(n951), .B(n952), .Z(n947) );
  ANDN U967 ( .B(n953), .A(n954), .Z(n951) );
  XNOR U968 ( .A(b[2034]), .B(n952), .Z(n953) );
  XNOR U969 ( .A(b[2034]), .B(n954), .Z(c[2034]) );
  XNOR U970 ( .A(a[2034]), .B(n955), .Z(n954) );
  IV U971 ( .A(n952), .Z(n955) );
  XOR U972 ( .A(n956), .B(n957), .Z(n952) );
  ANDN U973 ( .B(n958), .A(n959), .Z(n956) );
  XNOR U974 ( .A(b[2033]), .B(n957), .Z(n958) );
  XNOR U975 ( .A(b[2033]), .B(n959), .Z(c[2033]) );
  XNOR U976 ( .A(a[2033]), .B(n960), .Z(n959) );
  IV U977 ( .A(n957), .Z(n960) );
  XOR U978 ( .A(n961), .B(n962), .Z(n957) );
  ANDN U979 ( .B(n963), .A(n964), .Z(n961) );
  XNOR U980 ( .A(b[2032]), .B(n962), .Z(n963) );
  XNOR U981 ( .A(b[2032]), .B(n964), .Z(c[2032]) );
  XNOR U982 ( .A(a[2032]), .B(n965), .Z(n964) );
  IV U983 ( .A(n962), .Z(n965) );
  XOR U984 ( .A(n966), .B(n967), .Z(n962) );
  ANDN U985 ( .B(n968), .A(n969), .Z(n966) );
  XNOR U986 ( .A(b[2031]), .B(n967), .Z(n968) );
  XNOR U987 ( .A(b[2031]), .B(n969), .Z(c[2031]) );
  XNOR U988 ( .A(a[2031]), .B(n970), .Z(n969) );
  IV U989 ( .A(n967), .Z(n970) );
  XOR U990 ( .A(n971), .B(n972), .Z(n967) );
  ANDN U991 ( .B(n973), .A(n974), .Z(n971) );
  XNOR U992 ( .A(b[2030]), .B(n972), .Z(n973) );
  XNOR U993 ( .A(b[2030]), .B(n974), .Z(c[2030]) );
  XNOR U994 ( .A(a[2030]), .B(n975), .Z(n974) );
  IV U995 ( .A(n972), .Z(n975) );
  XOR U996 ( .A(n976), .B(n977), .Z(n972) );
  ANDN U997 ( .B(n978), .A(n979), .Z(n976) );
  XNOR U998 ( .A(b[2029]), .B(n977), .Z(n978) );
  XNOR U999 ( .A(b[202]), .B(n980), .Z(c[202]) );
  XNOR U1000 ( .A(b[2029]), .B(n979), .Z(c[2029]) );
  XNOR U1001 ( .A(a[2029]), .B(n981), .Z(n979) );
  IV U1002 ( .A(n977), .Z(n981) );
  XOR U1003 ( .A(n982), .B(n983), .Z(n977) );
  ANDN U1004 ( .B(n984), .A(n985), .Z(n982) );
  XNOR U1005 ( .A(b[2028]), .B(n983), .Z(n984) );
  XNOR U1006 ( .A(b[2028]), .B(n985), .Z(c[2028]) );
  XNOR U1007 ( .A(a[2028]), .B(n986), .Z(n985) );
  IV U1008 ( .A(n983), .Z(n986) );
  XOR U1009 ( .A(n987), .B(n988), .Z(n983) );
  ANDN U1010 ( .B(n989), .A(n990), .Z(n987) );
  XNOR U1011 ( .A(b[2027]), .B(n988), .Z(n989) );
  XNOR U1012 ( .A(b[2027]), .B(n990), .Z(c[2027]) );
  XNOR U1013 ( .A(a[2027]), .B(n991), .Z(n990) );
  IV U1014 ( .A(n988), .Z(n991) );
  XOR U1015 ( .A(n992), .B(n993), .Z(n988) );
  ANDN U1016 ( .B(n994), .A(n995), .Z(n992) );
  XNOR U1017 ( .A(b[2026]), .B(n993), .Z(n994) );
  XNOR U1018 ( .A(b[2026]), .B(n995), .Z(c[2026]) );
  XNOR U1019 ( .A(a[2026]), .B(n996), .Z(n995) );
  IV U1020 ( .A(n993), .Z(n996) );
  XOR U1021 ( .A(n997), .B(n998), .Z(n993) );
  ANDN U1022 ( .B(n999), .A(n1000), .Z(n997) );
  XNOR U1023 ( .A(b[2025]), .B(n998), .Z(n999) );
  XNOR U1024 ( .A(b[2025]), .B(n1000), .Z(c[2025]) );
  XNOR U1025 ( .A(a[2025]), .B(n1001), .Z(n1000) );
  IV U1026 ( .A(n998), .Z(n1001) );
  XOR U1027 ( .A(n1002), .B(n1003), .Z(n998) );
  ANDN U1028 ( .B(n1004), .A(n1005), .Z(n1002) );
  XNOR U1029 ( .A(b[2024]), .B(n1003), .Z(n1004) );
  XNOR U1030 ( .A(b[2024]), .B(n1005), .Z(c[2024]) );
  XNOR U1031 ( .A(a[2024]), .B(n1006), .Z(n1005) );
  IV U1032 ( .A(n1003), .Z(n1006) );
  XOR U1033 ( .A(n1007), .B(n1008), .Z(n1003) );
  ANDN U1034 ( .B(n1009), .A(n1010), .Z(n1007) );
  XNOR U1035 ( .A(b[2023]), .B(n1008), .Z(n1009) );
  XNOR U1036 ( .A(b[2023]), .B(n1010), .Z(c[2023]) );
  XNOR U1037 ( .A(a[2023]), .B(n1011), .Z(n1010) );
  IV U1038 ( .A(n1008), .Z(n1011) );
  XOR U1039 ( .A(n1012), .B(n1013), .Z(n1008) );
  ANDN U1040 ( .B(n1014), .A(n1015), .Z(n1012) );
  XNOR U1041 ( .A(b[2022]), .B(n1013), .Z(n1014) );
  XNOR U1042 ( .A(b[2022]), .B(n1015), .Z(c[2022]) );
  XNOR U1043 ( .A(a[2022]), .B(n1016), .Z(n1015) );
  IV U1044 ( .A(n1013), .Z(n1016) );
  XOR U1045 ( .A(n1017), .B(n1018), .Z(n1013) );
  ANDN U1046 ( .B(n1019), .A(n1020), .Z(n1017) );
  XNOR U1047 ( .A(b[2021]), .B(n1018), .Z(n1019) );
  XNOR U1048 ( .A(b[2021]), .B(n1020), .Z(c[2021]) );
  XNOR U1049 ( .A(a[2021]), .B(n1021), .Z(n1020) );
  IV U1050 ( .A(n1018), .Z(n1021) );
  XOR U1051 ( .A(n1022), .B(n1023), .Z(n1018) );
  ANDN U1052 ( .B(n1024), .A(n1025), .Z(n1022) );
  XNOR U1053 ( .A(b[2020]), .B(n1023), .Z(n1024) );
  XNOR U1054 ( .A(b[2020]), .B(n1025), .Z(c[2020]) );
  XNOR U1055 ( .A(a[2020]), .B(n1026), .Z(n1025) );
  IV U1056 ( .A(n1023), .Z(n1026) );
  XOR U1057 ( .A(n1027), .B(n1028), .Z(n1023) );
  ANDN U1058 ( .B(n1029), .A(n1030), .Z(n1027) );
  XNOR U1059 ( .A(b[2019]), .B(n1028), .Z(n1029) );
  XNOR U1060 ( .A(b[201]), .B(n1031), .Z(c[201]) );
  XNOR U1061 ( .A(b[2019]), .B(n1030), .Z(c[2019]) );
  XNOR U1062 ( .A(a[2019]), .B(n1032), .Z(n1030) );
  IV U1063 ( .A(n1028), .Z(n1032) );
  XOR U1064 ( .A(n1033), .B(n1034), .Z(n1028) );
  ANDN U1065 ( .B(n1035), .A(n1036), .Z(n1033) );
  XNOR U1066 ( .A(b[2018]), .B(n1034), .Z(n1035) );
  XNOR U1067 ( .A(b[2018]), .B(n1036), .Z(c[2018]) );
  XNOR U1068 ( .A(a[2018]), .B(n1037), .Z(n1036) );
  IV U1069 ( .A(n1034), .Z(n1037) );
  XOR U1070 ( .A(n1038), .B(n1039), .Z(n1034) );
  ANDN U1071 ( .B(n1040), .A(n1041), .Z(n1038) );
  XNOR U1072 ( .A(b[2017]), .B(n1039), .Z(n1040) );
  XNOR U1073 ( .A(b[2017]), .B(n1041), .Z(c[2017]) );
  XNOR U1074 ( .A(a[2017]), .B(n1042), .Z(n1041) );
  IV U1075 ( .A(n1039), .Z(n1042) );
  XOR U1076 ( .A(n1043), .B(n1044), .Z(n1039) );
  ANDN U1077 ( .B(n1045), .A(n1046), .Z(n1043) );
  XNOR U1078 ( .A(b[2016]), .B(n1044), .Z(n1045) );
  XNOR U1079 ( .A(b[2016]), .B(n1046), .Z(c[2016]) );
  XNOR U1080 ( .A(a[2016]), .B(n1047), .Z(n1046) );
  IV U1081 ( .A(n1044), .Z(n1047) );
  XOR U1082 ( .A(n1048), .B(n1049), .Z(n1044) );
  ANDN U1083 ( .B(n1050), .A(n1051), .Z(n1048) );
  XNOR U1084 ( .A(b[2015]), .B(n1049), .Z(n1050) );
  XNOR U1085 ( .A(b[2015]), .B(n1051), .Z(c[2015]) );
  XNOR U1086 ( .A(a[2015]), .B(n1052), .Z(n1051) );
  IV U1087 ( .A(n1049), .Z(n1052) );
  XOR U1088 ( .A(n1053), .B(n1054), .Z(n1049) );
  ANDN U1089 ( .B(n1055), .A(n1056), .Z(n1053) );
  XNOR U1090 ( .A(b[2014]), .B(n1054), .Z(n1055) );
  XNOR U1091 ( .A(b[2014]), .B(n1056), .Z(c[2014]) );
  XNOR U1092 ( .A(a[2014]), .B(n1057), .Z(n1056) );
  IV U1093 ( .A(n1054), .Z(n1057) );
  XOR U1094 ( .A(n1058), .B(n1059), .Z(n1054) );
  ANDN U1095 ( .B(n1060), .A(n1061), .Z(n1058) );
  XNOR U1096 ( .A(b[2013]), .B(n1059), .Z(n1060) );
  XNOR U1097 ( .A(b[2013]), .B(n1061), .Z(c[2013]) );
  XNOR U1098 ( .A(a[2013]), .B(n1062), .Z(n1061) );
  IV U1099 ( .A(n1059), .Z(n1062) );
  XOR U1100 ( .A(n1063), .B(n1064), .Z(n1059) );
  ANDN U1101 ( .B(n1065), .A(n1066), .Z(n1063) );
  XNOR U1102 ( .A(b[2012]), .B(n1064), .Z(n1065) );
  XNOR U1103 ( .A(b[2012]), .B(n1066), .Z(c[2012]) );
  XNOR U1104 ( .A(a[2012]), .B(n1067), .Z(n1066) );
  IV U1105 ( .A(n1064), .Z(n1067) );
  XOR U1106 ( .A(n1068), .B(n1069), .Z(n1064) );
  ANDN U1107 ( .B(n1070), .A(n1071), .Z(n1068) );
  XNOR U1108 ( .A(b[2011]), .B(n1069), .Z(n1070) );
  XNOR U1109 ( .A(b[2011]), .B(n1071), .Z(c[2011]) );
  XNOR U1110 ( .A(a[2011]), .B(n1072), .Z(n1071) );
  IV U1111 ( .A(n1069), .Z(n1072) );
  XOR U1112 ( .A(n1073), .B(n1074), .Z(n1069) );
  ANDN U1113 ( .B(n1075), .A(n1076), .Z(n1073) );
  XNOR U1114 ( .A(b[2010]), .B(n1074), .Z(n1075) );
  XNOR U1115 ( .A(b[2010]), .B(n1076), .Z(c[2010]) );
  XNOR U1116 ( .A(a[2010]), .B(n1077), .Z(n1076) );
  IV U1117 ( .A(n1074), .Z(n1077) );
  XOR U1118 ( .A(n1078), .B(n1079), .Z(n1074) );
  ANDN U1119 ( .B(n1080), .A(n1081), .Z(n1078) );
  XNOR U1120 ( .A(b[2009]), .B(n1079), .Z(n1080) );
  XNOR U1121 ( .A(b[200]), .B(n1082), .Z(c[200]) );
  XNOR U1122 ( .A(b[2009]), .B(n1081), .Z(c[2009]) );
  XNOR U1123 ( .A(a[2009]), .B(n1083), .Z(n1081) );
  IV U1124 ( .A(n1079), .Z(n1083) );
  XOR U1125 ( .A(n1084), .B(n1085), .Z(n1079) );
  ANDN U1126 ( .B(n1086), .A(n1087), .Z(n1084) );
  XNOR U1127 ( .A(b[2008]), .B(n1085), .Z(n1086) );
  XNOR U1128 ( .A(b[2008]), .B(n1087), .Z(c[2008]) );
  XNOR U1129 ( .A(a[2008]), .B(n1088), .Z(n1087) );
  IV U1130 ( .A(n1085), .Z(n1088) );
  XOR U1131 ( .A(n1089), .B(n1090), .Z(n1085) );
  ANDN U1132 ( .B(n1091), .A(n1092), .Z(n1089) );
  XNOR U1133 ( .A(b[2007]), .B(n1090), .Z(n1091) );
  XNOR U1134 ( .A(b[2007]), .B(n1092), .Z(c[2007]) );
  XNOR U1135 ( .A(a[2007]), .B(n1093), .Z(n1092) );
  IV U1136 ( .A(n1090), .Z(n1093) );
  XOR U1137 ( .A(n1094), .B(n1095), .Z(n1090) );
  ANDN U1138 ( .B(n1096), .A(n1097), .Z(n1094) );
  XNOR U1139 ( .A(b[2006]), .B(n1095), .Z(n1096) );
  XNOR U1140 ( .A(b[2006]), .B(n1097), .Z(c[2006]) );
  XNOR U1141 ( .A(a[2006]), .B(n1098), .Z(n1097) );
  IV U1142 ( .A(n1095), .Z(n1098) );
  XOR U1143 ( .A(n1099), .B(n1100), .Z(n1095) );
  ANDN U1144 ( .B(n1101), .A(n1102), .Z(n1099) );
  XNOR U1145 ( .A(b[2005]), .B(n1100), .Z(n1101) );
  XNOR U1146 ( .A(b[2005]), .B(n1102), .Z(c[2005]) );
  XNOR U1147 ( .A(a[2005]), .B(n1103), .Z(n1102) );
  IV U1148 ( .A(n1100), .Z(n1103) );
  XOR U1149 ( .A(n1104), .B(n1105), .Z(n1100) );
  ANDN U1150 ( .B(n1106), .A(n1107), .Z(n1104) );
  XNOR U1151 ( .A(b[2004]), .B(n1105), .Z(n1106) );
  XNOR U1152 ( .A(b[2004]), .B(n1107), .Z(c[2004]) );
  XNOR U1153 ( .A(a[2004]), .B(n1108), .Z(n1107) );
  IV U1154 ( .A(n1105), .Z(n1108) );
  XOR U1155 ( .A(n1109), .B(n1110), .Z(n1105) );
  ANDN U1156 ( .B(n1111), .A(n1112), .Z(n1109) );
  XNOR U1157 ( .A(b[2003]), .B(n1110), .Z(n1111) );
  XNOR U1158 ( .A(b[2003]), .B(n1112), .Z(c[2003]) );
  XNOR U1159 ( .A(a[2003]), .B(n1113), .Z(n1112) );
  IV U1160 ( .A(n1110), .Z(n1113) );
  XOR U1161 ( .A(n1114), .B(n1115), .Z(n1110) );
  ANDN U1162 ( .B(n1116), .A(n1117), .Z(n1114) );
  XNOR U1163 ( .A(b[2002]), .B(n1115), .Z(n1116) );
  XNOR U1164 ( .A(b[2002]), .B(n1117), .Z(c[2002]) );
  XNOR U1165 ( .A(a[2002]), .B(n1118), .Z(n1117) );
  IV U1166 ( .A(n1115), .Z(n1118) );
  XOR U1167 ( .A(n1119), .B(n1120), .Z(n1115) );
  ANDN U1168 ( .B(n1121), .A(n1122), .Z(n1119) );
  XNOR U1169 ( .A(b[2001]), .B(n1120), .Z(n1121) );
  XNOR U1170 ( .A(b[2001]), .B(n1122), .Z(c[2001]) );
  XNOR U1171 ( .A(a[2001]), .B(n1123), .Z(n1122) );
  IV U1172 ( .A(n1120), .Z(n1123) );
  XOR U1173 ( .A(n1124), .B(n1125), .Z(n1120) );
  ANDN U1174 ( .B(n1126), .A(n1127), .Z(n1124) );
  XNOR U1175 ( .A(b[2000]), .B(n1125), .Z(n1126) );
  XNOR U1176 ( .A(b[2000]), .B(n1127), .Z(c[2000]) );
  XNOR U1177 ( .A(a[2000]), .B(n1128), .Z(n1127) );
  IV U1178 ( .A(n1125), .Z(n1128) );
  XOR U1179 ( .A(n1129), .B(n1130), .Z(n1125) );
  ANDN U1180 ( .B(n1131), .A(n1132), .Z(n1129) );
  XNOR U1181 ( .A(b[1999]), .B(n1130), .Z(n1131) );
  XNOR U1182 ( .A(b[1]), .B(n1133), .Z(c[1]) );
  XNOR U1183 ( .A(b[19]), .B(n1134), .Z(c[19]) );
  XNOR U1184 ( .A(b[199]), .B(n1135), .Z(c[199]) );
  XNOR U1185 ( .A(b[1999]), .B(n1132), .Z(c[1999]) );
  XNOR U1186 ( .A(a[1999]), .B(n1136), .Z(n1132) );
  IV U1187 ( .A(n1130), .Z(n1136) );
  XOR U1188 ( .A(n1137), .B(n1138), .Z(n1130) );
  ANDN U1189 ( .B(n1139), .A(n1140), .Z(n1137) );
  XNOR U1190 ( .A(b[1998]), .B(n1138), .Z(n1139) );
  XNOR U1191 ( .A(b[1998]), .B(n1140), .Z(c[1998]) );
  XNOR U1192 ( .A(a[1998]), .B(n1141), .Z(n1140) );
  IV U1193 ( .A(n1138), .Z(n1141) );
  XOR U1194 ( .A(n1142), .B(n1143), .Z(n1138) );
  ANDN U1195 ( .B(n1144), .A(n1145), .Z(n1142) );
  XNOR U1196 ( .A(b[1997]), .B(n1143), .Z(n1144) );
  XNOR U1197 ( .A(b[1997]), .B(n1145), .Z(c[1997]) );
  XNOR U1198 ( .A(a[1997]), .B(n1146), .Z(n1145) );
  IV U1199 ( .A(n1143), .Z(n1146) );
  XOR U1200 ( .A(n1147), .B(n1148), .Z(n1143) );
  ANDN U1201 ( .B(n1149), .A(n1150), .Z(n1147) );
  XNOR U1202 ( .A(b[1996]), .B(n1148), .Z(n1149) );
  XNOR U1203 ( .A(b[1996]), .B(n1150), .Z(c[1996]) );
  XNOR U1204 ( .A(a[1996]), .B(n1151), .Z(n1150) );
  IV U1205 ( .A(n1148), .Z(n1151) );
  XOR U1206 ( .A(n1152), .B(n1153), .Z(n1148) );
  ANDN U1207 ( .B(n1154), .A(n1155), .Z(n1152) );
  XNOR U1208 ( .A(b[1995]), .B(n1153), .Z(n1154) );
  XNOR U1209 ( .A(b[1995]), .B(n1155), .Z(c[1995]) );
  XNOR U1210 ( .A(a[1995]), .B(n1156), .Z(n1155) );
  IV U1211 ( .A(n1153), .Z(n1156) );
  XOR U1212 ( .A(n1157), .B(n1158), .Z(n1153) );
  ANDN U1213 ( .B(n1159), .A(n1160), .Z(n1157) );
  XNOR U1214 ( .A(b[1994]), .B(n1158), .Z(n1159) );
  XNOR U1215 ( .A(b[1994]), .B(n1160), .Z(c[1994]) );
  XNOR U1216 ( .A(a[1994]), .B(n1161), .Z(n1160) );
  IV U1217 ( .A(n1158), .Z(n1161) );
  XOR U1218 ( .A(n1162), .B(n1163), .Z(n1158) );
  ANDN U1219 ( .B(n1164), .A(n1165), .Z(n1162) );
  XNOR U1220 ( .A(b[1993]), .B(n1163), .Z(n1164) );
  XNOR U1221 ( .A(b[1993]), .B(n1165), .Z(c[1993]) );
  XNOR U1222 ( .A(a[1993]), .B(n1166), .Z(n1165) );
  IV U1223 ( .A(n1163), .Z(n1166) );
  XOR U1224 ( .A(n1167), .B(n1168), .Z(n1163) );
  ANDN U1225 ( .B(n1169), .A(n1170), .Z(n1167) );
  XNOR U1226 ( .A(b[1992]), .B(n1168), .Z(n1169) );
  XNOR U1227 ( .A(b[1992]), .B(n1170), .Z(c[1992]) );
  XNOR U1228 ( .A(a[1992]), .B(n1171), .Z(n1170) );
  IV U1229 ( .A(n1168), .Z(n1171) );
  XOR U1230 ( .A(n1172), .B(n1173), .Z(n1168) );
  ANDN U1231 ( .B(n1174), .A(n1175), .Z(n1172) );
  XNOR U1232 ( .A(b[1991]), .B(n1173), .Z(n1174) );
  XNOR U1233 ( .A(b[1991]), .B(n1175), .Z(c[1991]) );
  XNOR U1234 ( .A(a[1991]), .B(n1176), .Z(n1175) );
  IV U1235 ( .A(n1173), .Z(n1176) );
  XOR U1236 ( .A(n1177), .B(n1178), .Z(n1173) );
  ANDN U1237 ( .B(n1179), .A(n1180), .Z(n1177) );
  XNOR U1238 ( .A(b[1990]), .B(n1178), .Z(n1179) );
  XNOR U1239 ( .A(b[1990]), .B(n1180), .Z(c[1990]) );
  XNOR U1240 ( .A(a[1990]), .B(n1181), .Z(n1180) );
  IV U1241 ( .A(n1178), .Z(n1181) );
  XOR U1242 ( .A(n1182), .B(n1183), .Z(n1178) );
  ANDN U1243 ( .B(n1184), .A(n1185), .Z(n1182) );
  XNOR U1244 ( .A(b[1989]), .B(n1183), .Z(n1184) );
  XNOR U1245 ( .A(b[198]), .B(n1186), .Z(c[198]) );
  XNOR U1246 ( .A(b[1989]), .B(n1185), .Z(c[1989]) );
  XNOR U1247 ( .A(a[1989]), .B(n1187), .Z(n1185) );
  IV U1248 ( .A(n1183), .Z(n1187) );
  XOR U1249 ( .A(n1188), .B(n1189), .Z(n1183) );
  ANDN U1250 ( .B(n1190), .A(n1191), .Z(n1188) );
  XNOR U1251 ( .A(b[1988]), .B(n1189), .Z(n1190) );
  XNOR U1252 ( .A(b[1988]), .B(n1191), .Z(c[1988]) );
  XNOR U1253 ( .A(a[1988]), .B(n1192), .Z(n1191) );
  IV U1254 ( .A(n1189), .Z(n1192) );
  XOR U1255 ( .A(n1193), .B(n1194), .Z(n1189) );
  ANDN U1256 ( .B(n1195), .A(n1196), .Z(n1193) );
  XNOR U1257 ( .A(b[1987]), .B(n1194), .Z(n1195) );
  XNOR U1258 ( .A(b[1987]), .B(n1196), .Z(c[1987]) );
  XNOR U1259 ( .A(a[1987]), .B(n1197), .Z(n1196) );
  IV U1260 ( .A(n1194), .Z(n1197) );
  XOR U1261 ( .A(n1198), .B(n1199), .Z(n1194) );
  ANDN U1262 ( .B(n1200), .A(n1201), .Z(n1198) );
  XNOR U1263 ( .A(b[1986]), .B(n1199), .Z(n1200) );
  XNOR U1264 ( .A(b[1986]), .B(n1201), .Z(c[1986]) );
  XNOR U1265 ( .A(a[1986]), .B(n1202), .Z(n1201) );
  IV U1266 ( .A(n1199), .Z(n1202) );
  XOR U1267 ( .A(n1203), .B(n1204), .Z(n1199) );
  ANDN U1268 ( .B(n1205), .A(n1206), .Z(n1203) );
  XNOR U1269 ( .A(b[1985]), .B(n1204), .Z(n1205) );
  XNOR U1270 ( .A(b[1985]), .B(n1206), .Z(c[1985]) );
  XNOR U1271 ( .A(a[1985]), .B(n1207), .Z(n1206) );
  IV U1272 ( .A(n1204), .Z(n1207) );
  XOR U1273 ( .A(n1208), .B(n1209), .Z(n1204) );
  ANDN U1274 ( .B(n1210), .A(n1211), .Z(n1208) );
  XNOR U1275 ( .A(b[1984]), .B(n1209), .Z(n1210) );
  XNOR U1276 ( .A(b[1984]), .B(n1211), .Z(c[1984]) );
  XNOR U1277 ( .A(a[1984]), .B(n1212), .Z(n1211) );
  IV U1278 ( .A(n1209), .Z(n1212) );
  XOR U1279 ( .A(n1213), .B(n1214), .Z(n1209) );
  ANDN U1280 ( .B(n1215), .A(n1216), .Z(n1213) );
  XNOR U1281 ( .A(b[1983]), .B(n1214), .Z(n1215) );
  XNOR U1282 ( .A(b[1983]), .B(n1216), .Z(c[1983]) );
  XNOR U1283 ( .A(a[1983]), .B(n1217), .Z(n1216) );
  IV U1284 ( .A(n1214), .Z(n1217) );
  XOR U1285 ( .A(n1218), .B(n1219), .Z(n1214) );
  ANDN U1286 ( .B(n1220), .A(n1221), .Z(n1218) );
  XNOR U1287 ( .A(b[1982]), .B(n1219), .Z(n1220) );
  XNOR U1288 ( .A(b[1982]), .B(n1221), .Z(c[1982]) );
  XNOR U1289 ( .A(a[1982]), .B(n1222), .Z(n1221) );
  IV U1290 ( .A(n1219), .Z(n1222) );
  XOR U1291 ( .A(n1223), .B(n1224), .Z(n1219) );
  ANDN U1292 ( .B(n1225), .A(n1226), .Z(n1223) );
  XNOR U1293 ( .A(b[1981]), .B(n1224), .Z(n1225) );
  XNOR U1294 ( .A(b[1981]), .B(n1226), .Z(c[1981]) );
  XNOR U1295 ( .A(a[1981]), .B(n1227), .Z(n1226) );
  IV U1296 ( .A(n1224), .Z(n1227) );
  XOR U1297 ( .A(n1228), .B(n1229), .Z(n1224) );
  ANDN U1298 ( .B(n1230), .A(n1231), .Z(n1228) );
  XNOR U1299 ( .A(b[1980]), .B(n1229), .Z(n1230) );
  XNOR U1300 ( .A(b[1980]), .B(n1231), .Z(c[1980]) );
  XNOR U1301 ( .A(a[1980]), .B(n1232), .Z(n1231) );
  IV U1302 ( .A(n1229), .Z(n1232) );
  XOR U1303 ( .A(n1233), .B(n1234), .Z(n1229) );
  ANDN U1304 ( .B(n1235), .A(n1236), .Z(n1233) );
  XNOR U1305 ( .A(b[1979]), .B(n1234), .Z(n1235) );
  XNOR U1306 ( .A(b[197]), .B(n1237), .Z(c[197]) );
  XNOR U1307 ( .A(b[1979]), .B(n1236), .Z(c[1979]) );
  XNOR U1308 ( .A(a[1979]), .B(n1238), .Z(n1236) );
  IV U1309 ( .A(n1234), .Z(n1238) );
  XOR U1310 ( .A(n1239), .B(n1240), .Z(n1234) );
  ANDN U1311 ( .B(n1241), .A(n1242), .Z(n1239) );
  XNOR U1312 ( .A(b[1978]), .B(n1240), .Z(n1241) );
  XNOR U1313 ( .A(b[1978]), .B(n1242), .Z(c[1978]) );
  XNOR U1314 ( .A(a[1978]), .B(n1243), .Z(n1242) );
  IV U1315 ( .A(n1240), .Z(n1243) );
  XOR U1316 ( .A(n1244), .B(n1245), .Z(n1240) );
  ANDN U1317 ( .B(n1246), .A(n1247), .Z(n1244) );
  XNOR U1318 ( .A(b[1977]), .B(n1245), .Z(n1246) );
  XNOR U1319 ( .A(b[1977]), .B(n1247), .Z(c[1977]) );
  XNOR U1320 ( .A(a[1977]), .B(n1248), .Z(n1247) );
  IV U1321 ( .A(n1245), .Z(n1248) );
  XOR U1322 ( .A(n1249), .B(n1250), .Z(n1245) );
  ANDN U1323 ( .B(n1251), .A(n1252), .Z(n1249) );
  XNOR U1324 ( .A(b[1976]), .B(n1250), .Z(n1251) );
  XNOR U1325 ( .A(b[1976]), .B(n1252), .Z(c[1976]) );
  XNOR U1326 ( .A(a[1976]), .B(n1253), .Z(n1252) );
  IV U1327 ( .A(n1250), .Z(n1253) );
  XOR U1328 ( .A(n1254), .B(n1255), .Z(n1250) );
  ANDN U1329 ( .B(n1256), .A(n1257), .Z(n1254) );
  XNOR U1330 ( .A(b[1975]), .B(n1255), .Z(n1256) );
  XNOR U1331 ( .A(b[1975]), .B(n1257), .Z(c[1975]) );
  XNOR U1332 ( .A(a[1975]), .B(n1258), .Z(n1257) );
  IV U1333 ( .A(n1255), .Z(n1258) );
  XOR U1334 ( .A(n1259), .B(n1260), .Z(n1255) );
  ANDN U1335 ( .B(n1261), .A(n1262), .Z(n1259) );
  XNOR U1336 ( .A(b[1974]), .B(n1260), .Z(n1261) );
  XNOR U1337 ( .A(b[1974]), .B(n1262), .Z(c[1974]) );
  XNOR U1338 ( .A(a[1974]), .B(n1263), .Z(n1262) );
  IV U1339 ( .A(n1260), .Z(n1263) );
  XOR U1340 ( .A(n1264), .B(n1265), .Z(n1260) );
  ANDN U1341 ( .B(n1266), .A(n1267), .Z(n1264) );
  XNOR U1342 ( .A(b[1973]), .B(n1265), .Z(n1266) );
  XNOR U1343 ( .A(b[1973]), .B(n1267), .Z(c[1973]) );
  XNOR U1344 ( .A(a[1973]), .B(n1268), .Z(n1267) );
  IV U1345 ( .A(n1265), .Z(n1268) );
  XOR U1346 ( .A(n1269), .B(n1270), .Z(n1265) );
  ANDN U1347 ( .B(n1271), .A(n1272), .Z(n1269) );
  XNOR U1348 ( .A(b[1972]), .B(n1270), .Z(n1271) );
  XNOR U1349 ( .A(b[1972]), .B(n1272), .Z(c[1972]) );
  XNOR U1350 ( .A(a[1972]), .B(n1273), .Z(n1272) );
  IV U1351 ( .A(n1270), .Z(n1273) );
  XOR U1352 ( .A(n1274), .B(n1275), .Z(n1270) );
  ANDN U1353 ( .B(n1276), .A(n1277), .Z(n1274) );
  XNOR U1354 ( .A(b[1971]), .B(n1275), .Z(n1276) );
  XNOR U1355 ( .A(b[1971]), .B(n1277), .Z(c[1971]) );
  XNOR U1356 ( .A(a[1971]), .B(n1278), .Z(n1277) );
  IV U1357 ( .A(n1275), .Z(n1278) );
  XOR U1358 ( .A(n1279), .B(n1280), .Z(n1275) );
  ANDN U1359 ( .B(n1281), .A(n1282), .Z(n1279) );
  XNOR U1360 ( .A(b[1970]), .B(n1280), .Z(n1281) );
  XNOR U1361 ( .A(b[1970]), .B(n1282), .Z(c[1970]) );
  XNOR U1362 ( .A(a[1970]), .B(n1283), .Z(n1282) );
  IV U1363 ( .A(n1280), .Z(n1283) );
  XOR U1364 ( .A(n1284), .B(n1285), .Z(n1280) );
  ANDN U1365 ( .B(n1286), .A(n1287), .Z(n1284) );
  XNOR U1366 ( .A(b[1969]), .B(n1285), .Z(n1286) );
  XNOR U1367 ( .A(b[196]), .B(n1288), .Z(c[196]) );
  XNOR U1368 ( .A(b[1969]), .B(n1287), .Z(c[1969]) );
  XNOR U1369 ( .A(a[1969]), .B(n1289), .Z(n1287) );
  IV U1370 ( .A(n1285), .Z(n1289) );
  XOR U1371 ( .A(n1290), .B(n1291), .Z(n1285) );
  ANDN U1372 ( .B(n1292), .A(n1293), .Z(n1290) );
  XNOR U1373 ( .A(b[1968]), .B(n1291), .Z(n1292) );
  XNOR U1374 ( .A(b[1968]), .B(n1293), .Z(c[1968]) );
  XNOR U1375 ( .A(a[1968]), .B(n1294), .Z(n1293) );
  IV U1376 ( .A(n1291), .Z(n1294) );
  XOR U1377 ( .A(n1295), .B(n1296), .Z(n1291) );
  ANDN U1378 ( .B(n1297), .A(n1298), .Z(n1295) );
  XNOR U1379 ( .A(b[1967]), .B(n1296), .Z(n1297) );
  XNOR U1380 ( .A(b[1967]), .B(n1298), .Z(c[1967]) );
  XNOR U1381 ( .A(a[1967]), .B(n1299), .Z(n1298) );
  IV U1382 ( .A(n1296), .Z(n1299) );
  XOR U1383 ( .A(n1300), .B(n1301), .Z(n1296) );
  ANDN U1384 ( .B(n1302), .A(n1303), .Z(n1300) );
  XNOR U1385 ( .A(b[1966]), .B(n1301), .Z(n1302) );
  XNOR U1386 ( .A(b[1966]), .B(n1303), .Z(c[1966]) );
  XNOR U1387 ( .A(a[1966]), .B(n1304), .Z(n1303) );
  IV U1388 ( .A(n1301), .Z(n1304) );
  XOR U1389 ( .A(n1305), .B(n1306), .Z(n1301) );
  ANDN U1390 ( .B(n1307), .A(n1308), .Z(n1305) );
  XNOR U1391 ( .A(b[1965]), .B(n1306), .Z(n1307) );
  XNOR U1392 ( .A(b[1965]), .B(n1308), .Z(c[1965]) );
  XNOR U1393 ( .A(a[1965]), .B(n1309), .Z(n1308) );
  IV U1394 ( .A(n1306), .Z(n1309) );
  XOR U1395 ( .A(n1310), .B(n1311), .Z(n1306) );
  ANDN U1396 ( .B(n1312), .A(n1313), .Z(n1310) );
  XNOR U1397 ( .A(b[1964]), .B(n1311), .Z(n1312) );
  XNOR U1398 ( .A(b[1964]), .B(n1313), .Z(c[1964]) );
  XNOR U1399 ( .A(a[1964]), .B(n1314), .Z(n1313) );
  IV U1400 ( .A(n1311), .Z(n1314) );
  XOR U1401 ( .A(n1315), .B(n1316), .Z(n1311) );
  ANDN U1402 ( .B(n1317), .A(n1318), .Z(n1315) );
  XNOR U1403 ( .A(b[1963]), .B(n1316), .Z(n1317) );
  XNOR U1404 ( .A(b[1963]), .B(n1318), .Z(c[1963]) );
  XNOR U1405 ( .A(a[1963]), .B(n1319), .Z(n1318) );
  IV U1406 ( .A(n1316), .Z(n1319) );
  XOR U1407 ( .A(n1320), .B(n1321), .Z(n1316) );
  ANDN U1408 ( .B(n1322), .A(n1323), .Z(n1320) );
  XNOR U1409 ( .A(b[1962]), .B(n1321), .Z(n1322) );
  XNOR U1410 ( .A(b[1962]), .B(n1323), .Z(c[1962]) );
  XNOR U1411 ( .A(a[1962]), .B(n1324), .Z(n1323) );
  IV U1412 ( .A(n1321), .Z(n1324) );
  XOR U1413 ( .A(n1325), .B(n1326), .Z(n1321) );
  ANDN U1414 ( .B(n1327), .A(n1328), .Z(n1325) );
  XNOR U1415 ( .A(b[1961]), .B(n1326), .Z(n1327) );
  XNOR U1416 ( .A(b[1961]), .B(n1328), .Z(c[1961]) );
  XNOR U1417 ( .A(a[1961]), .B(n1329), .Z(n1328) );
  IV U1418 ( .A(n1326), .Z(n1329) );
  XOR U1419 ( .A(n1330), .B(n1331), .Z(n1326) );
  ANDN U1420 ( .B(n1332), .A(n1333), .Z(n1330) );
  XNOR U1421 ( .A(b[1960]), .B(n1331), .Z(n1332) );
  XNOR U1422 ( .A(b[1960]), .B(n1333), .Z(c[1960]) );
  XNOR U1423 ( .A(a[1960]), .B(n1334), .Z(n1333) );
  IV U1424 ( .A(n1331), .Z(n1334) );
  XOR U1425 ( .A(n1335), .B(n1336), .Z(n1331) );
  ANDN U1426 ( .B(n1337), .A(n1338), .Z(n1335) );
  XNOR U1427 ( .A(b[1959]), .B(n1336), .Z(n1337) );
  XNOR U1428 ( .A(b[195]), .B(n1339), .Z(c[195]) );
  XNOR U1429 ( .A(b[1959]), .B(n1338), .Z(c[1959]) );
  XNOR U1430 ( .A(a[1959]), .B(n1340), .Z(n1338) );
  IV U1431 ( .A(n1336), .Z(n1340) );
  XOR U1432 ( .A(n1341), .B(n1342), .Z(n1336) );
  ANDN U1433 ( .B(n1343), .A(n1344), .Z(n1341) );
  XNOR U1434 ( .A(b[1958]), .B(n1342), .Z(n1343) );
  XNOR U1435 ( .A(b[1958]), .B(n1344), .Z(c[1958]) );
  XNOR U1436 ( .A(a[1958]), .B(n1345), .Z(n1344) );
  IV U1437 ( .A(n1342), .Z(n1345) );
  XOR U1438 ( .A(n1346), .B(n1347), .Z(n1342) );
  ANDN U1439 ( .B(n1348), .A(n1349), .Z(n1346) );
  XNOR U1440 ( .A(b[1957]), .B(n1347), .Z(n1348) );
  XNOR U1441 ( .A(b[1957]), .B(n1349), .Z(c[1957]) );
  XNOR U1442 ( .A(a[1957]), .B(n1350), .Z(n1349) );
  IV U1443 ( .A(n1347), .Z(n1350) );
  XOR U1444 ( .A(n1351), .B(n1352), .Z(n1347) );
  ANDN U1445 ( .B(n1353), .A(n1354), .Z(n1351) );
  XNOR U1446 ( .A(b[1956]), .B(n1352), .Z(n1353) );
  XNOR U1447 ( .A(b[1956]), .B(n1354), .Z(c[1956]) );
  XNOR U1448 ( .A(a[1956]), .B(n1355), .Z(n1354) );
  IV U1449 ( .A(n1352), .Z(n1355) );
  XOR U1450 ( .A(n1356), .B(n1357), .Z(n1352) );
  ANDN U1451 ( .B(n1358), .A(n1359), .Z(n1356) );
  XNOR U1452 ( .A(b[1955]), .B(n1357), .Z(n1358) );
  XNOR U1453 ( .A(b[1955]), .B(n1359), .Z(c[1955]) );
  XNOR U1454 ( .A(a[1955]), .B(n1360), .Z(n1359) );
  IV U1455 ( .A(n1357), .Z(n1360) );
  XOR U1456 ( .A(n1361), .B(n1362), .Z(n1357) );
  ANDN U1457 ( .B(n1363), .A(n1364), .Z(n1361) );
  XNOR U1458 ( .A(b[1954]), .B(n1362), .Z(n1363) );
  XNOR U1459 ( .A(b[1954]), .B(n1364), .Z(c[1954]) );
  XNOR U1460 ( .A(a[1954]), .B(n1365), .Z(n1364) );
  IV U1461 ( .A(n1362), .Z(n1365) );
  XOR U1462 ( .A(n1366), .B(n1367), .Z(n1362) );
  ANDN U1463 ( .B(n1368), .A(n1369), .Z(n1366) );
  XNOR U1464 ( .A(b[1953]), .B(n1367), .Z(n1368) );
  XNOR U1465 ( .A(b[1953]), .B(n1369), .Z(c[1953]) );
  XNOR U1466 ( .A(a[1953]), .B(n1370), .Z(n1369) );
  IV U1467 ( .A(n1367), .Z(n1370) );
  XOR U1468 ( .A(n1371), .B(n1372), .Z(n1367) );
  ANDN U1469 ( .B(n1373), .A(n1374), .Z(n1371) );
  XNOR U1470 ( .A(b[1952]), .B(n1372), .Z(n1373) );
  XNOR U1471 ( .A(b[1952]), .B(n1374), .Z(c[1952]) );
  XNOR U1472 ( .A(a[1952]), .B(n1375), .Z(n1374) );
  IV U1473 ( .A(n1372), .Z(n1375) );
  XOR U1474 ( .A(n1376), .B(n1377), .Z(n1372) );
  ANDN U1475 ( .B(n1378), .A(n1379), .Z(n1376) );
  XNOR U1476 ( .A(b[1951]), .B(n1377), .Z(n1378) );
  XNOR U1477 ( .A(b[1951]), .B(n1379), .Z(c[1951]) );
  XNOR U1478 ( .A(a[1951]), .B(n1380), .Z(n1379) );
  IV U1479 ( .A(n1377), .Z(n1380) );
  XOR U1480 ( .A(n1381), .B(n1382), .Z(n1377) );
  ANDN U1481 ( .B(n1383), .A(n1384), .Z(n1381) );
  XNOR U1482 ( .A(b[1950]), .B(n1382), .Z(n1383) );
  XNOR U1483 ( .A(b[1950]), .B(n1384), .Z(c[1950]) );
  XNOR U1484 ( .A(a[1950]), .B(n1385), .Z(n1384) );
  IV U1485 ( .A(n1382), .Z(n1385) );
  XOR U1486 ( .A(n1386), .B(n1387), .Z(n1382) );
  ANDN U1487 ( .B(n1388), .A(n1389), .Z(n1386) );
  XNOR U1488 ( .A(b[1949]), .B(n1387), .Z(n1388) );
  XNOR U1489 ( .A(b[194]), .B(n1390), .Z(c[194]) );
  XNOR U1490 ( .A(b[1949]), .B(n1389), .Z(c[1949]) );
  XNOR U1491 ( .A(a[1949]), .B(n1391), .Z(n1389) );
  IV U1492 ( .A(n1387), .Z(n1391) );
  XOR U1493 ( .A(n1392), .B(n1393), .Z(n1387) );
  ANDN U1494 ( .B(n1394), .A(n1395), .Z(n1392) );
  XNOR U1495 ( .A(b[1948]), .B(n1393), .Z(n1394) );
  XNOR U1496 ( .A(b[1948]), .B(n1395), .Z(c[1948]) );
  XNOR U1497 ( .A(a[1948]), .B(n1396), .Z(n1395) );
  IV U1498 ( .A(n1393), .Z(n1396) );
  XOR U1499 ( .A(n1397), .B(n1398), .Z(n1393) );
  ANDN U1500 ( .B(n1399), .A(n1400), .Z(n1397) );
  XNOR U1501 ( .A(b[1947]), .B(n1398), .Z(n1399) );
  XNOR U1502 ( .A(b[1947]), .B(n1400), .Z(c[1947]) );
  XNOR U1503 ( .A(a[1947]), .B(n1401), .Z(n1400) );
  IV U1504 ( .A(n1398), .Z(n1401) );
  XOR U1505 ( .A(n1402), .B(n1403), .Z(n1398) );
  ANDN U1506 ( .B(n1404), .A(n1405), .Z(n1402) );
  XNOR U1507 ( .A(b[1946]), .B(n1403), .Z(n1404) );
  XNOR U1508 ( .A(b[1946]), .B(n1405), .Z(c[1946]) );
  XNOR U1509 ( .A(a[1946]), .B(n1406), .Z(n1405) );
  IV U1510 ( .A(n1403), .Z(n1406) );
  XOR U1511 ( .A(n1407), .B(n1408), .Z(n1403) );
  ANDN U1512 ( .B(n1409), .A(n1410), .Z(n1407) );
  XNOR U1513 ( .A(b[1945]), .B(n1408), .Z(n1409) );
  XNOR U1514 ( .A(b[1945]), .B(n1410), .Z(c[1945]) );
  XNOR U1515 ( .A(a[1945]), .B(n1411), .Z(n1410) );
  IV U1516 ( .A(n1408), .Z(n1411) );
  XOR U1517 ( .A(n1412), .B(n1413), .Z(n1408) );
  ANDN U1518 ( .B(n1414), .A(n1415), .Z(n1412) );
  XNOR U1519 ( .A(b[1944]), .B(n1413), .Z(n1414) );
  XNOR U1520 ( .A(b[1944]), .B(n1415), .Z(c[1944]) );
  XNOR U1521 ( .A(a[1944]), .B(n1416), .Z(n1415) );
  IV U1522 ( .A(n1413), .Z(n1416) );
  XOR U1523 ( .A(n1417), .B(n1418), .Z(n1413) );
  ANDN U1524 ( .B(n1419), .A(n1420), .Z(n1417) );
  XNOR U1525 ( .A(b[1943]), .B(n1418), .Z(n1419) );
  XNOR U1526 ( .A(b[1943]), .B(n1420), .Z(c[1943]) );
  XNOR U1527 ( .A(a[1943]), .B(n1421), .Z(n1420) );
  IV U1528 ( .A(n1418), .Z(n1421) );
  XOR U1529 ( .A(n1422), .B(n1423), .Z(n1418) );
  ANDN U1530 ( .B(n1424), .A(n1425), .Z(n1422) );
  XNOR U1531 ( .A(b[1942]), .B(n1423), .Z(n1424) );
  XNOR U1532 ( .A(b[1942]), .B(n1425), .Z(c[1942]) );
  XNOR U1533 ( .A(a[1942]), .B(n1426), .Z(n1425) );
  IV U1534 ( .A(n1423), .Z(n1426) );
  XOR U1535 ( .A(n1427), .B(n1428), .Z(n1423) );
  ANDN U1536 ( .B(n1429), .A(n1430), .Z(n1427) );
  XNOR U1537 ( .A(b[1941]), .B(n1428), .Z(n1429) );
  XNOR U1538 ( .A(b[1941]), .B(n1430), .Z(c[1941]) );
  XNOR U1539 ( .A(a[1941]), .B(n1431), .Z(n1430) );
  IV U1540 ( .A(n1428), .Z(n1431) );
  XOR U1541 ( .A(n1432), .B(n1433), .Z(n1428) );
  ANDN U1542 ( .B(n1434), .A(n1435), .Z(n1432) );
  XNOR U1543 ( .A(b[1940]), .B(n1433), .Z(n1434) );
  XNOR U1544 ( .A(b[1940]), .B(n1435), .Z(c[1940]) );
  XNOR U1545 ( .A(a[1940]), .B(n1436), .Z(n1435) );
  IV U1546 ( .A(n1433), .Z(n1436) );
  XOR U1547 ( .A(n1437), .B(n1438), .Z(n1433) );
  ANDN U1548 ( .B(n1439), .A(n1440), .Z(n1437) );
  XNOR U1549 ( .A(b[1939]), .B(n1438), .Z(n1439) );
  XNOR U1550 ( .A(b[193]), .B(n1441), .Z(c[193]) );
  XNOR U1551 ( .A(b[1939]), .B(n1440), .Z(c[1939]) );
  XNOR U1552 ( .A(a[1939]), .B(n1442), .Z(n1440) );
  IV U1553 ( .A(n1438), .Z(n1442) );
  XOR U1554 ( .A(n1443), .B(n1444), .Z(n1438) );
  ANDN U1555 ( .B(n1445), .A(n1446), .Z(n1443) );
  XNOR U1556 ( .A(b[1938]), .B(n1444), .Z(n1445) );
  XNOR U1557 ( .A(b[1938]), .B(n1446), .Z(c[1938]) );
  XNOR U1558 ( .A(a[1938]), .B(n1447), .Z(n1446) );
  IV U1559 ( .A(n1444), .Z(n1447) );
  XOR U1560 ( .A(n1448), .B(n1449), .Z(n1444) );
  ANDN U1561 ( .B(n1450), .A(n1451), .Z(n1448) );
  XNOR U1562 ( .A(b[1937]), .B(n1449), .Z(n1450) );
  XNOR U1563 ( .A(b[1937]), .B(n1451), .Z(c[1937]) );
  XNOR U1564 ( .A(a[1937]), .B(n1452), .Z(n1451) );
  IV U1565 ( .A(n1449), .Z(n1452) );
  XOR U1566 ( .A(n1453), .B(n1454), .Z(n1449) );
  ANDN U1567 ( .B(n1455), .A(n1456), .Z(n1453) );
  XNOR U1568 ( .A(b[1936]), .B(n1454), .Z(n1455) );
  XNOR U1569 ( .A(b[1936]), .B(n1456), .Z(c[1936]) );
  XNOR U1570 ( .A(a[1936]), .B(n1457), .Z(n1456) );
  IV U1571 ( .A(n1454), .Z(n1457) );
  XOR U1572 ( .A(n1458), .B(n1459), .Z(n1454) );
  ANDN U1573 ( .B(n1460), .A(n1461), .Z(n1458) );
  XNOR U1574 ( .A(b[1935]), .B(n1459), .Z(n1460) );
  XNOR U1575 ( .A(b[1935]), .B(n1461), .Z(c[1935]) );
  XNOR U1576 ( .A(a[1935]), .B(n1462), .Z(n1461) );
  IV U1577 ( .A(n1459), .Z(n1462) );
  XOR U1578 ( .A(n1463), .B(n1464), .Z(n1459) );
  ANDN U1579 ( .B(n1465), .A(n1466), .Z(n1463) );
  XNOR U1580 ( .A(b[1934]), .B(n1464), .Z(n1465) );
  XNOR U1581 ( .A(b[1934]), .B(n1466), .Z(c[1934]) );
  XNOR U1582 ( .A(a[1934]), .B(n1467), .Z(n1466) );
  IV U1583 ( .A(n1464), .Z(n1467) );
  XOR U1584 ( .A(n1468), .B(n1469), .Z(n1464) );
  ANDN U1585 ( .B(n1470), .A(n1471), .Z(n1468) );
  XNOR U1586 ( .A(b[1933]), .B(n1469), .Z(n1470) );
  XNOR U1587 ( .A(b[1933]), .B(n1471), .Z(c[1933]) );
  XNOR U1588 ( .A(a[1933]), .B(n1472), .Z(n1471) );
  IV U1589 ( .A(n1469), .Z(n1472) );
  XOR U1590 ( .A(n1473), .B(n1474), .Z(n1469) );
  ANDN U1591 ( .B(n1475), .A(n1476), .Z(n1473) );
  XNOR U1592 ( .A(b[1932]), .B(n1474), .Z(n1475) );
  XNOR U1593 ( .A(b[1932]), .B(n1476), .Z(c[1932]) );
  XNOR U1594 ( .A(a[1932]), .B(n1477), .Z(n1476) );
  IV U1595 ( .A(n1474), .Z(n1477) );
  XOR U1596 ( .A(n1478), .B(n1479), .Z(n1474) );
  ANDN U1597 ( .B(n1480), .A(n1481), .Z(n1478) );
  XNOR U1598 ( .A(b[1931]), .B(n1479), .Z(n1480) );
  XNOR U1599 ( .A(b[1931]), .B(n1481), .Z(c[1931]) );
  XNOR U1600 ( .A(a[1931]), .B(n1482), .Z(n1481) );
  IV U1601 ( .A(n1479), .Z(n1482) );
  XOR U1602 ( .A(n1483), .B(n1484), .Z(n1479) );
  ANDN U1603 ( .B(n1485), .A(n1486), .Z(n1483) );
  XNOR U1604 ( .A(b[1930]), .B(n1484), .Z(n1485) );
  XNOR U1605 ( .A(b[1930]), .B(n1486), .Z(c[1930]) );
  XNOR U1606 ( .A(a[1930]), .B(n1487), .Z(n1486) );
  IV U1607 ( .A(n1484), .Z(n1487) );
  XOR U1608 ( .A(n1488), .B(n1489), .Z(n1484) );
  ANDN U1609 ( .B(n1490), .A(n1491), .Z(n1488) );
  XNOR U1610 ( .A(b[1929]), .B(n1489), .Z(n1490) );
  XNOR U1611 ( .A(b[192]), .B(n1492), .Z(c[192]) );
  XNOR U1612 ( .A(b[1929]), .B(n1491), .Z(c[1929]) );
  XNOR U1613 ( .A(a[1929]), .B(n1493), .Z(n1491) );
  IV U1614 ( .A(n1489), .Z(n1493) );
  XOR U1615 ( .A(n1494), .B(n1495), .Z(n1489) );
  ANDN U1616 ( .B(n1496), .A(n1497), .Z(n1494) );
  XNOR U1617 ( .A(b[1928]), .B(n1495), .Z(n1496) );
  XNOR U1618 ( .A(b[1928]), .B(n1497), .Z(c[1928]) );
  XNOR U1619 ( .A(a[1928]), .B(n1498), .Z(n1497) );
  IV U1620 ( .A(n1495), .Z(n1498) );
  XOR U1621 ( .A(n1499), .B(n1500), .Z(n1495) );
  ANDN U1622 ( .B(n1501), .A(n1502), .Z(n1499) );
  XNOR U1623 ( .A(b[1927]), .B(n1500), .Z(n1501) );
  XNOR U1624 ( .A(b[1927]), .B(n1502), .Z(c[1927]) );
  XNOR U1625 ( .A(a[1927]), .B(n1503), .Z(n1502) );
  IV U1626 ( .A(n1500), .Z(n1503) );
  XOR U1627 ( .A(n1504), .B(n1505), .Z(n1500) );
  ANDN U1628 ( .B(n1506), .A(n1507), .Z(n1504) );
  XNOR U1629 ( .A(b[1926]), .B(n1505), .Z(n1506) );
  XNOR U1630 ( .A(b[1926]), .B(n1507), .Z(c[1926]) );
  XNOR U1631 ( .A(a[1926]), .B(n1508), .Z(n1507) );
  IV U1632 ( .A(n1505), .Z(n1508) );
  XOR U1633 ( .A(n1509), .B(n1510), .Z(n1505) );
  ANDN U1634 ( .B(n1511), .A(n1512), .Z(n1509) );
  XNOR U1635 ( .A(b[1925]), .B(n1510), .Z(n1511) );
  XNOR U1636 ( .A(b[1925]), .B(n1512), .Z(c[1925]) );
  XNOR U1637 ( .A(a[1925]), .B(n1513), .Z(n1512) );
  IV U1638 ( .A(n1510), .Z(n1513) );
  XOR U1639 ( .A(n1514), .B(n1515), .Z(n1510) );
  ANDN U1640 ( .B(n1516), .A(n1517), .Z(n1514) );
  XNOR U1641 ( .A(b[1924]), .B(n1515), .Z(n1516) );
  XNOR U1642 ( .A(b[1924]), .B(n1517), .Z(c[1924]) );
  XNOR U1643 ( .A(a[1924]), .B(n1518), .Z(n1517) );
  IV U1644 ( .A(n1515), .Z(n1518) );
  XOR U1645 ( .A(n1519), .B(n1520), .Z(n1515) );
  ANDN U1646 ( .B(n1521), .A(n1522), .Z(n1519) );
  XNOR U1647 ( .A(b[1923]), .B(n1520), .Z(n1521) );
  XNOR U1648 ( .A(b[1923]), .B(n1522), .Z(c[1923]) );
  XNOR U1649 ( .A(a[1923]), .B(n1523), .Z(n1522) );
  IV U1650 ( .A(n1520), .Z(n1523) );
  XOR U1651 ( .A(n1524), .B(n1525), .Z(n1520) );
  ANDN U1652 ( .B(n1526), .A(n1527), .Z(n1524) );
  XNOR U1653 ( .A(b[1922]), .B(n1525), .Z(n1526) );
  XNOR U1654 ( .A(b[1922]), .B(n1527), .Z(c[1922]) );
  XNOR U1655 ( .A(a[1922]), .B(n1528), .Z(n1527) );
  IV U1656 ( .A(n1525), .Z(n1528) );
  XOR U1657 ( .A(n1529), .B(n1530), .Z(n1525) );
  ANDN U1658 ( .B(n1531), .A(n1532), .Z(n1529) );
  XNOR U1659 ( .A(b[1921]), .B(n1530), .Z(n1531) );
  XNOR U1660 ( .A(b[1921]), .B(n1532), .Z(c[1921]) );
  XNOR U1661 ( .A(a[1921]), .B(n1533), .Z(n1532) );
  IV U1662 ( .A(n1530), .Z(n1533) );
  XOR U1663 ( .A(n1534), .B(n1535), .Z(n1530) );
  ANDN U1664 ( .B(n1536), .A(n1537), .Z(n1534) );
  XNOR U1665 ( .A(b[1920]), .B(n1535), .Z(n1536) );
  XNOR U1666 ( .A(b[1920]), .B(n1537), .Z(c[1920]) );
  XNOR U1667 ( .A(a[1920]), .B(n1538), .Z(n1537) );
  IV U1668 ( .A(n1535), .Z(n1538) );
  XOR U1669 ( .A(n1539), .B(n1540), .Z(n1535) );
  ANDN U1670 ( .B(n1541), .A(n1542), .Z(n1539) );
  XNOR U1671 ( .A(b[1919]), .B(n1540), .Z(n1541) );
  XNOR U1672 ( .A(b[191]), .B(n1543), .Z(c[191]) );
  XNOR U1673 ( .A(b[1919]), .B(n1542), .Z(c[1919]) );
  XNOR U1674 ( .A(a[1919]), .B(n1544), .Z(n1542) );
  IV U1675 ( .A(n1540), .Z(n1544) );
  XOR U1676 ( .A(n1545), .B(n1546), .Z(n1540) );
  ANDN U1677 ( .B(n1547), .A(n1548), .Z(n1545) );
  XNOR U1678 ( .A(b[1918]), .B(n1546), .Z(n1547) );
  XNOR U1679 ( .A(b[1918]), .B(n1548), .Z(c[1918]) );
  XNOR U1680 ( .A(a[1918]), .B(n1549), .Z(n1548) );
  IV U1681 ( .A(n1546), .Z(n1549) );
  XOR U1682 ( .A(n1550), .B(n1551), .Z(n1546) );
  ANDN U1683 ( .B(n1552), .A(n1553), .Z(n1550) );
  XNOR U1684 ( .A(b[1917]), .B(n1551), .Z(n1552) );
  XNOR U1685 ( .A(b[1917]), .B(n1553), .Z(c[1917]) );
  XNOR U1686 ( .A(a[1917]), .B(n1554), .Z(n1553) );
  IV U1687 ( .A(n1551), .Z(n1554) );
  XOR U1688 ( .A(n1555), .B(n1556), .Z(n1551) );
  ANDN U1689 ( .B(n1557), .A(n1558), .Z(n1555) );
  XNOR U1690 ( .A(b[1916]), .B(n1556), .Z(n1557) );
  XNOR U1691 ( .A(b[1916]), .B(n1558), .Z(c[1916]) );
  XNOR U1692 ( .A(a[1916]), .B(n1559), .Z(n1558) );
  IV U1693 ( .A(n1556), .Z(n1559) );
  XOR U1694 ( .A(n1560), .B(n1561), .Z(n1556) );
  ANDN U1695 ( .B(n1562), .A(n1563), .Z(n1560) );
  XNOR U1696 ( .A(b[1915]), .B(n1561), .Z(n1562) );
  XNOR U1697 ( .A(b[1915]), .B(n1563), .Z(c[1915]) );
  XNOR U1698 ( .A(a[1915]), .B(n1564), .Z(n1563) );
  IV U1699 ( .A(n1561), .Z(n1564) );
  XOR U1700 ( .A(n1565), .B(n1566), .Z(n1561) );
  ANDN U1701 ( .B(n1567), .A(n1568), .Z(n1565) );
  XNOR U1702 ( .A(b[1914]), .B(n1566), .Z(n1567) );
  XNOR U1703 ( .A(b[1914]), .B(n1568), .Z(c[1914]) );
  XNOR U1704 ( .A(a[1914]), .B(n1569), .Z(n1568) );
  IV U1705 ( .A(n1566), .Z(n1569) );
  XOR U1706 ( .A(n1570), .B(n1571), .Z(n1566) );
  ANDN U1707 ( .B(n1572), .A(n1573), .Z(n1570) );
  XNOR U1708 ( .A(b[1913]), .B(n1571), .Z(n1572) );
  XNOR U1709 ( .A(b[1913]), .B(n1573), .Z(c[1913]) );
  XNOR U1710 ( .A(a[1913]), .B(n1574), .Z(n1573) );
  IV U1711 ( .A(n1571), .Z(n1574) );
  XOR U1712 ( .A(n1575), .B(n1576), .Z(n1571) );
  ANDN U1713 ( .B(n1577), .A(n1578), .Z(n1575) );
  XNOR U1714 ( .A(b[1912]), .B(n1576), .Z(n1577) );
  XNOR U1715 ( .A(b[1912]), .B(n1578), .Z(c[1912]) );
  XNOR U1716 ( .A(a[1912]), .B(n1579), .Z(n1578) );
  IV U1717 ( .A(n1576), .Z(n1579) );
  XOR U1718 ( .A(n1580), .B(n1581), .Z(n1576) );
  ANDN U1719 ( .B(n1582), .A(n1583), .Z(n1580) );
  XNOR U1720 ( .A(b[1911]), .B(n1581), .Z(n1582) );
  XNOR U1721 ( .A(b[1911]), .B(n1583), .Z(c[1911]) );
  XNOR U1722 ( .A(a[1911]), .B(n1584), .Z(n1583) );
  IV U1723 ( .A(n1581), .Z(n1584) );
  XOR U1724 ( .A(n1585), .B(n1586), .Z(n1581) );
  ANDN U1725 ( .B(n1587), .A(n1588), .Z(n1585) );
  XNOR U1726 ( .A(b[1910]), .B(n1586), .Z(n1587) );
  XNOR U1727 ( .A(b[1910]), .B(n1588), .Z(c[1910]) );
  XNOR U1728 ( .A(a[1910]), .B(n1589), .Z(n1588) );
  IV U1729 ( .A(n1586), .Z(n1589) );
  XOR U1730 ( .A(n1590), .B(n1591), .Z(n1586) );
  ANDN U1731 ( .B(n1592), .A(n1593), .Z(n1590) );
  XNOR U1732 ( .A(b[1909]), .B(n1591), .Z(n1592) );
  XNOR U1733 ( .A(b[190]), .B(n1594), .Z(c[190]) );
  XNOR U1734 ( .A(b[1909]), .B(n1593), .Z(c[1909]) );
  XNOR U1735 ( .A(a[1909]), .B(n1595), .Z(n1593) );
  IV U1736 ( .A(n1591), .Z(n1595) );
  XOR U1737 ( .A(n1596), .B(n1597), .Z(n1591) );
  ANDN U1738 ( .B(n1598), .A(n1599), .Z(n1596) );
  XNOR U1739 ( .A(b[1908]), .B(n1597), .Z(n1598) );
  XNOR U1740 ( .A(b[1908]), .B(n1599), .Z(c[1908]) );
  XNOR U1741 ( .A(a[1908]), .B(n1600), .Z(n1599) );
  IV U1742 ( .A(n1597), .Z(n1600) );
  XOR U1743 ( .A(n1601), .B(n1602), .Z(n1597) );
  ANDN U1744 ( .B(n1603), .A(n1604), .Z(n1601) );
  XNOR U1745 ( .A(b[1907]), .B(n1602), .Z(n1603) );
  XNOR U1746 ( .A(b[1907]), .B(n1604), .Z(c[1907]) );
  XNOR U1747 ( .A(a[1907]), .B(n1605), .Z(n1604) );
  IV U1748 ( .A(n1602), .Z(n1605) );
  XOR U1749 ( .A(n1606), .B(n1607), .Z(n1602) );
  ANDN U1750 ( .B(n1608), .A(n1609), .Z(n1606) );
  XNOR U1751 ( .A(b[1906]), .B(n1607), .Z(n1608) );
  XNOR U1752 ( .A(b[1906]), .B(n1609), .Z(c[1906]) );
  XNOR U1753 ( .A(a[1906]), .B(n1610), .Z(n1609) );
  IV U1754 ( .A(n1607), .Z(n1610) );
  XOR U1755 ( .A(n1611), .B(n1612), .Z(n1607) );
  ANDN U1756 ( .B(n1613), .A(n1614), .Z(n1611) );
  XNOR U1757 ( .A(b[1905]), .B(n1612), .Z(n1613) );
  XNOR U1758 ( .A(b[1905]), .B(n1614), .Z(c[1905]) );
  XNOR U1759 ( .A(a[1905]), .B(n1615), .Z(n1614) );
  IV U1760 ( .A(n1612), .Z(n1615) );
  XOR U1761 ( .A(n1616), .B(n1617), .Z(n1612) );
  ANDN U1762 ( .B(n1618), .A(n1619), .Z(n1616) );
  XNOR U1763 ( .A(b[1904]), .B(n1617), .Z(n1618) );
  XNOR U1764 ( .A(b[1904]), .B(n1619), .Z(c[1904]) );
  XNOR U1765 ( .A(a[1904]), .B(n1620), .Z(n1619) );
  IV U1766 ( .A(n1617), .Z(n1620) );
  XOR U1767 ( .A(n1621), .B(n1622), .Z(n1617) );
  ANDN U1768 ( .B(n1623), .A(n1624), .Z(n1621) );
  XNOR U1769 ( .A(b[1903]), .B(n1622), .Z(n1623) );
  XNOR U1770 ( .A(b[1903]), .B(n1624), .Z(c[1903]) );
  XNOR U1771 ( .A(a[1903]), .B(n1625), .Z(n1624) );
  IV U1772 ( .A(n1622), .Z(n1625) );
  XOR U1773 ( .A(n1626), .B(n1627), .Z(n1622) );
  ANDN U1774 ( .B(n1628), .A(n1629), .Z(n1626) );
  XNOR U1775 ( .A(b[1902]), .B(n1627), .Z(n1628) );
  XNOR U1776 ( .A(b[1902]), .B(n1629), .Z(c[1902]) );
  XNOR U1777 ( .A(a[1902]), .B(n1630), .Z(n1629) );
  IV U1778 ( .A(n1627), .Z(n1630) );
  XOR U1779 ( .A(n1631), .B(n1632), .Z(n1627) );
  ANDN U1780 ( .B(n1633), .A(n1634), .Z(n1631) );
  XNOR U1781 ( .A(b[1901]), .B(n1632), .Z(n1633) );
  XNOR U1782 ( .A(b[1901]), .B(n1634), .Z(c[1901]) );
  XNOR U1783 ( .A(a[1901]), .B(n1635), .Z(n1634) );
  IV U1784 ( .A(n1632), .Z(n1635) );
  XOR U1785 ( .A(n1636), .B(n1637), .Z(n1632) );
  ANDN U1786 ( .B(n1638), .A(n1639), .Z(n1636) );
  XNOR U1787 ( .A(b[1900]), .B(n1637), .Z(n1638) );
  XNOR U1788 ( .A(b[1900]), .B(n1639), .Z(c[1900]) );
  XNOR U1789 ( .A(a[1900]), .B(n1640), .Z(n1639) );
  IV U1790 ( .A(n1637), .Z(n1640) );
  XOR U1791 ( .A(n1641), .B(n1642), .Z(n1637) );
  ANDN U1792 ( .B(n1643), .A(n1644), .Z(n1641) );
  XNOR U1793 ( .A(b[1899]), .B(n1642), .Z(n1643) );
  XNOR U1794 ( .A(b[18]), .B(n1645), .Z(c[18]) );
  XNOR U1795 ( .A(b[189]), .B(n1646), .Z(c[189]) );
  XNOR U1796 ( .A(b[1899]), .B(n1644), .Z(c[1899]) );
  XNOR U1797 ( .A(a[1899]), .B(n1647), .Z(n1644) );
  IV U1798 ( .A(n1642), .Z(n1647) );
  XOR U1799 ( .A(n1648), .B(n1649), .Z(n1642) );
  ANDN U1800 ( .B(n1650), .A(n1651), .Z(n1648) );
  XNOR U1801 ( .A(b[1898]), .B(n1649), .Z(n1650) );
  XNOR U1802 ( .A(b[1898]), .B(n1651), .Z(c[1898]) );
  XNOR U1803 ( .A(a[1898]), .B(n1652), .Z(n1651) );
  IV U1804 ( .A(n1649), .Z(n1652) );
  XOR U1805 ( .A(n1653), .B(n1654), .Z(n1649) );
  ANDN U1806 ( .B(n1655), .A(n1656), .Z(n1653) );
  XNOR U1807 ( .A(b[1897]), .B(n1654), .Z(n1655) );
  XNOR U1808 ( .A(b[1897]), .B(n1656), .Z(c[1897]) );
  XNOR U1809 ( .A(a[1897]), .B(n1657), .Z(n1656) );
  IV U1810 ( .A(n1654), .Z(n1657) );
  XOR U1811 ( .A(n1658), .B(n1659), .Z(n1654) );
  ANDN U1812 ( .B(n1660), .A(n1661), .Z(n1658) );
  XNOR U1813 ( .A(b[1896]), .B(n1659), .Z(n1660) );
  XNOR U1814 ( .A(b[1896]), .B(n1661), .Z(c[1896]) );
  XNOR U1815 ( .A(a[1896]), .B(n1662), .Z(n1661) );
  IV U1816 ( .A(n1659), .Z(n1662) );
  XOR U1817 ( .A(n1663), .B(n1664), .Z(n1659) );
  ANDN U1818 ( .B(n1665), .A(n1666), .Z(n1663) );
  XNOR U1819 ( .A(b[1895]), .B(n1664), .Z(n1665) );
  XNOR U1820 ( .A(b[1895]), .B(n1666), .Z(c[1895]) );
  XNOR U1821 ( .A(a[1895]), .B(n1667), .Z(n1666) );
  IV U1822 ( .A(n1664), .Z(n1667) );
  XOR U1823 ( .A(n1668), .B(n1669), .Z(n1664) );
  ANDN U1824 ( .B(n1670), .A(n1671), .Z(n1668) );
  XNOR U1825 ( .A(b[1894]), .B(n1669), .Z(n1670) );
  XNOR U1826 ( .A(b[1894]), .B(n1671), .Z(c[1894]) );
  XNOR U1827 ( .A(a[1894]), .B(n1672), .Z(n1671) );
  IV U1828 ( .A(n1669), .Z(n1672) );
  XOR U1829 ( .A(n1673), .B(n1674), .Z(n1669) );
  ANDN U1830 ( .B(n1675), .A(n1676), .Z(n1673) );
  XNOR U1831 ( .A(b[1893]), .B(n1674), .Z(n1675) );
  XNOR U1832 ( .A(b[1893]), .B(n1676), .Z(c[1893]) );
  XNOR U1833 ( .A(a[1893]), .B(n1677), .Z(n1676) );
  IV U1834 ( .A(n1674), .Z(n1677) );
  XOR U1835 ( .A(n1678), .B(n1679), .Z(n1674) );
  ANDN U1836 ( .B(n1680), .A(n1681), .Z(n1678) );
  XNOR U1837 ( .A(b[1892]), .B(n1679), .Z(n1680) );
  XNOR U1838 ( .A(b[1892]), .B(n1681), .Z(c[1892]) );
  XNOR U1839 ( .A(a[1892]), .B(n1682), .Z(n1681) );
  IV U1840 ( .A(n1679), .Z(n1682) );
  XOR U1841 ( .A(n1683), .B(n1684), .Z(n1679) );
  ANDN U1842 ( .B(n1685), .A(n1686), .Z(n1683) );
  XNOR U1843 ( .A(b[1891]), .B(n1684), .Z(n1685) );
  XNOR U1844 ( .A(b[1891]), .B(n1686), .Z(c[1891]) );
  XNOR U1845 ( .A(a[1891]), .B(n1687), .Z(n1686) );
  IV U1846 ( .A(n1684), .Z(n1687) );
  XOR U1847 ( .A(n1688), .B(n1689), .Z(n1684) );
  ANDN U1848 ( .B(n1690), .A(n1691), .Z(n1688) );
  XNOR U1849 ( .A(b[1890]), .B(n1689), .Z(n1690) );
  XNOR U1850 ( .A(b[1890]), .B(n1691), .Z(c[1890]) );
  XNOR U1851 ( .A(a[1890]), .B(n1692), .Z(n1691) );
  IV U1852 ( .A(n1689), .Z(n1692) );
  XOR U1853 ( .A(n1693), .B(n1694), .Z(n1689) );
  ANDN U1854 ( .B(n1695), .A(n1696), .Z(n1693) );
  XNOR U1855 ( .A(b[1889]), .B(n1694), .Z(n1695) );
  XNOR U1856 ( .A(b[188]), .B(n1697), .Z(c[188]) );
  XNOR U1857 ( .A(b[1889]), .B(n1696), .Z(c[1889]) );
  XNOR U1858 ( .A(a[1889]), .B(n1698), .Z(n1696) );
  IV U1859 ( .A(n1694), .Z(n1698) );
  XOR U1860 ( .A(n1699), .B(n1700), .Z(n1694) );
  ANDN U1861 ( .B(n1701), .A(n1702), .Z(n1699) );
  XNOR U1862 ( .A(b[1888]), .B(n1700), .Z(n1701) );
  XNOR U1863 ( .A(b[1888]), .B(n1702), .Z(c[1888]) );
  XNOR U1864 ( .A(a[1888]), .B(n1703), .Z(n1702) );
  IV U1865 ( .A(n1700), .Z(n1703) );
  XOR U1866 ( .A(n1704), .B(n1705), .Z(n1700) );
  ANDN U1867 ( .B(n1706), .A(n1707), .Z(n1704) );
  XNOR U1868 ( .A(b[1887]), .B(n1705), .Z(n1706) );
  XNOR U1869 ( .A(b[1887]), .B(n1707), .Z(c[1887]) );
  XNOR U1870 ( .A(a[1887]), .B(n1708), .Z(n1707) );
  IV U1871 ( .A(n1705), .Z(n1708) );
  XOR U1872 ( .A(n1709), .B(n1710), .Z(n1705) );
  ANDN U1873 ( .B(n1711), .A(n1712), .Z(n1709) );
  XNOR U1874 ( .A(b[1886]), .B(n1710), .Z(n1711) );
  XNOR U1875 ( .A(b[1886]), .B(n1712), .Z(c[1886]) );
  XNOR U1876 ( .A(a[1886]), .B(n1713), .Z(n1712) );
  IV U1877 ( .A(n1710), .Z(n1713) );
  XOR U1878 ( .A(n1714), .B(n1715), .Z(n1710) );
  ANDN U1879 ( .B(n1716), .A(n1717), .Z(n1714) );
  XNOR U1880 ( .A(b[1885]), .B(n1715), .Z(n1716) );
  XNOR U1881 ( .A(b[1885]), .B(n1717), .Z(c[1885]) );
  XNOR U1882 ( .A(a[1885]), .B(n1718), .Z(n1717) );
  IV U1883 ( .A(n1715), .Z(n1718) );
  XOR U1884 ( .A(n1719), .B(n1720), .Z(n1715) );
  ANDN U1885 ( .B(n1721), .A(n1722), .Z(n1719) );
  XNOR U1886 ( .A(b[1884]), .B(n1720), .Z(n1721) );
  XNOR U1887 ( .A(b[1884]), .B(n1722), .Z(c[1884]) );
  XNOR U1888 ( .A(a[1884]), .B(n1723), .Z(n1722) );
  IV U1889 ( .A(n1720), .Z(n1723) );
  XOR U1890 ( .A(n1724), .B(n1725), .Z(n1720) );
  ANDN U1891 ( .B(n1726), .A(n1727), .Z(n1724) );
  XNOR U1892 ( .A(b[1883]), .B(n1725), .Z(n1726) );
  XNOR U1893 ( .A(b[1883]), .B(n1727), .Z(c[1883]) );
  XNOR U1894 ( .A(a[1883]), .B(n1728), .Z(n1727) );
  IV U1895 ( .A(n1725), .Z(n1728) );
  XOR U1896 ( .A(n1729), .B(n1730), .Z(n1725) );
  ANDN U1897 ( .B(n1731), .A(n1732), .Z(n1729) );
  XNOR U1898 ( .A(b[1882]), .B(n1730), .Z(n1731) );
  XNOR U1899 ( .A(b[1882]), .B(n1732), .Z(c[1882]) );
  XNOR U1900 ( .A(a[1882]), .B(n1733), .Z(n1732) );
  IV U1901 ( .A(n1730), .Z(n1733) );
  XOR U1902 ( .A(n1734), .B(n1735), .Z(n1730) );
  ANDN U1903 ( .B(n1736), .A(n1737), .Z(n1734) );
  XNOR U1904 ( .A(b[1881]), .B(n1735), .Z(n1736) );
  XNOR U1905 ( .A(b[1881]), .B(n1737), .Z(c[1881]) );
  XNOR U1906 ( .A(a[1881]), .B(n1738), .Z(n1737) );
  IV U1907 ( .A(n1735), .Z(n1738) );
  XOR U1908 ( .A(n1739), .B(n1740), .Z(n1735) );
  ANDN U1909 ( .B(n1741), .A(n1742), .Z(n1739) );
  XNOR U1910 ( .A(b[1880]), .B(n1740), .Z(n1741) );
  XNOR U1911 ( .A(b[1880]), .B(n1742), .Z(c[1880]) );
  XNOR U1912 ( .A(a[1880]), .B(n1743), .Z(n1742) );
  IV U1913 ( .A(n1740), .Z(n1743) );
  XOR U1914 ( .A(n1744), .B(n1745), .Z(n1740) );
  ANDN U1915 ( .B(n1746), .A(n1747), .Z(n1744) );
  XNOR U1916 ( .A(b[1879]), .B(n1745), .Z(n1746) );
  XNOR U1917 ( .A(b[187]), .B(n1748), .Z(c[187]) );
  XNOR U1918 ( .A(b[1879]), .B(n1747), .Z(c[1879]) );
  XNOR U1919 ( .A(a[1879]), .B(n1749), .Z(n1747) );
  IV U1920 ( .A(n1745), .Z(n1749) );
  XOR U1921 ( .A(n1750), .B(n1751), .Z(n1745) );
  ANDN U1922 ( .B(n1752), .A(n1753), .Z(n1750) );
  XNOR U1923 ( .A(b[1878]), .B(n1751), .Z(n1752) );
  XNOR U1924 ( .A(b[1878]), .B(n1753), .Z(c[1878]) );
  XNOR U1925 ( .A(a[1878]), .B(n1754), .Z(n1753) );
  IV U1926 ( .A(n1751), .Z(n1754) );
  XOR U1927 ( .A(n1755), .B(n1756), .Z(n1751) );
  ANDN U1928 ( .B(n1757), .A(n1758), .Z(n1755) );
  XNOR U1929 ( .A(b[1877]), .B(n1756), .Z(n1757) );
  XNOR U1930 ( .A(b[1877]), .B(n1758), .Z(c[1877]) );
  XNOR U1931 ( .A(a[1877]), .B(n1759), .Z(n1758) );
  IV U1932 ( .A(n1756), .Z(n1759) );
  XOR U1933 ( .A(n1760), .B(n1761), .Z(n1756) );
  ANDN U1934 ( .B(n1762), .A(n1763), .Z(n1760) );
  XNOR U1935 ( .A(b[1876]), .B(n1761), .Z(n1762) );
  XNOR U1936 ( .A(b[1876]), .B(n1763), .Z(c[1876]) );
  XNOR U1937 ( .A(a[1876]), .B(n1764), .Z(n1763) );
  IV U1938 ( .A(n1761), .Z(n1764) );
  XOR U1939 ( .A(n1765), .B(n1766), .Z(n1761) );
  ANDN U1940 ( .B(n1767), .A(n1768), .Z(n1765) );
  XNOR U1941 ( .A(b[1875]), .B(n1766), .Z(n1767) );
  XNOR U1942 ( .A(b[1875]), .B(n1768), .Z(c[1875]) );
  XNOR U1943 ( .A(a[1875]), .B(n1769), .Z(n1768) );
  IV U1944 ( .A(n1766), .Z(n1769) );
  XOR U1945 ( .A(n1770), .B(n1771), .Z(n1766) );
  ANDN U1946 ( .B(n1772), .A(n1773), .Z(n1770) );
  XNOR U1947 ( .A(b[1874]), .B(n1771), .Z(n1772) );
  XNOR U1948 ( .A(b[1874]), .B(n1773), .Z(c[1874]) );
  XNOR U1949 ( .A(a[1874]), .B(n1774), .Z(n1773) );
  IV U1950 ( .A(n1771), .Z(n1774) );
  XOR U1951 ( .A(n1775), .B(n1776), .Z(n1771) );
  ANDN U1952 ( .B(n1777), .A(n1778), .Z(n1775) );
  XNOR U1953 ( .A(b[1873]), .B(n1776), .Z(n1777) );
  XNOR U1954 ( .A(b[1873]), .B(n1778), .Z(c[1873]) );
  XNOR U1955 ( .A(a[1873]), .B(n1779), .Z(n1778) );
  IV U1956 ( .A(n1776), .Z(n1779) );
  XOR U1957 ( .A(n1780), .B(n1781), .Z(n1776) );
  ANDN U1958 ( .B(n1782), .A(n1783), .Z(n1780) );
  XNOR U1959 ( .A(b[1872]), .B(n1781), .Z(n1782) );
  XNOR U1960 ( .A(b[1872]), .B(n1783), .Z(c[1872]) );
  XNOR U1961 ( .A(a[1872]), .B(n1784), .Z(n1783) );
  IV U1962 ( .A(n1781), .Z(n1784) );
  XOR U1963 ( .A(n1785), .B(n1786), .Z(n1781) );
  ANDN U1964 ( .B(n1787), .A(n1788), .Z(n1785) );
  XNOR U1965 ( .A(b[1871]), .B(n1786), .Z(n1787) );
  XNOR U1966 ( .A(b[1871]), .B(n1788), .Z(c[1871]) );
  XNOR U1967 ( .A(a[1871]), .B(n1789), .Z(n1788) );
  IV U1968 ( .A(n1786), .Z(n1789) );
  XOR U1969 ( .A(n1790), .B(n1791), .Z(n1786) );
  ANDN U1970 ( .B(n1792), .A(n1793), .Z(n1790) );
  XNOR U1971 ( .A(b[1870]), .B(n1791), .Z(n1792) );
  XNOR U1972 ( .A(b[1870]), .B(n1793), .Z(c[1870]) );
  XNOR U1973 ( .A(a[1870]), .B(n1794), .Z(n1793) );
  IV U1974 ( .A(n1791), .Z(n1794) );
  XOR U1975 ( .A(n1795), .B(n1796), .Z(n1791) );
  ANDN U1976 ( .B(n1797), .A(n1798), .Z(n1795) );
  XNOR U1977 ( .A(b[1869]), .B(n1796), .Z(n1797) );
  XNOR U1978 ( .A(b[186]), .B(n1799), .Z(c[186]) );
  XNOR U1979 ( .A(b[1869]), .B(n1798), .Z(c[1869]) );
  XNOR U1980 ( .A(a[1869]), .B(n1800), .Z(n1798) );
  IV U1981 ( .A(n1796), .Z(n1800) );
  XOR U1982 ( .A(n1801), .B(n1802), .Z(n1796) );
  ANDN U1983 ( .B(n1803), .A(n1804), .Z(n1801) );
  XNOR U1984 ( .A(b[1868]), .B(n1802), .Z(n1803) );
  XNOR U1985 ( .A(b[1868]), .B(n1804), .Z(c[1868]) );
  XNOR U1986 ( .A(a[1868]), .B(n1805), .Z(n1804) );
  IV U1987 ( .A(n1802), .Z(n1805) );
  XOR U1988 ( .A(n1806), .B(n1807), .Z(n1802) );
  ANDN U1989 ( .B(n1808), .A(n1809), .Z(n1806) );
  XNOR U1990 ( .A(b[1867]), .B(n1807), .Z(n1808) );
  XNOR U1991 ( .A(b[1867]), .B(n1809), .Z(c[1867]) );
  XNOR U1992 ( .A(a[1867]), .B(n1810), .Z(n1809) );
  IV U1993 ( .A(n1807), .Z(n1810) );
  XOR U1994 ( .A(n1811), .B(n1812), .Z(n1807) );
  ANDN U1995 ( .B(n1813), .A(n1814), .Z(n1811) );
  XNOR U1996 ( .A(b[1866]), .B(n1812), .Z(n1813) );
  XNOR U1997 ( .A(b[1866]), .B(n1814), .Z(c[1866]) );
  XNOR U1998 ( .A(a[1866]), .B(n1815), .Z(n1814) );
  IV U1999 ( .A(n1812), .Z(n1815) );
  XOR U2000 ( .A(n1816), .B(n1817), .Z(n1812) );
  ANDN U2001 ( .B(n1818), .A(n1819), .Z(n1816) );
  XNOR U2002 ( .A(b[1865]), .B(n1817), .Z(n1818) );
  XNOR U2003 ( .A(b[1865]), .B(n1819), .Z(c[1865]) );
  XNOR U2004 ( .A(a[1865]), .B(n1820), .Z(n1819) );
  IV U2005 ( .A(n1817), .Z(n1820) );
  XOR U2006 ( .A(n1821), .B(n1822), .Z(n1817) );
  ANDN U2007 ( .B(n1823), .A(n1824), .Z(n1821) );
  XNOR U2008 ( .A(b[1864]), .B(n1822), .Z(n1823) );
  XNOR U2009 ( .A(b[1864]), .B(n1824), .Z(c[1864]) );
  XNOR U2010 ( .A(a[1864]), .B(n1825), .Z(n1824) );
  IV U2011 ( .A(n1822), .Z(n1825) );
  XOR U2012 ( .A(n1826), .B(n1827), .Z(n1822) );
  ANDN U2013 ( .B(n1828), .A(n1829), .Z(n1826) );
  XNOR U2014 ( .A(b[1863]), .B(n1827), .Z(n1828) );
  XNOR U2015 ( .A(b[1863]), .B(n1829), .Z(c[1863]) );
  XNOR U2016 ( .A(a[1863]), .B(n1830), .Z(n1829) );
  IV U2017 ( .A(n1827), .Z(n1830) );
  XOR U2018 ( .A(n1831), .B(n1832), .Z(n1827) );
  ANDN U2019 ( .B(n1833), .A(n1834), .Z(n1831) );
  XNOR U2020 ( .A(b[1862]), .B(n1832), .Z(n1833) );
  XNOR U2021 ( .A(b[1862]), .B(n1834), .Z(c[1862]) );
  XNOR U2022 ( .A(a[1862]), .B(n1835), .Z(n1834) );
  IV U2023 ( .A(n1832), .Z(n1835) );
  XOR U2024 ( .A(n1836), .B(n1837), .Z(n1832) );
  ANDN U2025 ( .B(n1838), .A(n1839), .Z(n1836) );
  XNOR U2026 ( .A(b[1861]), .B(n1837), .Z(n1838) );
  XNOR U2027 ( .A(b[1861]), .B(n1839), .Z(c[1861]) );
  XNOR U2028 ( .A(a[1861]), .B(n1840), .Z(n1839) );
  IV U2029 ( .A(n1837), .Z(n1840) );
  XOR U2030 ( .A(n1841), .B(n1842), .Z(n1837) );
  ANDN U2031 ( .B(n1843), .A(n1844), .Z(n1841) );
  XNOR U2032 ( .A(b[1860]), .B(n1842), .Z(n1843) );
  XNOR U2033 ( .A(b[1860]), .B(n1844), .Z(c[1860]) );
  XNOR U2034 ( .A(a[1860]), .B(n1845), .Z(n1844) );
  IV U2035 ( .A(n1842), .Z(n1845) );
  XOR U2036 ( .A(n1846), .B(n1847), .Z(n1842) );
  ANDN U2037 ( .B(n1848), .A(n1849), .Z(n1846) );
  XNOR U2038 ( .A(b[1859]), .B(n1847), .Z(n1848) );
  XNOR U2039 ( .A(b[185]), .B(n1850), .Z(c[185]) );
  XNOR U2040 ( .A(b[1859]), .B(n1849), .Z(c[1859]) );
  XNOR U2041 ( .A(a[1859]), .B(n1851), .Z(n1849) );
  IV U2042 ( .A(n1847), .Z(n1851) );
  XOR U2043 ( .A(n1852), .B(n1853), .Z(n1847) );
  ANDN U2044 ( .B(n1854), .A(n1855), .Z(n1852) );
  XNOR U2045 ( .A(b[1858]), .B(n1853), .Z(n1854) );
  XNOR U2046 ( .A(b[1858]), .B(n1855), .Z(c[1858]) );
  XNOR U2047 ( .A(a[1858]), .B(n1856), .Z(n1855) );
  IV U2048 ( .A(n1853), .Z(n1856) );
  XOR U2049 ( .A(n1857), .B(n1858), .Z(n1853) );
  ANDN U2050 ( .B(n1859), .A(n1860), .Z(n1857) );
  XNOR U2051 ( .A(b[1857]), .B(n1858), .Z(n1859) );
  XNOR U2052 ( .A(b[1857]), .B(n1860), .Z(c[1857]) );
  XNOR U2053 ( .A(a[1857]), .B(n1861), .Z(n1860) );
  IV U2054 ( .A(n1858), .Z(n1861) );
  XOR U2055 ( .A(n1862), .B(n1863), .Z(n1858) );
  ANDN U2056 ( .B(n1864), .A(n1865), .Z(n1862) );
  XNOR U2057 ( .A(b[1856]), .B(n1863), .Z(n1864) );
  XNOR U2058 ( .A(b[1856]), .B(n1865), .Z(c[1856]) );
  XNOR U2059 ( .A(a[1856]), .B(n1866), .Z(n1865) );
  IV U2060 ( .A(n1863), .Z(n1866) );
  XOR U2061 ( .A(n1867), .B(n1868), .Z(n1863) );
  ANDN U2062 ( .B(n1869), .A(n1870), .Z(n1867) );
  XNOR U2063 ( .A(b[1855]), .B(n1868), .Z(n1869) );
  XNOR U2064 ( .A(b[1855]), .B(n1870), .Z(c[1855]) );
  XNOR U2065 ( .A(a[1855]), .B(n1871), .Z(n1870) );
  IV U2066 ( .A(n1868), .Z(n1871) );
  XOR U2067 ( .A(n1872), .B(n1873), .Z(n1868) );
  ANDN U2068 ( .B(n1874), .A(n1875), .Z(n1872) );
  XNOR U2069 ( .A(b[1854]), .B(n1873), .Z(n1874) );
  XNOR U2070 ( .A(b[1854]), .B(n1875), .Z(c[1854]) );
  XNOR U2071 ( .A(a[1854]), .B(n1876), .Z(n1875) );
  IV U2072 ( .A(n1873), .Z(n1876) );
  XOR U2073 ( .A(n1877), .B(n1878), .Z(n1873) );
  ANDN U2074 ( .B(n1879), .A(n1880), .Z(n1877) );
  XNOR U2075 ( .A(b[1853]), .B(n1878), .Z(n1879) );
  XNOR U2076 ( .A(b[1853]), .B(n1880), .Z(c[1853]) );
  XNOR U2077 ( .A(a[1853]), .B(n1881), .Z(n1880) );
  IV U2078 ( .A(n1878), .Z(n1881) );
  XOR U2079 ( .A(n1882), .B(n1883), .Z(n1878) );
  ANDN U2080 ( .B(n1884), .A(n1885), .Z(n1882) );
  XNOR U2081 ( .A(b[1852]), .B(n1883), .Z(n1884) );
  XNOR U2082 ( .A(b[1852]), .B(n1885), .Z(c[1852]) );
  XNOR U2083 ( .A(a[1852]), .B(n1886), .Z(n1885) );
  IV U2084 ( .A(n1883), .Z(n1886) );
  XOR U2085 ( .A(n1887), .B(n1888), .Z(n1883) );
  ANDN U2086 ( .B(n1889), .A(n1890), .Z(n1887) );
  XNOR U2087 ( .A(b[1851]), .B(n1888), .Z(n1889) );
  XNOR U2088 ( .A(b[1851]), .B(n1890), .Z(c[1851]) );
  XNOR U2089 ( .A(a[1851]), .B(n1891), .Z(n1890) );
  IV U2090 ( .A(n1888), .Z(n1891) );
  XOR U2091 ( .A(n1892), .B(n1893), .Z(n1888) );
  ANDN U2092 ( .B(n1894), .A(n1895), .Z(n1892) );
  XNOR U2093 ( .A(b[1850]), .B(n1893), .Z(n1894) );
  XNOR U2094 ( .A(b[1850]), .B(n1895), .Z(c[1850]) );
  XNOR U2095 ( .A(a[1850]), .B(n1896), .Z(n1895) );
  IV U2096 ( .A(n1893), .Z(n1896) );
  XOR U2097 ( .A(n1897), .B(n1898), .Z(n1893) );
  ANDN U2098 ( .B(n1899), .A(n1900), .Z(n1897) );
  XNOR U2099 ( .A(b[1849]), .B(n1898), .Z(n1899) );
  XNOR U2100 ( .A(b[184]), .B(n1901), .Z(c[184]) );
  XNOR U2101 ( .A(b[1849]), .B(n1900), .Z(c[1849]) );
  XNOR U2102 ( .A(a[1849]), .B(n1902), .Z(n1900) );
  IV U2103 ( .A(n1898), .Z(n1902) );
  XOR U2104 ( .A(n1903), .B(n1904), .Z(n1898) );
  ANDN U2105 ( .B(n1905), .A(n1906), .Z(n1903) );
  XNOR U2106 ( .A(b[1848]), .B(n1904), .Z(n1905) );
  XNOR U2107 ( .A(b[1848]), .B(n1906), .Z(c[1848]) );
  XNOR U2108 ( .A(a[1848]), .B(n1907), .Z(n1906) );
  IV U2109 ( .A(n1904), .Z(n1907) );
  XOR U2110 ( .A(n1908), .B(n1909), .Z(n1904) );
  ANDN U2111 ( .B(n1910), .A(n1911), .Z(n1908) );
  XNOR U2112 ( .A(b[1847]), .B(n1909), .Z(n1910) );
  XNOR U2113 ( .A(b[1847]), .B(n1911), .Z(c[1847]) );
  XNOR U2114 ( .A(a[1847]), .B(n1912), .Z(n1911) );
  IV U2115 ( .A(n1909), .Z(n1912) );
  XOR U2116 ( .A(n1913), .B(n1914), .Z(n1909) );
  ANDN U2117 ( .B(n1915), .A(n1916), .Z(n1913) );
  XNOR U2118 ( .A(b[1846]), .B(n1914), .Z(n1915) );
  XNOR U2119 ( .A(b[1846]), .B(n1916), .Z(c[1846]) );
  XNOR U2120 ( .A(a[1846]), .B(n1917), .Z(n1916) );
  IV U2121 ( .A(n1914), .Z(n1917) );
  XOR U2122 ( .A(n1918), .B(n1919), .Z(n1914) );
  ANDN U2123 ( .B(n1920), .A(n1921), .Z(n1918) );
  XNOR U2124 ( .A(b[1845]), .B(n1919), .Z(n1920) );
  XNOR U2125 ( .A(b[1845]), .B(n1921), .Z(c[1845]) );
  XNOR U2126 ( .A(a[1845]), .B(n1922), .Z(n1921) );
  IV U2127 ( .A(n1919), .Z(n1922) );
  XOR U2128 ( .A(n1923), .B(n1924), .Z(n1919) );
  ANDN U2129 ( .B(n1925), .A(n1926), .Z(n1923) );
  XNOR U2130 ( .A(b[1844]), .B(n1924), .Z(n1925) );
  XNOR U2131 ( .A(b[1844]), .B(n1926), .Z(c[1844]) );
  XNOR U2132 ( .A(a[1844]), .B(n1927), .Z(n1926) );
  IV U2133 ( .A(n1924), .Z(n1927) );
  XOR U2134 ( .A(n1928), .B(n1929), .Z(n1924) );
  ANDN U2135 ( .B(n1930), .A(n1931), .Z(n1928) );
  XNOR U2136 ( .A(b[1843]), .B(n1929), .Z(n1930) );
  XNOR U2137 ( .A(b[1843]), .B(n1931), .Z(c[1843]) );
  XNOR U2138 ( .A(a[1843]), .B(n1932), .Z(n1931) );
  IV U2139 ( .A(n1929), .Z(n1932) );
  XOR U2140 ( .A(n1933), .B(n1934), .Z(n1929) );
  ANDN U2141 ( .B(n1935), .A(n1936), .Z(n1933) );
  XNOR U2142 ( .A(b[1842]), .B(n1934), .Z(n1935) );
  XNOR U2143 ( .A(b[1842]), .B(n1936), .Z(c[1842]) );
  XNOR U2144 ( .A(a[1842]), .B(n1937), .Z(n1936) );
  IV U2145 ( .A(n1934), .Z(n1937) );
  XOR U2146 ( .A(n1938), .B(n1939), .Z(n1934) );
  ANDN U2147 ( .B(n1940), .A(n1941), .Z(n1938) );
  XNOR U2148 ( .A(b[1841]), .B(n1939), .Z(n1940) );
  XNOR U2149 ( .A(b[1841]), .B(n1941), .Z(c[1841]) );
  XNOR U2150 ( .A(a[1841]), .B(n1942), .Z(n1941) );
  IV U2151 ( .A(n1939), .Z(n1942) );
  XOR U2152 ( .A(n1943), .B(n1944), .Z(n1939) );
  ANDN U2153 ( .B(n1945), .A(n1946), .Z(n1943) );
  XNOR U2154 ( .A(b[1840]), .B(n1944), .Z(n1945) );
  XNOR U2155 ( .A(b[1840]), .B(n1946), .Z(c[1840]) );
  XNOR U2156 ( .A(a[1840]), .B(n1947), .Z(n1946) );
  IV U2157 ( .A(n1944), .Z(n1947) );
  XOR U2158 ( .A(n1948), .B(n1949), .Z(n1944) );
  ANDN U2159 ( .B(n1950), .A(n1951), .Z(n1948) );
  XNOR U2160 ( .A(b[1839]), .B(n1949), .Z(n1950) );
  XNOR U2161 ( .A(b[183]), .B(n1952), .Z(c[183]) );
  XNOR U2162 ( .A(b[1839]), .B(n1951), .Z(c[1839]) );
  XNOR U2163 ( .A(a[1839]), .B(n1953), .Z(n1951) );
  IV U2164 ( .A(n1949), .Z(n1953) );
  XOR U2165 ( .A(n1954), .B(n1955), .Z(n1949) );
  ANDN U2166 ( .B(n1956), .A(n1957), .Z(n1954) );
  XNOR U2167 ( .A(b[1838]), .B(n1955), .Z(n1956) );
  XNOR U2168 ( .A(b[1838]), .B(n1957), .Z(c[1838]) );
  XNOR U2169 ( .A(a[1838]), .B(n1958), .Z(n1957) );
  IV U2170 ( .A(n1955), .Z(n1958) );
  XOR U2171 ( .A(n1959), .B(n1960), .Z(n1955) );
  ANDN U2172 ( .B(n1961), .A(n1962), .Z(n1959) );
  XNOR U2173 ( .A(b[1837]), .B(n1960), .Z(n1961) );
  XNOR U2174 ( .A(b[1837]), .B(n1962), .Z(c[1837]) );
  XNOR U2175 ( .A(a[1837]), .B(n1963), .Z(n1962) );
  IV U2176 ( .A(n1960), .Z(n1963) );
  XOR U2177 ( .A(n1964), .B(n1965), .Z(n1960) );
  ANDN U2178 ( .B(n1966), .A(n1967), .Z(n1964) );
  XNOR U2179 ( .A(b[1836]), .B(n1965), .Z(n1966) );
  XNOR U2180 ( .A(b[1836]), .B(n1967), .Z(c[1836]) );
  XNOR U2181 ( .A(a[1836]), .B(n1968), .Z(n1967) );
  IV U2182 ( .A(n1965), .Z(n1968) );
  XOR U2183 ( .A(n1969), .B(n1970), .Z(n1965) );
  ANDN U2184 ( .B(n1971), .A(n1972), .Z(n1969) );
  XNOR U2185 ( .A(b[1835]), .B(n1970), .Z(n1971) );
  XNOR U2186 ( .A(b[1835]), .B(n1972), .Z(c[1835]) );
  XNOR U2187 ( .A(a[1835]), .B(n1973), .Z(n1972) );
  IV U2188 ( .A(n1970), .Z(n1973) );
  XOR U2189 ( .A(n1974), .B(n1975), .Z(n1970) );
  ANDN U2190 ( .B(n1976), .A(n1977), .Z(n1974) );
  XNOR U2191 ( .A(b[1834]), .B(n1975), .Z(n1976) );
  XNOR U2192 ( .A(b[1834]), .B(n1977), .Z(c[1834]) );
  XNOR U2193 ( .A(a[1834]), .B(n1978), .Z(n1977) );
  IV U2194 ( .A(n1975), .Z(n1978) );
  XOR U2195 ( .A(n1979), .B(n1980), .Z(n1975) );
  ANDN U2196 ( .B(n1981), .A(n1982), .Z(n1979) );
  XNOR U2197 ( .A(b[1833]), .B(n1980), .Z(n1981) );
  XNOR U2198 ( .A(b[1833]), .B(n1982), .Z(c[1833]) );
  XNOR U2199 ( .A(a[1833]), .B(n1983), .Z(n1982) );
  IV U2200 ( .A(n1980), .Z(n1983) );
  XOR U2201 ( .A(n1984), .B(n1985), .Z(n1980) );
  ANDN U2202 ( .B(n1986), .A(n1987), .Z(n1984) );
  XNOR U2203 ( .A(b[1832]), .B(n1985), .Z(n1986) );
  XNOR U2204 ( .A(b[1832]), .B(n1987), .Z(c[1832]) );
  XNOR U2205 ( .A(a[1832]), .B(n1988), .Z(n1987) );
  IV U2206 ( .A(n1985), .Z(n1988) );
  XOR U2207 ( .A(n1989), .B(n1990), .Z(n1985) );
  ANDN U2208 ( .B(n1991), .A(n1992), .Z(n1989) );
  XNOR U2209 ( .A(b[1831]), .B(n1990), .Z(n1991) );
  XNOR U2210 ( .A(b[1831]), .B(n1992), .Z(c[1831]) );
  XNOR U2211 ( .A(a[1831]), .B(n1993), .Z(n1992) );
  IV U2212 ( .A(n1990), .Z(n1993) );
  XOR U2213 ( .A(n1994), .B(n1995), .Z(n1990) );
  ANDN U2214 ( .B(n1996), .A(n1997), .Z(n1994) );
  XNOR U2215 ( .A(b[1830]), .B(n1995), .Z(n1996) );
  XNOR U2216 ( .A(b[1830]), .B(n1997), .Z(c[1830]) );
  XNOR U2217 ( .A(a[1830]), .B(n1998), .Z(n1997) );
  IV U2218 ( .A(n1995), .Z(n1998) );
  XOR U2219 ( .A(n1999), .B(n2000), .Z(n1995) );
  ANDN U2220 ( .B(n2001), .A(n2002), .Z(n1999) );
  XNOR U2221 ( .A(b[1829]), .B(n2000), .Z(n2001) );
  XNOR U2222 ( .A(b[182]), .B(n2003), .Z(c[182]) );
  XNOR U2223 ( .A(b[1829]), .B(n2002), .Z(c[1829]) );
  XNOR U2224 ( .A(a[1829]), .B(n2004), .Z(n2002) );
  IV U2225 ( .A(n2000), .Z(n2004) );
  XOR U2226 ( .A(n2005), .B(n2006), .Z(n2000) );
  ANDN U2227 ( .B(n2007), .A(n2008), .Z(n2005) );
  XNOR U2228 ( .A(b[1828]), .B(n2006), .Z(n2007) );
  XNOR U2229 ( .A(b[1828]), .B(n2008), .Z(c[1828]) );
  XNOR U2230 ( .A(a[1828]), .B(n2009), .Z(n2008) );
  IV U2231 ( .A(n2006), .Z(n2009) );
  XOR U2232 ( .A(n2010), .B(n2011), .Z(n2006) );
  ANDN U2233 ( .B(n2012), .A(n2013), .Z(n2010) );
  XNOR U2234 ( .A(b[1827]), .B(n2011), .Z(n2012) );
  XNOR U2235 ( .A(b[1827]), .B(n2013), .Z(c[1827]) );
  XNOR U2236 ( .A(a[1827]), .B(n2014), .Z(n2013) );
  IV U2237 ( .A(n2011), .Z(n2014) );
  XOR U2238 ( .A(n2015), .B(n2016), .Z(n2011) );
  ANDN U2239 ( .B(n2017), .A(n2018), .Z(n2015) );
  XNOR U2240 ( .A(b[1826]), .B(n2016), .Z(n2017) );
  XNOR U2241 ( .A(b[1826]), .B(n2018), .Z(c[1826]) );
  XNOR U2242 ( .A(a[1826]), .B(n2019), .Z(n2018) );
  IV U2243 ( .A(n2016), .Z(n2019) );
  XOR U2244 ( .A(n2020), .B(n2021), .Z(n2016) );
  ANDN U2245 ( .B(n2022), .A(n2023), .Z(n2020) );
  XNOR U2246 ( .A(b[1825]), .B(n2021), .Z(n2022) );
  XNOR U2247 ( .A(b[1825]), .B(n2023), .Z(c[1825]) );
  XNOR U2248 ( .A(a[1825]), .B(n2024), .Z(n2023) );
  IV U2249 ( .A(n2021), .Z(n2024) );
  XOR U2250 ( .A(n2025), .B(n2026), .Z(n2021) );
  ANDN U2251 ( .B(n2027), .A(n2028), .Z(n2025) );
  XNOR U2252 ( .A(b[1824]), .B(n2026), .Z(n2027) );
  XNOR U2253 ( .A(b[1824]), .B(n2028), .Z(c[1824]) );
  XNOR U2254 ( .A(a[1824]), .B(n2029), .Z(n2028) );
  IV U2255 ( .A(n2026), .Z(n2029) );
  XOR U2256 ( .A(n2030), .B(n2031), .Z(n2026) );
  ANDN U2257 ( .B(n2032), .A(n2033), .Z(n2030) );
  XNOR U2258 ( .A(b[1823]), .B(n2031), .Z(n2032) );
  XNOR U2259 ( .A(b[1823]), .B(n2033), .Z(c[1823]) );
  XNOR U2260 ( .A(a[1823]), .B(n2034), .Z(n2033) );
  IV U2261 ( .A(n2031), .Z(n2034) );
  XOR U2262 ( .A(n2035), .B(n2036), .Z(n2031) );
  ANDN U2263 ( .B(n2037), .A(n2038), .Z(n2035) );
  XNOR U2264 ( .A(b[1822]), .B(n2036), .Z(n2037) );
  XNOR U2265 ( .A(b[1822]), .B(n2038), .Z(c[1822]) );
  XNOR U2266 ( .A(a[1822]), .B(n2039), .Z(n2038) );
  IV U2267 ( .A(n2036), .Z(n2039) );
  XOR U2268 ( .A(n2040), .B(n2041), .Z(n2036) );
  ANDN U2269 ( .B(n2042), .A(n2043), .Z(n2040) );
  XNOR U2270 ( .A(b[1821]), .B(n2041), .Z(n2042) );
  XNOR U2271 ( .A(b[1821]), .B(n2043), .Z(c[1821]) );
  XNOR U2272 ( .A(a[1821]), .B(n2044), .Z(n2043) );
  IV U2273 ( .A(n2041), .Z(n2044) );
  XOR U2274 ( .A(n2045), .B(n2046), .Z(n2041) );
  ANDN U2275 ( .B(n2047), .A(n2048), .Z(n2045) );
  XNOR U2276 ( .A(b[1820]), .B(n2046), .Z(n2047) );
  XNOR U2277 ( .A(b[1820]), .B(n2048), .Z(c[1820]) );
  XNOR U2278 ( .A(a[1820]), .B(n2049), .Z(n2048) );
  IV U2279 ( .A(n2046), .Z(n2049) );
  XOR U2280 ( .A(n2050), .B(n2051), .Z(n2046) );
  ANDN U2281 ( .B(n2052), .A(n2053), .Z(n2050) );
  XNOR U2282 ( .A(b[1819]), .B(n2051), .Z(n2052) );
  XNOR U2283 ( .A(b[181]), .B(n2054), .Z(c[181]) );
  XNOR U2284 ( .A(b[1819]), .B(n2053), .Z(c[1819]) );
  XNOR U2285 ( .A(a[1819]), .B(n2055), .Z(n2053) );
  IV U2286 ( .A(n2051), .Z(n2055) );
  XOR U2287 ( .A(n2056), .B(n2057), .Z(n2051) );
  ANDN U2288 ( .B(n2058), .A(n2059), .Z(n2056) );
  XNOR U2289 ( .A(b[1818]), .B(n2057), .Z(n2058) );
  XNOR U2290 ( .A(b[1818]), .B(n2059), .Z(c[1818]) );
  XNOR U2291 ( .A(a[1818]), .B(n2060), .Z(n2059) );
  IV U2292 ( .A(n2057), .Z(n2060) );
  XOR U2293 ( .A(n2061), .B(n2062), .Z(n2057) );
  ANDN U2294 ( .B(n2063), .A(n2064), .Z(n2061) );
  XNOR U2295 ( .A(b[1817]), .B(n2062), .Z(n2063) );
  XNOR U2296 ( .A(b[1817]), .B(n2064), .Z(c[1817]) );
  XNOR U2297 ( .A(a[1817]), .B(n2065), .Z(n2064) );
  IV U2298 ( .A(n2062), .Z(n2065) );
  XOR U2299 ( .A(n2066), .B(n2067), .Z(n2062) );
  ANDN U2300 ( .B(n2068), .A(n2069), .Z(n2066) );
  XNOR U2301 ( .A(b[1816]), .B(n2067), .Z(n2068) );
  XNOR U2302 ( .A(b[1816]), .B(n2069), .Z(c[1816]) );
  XNOR U2303 ( .A(a[1816]), .B(n2070), .Z(n2069) );
  IV U2304 ( .A(n2067), .Z(n2070) );
  XOR U2305 ( .A(n2071), .B(n2072), .Z(n2067) );
  ANDN U2306 ( .B(n2073), .A(n2074), .Z(n2071) );
  XNOR U2307 ( .A(b[1815]), .B(n2072), .Z(n2073) );
  XNOR U2308 ( .A(b[1815]), .B(n2074), .Z(c[1815]) );
  XNOR U2309 ( .A(a[1815]), .B(n2075), .Z(n2074) );
  IV U2310 ( .A(n2072), .Z(n2075) );
  XOR U2311 ( .A(n2076), .B(n2077), .Z(n2072) );
  ANDN U2312 ( .B(n2078), .A(n2079), .Z(n2076) );
  XNOR U2313 ( .A(b[1814]), .B(n2077), .Z(n2078) );
  XNOR U2314 ( .A(b[1814]), .B(n2079), .Z(c[1814]) );
  XNOR U2315 ( .A(a[1814]), .B(n2080), .Z(n2079) );
  IV U2316 ( .A(n2077), .Z(n2080) );
  XOR U2317 ( .A(n2081), .B(n2082), .Z(n2077) );
  ANDN U2318 ( .B(n2083), .A(n2084), .Z(n2081) );
  XNOR U2319 ( .A(b[1813]), .B(n2082), .Z(n2083) );
  XNOR U2320 ( .A(b[1813]), .B(n2084), .Z(c[1813]) );
  XNOR U2321 ( .A(a[1813]), .B(n2085), .Z(n2084) );
  IV U2322 ( .A(n2082), .Z(n2085) );
  XOR U2323 ( .A(n2086), .B(n2087), .Z(n2082) );
  ANDN U2324 ( .B(n2088), .A(n2089), .Z(n2086) );
  XNOR U2325 ( .A(b[1812]), .B(n2087), .Z(n2088) );
  XNOR U2326 ( .A(b[1812]), .B(n2089), .Z(c[1812]) );
  XNOR U2327 ( .A(a[1812]), .B(n2090), .Z(n2089) );
  IV U2328 ( .A(n2087), .Z(n2090) );
  XOR U2329 ( .A(n2091), .B(n2092), .Z(n2087) );
  ANDN U2330 ( .B(n2093), .A(n2094), .Z(n2091) );
  XNOR U2331 ( .A(b[1811]), .B(n2092), .Z(n2093) );
  XNOR U2332 ( .A(b[1811]), .B(n2094), .Z(c[1811]) );
  XNOR U2333 ( .A(a[1811]), .B(n2095), .Z(n2094) );
  IV U2334 ( .A(n2092), .Z(n2095) );
  XOR U2335 ( .A(n2096), .B(n2097), .Z(n2092) );
  ANDN U2336 ( .B(n2098), .A(n2099), .Z(n2096) );
  XNOR U2337 ( .A(b[1810]), .B(n2097), .Z(n2098) );
  XNOR U2338 ( .A(b[1810]), .B(n2099), .Z(c[1810]) );
  XNOR U2339 ( .A(a[1810]), .B(n2100), .Z(n2099) );
  IV U2340 ( .A(n2097), .Z(n2100) );
  XOR U2341 ( .A(n2101), .B(n2102), .Z(n2097) );
  ANDN U2342 ( .B(n2103), .A(n2104), .Z(n2101) );
  XNOR U2343 ( .A(b[1809]), .B(n2102), .Z(n2103) );
  XNOR U2344 ( .A(b[180]), .B(n2105), .Z(c[180]) );
  XNOR U2345 ( .A(b[1809]), .B(n2104), .Z(c[1809]) );
  XNOR U2346 ( .A(a[1809]), .B(n2106), .Z(n2104) );
  IV U2347 ( .A(n2102), .Z(n2106) );
  XOR U2348 ( .A(n2107), .B(n2108), .Z(n2102) );
  ANDN U2349 ( .B(n2109), .A(n2110), .Z(n2107) );
  XNOR U2350 ( .A(b[1808]), .B(n2108), .Z(n2109) );
  XNOR U2351 ( .A(b[1808]), .B(n2110), .Z(c[1808]) );
  XNOR U2352 ( .A(a[1808]), .B(n2111), .Z(n2110) );
  IV U2353 ( .A(n2108), .Z(n2111) );
  XOR U2354 ( .A(n2112), .B(n2113), .Z(n2108) );
  ANDN U2355 ( .B(n2114), .A(n2115), .Z(n2112) );
  XNOR U2356 ( .A(b[1807]), .B(n2113), .Z(n2114) );
  XNOR U2357 ( .A(b[1807]), .B(n2115), .Z(c[1807]) );
  XNOR U2358 ( .A(a[1807]), .B(n2116), .Z(n2115) );
  IV U2359 ( .A(n2113), .Z(n2116) );
  XOR U2360 ( .A(n2117), .B(n2118), .Z(n2113) );
  ANDN U2361 ( .B(n2119), .A(n2120), .Z(n2117) );
  XNOR U2362 ( .A(b[1806]), .B(n2118), .Z(n2119) );
  XNOR U2363 ( .A(b[1806]), .B(n2120), .Z(c[1806]) );
  XNOR U2364 ( .A(a[1806]), .B(n2121), .Z(n2120) );
  IV U2365 ( .A(n2118), .Z(n2121) );
  XOR U2366 ( .A(n2122), .B(n2123), .Z(n2118) );
  ANDN U2367 ( .B(n2124), .A(n2125), .Z(n2122) );
  XNOR U2368 ( .A(b[1805]), .B(n2123), .Z(n2124) );
  XNOR U2369 ( .A(b[1805]), .B(n2125), .Z(c[1805]) );
  XNOR U2370 ( .A(a[1805]), .B(n2126), .Z(n2125) );
  IV U2371 ( .A(n2123), .Z(n2126) );
  XOR U2372 ( .A(n2127), .B(n2128), .Z(n2123) );
  ANDN U2373 ( .B(n2129), .A(n2130), .Z(n2127) );
  XNOR U2374 ( .A(b[1804]), .B(n2128), .Z(n2129) );
  XNOR U2375 ( .A(b[1804]), .B(n2130), .Z(c[1804]) );
  XNOR U2376 ( .A(a[1804]), .B(n2131), .Z(n2130) );
  IV U2377 ( .A(n2128), .Z(n2131) );
  XOR U2378 ( .A(n2132), .B(n2133), .Z(n2128) );
  ANDN U2379 ( .B(n2134), .A(n2135), .Z(n2132) );
  XNOR U2380 ( .A(b[1803]), .B(n2133), .Z(n2134) );
  XNOR U2381 ( .A(b[1803]), .B(n2135), .Z(c[1803]) );
  XNOR U2382 ( .A(a[1803]), .B(n2136), .Z(n2135) );
  IV U2383 ( .A(n2133), .Z(n2136) );
  XOR U2384 ( .A(n2137), .B(n2138), .Z(n2133) );
  ANDN U2385 ( .B(n2139), .A(n2140), .Z(n2137) );
  XNOR U2386 ( .A(b[1802]), .B(n2138), .Z(n2139) );
  XNOR U2387 ( .A(b[1802]), .B(n2140), .Z(c[1802]) );
  XNOR U2388 ( .A(a[1802]), .B(n2141), .Z(n2140) );
  IV U2389 ( .A(n2138), .Z(n2141) );
  XOR U2390 ( .A(n2142), .B(n2143), .Z(n2138) );
  ANDN U2391 ( .B(n2144), .A(n2145), .Z(n2142) );
  XNOR U2392 ( .A(b[1801]), .B(n2143), .Z(n2144) );
  XNOR U2393 ( .A(b[1801]), .B(n2145), .Z(c[1801]) );
  XNOR U2394 ( .A(a[1801]), .B(n2146), .Z(n2145) );
  IV U2395 ( .A(n2143), .Z(n2146) );
  XOR U2396 ( .A(n2147), .B(n2148), .Z(n2143) );
  ANDN U2397 ( .B(n2149), .A(n2150), .Z(n2147) );
  XNOR U2398 ( .A(b[1800]), .B(n2148), .Z(n2149) );
  XNOR U2399 ( .A(b[1800]), .B(n2150), .Z(c[1800]) );
  XNOR U2400 ( .A(a[1800]), .B(n2151), .Z(n2150) );
  IV U2401 ( .A(n2148), .Z(n2151) );
  XOR U2402 ( .A(n2152), .B(n2153), .Z(n2148) );
  ANDN U2403 ( .B(n2154), .A(n2155), .Z(n2152) );
  XNOR U2404 ( .A(b[1799]), .B(n2153), .Z(n2154) );
  XNOR U2405 ( .A(b[17]), .B(n2156), .Z(c[17]) );
  XNOR U2406 ( .A(b[179]), .B(n2157), .Z(c[179]) );
  XNOR U2407 ( .A(b[1799]), .B(n2155), .Z(c[1799]) );
  XNOR U2408 ( .A(a[1799]), .B(n2158), .Z(n2155) );
  IV U2409 ( .A(n2153), .Z(n2158) );
  XOR U2410 ( .A(n2159), .B(n2160), .Z(n2153) );
  ANDN U2411 ( .B(n2161), .A(n2162), .Z(n2159) );
  XNOR U2412 ( .A(b[1798]), .B(n2160), .Z(n2161) );
  XNOR U2413 ( .A(b[1798]), .B(n2162), .Z(c[1798]) );
  XNOR U2414 ( .A(a[1798]), .B(n2163), .Z(n2162) );
  IV U2415 ( .A(n2160), .Z(n2163) );
  XOR U2416 ( .A(n2164), .B(n2165), .Z(n2160) );
  ANDN U2417 ( .B(n2166), .A(n2167), .Z(n2164) );
  XNOR U2418 ( .A(b[1797]), .B(n2165), .Z(n2166) );
  XNOR U2419 ( .A(b[1797]), .B(n2167), .Z(c[1797]) );
  XNOR U2420 ( .A(a[1797]), .B(n2168), .Z(n2167) );
  IV U2421 ( .A(n2165), .Z(n2168) );
  XOR U2422 ( .A(n2169), .B(n2170), .Z(n2165) );
  ANDN U2423 ( .B(n2171), .A(n2172), .Z(n2169) );
  XNOR U2424 ( .A(b[1796]), .B(n2170), .Z(n2171) );
  XNOR U2425 ( .A(b[1796]), .B(n2172), .Z(c[1796]) );
  XNOR U2426 ( .A(a[1796]), .B(n2173), .Z(n2172) );
  IV U2427 ( .A(n2170), .Z(n2173) );
  XOR U2428 ( .A(n2174), .B(n2175), .Z(n2170) );
  ANDN U2429 ( .B(n2176), .A(n2177), .Z(n2174) );
  XNOR U2430 ( .A(b[1795]), .B(n2175), .Z(n2176) );
  XNOR U2431 ( .A(b[1795]), .B(n2177), .Z(c[1795]) );
  XNOR U2432 ( .A(a[1795]), .B(n2178), .Z(n2177) );
  IV U2433 ( .A(n2175), .Z(n2178) );
  XOR U2434 ( .A(n2179), .B(n2180), .Z(n2175) );
  ANDN U2435 ( .B(n2181), .A(n2182), .Z(n2179) );
  XNOR U2436 ( .A(b[1794]), .B(n2180), .Z(n2181) );
  XNOR U2437 ( .A(b[1794]), .B(n2182), .Z(c[1794]) );
  XNOR U2438 ( .A(a[1794]), .B(n2183), .Z(n2182) );
  IV U2439 ( .A(n2180), .Z(n2183) );
  XOR U2440 ( .A(n2184), .B(n2185), .Z(n2180) );
  ANDN U2441 ( .B(n2186), .A(n2187), .Z(n2184) );
  XNOR U2442 ( .A(b[1793]), .B(n2185), .Z(n2186) );
  XNOR U2443 ( .A(b[1793]), .B(n2187), .Z(c[1793]) );
  XNOR U2444 ( .A(a[1793]), .B(n2188), .Z(n2187) );
  IV U2445 ( .A(n2185), .Z(n2188) );
  XOR U2446 ( .A(n2189), .B(n2190), .Z(n2185) );
  ANDN U2447 ( .B(n2191), .A(n2192), .Z(n2189) );
  XNOR U2448 ( .A(b[1792]), .B(n2190), .Z(n2191) );
  XNOR U2449 ( .A(b[1792]), .B(n2192), .Z(c[1792]) );
  XNOR U2450 ( .A(a[1792]), .B(n2193), .Z(n2192) );
  IV U2451 ( .A(n2190), .Z(n2193) );
  XOR U2452 ( .A(n2194), .B(n2195), .Z(n2190) );
  ANDN U2453 ( .B(n2196), .A(n2197), .Z(n2194) );
  XNOR U2454 ( .A(b[1791]), .B(n2195), .Z(n2196) );
  XNOR U2455 ( .A(b[1791]), .B(n2197), .Z(c[1791]) );
  XNOR U2456 ( .A(a[1791]), .B(n2198), .Z(n2197) );
  IV U2457 ( .A(n2195), .Z(n2198) );
  XOR U2458 ( .A(n2199), .B(n2200), .Z(n2195) );
  ANDN U2459 ( .B(n2201), .A(n2202), .Z(n2199) );
  XNOR U2460 ( .A(b[1790]), .B(n2200), .Z(n2201) );
  XNOR U2461 ( .A(b[1790]), .B(n2202), .Z(c[1790]) );
  XNOR U2462 ( .A(a[1790]), .B(n2203), .Z(n2202) );
  IV U2463 ( .A(n2200), .Z(n2203) );
  XOR U2464 ( .A(n2204), .B(n2205), .Z(n2200) );
  ANDN U2465 ( .B(n2206), .A(n2207), .Z(n2204) );
  XNOR U2466 ( .A(b[1789]), .B(n2205), .Z(n2206) );
  XNOR U2467 ( .A(b[178]), .B(n2208), .Z(c[178]) );
  XNOR U2468 ( .A(b[1789]), .B(n2207), .Z(c[1789]) );
  XNOR U2469 ( .A(a[1789]), .B(n2209), .Z(n2207) );
  IV U2470 ( .A(n2205), .Z(n2209) );
  XOR U2471 ( .A(n2210), .B(n2211), .Z(n2205) );
  ANDN U2472 ( .B(n2212), .A(n2213), .Z(n2210) );
  XNOR U2473 ( .A(b[1788]), .B(n2211), .Z(n2212) );
  XNOR U2474 ( .A(b[1788]), .B(n2213), .Z(c[1788]) );
  XNOR U2475 ( .A(a[1788]), .B(n2214), .Z(n2213) );
  IV U2476 ( .A(n2211), .Z(n2214) );
  XOR U2477 ( .A(n2215), .B(n2216), .Z(n2211) );
  ANDN U2478 ( .B(n2217), .A(n2218), .Z(n2215) );
  XNOR U2479 ( .A(b[1787]), .B(n2216), .Z(n2217) );
  XNOR U2480 ( .A(b[1787]), .B(n2218), .Z(c[1787]) );
  XNOR U2481 ( .A(a[1787]), .B(n2219), .Z(n2218) );
  IV U2482 ( .A(n2216), .Z(n2219) );
  XOR U2483 ( .A(n2220), .B(n2221), .Z(n2216) );
  ANDN U2484 ( .B(n2222), .A(n2223), .Z(n2220) );
  XNOR U2485 ( .A(b[1786]), .B(n2221), .Z(n2222) );
  XNOR U2486 ( .A(b[1786]), .B(n2223), .Z(c[1786]) );
  XNOR U2487 ( .A(a[1786]), .B(n2224), .Z(n2223) );
  IV U2488 ( .A(n2221), .Z(n2224) );
  XOR U2489 ( .A(n2225), .B(n2226), .Z(n2221) );
  ANDN U2490 ( .B(n2227), .A(n2228), .Z(n2225) );
  XNOR U2491 ( .A(b[1785]), .B(n2226), .Z(n2227) );
  XNOR U2492 ( .A(b[1785]), .B(n2228), .Z(c[1785]) );
  XNOR U2493 ( .A(a[1785]), .B(n2229), .Z(n2228) );
  IV U2494 ( .A(n2226), .Z(n2229) );
  XOR U2495 ( .A(n2230), .B(n2231), .Z(n2226) );
  ANDN U2496 ( .B(n2232), .A(n2233), .Z(n2230) );
  XNOR U2497 ( .A(b[1784]), .B(n2231), .Z(n2232) );
  XNOR U2498 ( .A(b[1784]), .B(n2233), .Z(c[1784]) );
  XNOR U2499 ( .A(a[1784]), .B(n2234), .Z(n2233) );
  IV U2500 ( .A(n2231), .Z(n2234) );
  XOR U2501 ( .A(n2235), .B(n2236), .Z(n2231) );
  ANDN U2502 ( .B(n2237), .A(n2238), .Z(n2235) );
  XNOR U2503 ( .A(b[1783]), .B(n2236), .Z(n2237) );
  XNOR U2504 ( .A(b[1783]), .B(n2238), .Z(c[1783]) );
  XNOR U2505 ( .A(a[1783]), .B(n2239), .Z(n2238) );
  IV U2506 ( .A(n2236), .Z(n2239) );
  XOR U2507 ( .A(n2240), .B(n2241), .Z(n2236) );
  ANDN U2508 ( .B(n2242), .A(n2243), .Z(n2240) );
  XNOR U2509 ( .A(b[1782]), .B(n2241), .Z(n2242) );
  XNOR U2510 ( .A(b[1782]), .B(n2243), .Z(c[1782]) );
  XNOR U2511 ( .A(a[1782]), .B(n2244), .Z(n2243) );
  IV U2512 ( .A(n2241), .Z(n2244) );
  XOR U2513 ( .A(n2245), .B(n2246), .Z(n2241) );
  ANDN U2514 ( .B(n2247), .A(n2248), .Z(n2245) );
  XNOR U2515 ( .A(b[1781]), .B(n2246), .Z(n2247) );
  XNOR U2516 ( .A(b[1781]), .B(n2248), .Z(c[1781]) );
  XNOR U2517 ( .A(a[1781]), .B(n2249), .Z(n2248) );
  IV U2518 ( .A(n2246), .Z(n2249) );
  XOR U2519 ( .A(n2250), .B(n2251), .Z(n2246) );
  ANDN U2520 ( .B(n2252), .A(n2253), .Z(n2250) );
  XNOR U2521 ( .A(b[1780]), .B(n2251), .Z(n2252) );
  XNOR U2522 ( .A(b[1780]), .B(n2253), .Z(c[1780]) );
  XNOR U2523 ( .A(a[1780]), .B(n2254), .Z(n2253) );
  IV U2524 ( .A(n2251), .Z(n2254) );
  XOR U2525 ( .A(n2255), .B(n2256), .Z(n2251) );
  ANDN U2526 ( .B(n2257), .A(n2258), .Z(n2255) );
  XNOR U2527 ( .A(b[1779]), .B(n2256), .Z(n2257) );
  XNOR U2528 ( .A(b[177]), .B(n2259), .Z(c[177]) );
  XNOR U2529 ( .A(b[1779]), .B(n2258), .Z(c[1779]) );
  XNOR U2530 ( .A(a[1779]), .B(n2260), .Z(n2258) );
  IV U2531 ( .A(n2256), .Z(n2260) );
  XOR U2532 ( .A(n2261), .B(n2262), .Z(n2256) );
  ANDN U2533 ( .B(n2263), .A(n2264), .Z(n2261) );
  XNOR U2534 ( .A(b[1778]), .B(n2262), .Z(n2263) );
  XNOR U2535 ( .A(b[1778]), .B(n2264), .Z(c[1778]) );
  XNOR U2536 ( .A(a[1778]), .B(n2265), .Z(n2264) );
  IV U2537 ( .A(n2262), .Z(n2265) );
  XOR U2538 ( .A(n2266), .B(n2267), .Z(n2262) );
  ANDN U2539 ( .B(n2268), .A(n2269), .Z(n2266) );
  XNOR U2540 ( .A(b[1777]), .B(n2267), .Z(n2268) );
  XNOR U2541 ( .A(b[1777]), .B(n2269), .Z(c[1777]) );
  XNOR U2542 ( .A(a[1777]), .B(n2270), .Z(n2269) );
  IV U2543 ( .A(n2267), .Z(n2270) );
  XOR U2544 ( .A(n2271), .B(n2272), .Z(n2267) );
  ANDN U2545 ( .B(n2273), .A(n2274), .Z(n2271) );
  XNOR U2546 ( .A(b[1776]), .B(n2272), .Z(n2273) );
  XNOR U2547 ( .A(b[1776]), .B(n2274), .Z(c[1776]) );
  XNOR U2548 ( .A(a[1776]), .B(n2275), .Z(n2274) );
  IV U2549 ( .A(n2272), .Z(n2275) );
  XOR U2550 ( .A(n2276), .B(n2277), .Z(n2272) );
  ANDN U2551 ( .B(n2278), .A(n2279), .Z(n2276) );
  XNOR U2552 ( .A(b[1775]), .B(n2277), .Z(n2278) );
  XNOR U2553 ( .A(b[1775]), .B(n2279), .Z(c[1775]) );
  XNOR U2554 ( .A(a[1775]), .B(n2280), .Z(n2279) );
  IV U2555 ( .A(n2277), .Z(n2280) );
  XOR U2556 ( .A(n2281), .B(n2282), .Z(n2277) );
  ANDN U2557 ( .B(n2283), .A(n2284), .Z(n2281) );
  XNOR U2558 ( .A(b[1774]), .B(n2282), .Z(n2283) );
  XNOR U2559 ( .A(b[1774]), .B(n2284), .Z(c[1774]) );
  XNOR U2560 ( .A(a[1774]), .B(n2285), .Z(n2284) );
  IV U2561 ( .A(n2282), .Z(n2285) );
  XOR U2562 ( .A(n2286), .B(n2287), .Z(n2282) );
  ANDN U2563 ( .B(n2288), .A(n2289), .Z(n2286) );
  XNOR U2564 ( .A(b[1773]), .B(n2287), .Z(n2288) );
  XNOR U2565 ( .A(b[1773]), .B(n2289), .Z(c[1773]) );
  XNOR U2566 ( .A(a[1773]), .B(n2290), .Z(n2289) );
  IV U2567 ( .A(n2287), .Z(n2290) );
  XOR U2568 ( .A(n2291), .B(n2292), .Z(n2287) );
  ANDN U2569 ( .B(n2293), .A(n2294), .Z(n2291) );
  XNOR U2570 ( .A(b[1772]), .B(n2292), .Z(n2293) );
  XNOR U2571 ( .A(b[1772]), .B(n2294), .Z(c[1772]) );
  XNOR U2572 ( .A(a[1772]), .B(n2295), .Z(n2294) );
  IV U2573 ( .A(n2292), .Z(n2295) );
  XOR U2574 ( .A(n2296), .B(n2297), .Z(n2292) );
  ANDN U2575 ( .B(n2298), .A(n2299), .Z(n2296) );
  XNOR U2576 ( .A(b[1771]), .B(n2297), .Z(n2298) );
  XNOR U2577 ( .A(b[1771]), .B(n2299), .Z(c[1771]) );
  XNOR U2578 ( .A(a[1771]), .B(n2300), .Z(n2299) );
  IV U2579 ( .A(n2297), .Z(n2300) );
  XOR U2580 ( .A(n2301), .B(n2302), .Z(n2297) );
  ANDN U2581 ( .B(n2303), .A(n2304), .Z(n2301) );
  XNOR U2582 ( .A(b[1770]), .B(n2302), .Z(n2303) );
  XNOR U2583 ( .A(b[1770]), .B(n2304), .Z(c[1770]) );
  XNOR U2584 ( .A(a[1770]), .B(n2305), .Z(n2304) );
  IV U2585 ( .A(n2302), .Z(n2305) );
  XOR U2586 ( .A(n2306), .B(n2307), .Z(n2302) );
  ANDN U2587 ( .B(n2308), .A(n2309), .Z(n2306) );
  XNOR U2588 ( .A(b[1769]), .B(n2307), .Z(n2308) );
  XNOR U2589 ( .A(b[176]), .B(n2310), .Z(c[176]) );
  XNOR U2590 ( .A(b[1769]), .B(n2309), .Z(c[1769]) );
  XNOR U2591 ( .A(a[1769]), .B(n2311), .Z(n2309) );
  IV U2592 ( .A(n2307), .Z(n2311) );
  XOR U2593 ( .A(n2312), .B(n2313), .Z(n2307) );
  ANDN U2594 ( .B(n2314), .A(n2315), .Z(n2312) );
  XNOR U2595 ( .A(b[1768]), .B(n2313), .Z(n2314) );
  XNOR U2596 ( .A(b[1768]), .B(n2315), .Z(c[1768]) );
  XNOR U2597 ( .A(a[1768]), .B(n2316), .Z(n2315) );
  IV U2598 ( .A(n2313), .Z(n2316) );
  XOR U2599 ( .A(n2317), .B(n2318), .Z(n2313) );
  ANDN U2600 ( .B(n2319), .A(n2320), .Z(n2317) );
  XNOR U2601 ( .A(b[1767]), .B(n2318), .Z(n2319) );
  XNOR U2602 ( .A(b[1767]), .B(n2320), .Z(c[1767]) );
  XNOR U2603 ( .A(a[1767]), .B(n2321), .Z(n2320) );
  IV U2604 ( .A(n2318), .Z(n2321) );
  XOR U2605 ( .A(n2322), .B(n2323), .Z(n2318) );
  ANDN U2606 ( .B(n2324), .A(n2325), .Z(n2322) );
  XNOR U2607 ( .A(b[1766]), .B(n2323), .Z(n2324) );
  XNOR U2608 ( .A(b[1766]), .B(n2325), .Z(c[1766]) );
  XNOR U2609 ( .A(a[1766]), .B(n2326), .Z(n2325) );
  IV U2610 ( .A(n2323), .Z(n2326) );
  XOR U2611 ( .A(n2327), .B(n2328), .Z(n2323) );
  ANDN U2612 ( .B(n2329), .A(n2330), .Z(n2327) );
  XNOR U2613 ( .A(b[1765]), .B(n2328), .Z(n2329) );
  XNOR U2614 ( .A(b[1765]), .B(n2330), .Z(c[1765]) );
  XNOR U2615 ( .A(a[1765]), .B(n2331), .Z(n2330) );
  IV U2616 ( .A(n2328), .Z(n2331) );
  XOR U2617 ( .A(n2332), .B(n2333), .Z(n2328) );
  ANDN U2618 ( .B(n2334), .A(n2335), .Z(n2332) );
  XNOR U2619 ( .A(b[1764]), .B(n2333), .Z(n2334) );
  XNOR U2620 ( .A(b[1764]), .B(n2335), .Z(c[1764]) );
  XNOR U2621 ( .A(a[1764]), .B(n2336), .Z(n2335) );
  IV U2622 ( .A(n2333), .Z(n2336) );
  XOR U2623 ( .A(n2337), .B(n2338), .Z(n2333) );
  ANDN U2624 ( .B(n2339), .A(n2340), .Z(n2337) );
  XNOR U2625 ( .A(b[1763]), .B(n2338), .Z(n2339) );
  XNOR U2626 ( .A(b[1763]), .B(n2340), .Z(c[1763]) );
  XNOR U2627 ( .A(a[1763]), .B(n2341), .Z(n2340) );
  IV U2628 ( .A(n2338), .Z(n2341) );
  XOR U2629 ( .A(n2342), .B(n2343), .Z(n2338) );
  ANDN U2630 ( .B(n2344), .A(n2345), .Z(n2342) );
  XNOR U2631 ( .A(b[1762]), .B(n2343), .Z(n2344) );
  XNOR U2632 ( .A(b[1762]), .B(n2345), .Z(c[1762]) );
  XNOR U2633 ( .A(a[1762]), .B(n2346), .Z(n2345) );
  IV U2634 ( .A(n2343), .Z(n2346) );
  XOR U2635 ( .A(n2347), .B(n2348), .Z(n2343) );
  ANDN U2636 ( .B(n2349), .A(n2350), .Z(n2347) );
  XNOR U2637 ( .A(b[1761]), .B(n2348), .Z(n2349) );
  XNOR U2638 ( .A(b[1761]), .B(n2350), .Z(c[1761]) );
  XNOR U2639 ( .A(a[1761]), .B(n2351), .Z(n2350) );
  IV U2640 ( .A(n2348), .Z(n2351) );
  XOR U2641 ( .A(n2352), .B(n2353), .Z(n2348) );
  ANDN U2642 ( .B(n2354), .A(n2355), .Z(n2352) );
  XNOR U2643 ( .A(b[1760]), .B(n2353), .Z(n2354) );
  XNOR U2644 ( .A(b[1760]), .B(n2355), .Z(c[1760]) );
  XNOR U2645 ( .A(a[1760]), .B(n2356), .Z(n2355) );
  IV U2646 ( .A(n2353), .Z(n2356) );
  XOR U2647 ( .A(n2357), .B(n2358), .Z(n2353) );
  ANDN U2648 ( .B(n2359), .A(n2360), .Z(n2357) );
  XNOR U2649 ( .A(b[1759]), .B(n2358), .Z(n2359) );
  XNOR U2650 ( .A(b[175]), .B(n2361), .Z(c[175]) );
  XNOR U2651 ( .A(b[1759]), .B(n2360), .Z(c[1759]) );
  XNOR U2652 ( .A(a[1759]), .B(n2362), .Z(n2360) );
  IV U2653 ( .A(n2358), .Z(n2362) );
  XOR U2654 ( .A(n2363), .B(n2364), .Z(n2358) );
  ANDN U2655 ( .B(n2365), .A(n2366), .Z(n2363) );
  XNOR U2656 ( .A(b[1758]), .B(n2364), .Z(n2365) );
  XNOR U2657 ( .A(b[1758]), .B(n2366), .Z(c[1758]) );
  XNOR U2658 ( .A(a[1758]), .B(n2367), .Z(n2366) );
  IV U2659 ( .A(n2364), .Z(n2367) );
  XOR U2660 ( .A(n2368), .B(n2369), .Z(n2364) );
  ANDN U2661 ( .B(n2370), .A(n2371), .Z(n2368) );
  XNOR U2662 ( .A(b[1757]), .B(n2369), .Z(n2370) );
  XNOR U2663 ( .A(b[1757]), .B(n2371), .Z(c[1757]) );
  XNOR U2664 ( .A(a[1757]), .B(n2372), .Z(n2371) );
  IV U2665 ( .A(n2369), .Z(n2372) );
  XOR U2666 ( .A(n2373), .B(n2374), .Z(n2369) );
  ANDN U2667 ( .B(n2375), .A(n2376), .Z(n2373) );
  XNOR U2668 ( .A(b[1756]), .B(n2374), .Z(n2375) );
  XNOR U2669 ( .A(b[1756]), .B(n2376), .Z(c[1756]) );
  XNOR U2670 ( .A(a[1756]), .B(n2377), .Z(n2376) );
  IV U2671 ( .A(n2374), .Z(n2377) );
  XOR U2672 ( .A(n2378), .B(n2379), .Z(n2374) );
  ANDN U2673 ( .B(n2380), .A(n2381), .Z(n2378) );
  XNOR U2674 ( .A(b[1755]), .B(n2379), .Z(n2380) );
  XNOR U2675 ( .A(b[1755]), .B(n2381), .Z(c[1755]) );
  XNOR U2676 ( .A(a[1755]), .B(n2382), .Z(n2381) );
  IV U2677 ( .A(n2379), .Z(n2382) );
  XOR U2678 ( .A(n2383), .B(n2384), .Z(n2379) );
  ANDN U2679 ( .B(n2385), .A(n2386), .Z(n2383) );
  XNOR U2680 ( .A(b[1754]), .B(n2384), .Z(n2385) );
  XNOR U2681 ( .A(b[1754]), .B(n2386), .Z(c[1754]) );
  XNOR U2682 ( .A(a[1754]), .B(n2387), .Z(n2386) );
  IV U2683 ( .A(n2384), .Z(n2387) );
  XOR U2684 ( .A(n2388), .B(n2389), .Z(n2384) );
  ANDN U2685 ( .B(n2390), .A(n2391), .Z(n2388) );
  XNOR U2686 ( .A(b[1753]), .B(n2389), .Z(n2390) );
  XNOR U2687 ( .A(b[1753]), .B(n2391), .Z(c[1753]) );
  XNOR U2688 ( .A(a[1753]), .B(n2392), .Z(n2391) );
  IV U2689 ( .A(n2389), .Z(n2392) );
  XOR U2690 ( .A(n2393), .B(n2394), .Z(n2389) );
  ANDN U2691 ( .B(n2395), .A(n2396), .Z(n2393) );
  XNOR U2692 ( .A(b[1752]), .B(n2394), .Z(n2395) );
  XNOR U2693 ( .A(b[1752]), .B(n2396), .Z(c[1752]) );
  XNOR U2694 ( .A(a[1752]), .B(n2397), .Z(n2396) );
  IV U2695 ( .A(n2394), .Z(n2397) );
  XOR U2696 ( .A(n2398), .B(n2399), .Z(n2394) );
  ANDN U2697 ( .B(n2400), .A(n2401), .Z(n2398) );
  XNOR U2698 ( .A(b[1751]), .B(n2399), .Z(n2400) );
  XNOR U2699 ( .A(b[1751]), .B(n2401), .Z(c[1751]) );
  XNOR U2700 ( .A(a[1751]), .B(n2402), .Z(n2401) );
  IV U2701 ( .A(n2399), .Z(n2402) );
  XOR U2702 ( .A(n2403), .B(n2404), .Z(n2399) );
  ANDN U2703 ( .B(n2405), .A(n2406), .Z(n2403) );
  XNOR U2704 ( .A(b[1750]), .B(n2404), .Z(n2405) );
  XNOR U2705 ( .A(b[1750]), .B(n2406), .Z(c[1750]) );
  XNOR U2706 ( .A(a[1750]), .B(n2407), .Z(n2406) );
  IV U2707 ( .A(n2404), .Z(n2407) );
  XOR U2708 ( .A(n2408), .B(n2409), .Z(n2404) );
  ANDN U2709 ( .B(n2410), .A(n2411), .Z(n2408) );
  XNOR U2710 ( .A(b[1749]), .B(n2409), .Z(n2410) );
  XNOR U2711 ( .A(b[174]), .B(n2412), .Z(c[174]) );
  XNOR U2712 ( .A(b[1749]), .B(n2411), .Z(c[1749]) );
  XNOR U2713 ( .A(a[1749]), .B(n2413), .Z(n2411) );
  IV U2714 ( .A(n2409), .Z(n2413) );
  XOR U2715 ( .A(n2414), .B(n2415), .Z(n2409) );
  ANDN U2716 ( .B(n2416), .A(n2417), .Z(n2414) );
  XNOR U2717 ( .A(b[1748]), .B(n2415), .Z(n2416) );
  XNOR U2718 ( .A(b[1748]), .B(n2417), .Z(c[1748]) );
  XNOR U2719 ( .A(a[1748]), .B(n2418), .Z(n2417) );
  IV U2720 ( .A(n2415), .Z(n2418) );
  XOR U2721 ( .A(n2419), .B(n2420), .Z(n2415) );
  ANDN U2722 ( .B(n2421), .A(n2422), .Z(n2419) );
  XNOR U2723 ( .A(b[1747]), .B(n2420), .Z(n2421) );
  XNOR U2724 ( .A(b[1747]), .B(n2422), .Z(c[1747]) );
  XNOR U2725 ( .A(a[1747]), .B(n2423), .Z(n2422) );
  IV U2726 ( .A(n2420), .Z(n2423) );
  XOR U2727 ( .A(n2424), .B(n2425), .Z(n2420) );
  ANDN U2728 ( .B(n2426), .A(n2427), .Z(n2424) );
  XNOR U2729 ( .A(b[1746]), .B(n2425), .Z(n2426) );
  XNOR U2730 ( .A(b[1746]), .B(n2427), .Z(c[1746]) );
  XNOR U2731 ( .A(a[1746]), .B(n2428), .Z(n2427) );
  IV U2732 ( .A(n2425), .Z(n2428) );
  XOR U2733 ( .A(n2429), .B(n2430), .Z(n2425) );
  ANDN U2734 ( .B(n2431), .A(n2432), .Z(n2429) );
  XNOR U2735 ( .A(b[1745]), .B(n2430), .Z(n2431) );
  XNOR U2736 ( .A(b[1745]), .B(n2432), .Z(c[1745]) );
  XNOR U2737 ( .A(a[1745]), .B(n2433), .Z(n2432) );
  IV U2738 ( .A(n2430), .Z(n2433) );
  XOR U2739 ( .A(n2434), .B(n2435), .Z(n2430) );
  ANDN U2740 ( .B(n2436), .A(n2437), .Z(n2434) );
  XNOR U2741 ( .A(b[1744]), .B(n2435), .Z(n2436) );
  XNOR U2742 ( .A(b[1744]), .B(n2437), .Z(c[1744]) );
  XNOR U2743 ( .A(a[1744]), .B(n2438), .Z(n2437) );
  IV U2744 ( .A(n2435), .Z(n2438) );
  XOR U2745 ( .A(n2439), .B(n2440), .Z(n2435) );
  ANDN U2746 ( .B(n2441), .A(n2442), .Z(n2439) );
  XNOR U2747 ( .A(b[1743]), .B(n2440), .Z(n2441) );
  XNOR U2748 ( .A(b[1743]), .B(n2442), .Z(c[1743]) );
  XNOR U2749 ( .A(a[1743]), .B(n2443), .Z(n2442) );
  IV U2750 ( .A(n2440), .Z(n2443) );
  XOR U2751 ( .A(n2444), .B(n2445), .Z(n2440) );
  ANDN U2752 ( .B(n2446), .A(n2447), .Z(n2444) );
  XNOR U2753 ( .A(b[1742]), .B(n2445), .Z(n2446) );
  XNOR U2754 ( .A(b[1742]), .B(n2447), .Z(c[1742]) );
  XNOR U2755 ( .A(a[1742]), .B(n2448), .Z(n2447) );
  IV U2756 ( .A(n2445), .Z(n2448) );
  XOR U2757 ( .A(n2449), .B(n2450), .Z(n2445) );
  ANDN U2758 ( .B(n2451), .A(n2452), .Z(n2449) );
  XNOR U2759 ( .A(b[1741]), .B(n2450), .Z(n2451) );
  XNOR U2760 ( .A(b[1741]), .B(n2452), .Z(c[1741]) );
  XNOR U2761 ( .A(a[1741]), .B(n2453), .Z(n2452) );
  IV U2762 ( .A(n2450), .Z(n2453) );
  XOR U2763 ( .A(n2454), .B(n2455), .Z(n2450) );
  ANDN U2764 ( .B(n2456), .A(n2457), .Z(n2454) );
  XNOR U2765 ( .A(b[1740]), .B(n2455), .Z(n2456) );
  XNOR U2766 ( .A(b[1740]), .B(n2457), .Z(c[1740]) );
  XNOR U2767 ( .A(a[1740]), .B(n2458), .Z(n2457) );
  IV U2768 ( .A(n2455), .Z(n2458) );
  XOR U2769 ( .A(n2459), .B(n2460), .Z(n2455) );
  ANDN U2770 ( .B(n2461), .A(n2462), .Z(n2459) );
  XNOR U2771 ( .A(b[1739]), .B(n2460), .Z(n2461) );
  XNOR U2772 ( .A(b[173]), .B(n2463), .Z(c[173]) );
  XNOR U2773 ( .A(b[1739]), .B(n2462), .Z(c[1739]) );
  XNOR U2774 ( .A(a[1739]), .B(n2464), .Z(n2462) );
  IV U2775 ( .A(n2460), .Z(n2464) );
  XOR U2776 ( .A(n2465), .B(n2466), .Z(n2460) );
  ANDN U2777 ( .B(n2467), .A(n2468), .Z(n2465) );
  XNOR U2778 ( .A(b[1738]), .B(n2466), .Z(n2467) );
  XNOR U2779 ( .A(b[1738]), .B(n2468), .Z(c[1738]) );
  XNOR U2780 ( .A(a[1738]), .B(n2469), .Z(n2468) );
  IV U2781 ( .A(n2466), .Z(n2469) );
  XOR U2782 ( .A(n2470), .B(n2471), .Z(n2466) );
  ANDN U2783 ( .B(n2472), .A(n2473), .Z(n2470) );
  XNOR U2784 ( .A(b[1737]), .B(n2471), .Z(n2472) );
  XNOR U2785 ( .A(b[1737]), .B(n2473), .Z(c[1737]) );
  XNOR U2786 ( .A(a[1737]), .B(n2474), .Z(n2473) );
  IV U2787 ( .A(n2471), .Z(n2474) );
  XOR U2788 ( .A(n2475), .B(n2476), .Z(n2471) );
  ANDN U2789 ( .B(n2477), .A(n2478), .Z(n2475) );
  XNOR U2790 ( .A(b[1736]), .B(n2476), .Z(n2477) );
  XNOR U2791 ( .A(b[1736]), .B(n2478), .Z(c[1736]) );
  XNOR U2792 ( .A(a[1736]), .B(n2479), .Z(n2478) );
  IV U2793 ( .A(n2476), .Z(n2479) );
  XOR U2794 ( .A(n2480), .B(n2481), .Z(n2476) );
  ANDN U2795 ( .B(n2482), .A(n2483), .Z(n2480) );
  XNOR U2796 ( .A(b[1735]), .B(n2481), .Z(n2482) );
  XNOR U2797 ( .A(b[1735]), .B(n2483), .Z(c[1735]) );
  XNOR U2798 ( .A(a[1735]), .B(n2484), .Z(n2483) );
  IV U2799 ( .A(n2481), .Z(n2484) );
  XOR U2800 ( .A(n2485), .B(n2486), .Z(n2481) );
  ANDN U2801 ( .B(n2487), .A(n2488), .Z(n2485) );
  XNOR U2802 ( .A(b[1734]), .B(n2486), .Z(n2487) );
  XNOR U2803 ( .A(b[1734]), .B(n2488), .Z(c[1734]) );
  XNOR U2804 ( .A(a[1734]), .B(n2489), .Z(n2488) );
  IV U2805 ( .A(n2486), .Z(n2489) );
  XOR U2806 ( .A(n2490), .B(n2491), .Z(n2486) );
  ANDN U2807 ( .B(n2492), .A(n2493), .Z(n2490) );
  XNOR U2808 ( .A(b[1733]), .B(n2491), .Z(n2492) );
  XNOR U2809 ( .A(b[1733]), .B(n2493), .Z(c[1733]) );
  XNOR U2810 ( .A(a[1733]), .B(n2494), .Z(n2493) );
  IV U2811 ( .A(n2491), .Z(n2494) );
  XOR U2812 ( .A(n2495), .B(n2496), .Z(n2491) );
  ANDN U2813 ( .B(n2497), .A(n2498), .Z(n2495) );
  XNOR U2814 ( .A(b[1732]), .B(n2496), .Z(n2497) );
  XNOR U2815 ( .A(b[1732]), .B(n2498), .Z(c[1732]) );
  XNOR U2816 ( .A(a[1732]), .B(n2499), .Z(n2498) );
  IV U2817 ( .A(n2496), .Z(n2499) );
  XOR U2818 ( .A(n2500), .B(n2501), .Z(n2496) );
  ANDN U2819 ( .B(n2502), .A(n2503), .Z(n2500) );
  XNOR U2820 ( .A(b[1731]), .B(n2501), .Z(n2502) );
  XNOR U2821 ( .A(b[1731]), .B(n2503), .Z(c[1731]) );
  XNOR U2822 ( .A(a[1731]), .B(n2504), .Z(n2503) );
  IV U2823 ( .A(n2501), .Z(n2504) );
  XOR U2824 ( .A(n2505), .B(n2506), .Z(n2501) );
  ANDN U2825 ( .B(n2507), .A(n2508), .Z(n2505) );
  XNOR U2826 ( .A(b[1730]), .B(n2506), .Z(n2507) );
  XNOR U2827 ( .A(b[1730]), .B(n2508), .Z(c[1730]) );
  XNOR U2828 ( .A(a[1730]), .B(n2509), .Z(n2508) );
  IV U2829 ( .A(n2506), .Z(n2509) );
  XOR U2830 ( .A(n2510), .B(n2511), .Z(n2506) );
  ANDN U2831 ( .B(n2512), .A(n2513), .Z(n2510) );
  XNOR U2832 ( .A(b[1729]), .B(n2511), .Z(n2512) );
  XNOR U2833 ( .A(b[172]), .B(n2514), .Z(c[172]) );
  XNOR U2834 ( .A(b[1729]), .B(n2513), .Z(c[1729]) );
  XNOR U2835 ( .A(a[1729]), .B(n2515), .Z(n2513) );
  IV U2836 ( .A(n2511), .Z(n2515) );
  XOR U2837 ( .A(n2516), .B(n2517), .Z(n2511) );
  ANDN U2838 ( .B(n2518), .A(n2519), .Z(n2516) );
  XNOR U2839 ( .A(b[1728]), .B(n2517), .Z(n2518) );
  XNOR U2840 ( .A(b[1728]), .B(n2519), .Z(c[1728]) );
  XNOR U2841 ( .A(a[1728]), .B(n2520), .Z(n2519) );
  IV U2842 ( .A(n2517), .Z(n2520) );
  XOR U2843 ( .A(n2521), .B(n2522), .Z(n2517) );
  ANDN U2844 ( .B(n2523), .A(n2524), .Z(n2521) );
  XNOR U2845 ( .A(b[1727]), .B(n2522), .Z(n2523) );
  XNOR U2846 ( .A(b[1727]), .B(n2524), .Z(c[1727]) );
  XNOR U2847 ( .A(a[1727]), .B(n2525), .Z(n2524) );
  IV U2848 ( .A(n2522), .Z(n2525) );
  XOR U2849 ( .A(n2526), .B(n2527), .Z(n2522) );
  ANDN U2850 ( .B(n2528), .A(n2529), .Z(n2526) );
  XNOR U2851 ( .A(b[1726]), .B(n2527), .Z(n2528) );
  XNOR U2852 ( .A(b[1726]), .B(n2529), .Z(c[1726]) );
  XNOR U2853 ( .A(a[1726]), .B(n2530), .Z(n2529) );
  IV U2854 ( .A(n2527), .Z(n2530) );
  XOR U2855 ( .A(n2531), .B(n2532), .Z(n2527) );
  ANDN U2856 ( .B(n2533), .A(n2534), .Z(n2531) );
  XNOR U2857 ( .A(b[1725]), .B(n2532), .Z(n2533) );
  XNOR U2858 ( .A(b[1725]), .B(n2534), .Z(c[1725]) );
  XNOR U2859 ( .A(a[1725]), .B(n2535), .Z(n2534) );
  IV U2860 ( .A(n2532), .Z(n2535) );
  XOR U2861 ( .A(n2536), .B(n2537), .Z(n2532) );
  ANDN U2862 ( .B(n2538), .A(n2539), .Z(n2536) );
  XNOR U2863 ( .A(b[1724]), .B(n2537), .Z(n2538) );
  XNOR U2864 ( .A(b[1724]), .B(n2539), .Z(c[1724]) );
  XNOR U2865 ( .A(a[1724]), .B(n2540), .Z(n2539) );
  IV U2866 ( .A(n2537), .Z(n2540) );
  XOR U2867 ( .A(n2541), .B(n2542), .Z(n2537) );
  ANDN U2868 ( .B(n2543), .A(n2544), .Z(n2541) );
  XNOR U2869 ( .A(b[1723]), .B(n2542), .Z(n2543) );
  XNOR U2870 ( .A(b[1723]), .B(n2544), .Z(c[1723]) );
  XNOR U2871 ( .A(a[1723]), .B(n2545), .Z(n2544) );
  IV U2872 ( .A(n2542), .Z(n2545) );
  XOR U2873 ( .A(n2546), .B(n2547), .Z(n2542) );
  ANDN U2874 ( .B(n2548), .A(n2549), .Z(n2546) );
  XNOR U2875 ( .A(b[1722]), .B(n2547), .Z(n2548) );
  XNOR U2876 ( .A(b[1722]), .B(n2549), .Z(c[1722]) );
  XNOR U2877 ( .A(a[1722]), .B(n2550), .Z(n2549) );
  IV U2878 ( .A(n2547), .Z(n2550) );
  XOR U2879 ( .A(n2551), .B(n2552), .Z(n2547) );
  ANDN U2880 ( .B(n2553), .A(n2554), .Z(n2551) );
  XNOR U2881 ( .A(b[1721]), .B(n2552), .Z(n2553) );
  XNOR U2882 ( .A(b[1721]), .B(n2554), .Z(c[1721]) );
  XNOR U2883 ( .A(a[1721]), .B(n2555), .Z(n2554) );
  IV U2884 ( .A(n2552), .Z(n2555) );
  XOR U2885 ( .A(n2556), .B(n2557), .Z(n2552) );
  ANDN U2886 ( .B(n2558), .A(n2559), .Z(n2556) );
  XNOR U2887 ( .A(b[1720]), .B(n2557), .Z(n2558) );
  XNOR U2888 ( .A(b[1720]), .B(n2559), .Z(c[1720]) );
  XNOR U2889 ( .A(a[1720]), .B(n2560), .Z(n2559) );
  IV U2890 ( .A(n2557), .Z(n2560) );
  XOR U2891 ( .A(n2561), .B(n2562), .Z(n2557) );
  ANDN U2892 ( .B(n2563), .A(n2564), .Z(n2561) );
  XNOR U2893 ( .A(b[1719]), .B(n2562), .Z(n2563) );
  XNOR U2894 ( .A(b[171]), .B(n2565), .Z(c[171]) );
  XNOR U2895 ( .A(b[1719]), .B(n2564), .Z(c[1719]) );
  XNOR U2896 ( .A(a[1719]), .B(n2566), .Z(n2564) );
  IV U2897 ( .A(n2562), .Z(n2566) );
  XOR U2898 ( .A(n2567), .B(n2568), .Z(n2562) );
  ANDN U2899 ( .B(n2569), .A(n2570), .Z(n2567) );
  XNOR U2900 ( .A(b[1718]), .B(n2568), .Z(n2569) );
  XNOR U2901 ( .A(b[1718]), .B(n2570), .Z(c[1718]) );
  XNOR U2902 ( .A(a[1718]), .B(n2571), .Z(n2570) );
  IV U2903 ( .A(n2568), .Z(n2571) );
  XOR U2904 ( .A(n2572), .B(n2573), .Z(n2568) );
  ANDN U2905 ( .B(n2574), .A(n2575), .Z(n2572) );
  XNOR U2906 ( .A(b[1717]), .B(n2573), .Z(n2574) );
  XNOR U2907 ( .A(b[1717]), .B(n2575), .Z(c[1717]) );
  XNOR U2908 ( .A(a[1717]), .B(n2576), .Z(n2575) );
  IV U2909 ( .A(n2573), .Z(n2576) );
  XOR U2910 ( .A(n2577), .B(n2578), .Z(n2573) );
  ANDN U2911 ( .B(n2579), .A(n2580), .Z(n2577) );
  XNOR U2912 ( .A(b[1716]), .B(n2578), .Z(n2579) );
  XNOR U2913 ( .A(b[1716]), .B(n2580), .Z(c[1716]) );
  XNOR U2914 ( .A(a[1716]), .B(n2581), .Z(n2580) );
  IV U2915 ( .A(n2578), .Z(n2581) );
  XOR U2916 ( .A(n2582), .B(n2583), .Z(n2578) );
  ANDN U2917 ( .B(n2584), .A(n2585), .Z(n2582) );
  XNOR U2918 ( .A(b[1715]), .B(n2583), .Z(n2584) );
  XNOR U2919 ( .A(b[1715]), .B(n2585), .Z(c[1715]) );
  XNOR U2920 ( .A(a[1715]), .B(n2586), .Z(n2585) );
  IV U2921 ( .A(n2583), .Z(n2586) );
  XOR U2922 ( .A(n2587), .B(n2588), .Z(n2583) );
  ANDN U2923 ( .B(n2589), .A(n2590), .Z(n2587) );
  XNOR U2924 ( .A(b[1714]), .B(n2588), .Z(n2589) );
  XNOR U2925 ( .A(b[1714]), .B(n2590), .Z(c[1714]) );
  XNOR U2926 ( .A(a[1714]), .B(n2591), .Z(n2590) );
  IV U2927 ( .A(n2588), .Z(n2591) );
  XOR U2928 ( .A(n2592), .B(n2593), .Z(n2588) );
  ANDN U2929 ( .B(n2594), .A(n2595), .Z(n2592) );
  XNOR U2930 ( .A(b[1713]), .B(n2593), .Z(n2594) );
  XNOR U2931 ( .A(b[1713]), .B(n2595), .Z(c[1713]) );
  XNOR U2932 ( .A(a[1713]), .B(n2596), .Z(n2595) );
  IV U2933 ( .A(n2593), .Z(n2596) );
  XOR U2934 ( .A(n2597), .B(n2598), .Z(n2593) );
  ANDN U2935 ( .B(n2599), .A(n2600), .Z(n2597) );
  XNOR U2936 ( .A(b[1712]), .B(n2598), .Z(n2599) );
  XNOR U2937 ( .A(b[1712]), .B(n2600), .Z(c[1712]) );
  XNOR U2938 ( .A(a[1712]), .B(n2601), .Z(n2600) );
  IV U2939 ( .A(n2598), .Z(n2601) );
  XOR U2940 ( .A(n2602), .B(n2603), .Z(n2598) );
  ANDN U2941 ( .B(n2604), .A(n2605), .Z(n2602) );
  XNOR U2942 ( .A(b[1711]), .B(n2603), .Z(n2604) );
  XNOR U2943 ( .A(b[1711]), .B(n2605), .Z(c[1711]) );
  XNOR U2944 ( .A(a[1711]), .B(n2606), .Z(n2605) );
  IV U2945 ( .A(n2603), .Z(n2606) );
  XOR U2946 ( .A(n2607), .B(n2608), .Z(n2603) );
  ANDN U2947 ( .B(n2609), .A(n2610), .Z(n2607) );
  XNOR U2948 ( .A(b[1710]), .B(n2608), .Z(n2609) );
  XNOR U2949 ( .A(b[1710]), .B(n2610), .Z(c[1710]) );
  XNOR U2950 ( .A(a[1710]), .B(n2611), .Z(n2610) );
  IV U2951 ( .A(n2608), .Z(n2611) );
  XOR U2952 ( .A(n2612), .B(n2613), .Z(n2608) );
  ANDN U2953 ( .B(n2614), .A(n2615), .Z(n2612) );
  XNOR U2954 ( .A(b[1709]), .B(n2613), .Z(n2614) );
  XNOR U2955 ( .A(b[170]), .B(n2616), .Z(c[170]) );
  XNOR U2956 ( .A(b[1709]), .B(n2615), .Z(c[1709]) );
  XNOR U2957 ( .A(a[1709]), .B(n2617), .Z(n2615) );
  IV U2958 ( .A(n2613), .Z(n2617) );
  XOR U2959 ( .A(n2618), .B(n2619), .Z(n2613) );
  ANDN U2960 ( .B(n2620), .A(n2621), .Z(n2618) );
  XNOR U2961 ( .A(b[1708]), .B(n2619), .Z(n2620) );
  XNOR U2962 ( .A(b[1708]), .B(n2621), .Z(c[1708]) );
  XNOR U2963 ( .A(a[1708]), .B(n2622), .Z(n2621) );
  IV U2964 ( .A(n2619), .Z(n2622) );
  XOR U2965 ( .A(n2623), .B(n2624), .Z(n2619) );
  ANDN U2966 ( .B(n2625), .A(n2626), .Z(n2623) );
  XNOR U2967 ( .A(b[1707]), .B(n2624), .Z(n2625) );
  XNOR U2968 ( .A(b[1707]), .B(n2626), .Z(c[1707]) );
  XNOR U2969 ( .A(a[1707]), .B(n2627), .Z(n2626) );
  IV U2970 ( .A(n2624), .Z(n2627) );
  XOR U2971 ( .A(n2628), .B(n2629), .Z(n2624) );
  ANDN U2972 ( .B(n2630), .A(n2631), .Z(n2628) );
  XNOR U2973 ( .A(b[1706]), .B(n2629), .Z(n2630) );
  XNOR U2974 ( .A(b[1706]), .B(n2631), .Z(c[1706]) );
  XNOR U2975 ( .A(a[1706]), .B(n2632), .Z(n2631) );
  IV U2976 ( .A(n2629), .Z(n2632) );
  XOR U2977 ( .A(n2633), .B(n2634), .Z(n2629) );
  ANDN U2978 ( .B(n2635), .A(n2636), .Z(n2633) );
  XNOR U2979 ( .A(b[1705]), .B(n2634), .Z(n2635) );
  XNOR U2980 ( .A(b[1705]), .B(n2636), .Z(c[1705]) );
  XNOR U2981 ( .A(a[1705]), .B(n2637), .Z(n2636) );
  IV U2982 ( .A(n2634), .Z(n2637) );
  XOR U2983 ( .A(n2638), .B(n2639), .Z(n2634) );
  ANDN U2984 ( .B(n2640), .A(n2641), .Z(n2638) );
  XNOR U2985 ( .A(b[1704]), .B(n2639), .Z(n2640) );
  XNOR U2986 ( .A(b[1704]), .B(n2641), .Z(c[1704]) );
  XNOR U2987 ( .A(a[1704]), .B(n2642), .Z(n2641) );
  IV U2988 ( .A(n2639), .Z(n2642) );
  XOR U2989 ( .A(n2643), .B(n2644), .Z(n2639) );
  ANDN U2990 ( .B(n2645), .A(n2646), .Z(n2643) );
  XNOR U2991 ( .A(b[1703]), .B(n2644), .Z(n2645) );
  XNOR U2992 ( .A(b[1703]), .B(n2646), .Z(c[1703]) );
  XNOR U2993 ( .A(a[1703]), .B(n2647), .Z(n2646) );
  IV U2994 ( .A(n2644), .Z(n2647) );
  XOR U2995 ( .A(n2648), .B(n2649), .Z(n2644) );
  ANDN U2996 ( .B(n2650), .A(n2651), .Z(n2648) );
  XNOR U2997 ( .A(b[1702]), .B(n2649), .Z(n2650) );
  XNOR U2998 ( .A(b[1702]), .B(n2651), .Z(c[1702]) );
  XNOR U2999 ( .A(a[1702]), .B(n2652), .Z(n2651) );
  IV U3000 ( .A(n2649), .Z(n2652) );
  XOR U3001 ( .A(n2653), .B(n2654), .Z(n2649) );
  ANDN U3002 ( .B(n2655), .A(n2656), .Z(n2653) );
  XNOR U3003 ( .A(b[1701]), .B(n2654), .Z(n2655) );
  XNOR U3004 ( .A(b[1701]), .B(n2656), .Z(c[1701]) );
  XNOR U3005 ( .A(a[1701]), .B(n2657), .Z(n2656) );
  IV U3006 ( .A(n2654), .Z(n2657) );
  XOR U3007 ( .A(n2658), .B(n2659), .Z(n2654) );
  ANDN U3008 ( .B(n2660), .A(n2661), .Z(n2658) );
  XNOR U3009 ( .A(b[1700]), .B(n2659), .Z(n2660) );
  XNOR U3010 ( .A(b[1700]), .B(n2661), .Z(c[1700]) );
  XNOR U3011 ( .A(a[1700]), .B(n2662), .Z(n2661) );
  IV U3012 ( .A(n2659), .Z(n2662) );
  XOR U3013 ( .A(n2663), .B(n2664), .Z(n2659) );
  ANDN U3014 ( .B(n2665), .A(n2666), .Z(n2663) );
  XNOR U3015 ( .A(b[1699]), .B(n2664), .Z(n2665) );
  XNOR U3016 ( .A(b[16]), .B(n2667), .Z(c[16]) );
  XNOR U3017 ( .A(b[169]), .B(n2668), .Z(c[169]) );
  XNOR U3018 ( .A(b[1699]), .B(n2666), .Z(c[1699]) );
  XNOR U3019 ( .A(a[1699]), .B(n2669), .Z(n2666) );
  IV U3020 ( .A(n2664), .Z(n2669) );
  XOR U3021 ( .A(n2670), .B(n2671), .Z(n2664) );
  ANDN U3022 ( .B(n2672), .A(n2673), .Z(n2670) );
  XNOR U3023 ( .A(b[1698]), .B(n2671), .Z(n2672) );
  XNOR U3024 ( .A(b[1698]), .B(n2673), .Z(c[1698]) );
  XNOR U3025 ( .A(a[1698]), .B(n2674), .Z(n2673) );
  IV U3026 ( .A(n2671), .Z(n2674) );
  XOR U3027 ( .A(n2675), .B(n2676), .Z(n2671) );
  ANDN U3028 ( .B(n2677), .A(n2678), .Z(n2675) );
  XNOR U3029 ( .A(b[1697]), .B(n2676), .Z(n2677) );
  XNOR U3030 ( .A(b[1697]), .B(n2678), .Z(c[1697]) );
  XNOR U3031 ( .A(a[1697]), .B(n2679), .Z(n2678) );
  IV U3032 ( .A(n2676), .Z(n2679) );
  XOR U3033 ( .A(n2680), .B(n2681), .Z(n2676) );
  ANDN U3034 ( .B(n2682), .A(n2683), .Z(n2680) );
  XNOR U3035 ( .A(b[1696]), .B(n2681), .Z(n2682) );
  XNOR U3036 ( .A(b[1696]), .B(n2683), .Z(c[1696]) );
  XNOR U3037 ( .A(a[1696]), .B(n2684), .Z(n2683) );
  IV U3038 ( .A(n2681), .Z(n2684) );
  XOR U3039 ( .A(n2685), .B(n2686), .Z(n2681) );
  ANDN U3040 ( .B(n2687), .A(n2688), .Z(n2685) );
  XNOR U3041 ( .A(b[1695]), .B(n2686), .Z(n2687) );
  XNOR U3042 ( .A(b[1695]), .B(n2688), .Z(c[1695]) );
  XNOR U3043 ( .A(a[1695]), .B(n2689), .Z(n2688) );
  IV U3044 ( .A(n2686), .Z(n2689) );
  XOR U3045 ( .A(n2690), .B(n2691), .Z(n2686) );
  ANDN U3046 ( .B(n2692), .A(n2693), .Z(n2690) );
  XNOR U3047 ( .A(b[1694]), .B(n2691), .Z(n2692) );
  XNOR U3048 ( .A(b[1694]), .B(n2693), .Z(c[1694]) );
  XNOR U3049 ( .A(a[1694]), .B(n2694), .Z(n2693) );
  IV U3050 ( .A(n2691), .Z(n2694) );
  XOR U3051 ( .A(n2695), .B(n2696), .Z(n2691) );
  ANDN U3052 ( .B(n2697), .A(n2698), .Z(n2695) );
  XNOR U3053 ( .A(b[1693]), .B(n2696), .Z(n2697) );
  XNOR U3054 ( .A(b[1693]), .B(n2698), .Z(c[1693]) );
  XNOR U3055 ( .A(a[1693]), .B(n2699), .Z(n2698) );
  IV U3056 ( .A(n2696), .Z(n2699) );
  XOR U3057 ( .A(n2700), .B(n2701), .Z(n2696) );
  ANDN U3058 ( .B(n2702), .A(n2703), .Z(n2700) );
  XNOR U3059 ( .A(b[1692]), .B(n2701), .Z(n2702) );
  XNOR U3060 ( .A(b[1692]), .B(n2703), .Z(c[1692]) );
  XNOR U3061 ( .A(a[1692]), .B(n2704), .Z(n2703) );
  IV U3062 ( .A(n2701), .Z(n2704) );
  XOR U3063 ( .A(n2705), .B(n2706), .Z(n2701) );
  ANDN U3064 ( .B(n2707), .A(n2708), .Z(n2705) );
  XNOR U3065 ( .A(b[1691]), .B(n2706), .Z(n2707) );
  XNOR U3066 ( .A(b[1691]), .B(n2708), .Z(c[1691]) );
  XNOR U3067 ( .A(a[1691]), .B(n2709), .Z(n2708) );
  IV U3068 ( .A(n2706), .Z(n2709) );
  XOR U3069 ( .A(n2710), .B(n2711), .Z(n2706) );
  ANDN U3070 ( .B(n2712), .A(n2713), .Z(n2710) );
  XNOR U3071 ( .A(b[1690]), .B(n2711), .Z(n2712) );
  XNOR U3072 ( .A(b[1690]), .B(n2713), .Z(c[1690]) );
  XNOR U3073 ( .A(a[1690]), .B(n2714), .Z(n2713) );
  IV U3074 ( .A(n2711), .Z(n2714) );
  XOR U3075 ( .A(n2715), .B(n2716), .Z(n2711) );
  ANDN U3076 ( .B(n2717), .A(n2718), .Z(n2715) );
  XNOR U3077 ( .A(b[1689]), .B(n2716), .Z(n2717) );
  XNOR U3078 ( .A(b[168]), .B(n2719), .Z(c[168]) );
  XNOR U3079 ( .A(b[1689]), .B(n2718), .Z(c[1689]) );
  XNOR U3080 ( .A(a[1689]), .B(n2720), .Z(n2718) );
  IV U3081 ( .A(n2716), .Z(n2720) );
  XOR U3082 ( .A(n2721), .B(n2722), .Z(n2716) );
  ANDN U3083 ( .B(n2723), .A(n2724), .Z(n2721) );
  XNOR U3084 ( .A(b[1688]), .B(n2722), .Z(n2723) );
  XNOR U3085 ( .A(b[1688]), .B(n2724), .Z(c[1688]) );
  XNOR U3086 ( .A(a[1688]), .B(n2725), .Z(n2724) );
  IV U3087 ( .A(n2722), .Z(n2725) );
  XOR U3088 ( .A(n2726), .B(n2727), .Z(n2722) );
  ANDN U3089 ( .B(n2728), .A(n2729), .Z(n2726) );
  XNOR U3090 ( .A(b[1687]), .B(n2727), .Z(n2728) );
  XNOR U3091 ( .A(b[1687]), .B(n2729), .Z(c[1687]) );
  XNOR U3092 ( .A(a[1687]), .B(n2730), .Z(n2729) );
  IV U3093 ( .A(n2727), .Z(n2730) );
  XOR U3094 ( .A(n2731), .B(n2732), .Z(n2727) );
  ANDN U3095 ( .B(n2733), .A(n2734), .Z(n2731) );
  XNOR U3096 ( .A(b[1686]), .B(n2732), .Z(n2733) );
  XNOR U3097 ( .A(b[1686]), .B(n2734), .Z(c[1686]) );
  XNOR U3098 ( .A(a[1686]), .B(n2735), .Z(n2734) );
  IV U3099 ( .A(n2732), .Z(n2735) );
  XOR U3100 ( .A(n2736), .B(n2737), .Z(n2732) );
  ANDN U3101 ( .B(n2738), .A(n2739), .Z(n2736) );
  XNOR U3102 ( .A(b[1685]), .B(n2737), .Z(n2738) );
  XNOR U3103 ( .A(b[1685]), .B(n2739), .Z(c[1685]) );
  XNOR U3104 ( .A(a[1685]), .B(n2740), .Z(n2739) );
  IV U3105 ( .A(n2737), .Z(n2740) );
  XOR U3106 ( .A(n2741), .B(n2742), .Z(n2737) );
  ANDN U3107 ( .B(n2743), .A(n2744), .Z(n2741) );
  XNOR U3108 ( .A(b[1684]), .B(n2742), .Z(n2743) );
  XNOR U3109 ( .A(b[1684]), .B(n2744), .Z(c[1684]) );
  XNOR U3110 ( .A(a[1684]), .B(n2745), .Z(n2744) );
  IV U3111 ( .A(n2742), .Z(n2745) );
  XOR U3112 ( .A(n2746), .B(n2747), .Z(n2742) );
  ANDN U3113 ( .B(n2748), .A(n2749), .Z(n2746) );
  XNOR U3114 ( .A(b[1683]), .B(n2747), .Z(n2748) );
  XNOR U3115 ( .A(b[1683]), .B(n2749), .Z(c[1683]) );
  XNOR U3116 ( .A(a[1683]), .B(n2750), .Z(n2749) );
  IV U3117 ( .A(n2747), .Z(n2750) );
  XOR U3118 ( .A(n2751), .B(n2752), .Z(n2747) );
  ANDN U3119 ( .B(n2753), .A(n2754), .Z(n2751) );
  XNOR U3120 ( .A(b[1682]), .B(n2752), .Z(n2753) );
  XNOR U3121 ( .A(b[1682]), .B(n2754), .Z(c[1682]) );
  XNOR U3122 ( .A(a[1682]), .B(n2755), .Z(n2754) );
  IV U3123 ( .A(n2752), .Z(n2755) );
  XOR U3124 ( .A(n2756), .B(n2757), .Z(n2752) );
  ANDN U3125 ( .B(n2758), .A(n2759), .Z(n2756) );
  XNOR U3126 ( .A(b[1681]), .B(n2757), .Z(n2758) );
  XNOR U3127 ( .A(b[1681]), .B(n2759), .Z(c[1681]) );
  XNOR U3128 ( .A(a[1681]), .B(n2760), .Z(n2759) );
  IV U3129 ( .A(n2757), .Z(n2760) );
  XOR U3130 ( .A(n2761), .B(n2762), .Z(n2757) );
  ANDN U3131 ( .B(n2763), .A(n2764), .Z(n2761) );
  XNOR U3132 ( .A(b[1680]), .B(n2762), .Z(n2763) );
  XNOR U3133 ( .A(b[1680]), .B(n2764), .Z(c[1680]) );
  XNOR U3134 ( .A(a[1680]), .B(n2765), .Z(n2764) );
  IV U3135 ( .A(n2762), .Z(n2765) );
  XOR U3136 ( .A(n2766), .B(n2767), .Z(n2762) );
  ANDN U3137 ( .B(n2768), .A(n2769), .Z(n2766) );
  XNOR U3138 ( .A(b[1679]), .B(n2767), .Z(n2768) );
  XNOR U3139 ( .A(b[167]), .B(n2770), .Z(c[167]) );
  XNOR U3140 ( .A(b[1679]), .B(n2769), .Z(c[1679]) );
  XNOR U3141 ( .A(a[1679]), .B(n2771), .Z(n2769) );
  IV U3142 ( .A(n2767), .Z(n2771) );
  XOR U3143 ( .A(n2772), .B(n2773), .Z(n2767) );
  ANDN U3144 ( .B(n2774), .A(n2775), .Z(n2772) );
  XNOR U3145 ( .A(b[1678]), .B(n2773), .Z(n2774) );
  XNOR U3146 ( .A(b[1678]), .B(n2775), .Z(c[1678]) );
  XNOR U3147 ( .A(a[1678]), .B(n2776), .Z(n2775) );
  IV U3148 ( .A(n2773), .Z(n2776) );
  XOR U3149 ( .A(n2777), .B(n2778), .Z(n2773) );
  ANDN U3150 ( .B(n2779), .A(n2780), .Z(n2777) );
  XNOR U3151 ( .A(b[1677]), .B(n2778), .Z(n2779) );
  XNOR U3152 ( .A(b[1677]), .B(n2780), .Z(c[1677]) );
  XNOR U3153 ( .A(a[1677]), .B(n2781), .Z(n2780) );
  IV U3154 ( .A(n2778), .Z(n2781) );
  XOR U3155 ( .A(n2782), .B(n2783), .Z(n2778) );
  ANDN U3156 ( .B(n2784), .A(n2785), .Z(n2782) );
  XNOR U3157 ( .A(b[1676]), .B(n2783), .Z(n2784) );
  XNOR U3158 ( .A(b[1676]), .B(n2785), .Z(c[1676]) );
  XNOR U3159 ( .A(a[1676]), .B(n2786), .Z(n2785) );
  IV U3160 ( .A(n2783), .Z(n2786) );
  XOR U3161 ( .A(n2787), .B(n2788), .Z(n2783) );
  ANDN U3162 ( .B(n2789), .A(n2790), .Z(n2787) );
  XNOR U3163 ( .A(b[1675]), .B(n2788), .Z(n2789) );
  XNOR U3164 ( .A(b[1675]), .B(n2790), .Z(c[1675]) );
  XNOR U3165 ( .A(a[1675]), .B(n2791), .Z(n2790) );
  IV U3166 ( .A(n2788), .Z(n2791) );
  XOR U3167 ( .A(n2792), .B(n2793), .Z(n2788) );
  ANDN U3168 ( .B(n2794), .A(n2795), .Z(n2792) );
  XNOR U3169 ( .A(b[1674]), .B(n2793), .Z(n2794) );
  XNOR U3170 ( .A(b[1674]), .B(n2795), .Z(c[1674]) );
  XNOR U3171 ( .A(a[1674]), .B(n2796), .Z(n2795) );
  IV U3172 ( .A(n2793), .Z(n2796) );
  XOR U3173 ( .A(n2797), .B(n2798), .Z(n2793) );
  ANDN U3174 ( .B(n2799), .A(n2800), .Z(n2797) );
  XNOR U3175 ( .A(b[1673]), .B(n2798), .Z(n2799) );
  XNOR U3176 ( .A(b[1673]), .B(n2800), .Z(c[1673]) );
  XNOR U3177 ( .A(a[1673]), .B(n2801), .Z(n2800) );
  IV U3178 ( .A(n2798), .Z(n2801) );
  XOR U3179 ( .A(n2802), .B(n2803), .Z(n2798) );
  ANDN U3180 ( .B(n2804), .A(n2805), .Z(n2802) );
  XNOR U3181 ( .A(b[1672]), .B(n2803), .Z(n2804) );
  XNOR U3182 ( .A(b[1672]), .B(n2805), .Z(c[1672]) );
  XNOR U3183 ( .A(a[1672]), .B(n2806), .Z(n2805) );
  IV U3184 ( .A(n2803), .Z(n2806) );
  XOR U3185 ( .A(n2807), .B(n2808), .Z(n2803) );
  ANDN U3186 ( .B(n2809), .A(n2810), .Z(n2807) );
  XNOR U3187 ( .A(b[1671]), .B(n2808), .Z(n2809) );
  XNOR U3188 ( .A(b[1671]), .B(n2810), .Z(c[1671]) );
  XNOR U3189 ( .A(a[1671]), .B(n2811), .Z(n2810) );
  IV U3190 ( .A(n2808), .Z(n2811) );
  XOR U3191 ( .A(n2812), .B(n2813), .Z(n2808) );
  ANDN U3192 ( .B(n2814), .A(n2815), .Z(n2812) );
  XNOR U3193 ( .A(b[1670]), .B(n2813), .Z(n2814) );
  XNOR U3194 ( .A(b[1670]), .B(n2815), .Z(c[1670]) );
  XNOR U3195 ( .A(a[1670]), .B(n2816), .Z(n2815) );
  IV U3196 ( .A(n2813), .Z(n2816) );
  XOR U3197 ( .A(n2817), .B(n2818), .Z(n2813) );
  ANDN U3198 ( .B(n2819), .A(n2820), .Z(n2817) );
  XNOR U3199 ( .A(b[1669]), .B(n2818), .Z(n2819) );
  XNOR U3200 ( .A(b[166]), .B(n2821), .Z(c[166]) );
  XNOR U3201 ( .A(b[1669]), .B(n2820), .Z(c[1669]) );
  XNOR U3202 ( .A(a[1669]), .B(n2822), .Z(n2820) );
  IV U3203 ( .A(n2818), .Z(n2822) );
  XOR U3204 ( .A(n2823), .B(n2824), .Z(n2818) );
  ANDN U3205 ( .B(n2825), .A(n2826), .Z(n2823) );
  XNOR U3206 ( .A(b[1668]), .B(n2824), .Z(n2825) );
  XNOR U3207 ( .A(b[1668]), .B(n2826), .Z(c[1668]) );
  XNOR U3208 ( .A(a[1668]), .B(n2827), .Z(n2826) );
  IV U3209 ( .A(n2824), .Z(n2827) );
  XOR U3210 ( .A(n2828), .B(n2829), .Z(n2824) );
  ANDN U3211 ( .B(n2830), .A(n2831), .Z(n2828) );
  XNOR U3212 ( .A(b[1667]), .B(n2829), .Z(n2830) );
  XNOR U3213 ( .A(b[1667]), .B(n2831), .Z(c[1667]) );
  XNOR U3214 ( .A(a[1667]), .B(n2832), .Z(n2831) );
  IV U3215 ( .A(n2829), .Z(n2832) );
  XOR U3216 ( .A(n2833), .B(n2834), .Z(n2829) );
  ANDN U3217 ( .B(n2835), .A(n2836), .Z(n2833) );
  XNOR U3218 ( .A(b[1666]), .B(n2834), .Z(n2835) );
  XNOR U3219 ( .A(b[1666]), .B(n2836), .Z(c[1666]) );
  XNOR U3220 ( .A(a[1666]), .B(n2837), .Z(n2836) );
  IV U3221 ( .A(n2834), .Z(n2837) );
  XOR U3222 ( .A(n2838), .B(n2839), .Z(n2834) );
  ANDN U3223 ( .B(n2840), .A(n2841), .Z(n2838) );
  XNOR U3224 ( .A(b[1665]), .B(n2839), .Z(n2840) );
  XNOR U3225 ( .A(b[1665]), .B(n2841), .Z(c[1665]) );
  XNOR U3226 ( .A(a[1665]), .B(n2842), .Z(n2841) );
  IV U3227 ( .A(n2839), .Z(n2842) );
  XOR U3228 ( .A(n2843), .B(n2844), .Z(n2839) );
  ANDN U3229 ( .B(n2845), .A(n2846), .Z(n2843) );
  XNOR U3230 ( .A(b[1664]), .B(n2844), .Z(n2845) );
  XNOR U3231 ( .A(b[1664]), .B(n2846), .Z(c[1664]) );
  XNOR U3232 ( .A(a[1664]), .B(n2847), .Z(n2846) );
  IV U3233 ( .A(n2844), .Z(n2847) );
  XOR U3234 ( .A(n2848), .B(n2849), .Z(n2844) );
  ANDN U3235 ( .B(n2850), .A(n2851), .Z(n2848) );
  XNOR U3236 ( .A(b[1663]), .B(n2849), .Z(n2850) );
  XNOR U3237 ( .A(b[1663]), .B(n2851), .Z(c[1663]) );
  XNOR U3238 ( .A(a[1663]), .B(n2852), .Z(n2851) );
  IV U3239 ( .A(n2849), .Z(n2852) );
  XOR U3240 ( .A(n2853), .B(n2854), .Z(n2849) );
  ANDN U3241 ( .B(n2855), .A(n2856), .Z(n2853) );
  XNOR U3242 ( .A(b[1662]), .B(n2854), .Z(n2855) );
  XNOR U3243 ( .A(b[1662]), .B(n2856), .Z(c[1662]) );
  XNOR U3244 ( .A(a[1662]), .B(n2857), .Z(n2856) );
  IV U3245 ( .A(n2854), .Z(n2857) );
  XOR U3246 ( .A(n2858), .B(n2859), .Z(n2854) );
  ANDN U3247 ( .B(n2860), .A(n2861), .Z(n2858) );
  XNOR U3248 ( .A(b[1661]), .B(n2859), .Z(n2860) );
  XNOR U3249 ( .A(b[1661]), .B(n2861), .Z(c[1661]) );
  XNOR U3250 ( .A(a[1661]), .B(n2862), .Z(n2861) );
  IV U3251 ( .A(n2859), .Z(n2862) );
  XOR U3252 ( .A(n2863), .B(n2864), .Z(n2859) );
  ANDN U3253 ( .B(n2865), .A(n2866), .Z(n2863) );
  XNOR U3254 ( .A(b[1660]), .B(n2864), .Z(n2865) );
  XNOR U3255 ( .A(b[1660]), .B(n2866), .Z(c[1660]) );
  XNOR U3256 ( .A(a[1660]), .B(n2867), .Z(n2866) );
  IV U3257 ( .A(n2864), .Z(n2867) );
  XOR U3258 ( .A(n2868), .B(n2869), .Z(n2864) );
  ANDN U3259 ( .B(n2870), .A(n2871), .Z(n2868) );
  XNOR U3260 ( .A(b[1659]), .B(n2869), .Z(n2870) );
  XNOR U3261 ( .A(b[165]), .B(n2872), .Z(c[165]) );
  XNOR U3262 ( .A(b[1659]), .B(n2871), .Z(c[1659]) );
  XNOR U3263 ( .A(a[1659]), .B(n2873), .Z(n2871) );
  IV U3264 ( .A(n2869), .Z(n2873) );
  XOR U3265 ( .A(n2874), .B(n2875), .Z(n2869) );
  ANDN U3266 ( .B(n2876), .A(n2877), .Z(n2874) );
  XNOR U3267 ( .A(b[1658]), .B(n2875), .Z(n2876) );
  XNOR U3268 ( .A(b[1658]), .B(n2877), .Z(c[1658]) );
  XNOR U3269 ( .A(a[1658]), .B(n2878), .Z(n2877) );
  IV U3270 ( .A(n2875), .Z(n2878) );
  XOR U3271 ( .A(n2879), .B(n2880), .Z(n2875) );
  ANDN U3272 ( .B(n2881), .A(n2882), .Z(n2879) );
  XNOR U3273 ( .A(b[1657]), .B(n2880), .Z(n2881) );
  XNOR U3274 ( .A(b[1657]), .B(n2882), .Z(c[1657]) );
  XNOR U3275 ( .A(a[1657]), .B(n2883), .Z(n2882) );
  IV U3276 ( .A(n2880), .Z(n2883) );
  XOR U3277 ( .A(n2884), .B(n2885), .Z(n2880) );
  ANDN U3278 ( .B(n2886), .A(n2887), .Z(n2884) );
  XNOR U3279 ( .A(b[1656]), .B(n2885), .Z(n2886) );
  XNOR U3280 ( .A(b[1656]), .B(n2887), .Z(c[1656]) );
  XNOR U3281 ( .A(a[1656]), .B(n2888), .Z(n2887) );
  IV U3282 ( .A(n2885), .Z(n2888) );
  XOR U3283 ( .A(n2889), .B(n2890), .Z(n2885) );
  ANDN U3284 ( .B(n2891), .A(n2892), .Z(n2889) );
  XNOR U3285 ( .A(b[1655]), .B(n2890), .Z(n2891) );
  XNOR U3286 ( .A(b[1655]), .B(n2892), .Z(c[1655]) );
  XNOR U3287 ( .A(a[1655]), .B(n2893), .Z(n2892) );
  IV U3288 ( .A(n2890), .Z(n2893) );
  XOR U3289 ( .A(n2894), .B(n2895), .Z(n2890) );
  ANDN U3290 ( .B(n2896), .A(n2897), .Z(n2894) );
  XNOR U3291 ( .A(b[1654]), .B(n2895), .Z(n2896) );
  XNOR U3292 ( .A(b[1654]), .B(n2897), .Z(c[1654]) );
  XNOR U3293 ( .A(a[1654]), .B(n2898), .Z(n2897) );
  IV U3294 ( .A(n2895), .Z(n2898) );
  XOR U3295 ( .A(n2899), .B(n2900), .Z(n2895) );
  ANDN U3296 ( .B(n2901), .A(n2902), .Z(n2899) );
  XNOR U3297 ( .A(b[1653]), .B(n2900), .Z(n2901) );
  XNOR U3298 ( .A(b[1653]), .B(n2902), .Z(c[1653]) );
  XNOR U3299 ( .A(a[1653]), .B(n2903), .Z(n2902) );
  IV U3300 ( .A(n2900), .Z(n2903) );
  XOR U3301 ( .A(n2904), .B(n2905), .Z(n2900) );
  ANDN U3302 ( .B(n2906), .A(n2907), .Z(n2904) );
  XNOR U3303 ( .A(b[1652]), .B(n2905), .Z(n2906) );
  XNOR U3304 ( .A(b[1652]), .B(n2907), .Z(c[1652]) );
  XNOR U3305 ( .A(a[1652]), .B(n2908), .Z(n2907) );
  IV U3306 ( .A(n2905), .Z(n2908) );
  XOR U3307 ( .A(n2909), .B(n2910), .Z(n2905) );
  ANDN U3308 ( .B(n2911), .A(n2912), .Z(n2909) );
  XNOR U3309 ( .A(b[1651]), .B(n2910), .Z(n2911) );
  XNOR U3310 ( .A(b[1651]), .B(n2912), .Z(c[1651]) );
  XNOR U3311 ( .A(a[1651]), .B(n2913), .Z(n2912) );
  IV U3312 ( .A(n2910), .Z(n2913) );
  XOR U3313 ( .A(n2914), .B(n2915), .Z(n2910) );
  ANDN U3314 ( .B(n2916), .A(n2917), .Z(n2914) );
  XNOR U3315 ( .A(b[1650]), .B(n2915), .Z(n2916) );
  XNOR U3316 ( .A(b[1650]), .B(n2917), .Z(c[1650]) );
  XNOR U3317 ( .A(a[1650]), .B(n2918), .Z(n2917) );
  IV U3318 ( .A(n2915), .Z(n2918) );
  XOR U3319 ( .A(n2919), .B(n2920), .Z(n2915) );
  ANDN U3320 ( .B(n2921), .A(n2922), .Z(n2919) );
  XNOR U3321 ( .A(b[1649]), .B(n2920), .Z(n2921) );
  XNOR U3322 ( .A(b[164]), .B(n2923), .Z(c[164]) );
  XNOR U3323 ( .A(b[1649]), .B(n2922), .Z(c[1649]) );
  XNOR U3324 ( .A(a[1649]), .B(n2924), .Z(n2922) );
  IV U3325 ( .A(n2920), .Z(n2924) );
  XOR U3326 ( .A(n2925), .B(n2926), .Z(n2920) );
  ANDN U3327 ( .B(n2927), .A(n2928), .Z(n2925) );
  XNOR U3328 ( .A(b[1648]), .B(n2926), .Z(n2927) );
  XNOR U3329 ( .A(b[1648]), .B(n2928), .Z(c[1648]) );
  XNOR U3330 ( .A(a[1648]), .B(n2929), .Z(n2928) );
  IV U3331 ( .A(n2926), .Z(n2929) );
  XOR U3332 ( .A(n2930), .B(n2931), .Z(n2926) );
  ANDN U3333 ( .B(n2932), .A(n2933), .Z(n2930) );
  XNOR U3334 ( .A(b[1647]), .B(n2931), .Z(n2932) );
  XNOR U3335 ( .A(b[1647]), .B(n2933), .Z(c[1647]) );
  XNOR U3336 ( .A(a[1647]), .B(n2934), .Z(n2933) );
  IV U3337 ( .A(n2931), .Z(n2934) );
  XOR U3338 ( .A(n2935), .B(n2936), .Z(n2931) );
  ANDN U3339 ( .B(n2937), .A(n2938), .Z(n2935) );
  XNOR U3340 ( .A(b[1646]), .B(n2936), .Z(n2937) );
  XNOR U3341 ( .A(b[1646]), .B(n2938), .Z(c[1646]) );
  XNOR U3342 ( .A(a[1646]), .B(n2939), .Z(n2938) );
  IV U3343 ( .A(n2936), .Z(n2939) );
  XOR U3344 ( .A(n2940), .B(n2941), .Z(n2936) );
  ANDN U3345 ( .B(n2942), .A(n2943), .Z(n2940) );
  XNOR U3346 ( .A(b[1645]), .B(n2941), .Z(n2942) );
  XNOR U3347 ( .A(b[1645]), .B(n2943), .Z(c[1645]) );
  XNOR U3348 ( .A(a[1645]), .B(n2944), .Z(n2943) );
  IV U3349 ( .A(n2941), .Z(n2944) );
  XOR U3350 ( .A(n2945), .B(n2946), .Z(n2941) );
  ANDN U3351 ( .B(n2947), .A(n2948), .Z(n2945) );
  XNOR U3352 ( .A(b[1644]), .B(n2946), .Z(n2947) );
  XNOR U3353 ( .A(b[1644]), .B(n2948), .Z(c[1644]) );
  XNOR U3354 ( .A(a[1644]), .B(n2949), .Z(n2948) );
  IV U3355 ( .A(n2946), .Z(n2949) );
  XOR U3356 ( .A(n2950), .B(n2951), .Z(n2946) );
  ANDN U3357 ( .B(n2952), .A(n2953), .Z(n2950) );
  XNOR U3358 ( .A(b[1643]), .B(n2951), .Z(n2952) );
  XNOR U3359 ( .A(b[1643]), .B(n2953), .Z(c[1643]) );
  XNOR U3360 ( .A(a[1643]), .B(n2954), .Z(n2953) );
  IV U3361 ( .A(n2951), .Z(n2954) );
  XOR U3362 ( .A(n2955), .B(n2956), .Z(n2951) );
  ANDN U3363 ( .B(n2957), .A(n2958), .Z(n2955) );
  XNOR U3364 ( .A(b[1642]), .B(n2956), .Z(n2957) );
  XNOR U3365 ( .A(b[1642]), .B(n2958), .Z(c[1642]) );
  XNOR U3366 ( .A(a[1642]), .B(n2959), .Z(n2958) );
  IV U3367 ( .A(n2956), .Z(n2959) );
  XOR U3368 ( .A(n2960), .B(n2961), .Z(n2956) );
  ANDN U3369 ( .B(n2962), .A(n2963), .Z(n2960) );
  XNOR U3370 ( .A(b[1641]), .B(n2961), .Z(n2962) );
  XNOR U3371 ( .A(b[1641]), .B(n2963), .Z(c[1641]) );
  XNOR U3372 ( .A(a[1641]), .B(n2964), .Z(n2963) );
  IV U3373 ( .A(n2961), .Z(n2964) );
  XOR U3374 ( .A(n2965), .B(n2966), .Z(n2961) );
  ANDN U3375 ( .B(n2967), .A(n2968), .Z(n2965) );
  XNOR U3376 ( .A(b[1640]), .B(n2966), .Z(n2967) );
  XNOR U3377 ( .A(b[1640]), .B(n2968), .Z(c[1640]) );
  XNOR U3378 ( .A(a[1640]), .B(n2969), .Z(n2968) );
  IV U3379 ( .A(n2966), .Z(n2969) );
  XOR U3380 ( .A(n2970), .B(n2971), .Z(n2966) );
  ANDN U3381 ( .B(n2972), .A(n2973), .Z(n2970) );
  XNOR U3382 ( .A(b[1639]), .B(n2971), .Z(n2972) );
  XNOR U3383 ( .A(b[163]), .B(n2974), .Z(c[163]) );
  XNOR U3384 ( .A(b[1639]), .B(n2973), .Z(c[1639]) );
  XNOR U3385 ( .A(a[1639]), .B(n2975), .Z(n2973) );
  IV U3386 ( .A(n2971), .Z(n2975) );
  XOR U3387 ( .A(n2976), .B(n2977), .Z(n2971) );
  ANDN U3388 ( .B(n2978), .A(n2979), .Z(n2976) );
  XNOR U3389 ( .A(b[1638]), .B(n2977), .Z(n2978) );
  XNOR U3390 ( .A(b[1638]), .B(n2979), .Z(c[1638]) );
  XNOR U3391 ( .A(a[1638]), .B(n2980), .Z(n2979) );
  IV U3392 ( .A(n2977), .Z(n2980) );
  XOR U3393 ( .A(n2981), .B(n2982), .Z(n2977) );
  ANDN U3394 ( .B(n2983), .A(n2984), .Z(n2981) );
  XNOR U3395 ( .A(b[1637]), .B(n2982), .Z(n2983) );
  XNOR U3396 ( .A(b[1637]), .B(n2984), .Z(c[1637]) );
  XNOR U3397 ( .A(a[1637]), .B(n2985), .Z(n2984) );
  IV U3398 ( .A(n2982), .Z(n2985) );
  XOR U3399 ( .A(n2986), .B(n2987), .Z(n2982) );
  ANDN U3400 ( .B(n2988), .A(n2989), .Z(n2986) );
  XNOR U3401 ( .A(b[1636]), .B(n2987), .Z(n2988) );
  XNOR U3402 ( .A(b[1636]), .B(n2989), .Z(c[1636]) );
  XNOR U3403 ( .A(a[1636]), .B(n2990), .Z(n2989) );
  IV U3404 ( .A(n2987), .Z(n2990) );
  XOR U3405 ( .A(n2991), .B(n2992), .Z(n2987) );
  ANDN U3406 ( .B(n2993), .A(n2994), .Z(n2991) );
  XNOR U3407 ( .A(b[1635]), .B(n2992), .Z(n2993) );
  XNOR U3408 ( .A(b[1635]), .B(n2994), .Z(c[1635]) );
  XNOR U3409 ( .A(a[1635]), .B(n2995), .Z(n2994) );
  IV U3410 ( .A(n2992), .Z(n2995) );
  XOR U3411 ( .A(n2996), .B(n2997), .Z(n2992) );
  ANDN U3412 ( .B(n2998), .A(n2999), .Z(n2996) );
  XNOR U3413 ( .A(b[1634]), .B(n2997), .Z(n2998) );
  XNOR U3414 ( .A(b[1634]), .B(n2999), .Z(c[1634]) );
  XNOR U3415 ( .A(a[1634]), .B(n3000), .Z(n2999) );
  IV U3416 ( .A(n2997), .Z(n3000) );
  XOR U3417 ( .A(n3001), .B(n3002), .Z(n2997) );
  ANDN U3418 ( .B(n3003), .A(n3004), .Z(n3001) );
  XNOR U3419 ( .A(b[1633]), .B(n3002), .Z(n3003) );
  XNOR U3420 ( .A(b[1633]), .B(n3004), .Z(c[1633]) );
  XNOR U3421 ( .A(a[1633]), .B(n3005), .Z(n3004) );
  IV U3422 ( .A(n3002), .Z(n3005) );
  XOR U3423 ( .A(n3006), .B(n3007), .Z(n3002) );
  ANDN U3424 ( .B(n3008), .A(n3009), .Z(n3006) );
  XNOR U3425 ( .A(b[1632]), .B(n3007), .Z(n3008) );
  XNOR U3426 ( .A(b[1632]), .B(n3009), .Z(c[1632]) );
  XNOR U3427 ( .A(a[1632]), .B(n3010), .Z(n3009) );
  IV U3428 ( .A(n3007), .Z(n3010) );
  XOR U3429 ( .A(n3011), .B(n3012), .Z(n3007) );
  ANDN U3430 ( .B(n3013), .A(n3014), .Z(n3011) );
  XNOR U3431 ( .A(b[1631]), .B(n3012), .Z(n3013) );
  XNOR U3432 ( .A(b[1631]), .B(n3014), .Z(c[1631]) );
  XNOR U3433 ( .A(a[1631]), .B(n3015), .Z(n3014) );
  IV U3434 ( .A(n3012), .Z(n3015) );
  XOR U3435 ( .A(n3016), .B(n3017), .Z(n3012) );
  ANDN U3436 ( .B(n3018), .A(n3019), .Z(n3016) );
  XNOR U3437 ( .A(b[1630]), .B(n3017), .Z(n3018) );
  XNOR U3438 ( .A(b[1630]), .B(n3019), .Z(c[1630]) );
  XNOR U3439 ( .A(a[1630]), .B(n3020), .Z(n3019) );
  IV U3440 ( .A(n3017), .Z(n3020) );
  XOR U3441 ( .A(n3021), .B(n3022), .Z(n3017) );
  ANDN U3442 ( .B(n3023), .A(n3024), .Z(n3021) );
  XNOR U3443 ( .A(b[1629]), .B(n3022), .Z(n3023) );
  XNOR U3444 ( .A(b[162]), .B(n3025), .Z(c[162]) );
  XNOR U3445 ( .A(b[1629]), .B(n3024), .Z(c[1629]) );
  XNOR U3446 ( .A(a[1629]), .B(n3026), .Z(n3024) );
  IV U3447 ( .A(n3022), .Z(n3026) );
  XOR U3448 ( .A(n3027), .B(n3028), .Z(n3022) );
  ANDN U3449 ( .B(n3029), .A(n3030), .Z(n3027) );
  XNOR U3450 ( .A(b[1628]), .B(n3028), .Z(n3029) );
  XNOR U3451 ( .A(b[1628]), .B(n3030), .Z(c[1628]) );
  XNOR U3452 ( .A(a[1628]), .B(n3031), .Z(n3030) );
  IV U3453 ( .A(n3028), .Z(n3031) );
  XOR U3454 ( .A(n3032), .B(n3033), .Z(n3028) );
  ANDN U3455 ( .B(n3034), .A(n3035), .Z(n3032) );
  XNOR U3456 ( .A(b[1627]), .B(n3033), .Z(n3034) );
  XNOR U3457 ( .A(b[1627]), .B(n3035), .Z(c[1627]) );
  XNOR U3458 ( .A(a[1627]), .B(n3036), .Z(n3035) );
  IV U3459 ( .A(n3033), .Z(n3036) );
  XOR U3460 ( .A(n3037), .B(n3038), .Z(n3033) );
  ANDN U3461 ( .B(n3039), .A(n3040), .Z(n3037) );
  XNOR U3462 ( .A(b[1626]), .B(n3038), .Z(n3039) );
  XNOR U3463 ( .A(b[1626]), .B(n3040), .Z(c[1626]) );
  XNOR U3464 ( .A(a[1626]), .B(n3041), .Z(n3040) );
  IV U3465 ( .A(n3038), .Z(n3041) );
  XOR U3466 ( .A(n3042), .B(n3043), .Z(n3038) );
  ANDN U3467 ( .B(n3044), .A(n3045), .Z(n3042) );
  XNOR U3468 ( .A(b[1625]), .B(n3043), .Z(n3044) );
  XNOR U3469 ( .A(b[1625]), .B(n3045), .Z(c[1625]) );
  XNOR U3470 ( .A(a[1625]), .B(n3046), .Z(n3045) );
  IV U3471 ( .A(n3043), .Z(n3046) );
  XOR U3472 ( .A(n3047), .B(n3048), .Z(n3043) );
  ANDN U3473 ( .B(n3049), .A(n3050), .Z(n3047) );
  XNOR U3474 ( .A(b[1624]), .B(n3048), .Z(n3049) );
  XNOR U3475 ( .A(b[1624]), .B(n3050), .Z(c[1624]) );
  XNOR U3476 ( .A(a[1624]), .B(n3051), .Z(n3050) );
  IV U3477 ( .A(n3048), .Z(n3051) );
  XOR U3478 ( .A(n3052), .B(n3053), .Z(n3048) );
  ANDN U3479 ( .B(n3054), .A(n3055), .Z(n3052) );
  XNOR U3480 ( .A(b[1623]), .B(n3053), .Z(n3054) );
  XNOR U3481 ( .A(b[1623]), .B(n3055), .Z(c[1623]) );
  XNOR U3482 ( .A(a[1623]), .B(n3056), .Z(n3055) );
  IV U3483 ( .A(n3053), .Z(n3056) );
  XOR U3484 ( .A(n3057), .B(n3058), .Z(n3053) );
  ANDN U3485 ( .B(n3059), .A(n3060), .Z(n3057) );
  XNOR U3486 ( .A(b[1622]), .B(n3058), .Z(n3059) );
  XNOR U3487 ( .A(b[1622]), .B(n3060), .Z(c[1622]) );
  XNOR U3488 ( .A(a[1622]), .B(n3061), .Z(n3060) );
  IV U3489 ( .A(n3058), .Z(n3061) );
  XOR U3490 ( .A(n3062), .B(n3063), .Z(n3058) );
  ANDN U3491 ( .B(n3064), .A(n3065), .Z(n3062) );
  XNOR U3492 ( .A(b[1621]), .B(n3063), .Z(n3064) );
  XNOR U3493 ( .A(b[1621]), .B(n3065), .Z(c[1621]) );
  XNOR U3494 ( .A(a[1621]), .B(n3066), .Z(n3065) );
  IV U3495 ( .A(n3063), .Z(n3066) );
  XOR U3496 ( .A(n3067), .B(n3068), .Z(n3063) );
  ANDN U3497 ( .B(n3069), .A(n3070), .Z(n3067) );
  XNOR U3498 ( .A(b[1620]), .B(n3068), .Z(n3069) );
  XNOR U3499 ( .A(b[1620]), .B(n3070), .Z(c[1620]) );
  XNOR U3500 ( .A(a[1620]), .B(n3071), .Z(n3070) );
  IV U3501 ( .A(n3068), .Z(n3071) );
  XOR U3502 ( .A(n3072), .B(n3073), .Z(n3068) );
  ANDN U3503 ( .B(n3074), .A(n3075), .Z(n3072) );
  XNOR U3504 ( .A(b[1619]), .B(n3073), .Z(n3074) );
  XNOR U3505 ( .A(b[161]), .B(n3076), .Z(c[161]) );
  XNOR U3506 ( .A(b[1619]), .B(n3075), .Z(c[1619]) );
  XNOR U3507 ( .A(a[1619]), .B(n3077), .Z(n3075) );
  IV U3508 ( .A(n3073), .Z(n3077) );
  XOR U3509 ( .A(n3078), .B(n3079), .Z(n3073) );
  ANDN U3510 ( .B(n3080), .A(n3081), .Z(n3078) );
  XNOR U3511 ( .A(b[1618]), .B(n3079), .Z(n3080) );
  XNOR U3512 ( .A(b[1618]), .B(n3081), .Z(c[1618]) );
  XNOR U3513 ( .A(a[1618]), .B(n3082), .Z(n3081) );
  IV U3514 ( .A(n3079), .Z(n3082) );
  XOR U3515 ( .A(n3083), .B(n3084), .Z(n3079) );
  ANDN U3516 ( .B(n3085), .A(n3086), .Z(n3083) );
  XNOR U3517 ( .A(b[1617]), .B(n3084), .Z(n3085) );
  XNOR U3518 ( .A(b[1617]), .B(n3086), .Z(c[1617]) );
  XNOR U3519 ( .A(a[1617]), .B(n3087), .Z(n3086) );
  IV U3520 ( .A(n3084), .Z(n3087) );
  XOR U3521 ( .A(n3088), .B(n3089), .Z(n3084) );
  ANDN U3522 ( .B(n3090), .A(n3091), .Z(n3088) );
  XNOR U3523 ( .A(b[1616]), .B(n3089), .Z(n3090) );
  XNOR U3524 ( .A(b[1616]), .B(n3091), .Z(c[1616]) );
  XNOR U3525 ( .A(a[1616]), .B(n3092), .Z(n3091) );
  IV U3526 ( .A(n3089), .Z(n3092) );
  XOR U3527 ( .A(n3093), .B(n3094), .Z(n3089) );
  ANDN U3528 ( .B(n3095), .A(n3096), .Z(n3093) );
  XNOR U3529 ( .A(b[1615]), .B(n3094), .Z(n3095) );
  XNOR U3530 ( .A(b[1615]), .B(n3096), .Z(c[1615]) );
  XNOR U3531 ( .A(a[1615]), .B(n3097), .Z(n3096) );
  IV U3532 ( .A(n3094), .Z(n3097) );
  XOR U3533 ( .A(n3098), .B(n3099), .Z(n3094) );
  ANDN U3534 ( .B(n3100), .A(n3101), .Z(n3098) );
  XNOR U3535 ( .A(b[1614]), .B(n3099), .Z(n3100) );
  XNOR U3536 ( .A(b[1614]), .B(n3101), .Z(c[1614]) );
  XNOR U3537 ( .A(a[1614]), .B(n3102), .Z(n3101) );
  IV U3538 ( .A(n3099), .Z(n3102) );
  XOR U3539 ( .A(n3103), .B(n3104), .Z(n3099) );
  ANDN U3540 ( .B(n3105), .A(n3106), .Z(n3103) );
  XNOR U3541 ( .A(b[1613]), .B(n3104), .Z(n3105) );
  XNOR U3542 ( .A(b[1613]), .B(n3106), .Z(c[1613]) );
  XNOR U3543 ( .A(a[1613]), .B(n3107), .Z(n3106) );
  IV U3544 ( .A(n3104), .Z(n3107) );
  XOR U3545 ( .A(n3108), .B(n3109), .Z(n3104) );
  ANDN U3546 ( .B(n3110), .A(n3111), .Z(n3108) );
  XNOR U3547 ( .A(b[1612]), .B(n3109), .Z(n3110) );
  XNOR U3548 ( .A(b[1612]), .B(n3111), .Z(c[1612]) );
  XNOR U3549 ( .A(a[1612]), .B(n3112), .Z(n3111) );
  IV U3550 ( .A(n3109), .Z(n3112) );
  XOR U3551 ( .A(n3113), .B(n3114), .Z(n3109) );
  ANDN U3552 ( .B(n3115), .A(n3116), .Z(n3113) );
  XNOR U3553 ( .A(b[1611]), .B(n3114), .Z(n3115) );
  XNOR U3554 ( .A(b[1611]), .B(n3116), .Z(c[1611]) );
  XNOR U3555 ( .A(a[1611]), .B(n3117), .Z(n3116) );
  IV U3556 ( .A(n3114), .Z(n3117) );
  XOR U3557 ( .A(n3118), .B(n3119), .Z(n3114) );
  ANDN U3558 ( .B(n3120), .A(n3121), .Z(n3118) );
  XNOR U3559 ( .A(b[1610]), .B(n3119), .Z(n3120) );
  XNOR U3560 ( .A(b[1610]), .B(n3121), .Z(c[1610]) );
  XNOR U3561 ( .A(a[1610]), .B(n3122), .Z(n3121) );
  IV U3562 ( .A(n3119), .Z(n3122) );
  XOR U3563 ( .A(n3123), .B(n3124), .Z(n3119) );
  ANDN U3564 ( .B(n3125), .A(n3126), .Z(n3123) );
  XNOR U3565 ( .A(b[1609]), .B(n3124), .Z(n3125) );
  XNOR U3566 ( .A(b[160]), .B(n3127), .Z(c[160]) );
  XNOR U3567 ( .A(b[1609]), .B(n3126), .Z(c[1609]) );
  XNOR U3568 ( .A(a[1609]), .B(n3128), .Z(n3126) );
  IV U3569 ( .A(n3124), .Z(n3128) );
  XOR U3570 ( .A(n3129), .B(n3130), .Z(n3124) );
  ANDN U3571 ( .B(n3131), .A(n3132), .Z(n3129) );
  XNOR U3572 ( .A(b[1608]), .B(n3130), .Z(n3131) );
  XNOR U3573 ( .A(b[1608]), .B(n3132), .Z(c[1608]) );
  XNOR U3574 ( .A(a[1608]), .B(n3133), .Z(n3132) );
  IV U3575 ( .A(n3130), .Z(n3133) );
  XOR U3576 ( .A(n3134), .B(n3135), .Z(n3130) );
  ANDN U3577 ( .B(n3136), .A(n3137), .Z(n3134) );
  XNOR U3578 ( .A(b[1607]), .B(n3135), .Z(n3136) );
  XNOR U3579 ( .A(b[1607]), .B(n3137), .Z(c[1607]) );
  XNOR U3580 ( .A(a[1607]), .B(n3138), .Z(n3137) );
  IV U3581 ( .A(n3135), .Z(n3138) );
  XOR U3582 ( .A(n3139), .B(n3140), .Z(n3135) );
  ANDN U3583 ( .B(n3141), .A(n3142), .Z(n3139) );
  XNOR U3584 ( .A(b[1606]), .B(n3140), .Z(n3141) );
  XNOR U3585 ( .A(b[1606]), .B(n3142), .Z(c[1606]) );
  XNOR U3586 ( .A(a[1606]), .B(n3143), .Z(n3142) );
  IV U3587 ( .A(n3140), .Z(n3143) );
  XOR U3588 ( .A(n3144), .B(n3145), .Z(n3140) );
  ANDN U3589 ( .B(n3146), .A(n3147), .Z(n3144) );
  XNOR U3590 ( .A(b[1605]), .B(n3145), .Z(n3146) );
  XNOR U3591 ( .A(b[1605]), .B(n3147), .Z(c[1605]) );
  XNOR U3592 ( .A(a[1605]), .B(n3148), .Z(n3147) );
  IV U3593 ( .A(n3145), .Z(n3148) );
  XOR U3594 ( .A(n3149), .B(n3150), .Z(n3145) );
  ANDN U3595 ( .B(n3151), .A(n3152), .Z(n3149) );
  XNOR U3596 ( .A(b[1604]), .B(n3150), .Z(n3151) );
  XNOR U3597 ( .A(b[1604]), .B(n3152), .Z(c[1604]) );
  XNOR U3598 ( .A(a[1604]), .B(n3153), .Z(n3152) );
  IV U3599 ( .A(n3150), .Z(n3153) );
  XOR U3600 ( .A(n3154), .B(n3155), .Z(n3150) );
  ANDN U3601 ( .B(n3156), .A(n3157), .Z(n3154) );
  XNOR U3602 ( .A(b[1603]), .B(n3155), .Z(n3156) );
  XNOR U3603 ( .A(b[1603]), .B(n3157), .Z(c[1603]) );
  XNOR U3604 ( .A(a[1603]), .B(n3158), .Z(n3157) );
  IV U3605 ( .A(n3155), .Z(n3158) );
  XOR U3606 ( .A(n3159), .B(n3160), .Z(n3155) );
  ANDN U3607 ( .B(n3161), .A(n3162), .Z(n3159) );
  XNOR U3608 ( .A(b[1602]), .B(n3160), .Z(n3161) );
  XNOR U3609 ( .A(b[1602]), .B(n3162), .Z(c[1602]) );
  XNOR U3610 ( .A(a[1602]), .B(n3163), .Z(n3162) );
  IV U3611 ( .A(n3160), .Z(n3163) );
  XOR U3612 ( .A(n3164), .B(n3165), .Z(n3160) );
  ANDN U3613 ( .B(n3166), .A(n3167), .Z(n3164) );
  XNOR U3614 ( .A(b[1601]), .B(n3165), .Z(n3166) );
  XNOR U3615 ( .A(b[1601]), .B(n3167), .Z(c[1601]) );
  XNOR U3616 ( .A(a[1601]), .B(n3168), .Z(n3167) );
  IV U3617 ( .A(n3165), .Z(n3168) );
  XOR U3618 ( .A(n3169), .B(n3170), .Z(n3165) );
  ANDN U3619 ( .B(n3171), .A(n3172), .Z(n3169) );
  XNOR U3620 ( .A(b[1600]), .B(n3170), .Z(n3171) );
  XNOR U3621 ( .A(b[1600]), .B(n3172), .Z(c[1600]) );
  XNOR U3622 ( .A(a[1600]), .B(n3173), .Z(n3172) );
  IV U3623 ( .A(n3170), .Z(n3173) );
  XOR U3624 ( .A(n3174), .B(n3175), .Z(n3170) );
  ANDN U3625 ( .B(n3176), .A(n3177), .Z(n3174) );
  XNOR U3626 ( .A(b[1599]), .B(n3175), .Z(n3176) );
  XNOR U3627 ( .A(b[15]), .B(n3178), .Z(c[15]) );
  XNOR U3628 ( .A(b[159]), .B(n3179), .Z(c[159]) );
  XNOR U3629 ( .A(b[1599]), .B(n3177), .Z(c[1599]) );
  XNOR U3630 ( .A(a[1599]), .B(n3180), .Z(n3177) );
  IV U3631 ( .A(n3175), .Z(n3180) );
  XOR U3632 ( .A(n3181), .B(n3182), .Z(n3175) );
  ANDN U3633 ( .B(n3183), .A(n3184), .Z(n3181) );
  XNOR U3634 ( .A(b[1598]), .B(n3182), .Z(n3183) );
  XNOR U3635 ( .A(b[1598]), .B(n3184), .Z(c[1598]) );
  XNOR U3636 ( .A(a[1598]), .B(n3185), .Z(n3184) );
  IV U3637 ( .A(n3182), .Z(n3185) );
  XOR U3638 ( .A(n3186), .B(n3187), .Z(n3182) );
  ANDN U3639 ( .B(n3188), .A(n3189), .Z(n3186) );
  XNOR U3640 ( .A(b[1597]), .B(n3187), .Z(n3188) );
  XNOR U3641 ( .A(b[1597]), .B(n3189), .Z(c[1597]) );
  XNOR U3642 ( .A(a[1597]), .B(n3190), .Z(n3189) );
  IV U3643 ( .A(n3187), .Z(n3190) );
  XOR U3644 ( .A(n3191), .B(n3192), .Z(n3187) );
  ANDN U3645 ( .B(n3193), .A(n3194), .Z(n3191) );
  XNOR U3646 ( .A(b[1596]), .B(n3192), .Z(n3193) );
  XNOR U3647 ( .A(b[1596]), .B(n3194), .Z(c[1596]) );
  XNOR U3648 ( .A(a[1596]), .B(n3195), .Z(n3194) );
  IV U3649 ( .A(n3192), .Z(n3195) );
  XOR U3650 ( .A(n3196), .B(n3197), .Z(n3192) );
  ANDN U3651 ( .B(n3198), .A(n3199), .Z(n3196) );
  XNOR U3652 ( .A(b[1595]), .B(n3197), .Z(n3198) );
  XNOR U3653 ( .A(b[1595]), .B(n3199), .Z(c[1595]) );
  XNOR U3654 ( .A(a[1595]), .B(n3200), .Z(n3199) );
  IV U3655 ( .A(n3197), .Z(n3200) );
  XOR U3656 ( .A(n3201), .B(n3202), .Z(n3197) );
  ANDN U3657 ( .B(n3203), .A(n3204), .Z(n3201) );
  XNOR U3658 ( .A(b[1594]), .B(n3202), .Z(n3203) );
  XNOR U3659 ( .A(b[1594]), .B(n3204), .Z(c[1594]) );
  XNOR U3660 ( .A(a[1594]), .B(n3205), .Z(n3204) );
  IV U3661 ( .A(n3202), .Z(n3205) );
  XOR U3662 ( .A(n3206), .B(n3207), .Z(n3202) );
  ANDN U3663 ( .B(n3208), .A(n3209), .Z(n3206) );
  XNOR U3664 ( .A(b[1593]), .B(n3207), .Z(n3208) );
  XNOR U3665 ( .A(b[1593]), .B(n3209), .Z(c[1593]) );
  XNOR U3666 ( .A(a[1593]), .B(n3210), .Z(n3209) );
  IV U3667 ( .A(n3207), .Z(n3210) );
  XOR U3668 ( .A(n3211), .B(n3212), .Z(n3207) );
  ANDN U3669 ( .B(n3213), .A(n3214), .Z(n3211) );
  XNOR U3670 ( .A(b[1592]), .B(n3212), .Z(n3213) );
  XNOR U3671 ( .A(b[1592]), .B(n3214), .Z(c[1592]) );
  XNOR U3672 ( .A(a[1592]), .B(n3215), .Z(n3214) );
  IV U3673 ( .A(n3212), .Z(n3215) );
  XOR U3674 ( .A(n3216), .B(n3217), .Z(n3212) );
  ANDN U3675 ( .B(n3218), .A(n3219), .Z(n3216) );
  XNOR U3676 ( .A(b[1591]), .B(n3217), .Z(n3218) );
  XNOR U3677 ( .A(b[1591]), .B(n3219), .Z(c[1591]) );
  XNOR U3678 ( .A(a[1591]), .B(n3220), .Z(n3219) );
  IV U3679 ( .A(n3217), .Z(n3220) );
  XOR U3680 ( .A(n3221), .B(n3222), .Z(n3217) );
  ANDN U3681 ( .B(n3223), .A(n3224), .Z(n3221) );
  XNOR U3682 ( .A(b[1590]), .B(n3222), .Z(n3223) );
  XNOR U3683 ( .A(b[1590]), .B(n3224), .Z(c[1590]) );
  XNOR U3684 ( .A(a[1590]), .B(n3225), .Z(n3224) );
  IV U3685 ( .A(n3222), .Z(n3225) );
  XOR U3686 ( .A(n3226), .B(n3227), .Z(n3222) );
  ANDN U3687 ( .B(n3228), .A(n3229), .Z(n3226) );
  XNOR U3688 ( .A(b[1589]), .B(n3227), .Z(n3228) );
  XNOR U3689 ( .A(b[158]), .B(n3230), .Z(c[158]) );
  XNOR U3690 ( .A(b[1589]), .B(n3229), .Z(c[1589]) );
  XNOR U3691 ( .A(a[1589]), .B(n3231), .Z(n3229) );
  IV U3692 ( .A(n3227), .Z(n3231) );
  XOR U3693 ( .A(n3232), .B(n3233), .Z(n3227) );
  ANDN U3694 ( .B(n3234), .A(n3235), .Z(n3232) );
  XNOR U3695 ( .A(b[1588]), .B(n3233), .Z(n3234) );
  XNOR U3696 ( .A(b[1588]), .B(n3235), .Z(c[1588]) );
  XNOR U3697 ( .A(a[1588]), .B(n3236), .Z(n3235) );
  IV U3698 ( .A(n3233), .Z(n3236) );
  XOR U3699 ( .A(n3237), .B(n3238), .Z(n3233) );
  ANDN U3700 ( .B(n3239), .A(n3240), .Z(n3237) );
  XNOR U3701 ( .A(b[1587]), .B(n3238), .Z(n3239) );
  XNOR U3702 ( .A(b[1587]), .B(n3240), .Z(c[1587]) );
  XNOR U3703 ( .A(a[1587]), .B(n3241), .Z(n3240) );
  IV U3704 ( .A(n3238), .Z(n3241) );
  XOR U3705 ( .A(n3242), .B(n3243), .Z(n3238) );
  ANDN U3706 ( .B(n3244), .A(n3245), .Z(n3242) );
  XNOR U3707 ( .A(b[1586]), .B(n3243), .Z(n3244) );
  XNOR U3708 ( .A(b[1586]), .B(n3245), .Z(c[1586]) );
  XNOR U3709 ( .A(a[1586]), .B(n3246), .Z(n3245) );
  IV U3710 ( .A(n3243), .Z(n3246) );
  XOR U3711 ( .A(n3247), .B(n3248), .Z(n3243) );
  ANDN U3712 ( .B(n3249), .A(n3250), .Z(n3247) );
  XNOR U3713 ( .A(b[1585]), .B(n3248), .Z(n3249) );
  XNOR U3714 ( .A(b[1585]), .B(n3250), .Z(c[1585]) );
  XNOR U3715 ( .A(a[1585]), .B(n3251), .Z(n3250) );
  IV U3716 ( .A(n3248), .Z(n3251) );
  XOR U3717 ( .A(n3252), .B(n3253), .Z(n3248) );
  ANDN U3718 ( .B(n3254), .A(n3255), .Z(n3252) );
  XNOR U3719 ( .A(b[1584]), .B(n3253), .Z(n3254) );
  XNOR U3720 ( .A(b[1584]), .B(n3255), .Z(c[1584]) );
  XNOR U3721 ( .A(a[1584]), .B(n3256), .Z(n3255) );
  IV U3722 ( .A(n3253), .Z(n3256) );
  XOR U3723 ( .A(n3257), .B(n3258), .Z(n3253) );
  ANDN U3724 ( .B(n3259), .A(n3260), .Z(n3257) );
  XNOR U3725 ( .A(b[1583]), .B(n3258), .Z(n3259) );
  XNOR U3726 ( .A(b[1583]), .B(n3260), .Z(c[1583]) );
  XNOR U3727 ( .A(a[1583]), .B(n3261), .Z(n3260) );
  IV U3728 ( .A(n3258), .Z(n3261) );
  XOR U3729 ( .A(n3262), .B(n3263), .Z(n3258) );
  ANDN U3730 ( .B(n3264), .A(n3265), .Z(n3262) );
  XNOR U3731 ( .A(b[1582]), .B(n3263), .Z(n3264) );
  XNOR U3732 ( .A(b[1582]), .B(n3265), .Z(c[1582]) );
  XNOR U3733 ( .A(a[1582]), .B(n3266), .Z(n3265) );
  IV U3734 ( .A(n3263), .Z(n3266) );
  XOR U3735 ( .A(n3267), .B(n3268), .Z(n3263) );
  ANDN U3736 ( .B(n3269), .A(n3270), .Z(n3267) );
  XNOR U3737 ( .A(b[1581]), .B(n3268), .Z(n3269) );
  XNOR U3738 ( .A(b[1581]), .B(n3270), .Z(c[1581]) );
  XNOR U3739 ( .A(a[1581]), .B(n3271), .Z(n3270) );
  IV U3740 ( .A(n3268), .Z(n3271) );
  XOR U3741 ( .A(n3272), .B(n3273), .Z(n3268) );
  ANDN U3742 ( .B(n3274), .A(n3275), .Z(n3272) );
  XNOR U3743 ( .A(b[1580]), .B(n3273), .Z(n3274) );
  XNOR U3744 ( .A(b[1580]), .B(n3275), .Z(c[1580]) );
  XNOR U3745 ( .A(a[1580]), .B(n3276), .Z(n3275) );
  IV U3746 ( .A(n3273), .Z(n3276) );
  XOR U3747 ( .A(n3277), .B(n3278), .Z(n3273) );
  ANDN U3748 ( .B(n3279), .A(n3280), .Z(n3277) );
  XNOR U3749 ( .A(b[1579]), .B(n3278), .Z(n3279) );
  XNOR U3750 ( .A(b[157]), .B(n3281), .Z(c[157]) );
  XNOR U3751 ( .A(b[1579]), .B(n3280), .Z(c[1579]) );
  XNOR U3752 ( .A(a[1579]), .B(n3282), .Z(n3280) );
  IV U3753 ( .A(n3278), .Z(n3282) );
  XOR U3754 ( .A(n3283), .B(n3284), .Z(n3278) );
  ANDN U3755 ( .B(n3285), .A(n3286), .Z(n3283) );
  XNOR U3756 ( .A(b[1578]), .B(n3284), .Z(n3285) );
  XNOR U3757 ( .A(b[1578]), .B(n3286), .Z(c[1578]) );
  XNOR U3758 ( .A(a[1578]), .B(n3287), .Z(n3286) );
  IV U3759 ( .A(n3284), .Z(n3287) );
  XOR U3760 ( .A(n3288), .B(n3289), .Z(n3284) );
  ANDN U3761 ( .B(n3290), .A(n3291), .Z(n3288) );
  XNOR U3762 ( .A(b[1577]), .B(n3289), .Z(n3290) );
  XNOR U3763 ( .A(b[1577]), .B(n3291), .Z(c[1577]) );
  XNOR U3764 ( .A(a[1577]), .B(n3292), .Z(n3291) );
  IV U3765 ( .A(n3289), .Z(n3292) );
  XOR U3766 ( .A(n3293), .B(n3294), .Z(n3289) );
  ANDN U3767 ( .B(n3295), .A(n3296), .Z(n3293) );
  XNOR U3768 ( .A(b[1576]), .B(n3294), .Z(n3295) );
  XNOR U3769 ( .A(b[1576]), .B(n3296), .Z(c[1576]) );
  XNOR U3770 ( .A(a[1576]), .B(n3297), .Z(n3296) );
  IV U3771 ( .A(n3294), .Z(n3297) );
  XOR U3772 ( .A(n3298), .B(n3299), .Z(n3294) );
  ANDN U3773 ( .B(n3300), .A(n3301), .Z(n3298) );
  XNOR U3774 ( .A(b[1575]), .B(n3299), .Z(n3300) );
  XNOR U3775 ( .A(b[1575]), .B(n3301), .Z(c[1575]) );
  XNOR U3776 ( .A(a[1575]), .B(n3302), .Z(n3301) );
  IV U3777 ( .A(n3299), .Z(n3302) );
  XOR U3778 ( .A(n3303), .B(n3304), .Z(n3299) );
  ANDN U3779 ( .B(n3305), .A(n3306), .Z(n3303) );
  XNOR U3780 ( .A(b[1574]), .B(n3304), .Z(n3305) );
  XNOR U3781 ( .A(b[1574]), .B(n3306), .Z(c[1574]) );
  XNOR U3782 ( .A(a[1574]), .B(n3307), .Z(n3306) );
  IV U3783 ( .A(n3304), .Z(n3307) );
  XOR U3784 ( .A(n3308), .B(n3309), .Z(n3304) );
  ANDN U3785 ( .B(n3310), .A(n3311), .Z(n3308) );
  XNOR U3786 ( .A(b[1573]), .B(n3309), .Z(n3310) );
  XNOR U3787 ( .A(b[1573]), .B(n3311), .Z(c[1573]) );
  XNOR U3788 ( .A(a[1573]), .B(n3312), .Z(n3311) );
  IV U3789 ( .A(n3309), .Z(n3312) );
  XOR U3790 ( .A(n3313), .B(n3314), .Z(n3309) );
  ANDN U3791 ( .B(n3315), .A(n3316), .Z(n3313) );
  XNOR U3792 ( .A(b[1572]), .B(n3314), .Z(n3315) );
  XNOR U3793 ( .A(b[1572]), .B(n3316), .Z(c[1572]) );
  XNOR U3794 ( .A(a[1572]), .B(n3317), .Z(n3316) );
  IV U3795 ( .A(n3314), .Z(n3317) );
  XOR U3796 ( .A(n3318), .B(n3319), .Z(n3314) );
  ANDN U3797 ( .B(n3320), .A(n3321), .Z(n3318) );
  XNOR U3798 ( .A(b[1571]), .B(n3319), .Z(n3320) );
  XNOR U3799 ( .A(b[1571]), .B(n3321), .Z(c[1571]) );
  XNOR U3800 ( .A(a[1571]), .B(n3322), .Z(n3321) );
  IV U3801 ( .A(n3319), .Z(n3322) );
  XOR U3802 ( .A(n3323), .B(n3324), .Z(n3319) );
  ANDN U3803 ( .B(n3325), .A(n3326), .Z(n3323) );
  XNOR U3804 ( .A(b[1570]), .B(n3324), .Z(n3325) );
  XNOR U3805 ( .A(b[1570]), .B(n3326), .Z(c[1570]) );
  XNOR U3806 ( .A(a[1570]), .B(n3327), .Z(n3326) );
  IV U3807 ( .A(n3324), .Z(n3327) );
  XOR U3808 ( .A(n3328), .B(n3329), .Z(n3324) );
  ANDN U3809 ( .B(n3330), .A(n3331), .Z(n3328) );
  XNOR U3810 ( .A(b[1569]), .B(n3329), .Z(n3330) );
  XNOR U3811 ( .A(b[156]), .B(n3332), .Z(c[156]) );
  XNOR U3812 ( .A(b[1569]), .B(n3331), .Z(c[1569]) );
  XNOR U3813 ( .A(a[1569]), .B(n3333), .Z(n3331) );
  IV U3814 ( .A(n3329), .Z(n3333) );
  XOR U3815 ( .A(n3334), .B(n3335), .Z(n3329) );
  ANDN U3816 ( .B(n3336), .A(n3337), .Z(n3334) );
  XNOR U3817 ( .A(b[1568]), .B(n3335), .Z(n3336) );
  XNOR U3818 ( .A(b[1568]), .B(n3337), .Z(c[1568]) );
  XNOR U3819 ( .A(a[1568]), .B(n3338), .Z(n3337) );
  IV U3820 ( .A(n3335), .Z(n3338) );
  XOR U3821 ( .A(n3339), .B(n3340), .Z(n3335) );
  ANDN U3822 ( .B(n3341), .A(n3342), .Z(n3339) );
  XNOR U3823 ( .A(b[1567]), .B(n3340), .Z(n3341) );
  XNOR U3824 ( .A(b[1567]), .B(n3342), .Z(c[1567]) );
  XNOR U3825 ( .A(a[1567]), .B(n3343), .Z(n3342) );
  IV U3826 ( .A(n3340), .Z(n3343) );
  XOR U3827 ( .A(n3344), .B(n3345), .Z(n3340) );
  ANDN U3828 ( .B(n3346), .A(n3347), .Z(n3344) );
  XNOR U3829 ( .A(b[1566]), .B(n3345), .Z(n3346) );
  XNOR U3830 ( .A(b[1566]), .B(n3347), .Z(c[1566]) );
  XNOR U3831 ( .A(a[1566]), .B(n3348), .Z(n3347) );
  IV U3832 ( .A(n3345), .Z(n3348) );
  XOR U3833 ( .A(n3349), .B(n3350), .Z(n3345) );
  ANDN U3834 ( .B(n3351), .A(n3352), .Z(n3349) );
  XNOR U3835 ( .A(b[1565]), .B(n3350), .Z(n3351) );
  XNOR U3836 ( .A(b[1565]), .B(n3352), .Z(c[1565]) );
  XNOR U3837 ( .A(a[1565]), .B(n3353), .Z(n3352) );
  IV U3838 ( .A(n3350), .Z(n3353) );
  XOR U3839 ( .A(n3354), .B(n3355), .Z(n3350) );
  ANDN U3840 ( .B(n3356), .A(n3357), .Z(n3354) );
  XNOR U3841 ( .A(b[1564]), .B(n3355), .Z(n3356) );
  XNOR U3842 ( .A(b[1564]), .B(n3357), .Z(c[1564]) );
  XNOR U3843 ( .A(a[1564]), .B(n3358), .Z(n3357) );
  IV U3844 ( .A(n3355), .Z(n3358) );
  XOR U3845 ( .A(n3359), .B(n3360), .Z(n3355) );
  ANDN U3846 ( .B(n3361), .A(n3362), .Z(n3359) );
  XNOR U3847 ( .A(b[1563]), .B(n3360), .Z(n3361) );
  XNOR U3848 ( .A(b[1563]), .B(n3362), .Z(c[1563]) );
  XNOR U3849 ( .A(a[1563]), .B(n3363), .Z(n3362) );
  IV U3850 ( .A(n3360), .Z(n3363) );
  XOR U3851 ( .A(n3364), .B(n3365), .Z(n3360) );
  ANDN U3852 ( .B(n3366), .A(n3367), .Z(n3364) );
  XNOR U3853 ( .A(b[1562]), .B(n3365), .Z(n3366) );
  XNOR U3854 ( .A(b[1562]), .B(n3367), .Z(c[1562]) );
  XNOR U3855 ( .A(a[1562]), .B(n3368), .Z(n3367) );
  IV U3856 ( .A(n3365), .Z(n3368) );
  XOR U3857 ( .A(n3369), .B(n3370), .Z(n3365) );
  ANDN U3858 ( .B(n3371), .A(n3372), .Z(n3369) );
  XNOR U3859 ( .A(b[1561]), .B(n3370), .Z(n3371) );
  XNOR U3860 ( .A(b[1561]), .B(n3372), .Z(c[1561]) );
  XNOR U3861 ( .A(a[1561]), .B(n3373), .Z(n3372) );
  IV U3862 ( .A(n3370), .Z(n3373) );
  XOR U3863 ( .A(n3374), .B(n3375), .Z(n3370) );
  ANDN U3864 ( .B(n3376), .A(n3377), .Z(n3374) );
  XNOR U3865 ( .A(b[1560]), .B(n3375), .Z(n3376) );
  XNOR U3866 ( .A(b[1560]), .B(n3377), .Z(c[1560]) );
  XNOR U3867 ( .A(a[1560]), .B(n3378), .Z(n3377) );
  IV U3868 ( .A(n3375), .Z(n3378) );
  XOR U3869 ( .A(n3379), .B(n3380), .Z(n3375) );
  ANDN U3870 ( .B(n3381), .A(n3382), .Z(n3379) );
  XNOR U3871 ( .A(b[1559]), .B(n3380), .Z(n3381) );
  XNOR U3872 ( .A(b[155]), .B(n3383), .Z(c[155]) );
  XNOR U3873 ( .A(b[1559]), .B(n3382), .Z(c[1559]) );
  XNOR U3874 ( .A(a[1559]), .B(n3384), .Z(n3382) );
  IV U3875 ( .A(n3380), .Z(n3384) );
  XOR U3876 ( .A(n3385), .B(n3386), .Z(n3380) );
  ANDN U3877 ( .B(n3387), .A(n3388), .Z(n3385) );
  XNOR U3878 ( .A(b[1558]), .B(n3386), .Z(n3387) );
  XNOR U3879 ( .A(b[1558]), .B(n3388), .Z(c[1558]) );
  XNOR U3880 ( .A(a[1558]), .B(n3389), .Z(n3388) );
  IV U3881 ( .A(n3386), .Z(n3389) );
  XOR U3882 ( .A(n3390), .B(n3391), .Z(n3386) );
  ANDN U3883 ( .B(n3392), .A(n3393), .Z(n3390) );
  XNOR U3884 ( .A(b[1557]), .B(n3391), .Z(n3392) );
  XNOR U3885 ( .A(b[1557]), .B(n3393), .Z(c[1557]) );
  XNOR U3886 ( .A(a[1557]), .B(n3394), .Z(n3393) );
  IV U3887 ( .A(n3391), .Z(n3394) );
  XOR U3888 ( .A(n3395), .B(n3396), .Z(n3391) );
  ANDN U3889 ( .B(n3397), .A(n3398), .Z(n3395) );
  XNOR U3890 ( .A(b[1556]), .B(n3396), .Z(n3397) );
  XNOR U3891 ( .A(b[1556]), .B(n3398), .Z(c[1556]) );
  XNOR U3892 ( .A(a[1556]), .B(n3399), .Z(n3398) );
  IV U3893 ( .A(n3396), .Z(n3399) );
  XOR U3894 ( .A(n3400), .B(n3401), .Z(n3396) );
  ANDN U3895 ( .B(n3402), .A(n3403), .Z(n3400) );
  XNOR U3896 ( .A(b[1555]), .B(n3401), .Z(n3402) );
  XNOR U3897 ( .A(b[1555]), .B(n3403), .Z(c[1555]) );
  XNOR U3898 ( .A(a[1555]), .B(n3404), .Z(n3403) );
  IV U3899 ( .A(n3401), .Z(n3404) );
  XOR U3900 ( .A(n3405), .B(n3406), .Z(n3401) );
  ANDN U3901 ( .B(n3407), .A(n3408), .Z(n3405) );
  XNOR U3902 ( .A(b[1554]), .B(n3406), .Z(n3407) );
  XNOR U3903 ( .A(b[1554]), .B(n3408), .Z(c[1554]) );
  XNOR U3904 ( .A(a[1554]), .B(n3409), .Z(n3408) );
  IV U3905 ( .A(n3406), .Z(n3409) );
  XOR U3906 ( .A(n3410), .B(n3411), .Z(n3406) );
  ANDN U3907 ( .B(n3412), .A(n3413), .Z(n3410) );
  XNOR U3908 ( .A(b[1553]), .B(n3411), .Z(n3412) );
  XNOR U3909 ( .A(b[1553]), .B(n3413), .Z(c[1553]) );
  XNOR U3910 ( .A(a[1553]), .B(n3414), .Z(n3413) );
  IV U3911 ( .A(n3411), .Z(n3414) );
  XOR U3912 ( .A(n3415), .B(n3416), .Z(n3411) );
  ANDN U3913 ( .B(n3417), .A(n3418), .Z(n3415) );
  XNOR U3914 ( .A(b[1552]), .B(n3416), .Z(n3417) );
  XNOR U3915 ( .A(b[1552]), .B(n3418), .Z(c[1552]) );
  XNOR U3916 ( .A(a[1552]), .B(n3419), .Z(n3418) );
  IV U3917 ( .A(n3416), .Z(n3419) );
  XOR U3918 ( .A(n3420), .B(n3421), .Z(n3416) );
  ANDN U3919 ( .B(n3422), .A(n3423), .Z(n3420) );
  XNOR U3920 ( .A(b[1551]), .B(n3421), .Z(n3422) );
  XNOR U3921 ( .A(b[1551]), .B(n3423), .Z(c[1551]) );
  XNOR U3922 ( .A(a[1551]), .B(n3424), .Z(n3423) );
  IV U3923 ( .A(n3421), .Z(n3424) );
  XOR U3924 ( .A(n3425), .B(n3426), .Z(n3421) );
  ANDN U3925 ( .B(n3427), .A(n3428), .Z(n3425) );
  XNOR U3926 ( .A(b[1550]), .B(n3426), .Z(n3427) );
  XNOR U3927 ( .A(b[1550]), .B(n3428), .Z(c[1550]) );
  XNOR U3928 ( .A(a[1550]), .B(n3429), .Z(n3428) );
  IV U3929 ( .A(n3426), .Z(n3429) );
  XOR U3930 ( .A(n3430), .B(n3431), .Z(n3426) );
  ANDN U3931 ( .B(n3432), .A(n3433), .Z(n3430) );
  XNOR U3932 ( .A(b[1549]), .B(n3431), .Z(n3432) );
  XNOR U3933 ( .A(b[154]), .B(n3434), .Z(c[154]) );
  XNOR U3934 ( .A(b[1549]), .B(n3433), .Z(c[1549]) );
  XNOR U3935 ( .A(a[1549]), .B(n3435), .Z(n3433) );
  IV U3936 ( .A(n3431), .Z(n3435) );
  XOR U3937 ( .A(n3436), .B(n3437), .Z(n3431) );
  ANDN U3938 ( .B(n3438), .A(n3439), .Z(n3436) );
  XNOR U3939 ( .A(b[1548]), .B(n3437), .Z(n3438) );
  XNOR U3940 ( .A(b[1548]), .B(n3439), .Z(c[1548]) );
  XNOR U3941 ( .A(a[1548]), .B(n3440), .Z(n3439) );
  IV U3942 ( .A(n3437), .Z(n3440) );
  XOR U3943 ( .A(n3441), .B(n3442), .Z(n3437) );
  ANDN U3944 ( .B(n3443), .A(n3444), .Z(n3441) );
  XNOR U3945 ( .A(b[1547]), .B(n3442), .Z(n3443) );
  XNOR U3946 ( .A(b[1547]), .B(n3444), .Z(c[1547]) );
  XNOR U3947 ( .A(a[1547]), .B(n3445), .Z(n3444) );
  IV U3948 ( .A(n3442), .Z(n3445) );
  XOR U3949 ( .A(n3446), .B(n3447), .Z(n3442) );
  ANDN U3950 ( .B(n3448), .A(n3449), .Z(n3446) );
  XNOR U3951 ( .A(b[1546]), .B(n3447), .Z(n3448) );
  XNOR U3952 ( .A(b[1546]), .B(n3449), .Z(c[1546]) );
  XNOR U3953 ( .A(a[1546]), .B(n3450), .Z(n3449) );
  IV U3954 ( .A(n3447), .Z(n3450) );
  XOR U3955 ( .A(n3451), .B(n3452), .Z(n3447) );
  ANDN U3956 ( .B(n3453), .A(n3454), .Z(n3451) );
  XNOR U3957 ( .A(b[1545]), .B(n3452), .Z(n3453) );
  XNOR U3958 ( .A(b[1545]), .B(n3454), .Z(c[1545]) );
  XNOR U3959 ( .A(a[1545]), .B(n3455), .Z(n3454) );
  IV U3960 ( .A(n3452), .Z(n3455) );
  XOR U3961 ( .A(n3456), .B(n3457), .Z(n3452) );
  ANDN U3962 ( .B(n3458), .A(n3459), .Z(n3456) );
  XNOR U3963 ( .A(b[1544]), .B(n3457), .Z(n3458) );
  XNOR U3964 ( .A(b[1544]), .B(n3459), .Z(c[1544]) );
  XNOR U3965 ( .A(a[1544]), .B(n3460), .Z(n3459) );
  IV U3966 ( .A(n3457), .Z(n3460) );
  XOR U3967 ( .A(n3461), .B(n3462), .Z(n3457) );
  ANDN U3968 ( .B(n3463), .A(n3464), .Z(n3461) );
  XNOR U3969 ( .A(b[1543]), .B(n3462), .Z(n3463) );
  XNOR U3970 ( .A(b[1543]), .B(n3464), .Z(c[1543]) );
  XNOR U3971 ( .A(a[1543]), .B(n3465), .Z(n3464) );
  IV U3972 ( .A(n3462), .Z(n3465) );
  XOR U3973 ( .A(n3466), .B(n3467), .Z(n3462) );
  ANDN U3974 ( .B(n3468), .A(n3469), .Z(n3466) );
  XNOR U3975 ( .A(b[1542]), .B(n3467), .Z(n3468) );
  XNOR U3976 ( .A(b[1542]), .B(n3469), .Z(c[1542]) );
  XNOR U3977 ( .A(a[1542]), .B(n3470), .Z(n3469) );
  IV U3978 ( .A(n3467), .Z(n3470) );
  XOR U3979 ( .A(n3471), .B(n3472), .Z(n3467) );
  ANDN U3980 ( .B(n3473), .A(n3474), .Z(n3471) );
  XNOR U3981 ( .A(b[1541]), .B(n3472), .Z(n3473) );
  XNOR U3982 ( .A(b[1541]), .B(n3474), .Z(c[1541]) );
  XNOR U3983 ( .A(a[1541]), .B(n3475), .Z(n3474) );
  IV U3984 ( .A(n3472), .Z(n3475) );
  XOR U3985 ( .A(n3476), .B(n3477), .Z(n3472) );
  ANDN U3986 ( .B(n3478), .A(n3479), .Z(n3476) );
  XNOR U3987 ( .A(b[1540]), .B(n3477), .Z(n3478) );
  XNOR U3988 ( .A(b[1540]), .B(n3479), .Z(c[1540]) );
  XNOR U3989 ( .A(a[1540]), .B(n3480), .Z(n3479) );
  IV U3990 ( .A(n3477), .Z(n3480) );
  XOR U3991 ( .A(n3481), .B(n3482), .Z(n3477) );
  ANDN U3992 ( .B(n3483), .A(n3484), .Z(n3481) );
  XNOR U3993 ( .A(b[1539]), .B(n3482), .Z(n3483) );
  XNOR U3994 ( .A(b[153]), .B(n3485), .Z(c[153]) );
  XNOR U3995 ( .A(b[1539]), .B(n3484), .Z(c[1539]) );
  XNOR U3996 ( .A(a[1539]), .B(n3486), .Z(n3484) );
  IV U3997 ( .A(n3482), .Z(n3486) );
  XOR U3998 ( .A(n3487), .B(n3488), .Z(n3482) );
  ANDN U3999 ( .B(n3489), .A(n3490), .Z(n3487) );
  XNOR U4000 ( .A(b[1538]), .B(n3488), .Z(n3489) );
  XNOR U4001 ( .A(b[1538]), .B(n3490), .Z(c[1538]) );
  XNOR U4002 ( .A(a[1538]), .B(n3491), .Z(n3490) );
  IV U4003 ( .A(n3488), .Z(n3491) );
  XOR U4004 ( .A(n3492), .B(n3493), .Z(n3488) );
  ANDN U4005 ( .B(n3494), .A(n3495), .Z(n3492) );
  XNOR U4006 ( .A(b[1537]), .B(n3493), .Z(n3494) );
  XNOR U4007 ( .A(b[1537]), .B(n3495), .Z(c[1537]) );
  XNOR U4008 ( .A(a[1537]), .B(n3496), .Z(n3495) );
  IV U4009 ( .A(n3493), .Z(n3496) );
  XOR U4010 ( .A(n3497), .B(n3498), .Z(n3493) );
  ANDN U4011 ( .B(n3499), .A(n3500), .Z(n3497) );
  XNOR U4012 ( .A(b[1536]), .B(n3498), .Z(n3499) );
  XNOR U4013 ( .A(b[1536]), .B(n3500), .Z(c[1536]) );
  XNOR U4014 ( .A(a[1536]), .B(n3501), .Z(n3500) );
  IV U4015 ( .A(n3498), .Z(n3501) );
  XOR U4016 ( .A(n3502), .B(n3503), .Z(n3498) );
  ANDN U4017 ( .B(n3504), .A(n3505), .Z(n3502) );
  XNOR U4018 ( .A(b[1535]), .B(n3503), .Z(n3504) );
  XNOR U4019 ( .A(b[1535]), .B(n3505), .Z(c[1535]) );
  XNOR U4020 ( .A(a[1535]), .B(n3506), .Z(n3505) );
  IV U4021 ( .A(n3503), .Z(n3506) );
  XOR U4022 ( .A(n3507), .B(n3508), .Z(n3503) );
  ANDN U4023 ( .B(n3509), .A(n3510), .Z(n3507) );
  XNOR U4024 ( .A(b[1534]), .B(n3508), .Z(n3509) );
  XNOR U4025 ( .A(b[1534]), .B(n3510), .Z(c[1534]) );
  XNOR U4026 ( .A(a[1534]), .B(n3511), .Z(n3510) );
  IV U4027 ( .A(n3508), .Z(n3511) );
  XOR U4028 ( .A(n3512), .B(n3513), .Z(n3508) );
  ANDN U4029 ( .B(n3514), .A(n3515), .Z(n3512) );
  XNOR U4030 ( .A(b[1533]), .B(n3513), .Z(n3514) );
  XNOR U4031 ( .A(b[1533]), .B(n3515), .Z(c[1533]) );
  XNOR U4032 ( .A(a[1533]), .B(n3516), .Z(n3515) );
  IV U4033 ( .A(n3513), .Z(n3516) );
  XOR U4034 ( .A(n3517), .B(n3518), .Z(n3513) );
  ANDN U4035 ( .B(n3519), .A(n3520), .Z(n3517) );
  XNOR U4036 ( .A(b[1532]), .B(n3518), .Z(n3519) );
  XNOR U4037 ( .A(b[1532]), .B(n3520), .Z(c[1532]) );
  XNOR U4038 ( .A(a[1532]), .B(n3521), .Z(n3520) );
  IV U4039 ( .A(n3518), .Z(n3521) );
  XOR U4040 ( .A(n3522), .B(n3523), .Z(n3518) );
  ANDN U4041 ( .B(n3524), .A(n3525), .Z(n3522) );
  XNOR U4042 ( .A(b[1531]), .B(n3523), .Z(n3524) );
  XNOR U4043 ( .A(b[1531]), .B(n3525), .Z(c[1531]) );
  XNOR U4044 ( .A(a[1531]), .B(n3526), .Z(n3525) );
  IV U4045 ( .A(n3523), .Z(n3526) );
  XOR U4046 ( .A(n3527), .B(n3528), .Z(n3523) );
  ANDN U4047 ( .B(n3529), .A(n3530), .Z(n3527) );
  XNOR U4048 ( .A(b[1530]), .B(n3528), .Z(n3529) );
  XNOR U4049 ( .A(b[1530]), .B(n3530), .Z(c[1530]) );
  XNOR U4050 ( .A(a[1530]), .B(n3531), .Z(n3530) );
  IV U4051 ( .A(n3528), .Z(n3531) );
  XOR U4052 ( .A(n3532), .B(n3533), .Z(n3528) );
  ANDN U4053 ( .B(n3534), .A(n3535), .Z(n3532) );
  XNOR U4054 ( .A(b[1529]), .B(n3533), .Z(n3534) );
  XNOR U4055 ( .A(b[152]), .B(n3536), .Z(c[152]) );
  XNOR U4056 ( .A(b[1529]), .B(n3535), .Z(c[1529]) );
  XNOR U4057 ( .A(a[1529]), .B(n3537), .Z(n3535) );
  IV U4058 ( .A(n3533), .Z(n3537) );
  XOR U4059 ( .A(n3538), .B(n3539), .Z(n3533) );
  ANDN U4060 ( .B(n3540), .A(n3541), .Z(n3538) );
  XNOR U4061 ( .A(b[1528]), .B(n3539), .Z(n3540) );
  XNOR U4062 ( .A(b[1528]), .B(n3541), .Z(c[1528]) );
  XNOR U4063 ( .A(a[1528]), .B(n3542), .Z(n3541) );
  IV U4064 ( .A(n3539), .Z(n3542) );
  XOR U4065 ( .A(n3543), .B(n3544), .Z(n3539) );
  ANDN U4066 ( .B(n3545), .A(n3546), .Z(n3543) );
  XNOR U4067 ( .A(b[1527]), .B(n3544), .Z(n3545) );
  XNOR U4068 ( .A(b[1527]), .B(n3546), .Z(c[1527]) );
  XNOR U4069 ( .A(a[1527]), .B(n3547), .Z(n3546) );
  IV U4070 ( .A(n3544), .Z(n3547) );
  XOR U4071 ( .A(n3548), .B(n3549), .Z(n3544) );
  ANDN U4072 ( .B(n3550), .A(n3551), .Z(n3548) );
  XNOR U4073 ( .A(b[1526]), .B(n3549), .Z(n3550) );
  XNOR U4074 ( .A(b[1526]), .B(n3551), .Z(c[1526]) );
  XNOR U4075 ( .A(a[1526]), .B(n3552), .Z(n3551) );
  IV U4076 ( .A(n3549), .Z(n3552) );
  XOR U4077 ( .A(n3553), .B(n3554), .Z(n3549) );
  ANDN U4078 ( .B(n3555), .A(n3556), .Z(n3553) );
  XNOR U4079 ( .A(b[1525]), .B(n3554), .Z(n3555) );
  XNOR U4080 ( .A(b[1525]), .B(n3556), .Z(c[1525]) );
  XNOR U4081 ( .A(a[1525]), .B(n3557), .Z(n3556) );
  IV U4082 ( .A(n3554), .Z(n3557) );
  XOR U4083 ( .A(n3558), .B(n3559), .Z(n3554) );
  ANDN U4084 ( .B(n3560), .A(n3561), .Z(n3558) );
  XNOR U4085 ( .A(b[1524]), .B(n3559), .Z(n3560) );
  XNOR U4086 ( .A(b[1524]), .B(n3561), .Z(c[1524]) );
  XNOR U4087 ( .A(a[1524]), .B(n3562), .Z(n3561) );
  IV U4088 ( .A(n3559), .Z(n3562) );
  XOR U4089 ( .A(n3563), .B(n3564), .Z(n3559) );
  ANDN U4090 ( .B(n3565), .A(n3566), .Z(n3563) );
  XNOR U4091 ( .A(b[1523]), .B(n3564), .Z(n3565) );
  XNOR U4092 ( .A(b[1523]), .B(n3566), .Z(c[1523]) );
  XNOR U4093 ( .A(a[1523]), .B(n3567), .Z(n3566) );
  IV U4094 ( .A(n3564), .Z(n3567) );
  XOR U4095 ( .A(n3568), .B(n3569), .Z(n3564) );
  ANDN U4096 ( .B(n3570), .A(n3571), .Z(n3568) );
  XNOR U4097 ( .A(b[1522]), .B(n3569), .Z(n3570) );
  XNOR U4098 ( .A(b[1522]), .B(n3571), .Z(c[1522]) );
  XNOR U4099 ( .A(a[1522]), .B(n3572), .Z(n3571) );
  IV U4100 ( .A(n3569), .Z(n3572) );
  XOR U4101 ( .A(n3573), .B(n3574), .Z(n3569) );
  ANDN U4102 ( .B(n3575), .A(n3576), .Z(n3573) );
  XNOR U4103 ( .A(b[1521]), .B(n3574), .Z(n3575) );
  XNOR U4104 ( .A(b[1521]), .B(n3576), .Z(c[1521]) );
  XNOR U4105 ( .A(a[1521]), .B(n3577), .Z(n3576) );
  IV U4106 ( .A(n3574), .Z(n3577) );
  XOR U4107 ( .A(n3578), .B(n3579), .Z(n3574) );
  ANDN U4108 ( .B(n3580), .A(n3581), .Z(n3578) );
  XNOR U4109 ( .A(b[1520]), .B(n3579), .Z(n3580) );
  XNOR U4110 ( .A(b[1520]), .B(n3581), .Z(c[1520]) );
  XNOR U4111 ( .A(a[1520]), .B(n3582), .Z(n3581) );
  IV U4112 ( .A(n3579), .Z(n3582) );
  XOR U4113 ( .A(n3583), .B(n3584), .Z(n3579) );
  ANDN U4114 ( .B(n3585), .A(n3586), .Z(n3583) );
  XNOR U4115 ( .A(b[1519]), .B(n3584), .Z(n3585) );
  XNOR U4116 ( .A(b[151]), .B(n3587), .Z(c[151]) );
  XNOR U4117 ( .A(b[1519]), .B(n3586), .Z(c[1519]) );
  XNOR U4118 ( .A(a[1519]), .B(n3588), .Z(n3586) );
  IV U4119 ( .A(n3584), .Z(n3588) );
  XOR U4120 ( .A(n3589), .B(n3590), .Z(n3584) );
  ANDN U4121 ( .B(n3591), .A(n3592), .Z(n3589) );
  XNOR U4122 ( .A(b[1518]), .B(n3590), .Z(n3591) );
  XNOR U4123 ( .A(b[1518]), .B(n3592), .Z(c[1518]) );
  XNOR U4124 ( .A(a[1518]), .B(n3593), .Z(n3592) );
  IV U4125 ( .A(n3590), .Z(n3593) );
  XOR U4126 ( .A(n3594), .B(n3595), .Z(n3590) );
  ANDN U4127 ( .B(n3596), .A(n3597), .Z(n3594) );
  XNOR U4128 ( .A(b[1517]), .B(n3595), .Z(n3596) );
  XNOR U4129 ( .A(b[1517]), .B(n3597), .Z(c[1517]) );
  XNOR U4130 ( .A(a[1517]), .B(n3598), .Z(n3597) );
  IV U4131 ( .A(n3595), .Z(n3598) );
  XOR U4132 ( .A(n3599), .B(n3600), .Z(n3595) );
  ANDN U4133 ( .B(n3601), .A(n3602), .Z(n3599) );
  XNOR U4134 ( .A(b[1516]), .B(n3600), .Z(n3601) );
  XNOR U4135 ( .A(b[1516]), .B(n3602), .Z(c[1516]) );
  XNOR U4136 ( .A(a[1516]), .B(n3603), .Z(n3602) );
  IV U4137 ( .A(n3600), .Z(n3603) );
  XOR U4138 ( .A(n3604), .B(n3605), .Z(n3600) );
  ANDN U4139 ( .B(n3606), .A(n3607), .Z(n3604) );
  XNOR U4140 ( .A(b[1515]), .B(n3605), .Z(n3606) );
  XNOR U4141 ( .A(b[1515]), .B(n3607), .Z(c[1515]) );
  XNOR U4142 ( .A(a[1515]), .B(n3608), .Z(n3607) );
  IV U4143 ( .A(n3605), .Z(n3608) );
  XOR U4144 ( .A(n3609), .B(n3610), .Z(n3605) );
  ANDN U4145 ( .B(n3611), .A(n3612), .Z(n3609) );
  XNOR U4146 ( .A(b[1514]), .B(n3610), .Z(n3611) );
  XNOR U4147 ( .A(b[1514]), .B(n3612), .Z(c[1514]) );
  XNOR U4148 ( .A(a[1514]), .B(n3613), .Z(n3612) );
  IV U4149 ( .A(n3610), .Z(n3613) );
  XOR U4150 ( .A(n3614), .B(n3615), .Z(n3610) );
  ANDN U4151 ( .B(n3616), .A(n3617), .Z(n3614) );
  XNOR U4152 ( .A(b[1513]), .B(n3615), .Z(n3616) );
  XNOR U4153 ( .A(b[1513]), .B(n3617), .Z(c[1513]) );
  XNOR U4154 ( .A(a[1513]), .B(n3618), .Z(n3617) );
  IV U4155 ( .A(n3615), .Z(n3618) );
  XOR U4156 ( .A(n3619), .B(n3620), .Z(n3615) );
  ANDN U4157 ( .B(n3621), .A(n3622), .Z(n3619) );
  XNOR U4158 ( .A(b[1512]), .B(n3620), .Z(n3621) );
  XNOR U4159 ( .A(b[1512]), .B(n3622), .Z(c[1512]) );
  XNOR U4160 ( .A(a[1512]), .B(n3623), .Z(n3622) );
  IV U4161 ( .A(n3620), .Z(n3623) );
  XOR U4162 ( .A(n3624), .B(n3625), .Z(n3620) );
  ANDN U4163 ( .B(n3626), .A(n3627), .Z(n3624) );
  XNOR U4164 ( .A(b[1511]), .B(n3625), .Z(n3626) );
  XNOR U4165 ( .A(b[1511]), .B(n3627), .Z(c[1511]) );
  XNOR U4166 ( .A(a[1511]), .B(n3628), .Z(n3627) );
  IV U4167 ( .A(n3625), .Z(n3628) );
  XOR U4168 ( .A(n3629), .B(n3630), .Z(n3625) );
  ANDN U4169 ( .B(n3631), .A(n3632), .Z(n3629) );
  XNOR U4170 ( .A(b[1510]), .B(n3630), .Z(n3631) );
  XNOR U4171 ( .A(b[1510]), .B(n3632), .Z(c[1510]) );
  XNOR U4172 ( .A(a[1510]), .B(n3633), .Z(n3632) );
  IV U4173 ( .A(n3630), .Z(n3633) );
  XOR U4174 ( .A(n3634), .B(n3635), .Z(n3630) );
  ANDN U4175 ( .B(n3636), .A(n3637), .Z(n3634) );
  XNOR U4176 ( .A(b[1509]), .B(n3635), .Z(n3636) );
  XNOR U4177 ( .A(b[150]), .B(n3638), .Z(c[150]) );
  XNOR U4178 ( .A(b[1509]), .B(n3637), .Z(c[1509]) );
  XNOR U4179 ( .A(a[1509]), .B(n3639), .Z(n3637) );
  IV U4180 ( .A(n3635), .Z(n3639) );
  XOR U4181 ( .A(n3640), .B(n3641), .Z(n3635) );
  ANDN U4182 ( .B(n3642), .A(n3643), .Z(n3640) );
  XNOR U4183 ( .A(b[1508]), .B(n3641), .Z(n3642) );
  XNOR U4184 ( .A(b[1508]), .B(n3643), .Z(c[1508]) );
  XNOR U4185 ( .A(a[1508]), .B(n3644), .Z(n3643) );
  IV U4186 ( .A(n3641), .Z(n3644) );
  XOR U4187 ( .A(n3645), .B(n3646), .Z(n3641) );
  ANDN U4188 ( .B(n3647), .A(n3648), .Z(n3645) );
  XNOR U4189 ( .A(b[1507]), .B(n3646), .Z(n3647) );
  XNOR U4190 ( .A(b[1507]), .B(n3648), .Z(c[1507]) );
  XNOR U4191 ( .A(a[1507]), .B(n3649), .Z(n3648) );
  IV U4192 ( .A(n3646), .Z(n3649) );
  XOR U4193 ( .A(n3650), .B(n3651), .Z(n3646) );
  ANDN U4194 ( .B(n3652), .A(n3653), .Z(n3650) );
  XNOR U4195 ( .A(b[1506]), .B(n3651), .Z(n3652) );
  XNOR U4196 ( .A(b[1506]), .B(n3653), .Z(c[1506]) );
  XNOR U4197 ( .A(a[1506]), .B(n3654), .Z(n3653) );
  IV U4198 ( .A(n3651), .Z(n3654) );
  XOR U4199 ( .A(n3655), .B(n3656), .Z(n3651) );
  ANDN U4200 ( .B(n3657), .A(n3658), .Z(n3655) );
  XNOR U4201 ( .A(b[1505]), .B(n3656), .Z(n3657) );
  XNOR U4202 ( .A(b[1505]), .B(n3658), .Z(c[1505]) );
  XNOR U4203 ( .A(a[1505]), .B(n3659), .Z(n3658) );
  IV U4204 ( .A(n3656), .Z(n3659) );
  XOR U4205 ( .A(n3660), .B(n3661), .Z(n3656) );
  ANDN U4206 ( .B(n3662), .A(n3663), .Z(n3660) );
  XNOR U4207 ( .A(b[1504]), .B(n3661), .Z(n3662) );
  XNOR U4208 ( .A(b[1504]), .B(n3663), .Z(c[1504]) );
  XNOR U4209 ( .A(a[1504]), .B(n3664), .Z(n3663) );
  IV U4210 ( .A(n3661), .Z(n3664) );
  XOR U4211 ( .A(n3665), .B(n3666), .Z(n3661) );
  ANDN U4212 ( .B(n3667), .A(n3668), .Z(n3665) );
  XNOR U4213 ( .A(b[1503]), .B(n3666), .Z(n3667) );
  XNOR U4214 ( .A(b[1503]), .B(n3668), .Z(c[1503]) );
  XNOR U4215 ( .A(a[1503]), .B(n3669), .Z(n3668) );
  IV U4216 ( .A(n3666), .Z(n3669) );
  XOR U4217 ( .A(n3670), .B(n3671), .Z(n3666) );
  ANDN U4218 ( .B(n3672), .A(n3673), .Z(n3670) );
  XNOR U4219 ( .A(b[1502]), .B(n3671), .Z(n3672) );
  XNOR U4220 ( .A(b[1502]), .B(n3673), .Z(c[1502]) );
  XNOR U4221 ( .A(a[1502]), .B(n3674), .Z(n3673) );
  IV U4222 ( .A(n3671), .Z(n3674) );
  XOR U4223 ( .A(n3675), .B(n3676), .Z(n3671) );
  ANDN U4224 ( .B(n3677), .A(n3678), .Z(n3675) );
  XNOR U4225 ( .A(b[1501]), .B(n3676), .Z(n3677) );
  XNOR U4226 ( .A(b[1501]), .B(n3678), .Z(c[1501]) );
  XNOR U4227 ( .A(a[1501]), .B(n3679), .Z(n3678) );
  IV U4228 ( .A(n3676), .Z(n3679) );
  XOR U4229 ( .A(n3680), .B(n3681), .Z(n3676) );
  ANDN U4230 ( .B(n3682), .A(n3683), .Z(n3680) );
  XNOR U4231 ( .A(b[1500]), .B(n3681), .Z(n3682) );
  XNOR U4232 ( .A(b[1500]), .B(n3683), .Z(c[1500]) );
  XNOR U4233 ( .A(a[1500]), .B(n3684), .Z(n3683) );
  IV U4234 ( .A(n3681), .Z(n3684) );
  XOR U4235 ( .A(n3685), .B(n3686), .Z(n3681) );
  ANDN U4236 ( .B(n3687), .A(n3688), .Z(n3685) );
  XNOR U4237 ( .A(b[1499]), .B(n3686), .Z(n3687) );
  XNOR U4238 ( .A(b[14]), .B(n3689), .Z(c[14]) );
  XNOR U4239 ( .A(b[149]), .B(n3690), .Z(c[149]) );
  XNOR U4240 ( .A(b[1499]), .B(n3688), .Z(c[1499]) );
  XNOR U4241 ( .A(a[1499]), .B(n3691), .Z(n3688) );
  IV U4242 ( .A(n3686), .Z(n3691) );
  XOR U4243 ( .A(n3692), .B(n3693), .Z(n3686) );
  ANDN U4244 ( .B(n3694), .A(n3695), .Z(n3692) );
  XNOR U4245 ( .A(b[1498]), .B(n3693), .Z(n3694) );
  XNOR U4246 ( .A(b[1498]), .B(n3695), .Z(c[1498]) );
  XNOR U4247 ( .A(a[1498]), .B(n3696), .Z(n3695) );
  IV U4248 ( .A(n3693), .Z(n3696) );
  XOR U4249 ( .A(n3697), .B(n3698), .Z(n3693) );
  ANDN U4250 ( .B(n3699), .A(n3700), .Z(n3697) );
  XNOR U4251 ( .A(b[1497]), .B(n3698), .Z(n3699) );
  XNOR U4252 ( .A(b[1497]), .B(n3700), .Z(c[1497]) );
  XNOR U4253 ( .A(a[1497]), .B(n3701), .Z(n3700) );
  IV U4254 ( .A(n3698), .Z(n3701) );
  XOR U4255 ( .A(n3702), .B(n3703), .Z(n3698) );
  ANDN U4256 ( .B(n3704), .A(n3705), .Z(n3702) );
  XNOR U4257 ( .A(b[1496]), .B(n3703), .Z(n3704) );
  XNOR U4258 ( .A(b[1496]), .B(n3705), .Z(c[1496]) );
  XNOR U4259 ( .A(a[1496]), .B(n3706), .Z(n3705) );
  IV U4260 ( .A(n3703), .Z(n3706) );
  XOR U4261 ( .A(n3707), .B(n3708), .Z(n3703) );
  ANDN U4262 ( .B(n3709), .A(n3710), .Z(n3707) );
  XNOR U4263 ( .A(b[1495]), .B(n3708), .Z(n3709) );
  XNOR U4264 ( .A(b[1495]), .B(n3710), .Z(c[1495]) );
  XNOR U4265 ( .A(a[1495]), .B(n3711), .Z(n3710) );
  IV U4266 ( .A(n3708), .Z(n3711) );
  XOR U4267 ( .A(n3712), .B(n3713), .Z(n3708) );
  ANDN U4268 ( .B(n3714), .A(n3715), .Z(n3712) );
  XNOR U4269 ( .A(b[1494]), .B(n3713), .Z(n3714) );
  XNOR U4270 ( .A(b[1494]), .B(n3715), .Z(c[1494]) );
  XNOR U4271 ( .A(a[1494]), .B(n3716), .Z(n3715) );
  IV U4272 ( .A(n3713), .Z(n3716) );
  XOR U4273 ( .A(n3717), .B(n3718), .Z(n3713) );
  ANDN U4274 ( .B(n3719), .A(n3720), .Z(n3717) );
  XNOR U4275 ( .A(b[1493]), .B(n3718), .Z(n3719) );
  XNOR U4276 ( .A(b[1493]), .B(n3720), .Z(c[1493]) );
  XNOR U4277 ( .A(a[1493]), .B(n3721), .Z(n3720) );
  IV U4278 ( .A(n3718), .Z(n3721) );
  XOR U4279 ( .A(n3722), .B(n3723), .Z(n3718) );
  ANDN U4280 ( .B(n3724), .A(n3725), .Z(n3722) );
  XNOR U4281 ( .A(b[1492]), .B(n3723), .Z(n3724) );
  XNOR U4282 ( .A(b[1492]), .B(n3725), .Z(c[1492]) );
  XNOR U4283 ( .A(a[1492]), .B(n3726), .Z(n3725) );
  IV U4284 ( .A(n3723), .Z(n3726) );
  XOR U4285 ( .A(n3727), .B(n3728), .Z(n3723) );
  ANDN U4286 ( .B(n3729), .A(n3730), .Z(n3727) );
  XNOR U4287 ( .A(b[1491]), .B(n3728), .Z(n3729) );
  XNOR U4288 ( .A(b[1491]), .B(n3730), .Z(c[1491]) );
  XNOR U4289 ( .A(a[1491]), .B(n3731), .Z(n3730) );
  IV U4290 ( .A(n3728), .Z(n3731) );
  XOR U4291 ( .A(n3732), .B(n3733), .Z(n3728) );
  ANDN U4292 ( .B(n3734), .A(n3735), .Z(n3732) );
  XNOR U4293 ( .A(b[1490]), .B(n3733), .Z(n3734) );
  XNOR U4294 ( .A(b[1490]), .B(n3735), .Z(c[1490]) );
  XNOR U4295 ( .A(a[1490]), .B(n3736), .Z(n3735) );
  IV U4296 ( .A(n3733), .Z(n3736) );
  XOR U4297 ( .A(n3737), .B(n3738), .Z(n3733) );
  ANDN U4298 ( .B(n3739), .A(n3740), .Z(n3737) );
  XNOR U4299 ( .A(b[1489]), .B(n3738), .Z(n3739) );
  XNOR U4300 ( .A(b[148]), .B(n3741), .Z(c[148]) );
  XNOR U4301 ( .A(b[1489]), .B(n3740), .Z(c[1489]) );
  XNOR U4302 ( .A(a[1489]), .B(n3742), .Z(n3740) );
  IV U4303 ( .A(n3738), .Z(n3742) );
  XOR U4304 ( .A(n3743), .B(n3744), .Z(n3738) );
  ANDN U4305 ( .B(n3745), .A(n3746), .Z(n3743) );
  XNOR U4306 ( .A(b[1488]), .B(n3744), .Z(n3745) );
  XNOR U4307 ( .A(b[1488]), .B(n3746), .Z(c[1488]) );
  XNOR U4308 ( .A(a[1488]), .B(n3747), .Z(n3746) );
  IV U4309 ( .A(n3744), .Z(n3747) );
  XOR U4310 ( .A(n3748), .B(n3749), .Z(n3744) );
  ANDN U4311 ( .B(n3750), .A(n3751), .Z(n3748) );
  XNOR U4312 ( .A(b[1487]), .B(n3749), .Z(n3750) );
  XNOR U4313 ( .A(b[1487]), .B(n3751), .Z(c[1487]) );
  XNOR U4314 ( .A(a[1487]), .B(n3752), .Z(n3751) );
  IV U4315 ( .A(n3749), .Z(n3752) );
  XOR U4316 ( .A(n3753), .B(n3754), .Z(n3749) );
  ANDN U4317 ( .B(n3755), .A(n3756), .Z(n3753) );
  XNOR U4318 ( .A(b[1486]), .B(n3754), .Z(n3755) );
  XNOR U4319 ( .A(b[1486]), .B(n3756), .Z(c[1486]) );
  XNOR U4320 ( .A(a[1486]), .B(n3757), .Z(n3756) );
  IV U4321 ( .A(n3754), .Z(n3757) );
  XOR U4322 ( .A(n3758), .B(n3759), .Z(n3754) );
  ANDN U4323 ( .B(n3760), .A(n3761), .Z(n3758) );
  XNOR U4324 ( .A(b[1485]), .B(n3759), .Z(n3760) );
  XNOR U4325 ( .A(b[1485]), .B(n3761), .Z(c[1485]) );
  XNOR U4326 ( .A(a[1485]), .B(n3762), .Z(n3761) );
  IV U4327 ( .A(n3759), .Z(n3762) );
  XOR U4328 ( .A(n3763), .B(n3764), .Z(n3759) );
  ANDN U4329 ( .B(n3765), .A(n3766), .Z(n3763) );
  XNOR U4330 ( .A(b[1484]), .B(n3764), .Z(n3765) );
  XNOR U4331 ( .A(b[1484]), .B(n3766), .Z(c[1484]) );
  XNOR U4332 ( .A(a[1484]), .B(n3767), .Z(n3766) );
  IV U4333 ( .A(n3764), .Z(n3767) );
  XOR U4334 ( .A(n3768), .B(n3769), .Z(n3764) );
  ANDN U4335 ( .B(n3770), .A(n3771), .Z(n3768) );
  XNOR U4336 ( .A(b[1483]), .B(n3769), .Z(n3770) );
  XNOR U4337 ( .A(b[1483]), .B(n3771), .Z(c[1483]) );
  XNOR U4338 ( .A(a[1483]), .B(n3772), .Z(n3771) );
  IV U4339 ( .A(n3769), .Z(n3772) );
  XOR U4340 ( .A(n3773), .B(n3774), .Z(n3769) );
  ANDN U4341 ( .B(n3775), .A(n3776), .Z(n3773) );
  XNOR U4342 ( .A(b[1482]), .B(n3774), .Z(n3775) );
  XNOR U4343 ( .A(b[1482]), .B(n3776), .Z(c[1482]) );
  XNOR U4344 ( .A(a[1482]), .B(n3777), .Z(n3776) );
  IV U4345 ( .A(n3774), .Z(n3777) );
  XOR U4346 ( .A(n3778), .B(n3779), .Z(n3774) );
  ANDN U4347 ( .B(n3780), .A(n3781), .Z(n3778) );
  XNOR U4348 ( .A(b[1481]), .B(n3779), .Z(n3780) );
  XNOR U4349 ( .A(b[1481]), .B(n3781), .Z(c[1481]) );
  XNOR U4350 ( .A(a[1481]), .B(n3782), .Z(n3781) );
  IV U4351 ( .A(n3779), .Z(n3782) );
  XOR U4352 ( .A(n3783), .B(n3784), .Z(n3779) );
  ANDN U4353 ( .B(n3785), .A(n3786), .Z(n3783) );
  XNOR U4354 ( .A(b[1480]), .B(n3784), .Z(n3785) );
  XNOR U4355 ( .A(b[1480]), .B(n3786), .Z(c[1480]) );
  XNOR U4356 ( .A(a[1480]), .B(n3787), .Z(n3786) );
  IV U4357 ( .A(n3784), .Z(n3787) );
  XOR U4358 ( .A(n3788), .B(n3789), .Z(n3784) );
  ANDN U4359 ( .B(n3790), .A(n3791), .Z(n3788) );
  XNOR U4360 ( .A(b[1479]), .B(n3789), .Z(n3790) );
  XNOR U4361 ( .A(b[147]), .B(n3792), .Z(c[147]) );
  XNOR U4362 ( .A(b[1479]), .B(n3791), .Z(c[1479]) );
  XNOR U4363 ( .A(a[1479]), .B(n3793), .Z(n3791) );
  IV U4364 ( .A(n3789), .Z(n3793) );
  XOR U4365 ( .A(n3794), .B(n3795), .Z(n3789) );
  ANDN U4366 ( .B(n3796), .A(n3797), .Z(n3794) );
  XNOR U4367 ( .A(b[1478]), .B(n3795), .Z(n3796) );
  XNOR U4368 ( .A(b[1478]), .B(n3797), .Z(c[1478]) );
  XNOR U4369 ( .A(a[1478]), .B(n3798), .Z(n3797) );
  IV U4370 ( .A(n3795), .Z(n3798) );
  XOR U4371 ( .A(n3799), .B(n3800), .Z(n3795) );
  ANDN U4372 ( .B(n3801), .A(n3802), .Z(n3799) );
  XNOR U4373 ( .A(b[1477]), .B(n3800), .Z(n3801) );
  XNOR U4374 ( .A(b[1477]), .B(n3802), .Z(c[1477]) );
  XNOR U4375 ( .A(a[1477]), .B(n3803), .Z(n3802) );
  IV U4376 ( .A(n3800), .Z(n3803) );
  XOR U4377 ( .A(n3804), .B(n3805), .Z(n3800) );
  ANDN U4378 ( .B(n3806), .A(n3807), .Z(n3804) );
  XNOR U4379 ( .A(b[1476]), .B(n3805), .Z(n3806) );
  XNOR U4380 ( .A(b[1476]), .B(n3807), .Z(c[1476]) );
  XNOR U4381 ( .A(a[1476]), .B(n3808), .Z(n3807) );
  IV U4382 ( .A(n3805), .Z(n3808) );
  XOR U4383 ( .A(n3809), .B(n3810), .Z(n3805) );
  ANDN U4384 ( .B(n3811), .A(n3812), .Z(n3809) );
  XNOR U4385 ( .A(b[1475]), .B(n3810), .Z(n3811) );
  XNOR U4386 ( .A(b[1475]), .B(n3812), .Z(c[1475]) );
  XNOR U4387 ( .A(a[1475]), .B(n3813), .Z(n3812) );
  IV U4388 ( .A(n3810), .Z(n3813) );
  XOR U4389 ( .A(n3814), .B(n3815), .Z(n3810) );
  ANDN U4390 ( .B(n3816), .A(n3817), .Z(n3814) );
  XNOR U4391 ( .A(b[1474]), .B(n3815), .Z(n3816) );
  XNOR U4392 ( .A(b[1474]), .B(n3817), .Z(c[1474]) );
  XNOR U4393 ( .A(a[1474]), .B(n3818), .Z(n3817) );
  IV U4394 ( .A(n3815), .Z(n3818) );
  XOR U4395 ( .A(n3819), .B(n3820), .Z(n3815) );
  ANDN U4396 ( .B(n3821), .A(n3822), .Z(n3819) );
  XNOR U4397 ( .A(b[1473]), .B(n3820), .Z(n3821) );
  XNOR U4398 ( .A(b[1473]), .B(n3822), .Z(c[1473]) );
  XNOR U4399 ( .A(a[1473]), .B(n3823), .Z(n3822) );
  IV U4400 ( .A(n3820), .Z(n3823) );
  XOR U4401 ( .A(n3824), .B(n3825), .Z(n3820) );
  ANDN U4402 ( .B(n3826), .A(n3827), .Z(n3824) );
  XNOR U4403 ( .A(b[1472]), .B(n3825), .Z(n3826) );
  XNOR U4404 ( .A(b[1472]), .B(n3827), .Z(c[1472]) );
  XNOR U4405 ( .A(a[1472]), .B(n3828), .Z(n3827) );
  IV U4406 ( .A(n3825), .Z(n3828) );
  XOR U4407 ( .A(n3829), .B(n3830), .Z(n3825) );
  ANDN U4408 ( .B(n3831), .A(n3832), .Z(n3829) );
  XNOR U4409 ( .A(b[1471]), .B(n3830), .Z(n3831) );
  XNOR U4410 ( .A(b[1471]), .B(n3832), .Z(c[1471]) );
  XNOR U4411 ( .A(a[1471]), .B(n3833), .Z(n3832) );
  IV U4412 ( .A(n3830), .Z(n3833) );
  XOR U4413 ( .A(n3834), .B(n3835), .Z(n3830) );
  ANDN U4414 ( .B(n3836), .A(n3837), .Z(n3834) );
  XNOR U4415 ( .A(b[1470]), .B(n3835), .Z(n3836) );
  XNOR U4416 ( .A(b[1470]), .B(n3837), .Z(c[1470]) );
  XNOR U4417 ( .A(a[1470]), .B(n3838), .Z(n3837) );
  IV U4418 ( .A(n3835), .Z(n3838) );
  XOR U4419 ( .A(n3839), .B(n3840), .Z(n3835) );
  ANDN U4420 ( .B(n3841), .A(n3842), .Z(n3839) );
  XNOR U4421 ( .A(b[1469]), .B(n3840), .Z(n3841) );
  XNOR U4422 ( .A(b[146]), .B(n3843), .Z(c[146]) );
  XNOR U4423 ( .A(b[1469]), .B(n3842), .Z(c[1469]) );
  XNOR U4424 ( .A(a[1469]), .B(n3844), .Z(n3842) );
  IV U4425 ( .A(n3840), .Z(n3844) );
  XOR U4426 ( .A(n3845), .B(n3846), .Z(n3840) );
  ANDN U4427 ( .B(n3847), .A(n3848), .Z(n3845) );
  XNOR U4428 ( .A(b[1468]), .B(n3846), .Z(n3847) );
  XNOR U4429 ( .A(b[1468]), .B(n3848), .Z(c[1468]) );
  XNOR U4430 ( .A(a[1468]), .B(n3849), .Z(n3848) );
  IV U4431 ( .A(n3846), .Z(n3849) );
  XOR U4432 ( .A(n3850), .B(n3851), .Z(n3846) );
  ANDN U4433 ( .B(n3852), .A(n3853), .Z(n3850) );
  XNOR U4434 ( .A(b[1467]), .B(n3851), .Z(n3852) );
  XNOR U4435 ( .A(b[1467]), .B(n3853), .Z(c[1467]) );
  XNOR U4436 ( .A(a[1467]), .B(n3854), .Z(n3853) );
  IV U4437 ( .A(n3851), .Z(n3854) );
  XOR U4438 ( .A(n3855), .B(n3856), .Z(n3851) );
  ANDN U4439 ( .B(n3857), .A(n3858), .Z(n3855) );
  XNOR U4440 ( .A(b[1466]), .B(n3856), .Z(n3857) );
  XNOR U4441 ( .A(b[1466]), .B(n3858), .Z(c[1466]) );
  XNOR U4442 ( .A(a[1466]), .B(n3859), .Z(n3858) );
  IV U4443 ( .A(n3856), .Z(n3859) );
  XOR U4444 ( .A(n3860), .B(n3861), .Z(n3856) );
  ANDN U4445 ( .B(n3862), .A(n3863), .Z(n3860) );
  XNOR U4446 ( .A(b[1465]), .B(n3861), .Z(n3862) );
  XNOR U4447 ( .A(b[1465]), .B(n3863), .Z(c[1465]) );
  XNOR U4448 ( .A(a[1465]), .B(n3864), .Z(n3863) );
  IV U4449 ( .A(n3861), .Z(n3864) );
  XOR U4450 ( .A(n3865), .B(n3866), .Z(n3861) );
  ANDN U4451 ( .B(n3867), .A(n3868), .Z(n3865) );
  XNOR U4452 ( .A(b[1464]), .B(n3866), .Z(n3867) );
  XNOR U4453 ( .A(b[1464]), .B(n3868), .Z(c[1464]) );
  XNOR U4454 ( .A(a[1464]), .B(n3869), .Z(n3868) );
  IV U4455 ( .A(n3866), .Z(n3869) );
  XOR U4456 ( .A(n3870), .B(n3871), .Z(n3866) );
  ANDN U4457 ( .B(n3872), .A(n3873), .Z(n3870) );
  XNOR U4458 ( .A(b[1463]), .B(n3871), .Z(n3872) );
  XNOR U4459 ( .A(b[1463]), .B(n3873), .Z(c[1463]) );
  XNOR U4460 ( .A(a[1463]), .B(n3874), .Z(n3873) );
  IV U4461 ( .A(n3871), .Z(n3874) );
  XOR U4462 ( .A(n3875), .B(n3876), .Z(n3871) );
  ANDN U4463 ( .B(n3877), .A(n3878), .Z(n3875) );
  XNOR U4464 ( .A(b[1462]), .B(n3876), .Z(n3877) );
  XNOR U4465 ( .A(b[1462]), .B(n3878), .Z(c[1462]) );
  XNOR U4466 ( .A(a[1462]), .B(n3879), .Z(n3878) );
  IV U4467 ( .A(n3876), .Z(n3879) );
  XOR U4468 ( .A(n3880), .B(n3881), .Z(n3876) );
  ANDN U4469 ( .B(n3882), .A(n3883), .Z(n3880) );
  XNOR U4470 ( .A(b[1461]), .B(n3881), .Z(n3882) );
  XNOR U4471 ( .A(b[1461]), .B(n3883), .Z(c[1461]) );
  XNOR U4472 ( .A(a[1461]), .B(n3884), .Z(n3883) );
  IV U4473 ( .A(n3881), .Z(n3884) );
  XOR U4474 ( .A(n3885), .B(n3886), .Z(n3881) );
  ANDN U4475 ( .B(n3887), .A(n3888), .Z(n3885) );
  XNOR U4476 ( .A(b[1460]), .B(n3886), .Z(n3887) );
  XNOR U4477 ( .A(b[1460]), .B(n3888), .Z(c[1460]) );
  XNOR U4478 ( .A(a[1460]), .B(n3889), .Z(n3888) );
  IV U4479 ( .A(n3886), .Z(n3889) );
  XOR U4480 ( .A(n3890), .B(n3891), .Z(n3886) );
  ANDN U4481 ( .B(n3892), .A(n3893), .Z(n3890) );
  XNOR U4482 ( .A(b[1459]), .B(n3891), .Z(n3892) );
  XNOR U4483 ( .A(b[145]), .B(n3894), .Z(c[145]) );
  XNOR U4484 ( .A(b[1459]), .B(n3893), .Z(c[1459]) );
  XNOR U4485 ( .A(a[1459]), .B(n3895), .Z(n3893) );
  IV U4486 ( .A(n3891), .Z(n3895) );
  XOR U4487 ( .A(n3896), .B(n3897), .Z(n3891) );
  ANDN U4488 ( .B(n3898), .A(n3899), .Z(n3896) );
  XNOR U4489 ( .A(b[1458]), .B(n3897), .Z(n3898) );
  XNOR U4490 ( .A(b[1458]), .B(n3899), .Z(c[1458]) );
  XNOR U4491 ( .A(a[1458]), .B(n3900), .Z(n3899) );
  IV U4492 ( .A(n3897), .Z(n3900) );
  XOR U4493 ( .A(n3901), .B(n3902), .Z(n3897) );
  ANDN U4494 ( .B(n3903), .A(n3904), .Z(n3901) );
  XNOR U4495 ( .A(b[1457]), .B(n3902), .Z(n3903) );
  XNOR U4496 ( .A(b[1457]), .B(n3904), .Z(c[1457]) );
  XNOR U4497 ( .A(a[1457]), .B(n3905), .Z(n3904) );
  IV U4498 ( .A(n3902), .Z(n3905) );
  XOR U4499 ( .A(n3906), .B(n3907), .Z(n3902) );
  ANDN U4500 ( .B(n3908), .A(n3909), .Z(n3906) );
  XNOR U4501 ( .A(b[1456]), .B(n3907), .Z(n3908) );
  XNOR U4502 ( .A(b[1456]), .B(n3909), .Z(c[1456]) );
  XNOR U4503 ( .A(a[1456]), .B(n3910), .Z(n3909) );
  IV U4504 ( .A(n3907), .Z(n3910) );
  XOR U4505 ( .A(n3911), .B(n3912), .Z(n3907) );
  ANDN U4506 ( .B(n3913), .A(n3914), .Z(n3911) );
  XNOR U4507 ( .A(b[1455]), .B(n3912), .Z(n3913) );
  XNOR U4508 ( .A(b[1455]), .B(n3914), .Z(c[1455]) );
  XNOR U4509 ( .A(a[1455]), .B(n3915), .Z(n3914) );
  IV U4510 ( .A(n3912), .Z(n3915) );
  XOR U4511 ( .A(n3916), .B(n3917), .Z(n3912) );
  ANDN U4512 ( .B(n3918), .A(n3919), .Z(n3916) );
  XNOR U4513 ( .A(b[1454]), .B(n3917), .Z(n3918) );
  XNOR U4514 ( .A(b[1454]), .B(n3919), .Z(c[1454]) );
  XNOR U4515 ( .A(a[1454]), .B(n3920), .Z(n3919) );
  IV U4516 ( .A(n3917), .Z(n3920) );
  XOR U4517 ( .A(n3921), .B(n3922), .Z(n3917) );
  ANDN U4518 ( .B(n3923), .A(n3924), .Z(n3921) );
  XNOR U4519 ( .A(b[1453]), .B(n3922), .Z(n3923) );
  XNOR U4520 ( .A(b[1453]), .B(n3924), .Z(c[1453]) );
  XNOR U4521 ( .A(a[1453]), .B(n3925), .Z(n3924) );
  IV U4522 ( .A(n3922), .Z(n3925) );
  XOR U4523 ( .A(n3926), .B(n3927), .Z(n3922) );
  ANDN U4524 ( .B(n3928), .A(n3929), .Z(n3926) );
  XNOR U4525 ( .A(b[1452]), .B(n3927), .Z(n3928) );
  XNOR U4526 ( .A(b[1452]), .B(n3929), .Z(c[1452]) );
  XNOR U4527 ( .A(a[1452]), .B(n3930), .Z(n3929) );
  IV U4528 ( .A(n3927), .Z(n3930) );
  XOR U4529 ( .A(n3931), .B(n3932), .Z(n3927) );
  ANDN U4530 ( .B(n3933), .A(n3934), .Z(n3931) );
  XNOR U4531 ( .A(b[1451]), .B(n3932), .Z(n3933) );
  XNOR U4532 ( .A(b[1451]), .B(n3934), .Z(c[1451]) );
  XNOR U4533 ( .A(a[1451]), .B(n3935), .Z(n3934) );
  IV U4534 ( .A(n3932), .Z(n3935) );
  XOR U4535 ( .A(n3936), .B(n3937), .Z(n3932) );
  ANDN U4536 ( .B(n3938), .A(n3939), .Z(n3936) );
  XNOR U4537 ( .A(b[1450]), .B(n3937), .Z(n3938) );
  XNOR U4538 ( .A(b[1450]), .B(n3939), .Z(c[1450]) );
  XNOR U4539 ( .A(a[1450]), .B(n3940), .Z(n3939) );
  IV U4540 ( .A(n3937), .Z(n3940) );
  XOR U4541 ( .A(n3941), .B(n3942), .Z(n3937) );
  ANDN U4542 ( .B(n3943), .A(n3944), .Z(n3941) );
  XNOR U4543 ( .A(b[1449]), .B(n3942), .Z(n3943) );
  XNOR U4544 ( .A(b[144]), .B(n3945), .Z(c[144]) );
  XNOR U4545 ( .A(b[1449]), .B(n3944), .Z(c[1449]) );
  XNOR U4546 ( .A(a[1449]), .B(n3946), .Z(n3944) );
  IV U4547 ( .A(n3942), .Z(n3946) );
  XOR U4548 ( .A(n3947), .B(n3948), .Z(n3942) );
  ANDN U4549 ( .B(n3949), .A(n3950), .Z(n3947) );
  XNOR U4550 ( .A(b[1448]), .B(n3948), .Z(n3949) );
  XNOR U4551 ( .A(b[1448]), .B(n3950), .Z(c[1448]) );
  XNOR U4552 ( .A(a[1448]), .B(n3951), .Z(n3950) );
  IV U4553 ( .A(n3948), .Z(n3951) );
  XOR U4554 ( .A(n3952), .B(n3953), .Z(n3948) );
  ANDN U4555 ( .B(n3954), .A(n3955), .Z(n3952) );
  XNOR U4556 ( .A(b[1447]), .B(n3953), .Z(n3954) );
  XNOR U4557 ( .A(b[1447]), .B(n3955), .Z(c[1447]) );
  XNOR U4558 ( .A(a[1447]), .B(n3956), .Z(n3955) );
  IV U4559 ( .A(n3953), .Z(n3956) );
  XOR U4560 ( .A(n3957), .B(n3958), .Z(n3953) );
  ANDN U4561 ( .B(n3959), .A(n3960), .Z(n3957) );
  XNOR U4562 ( .A(b[1446]), .B(n3958), .Z(n3959) );
  XNOR U4563 ( .A(b[1446]), .B(n3960), .Z(c[1446]) );
  XNOR U4564 ( .A(a[1446]), .B(n3961), .Z(n3960) );
  IV U4565 ( .A(n3958), .Z(n3961) );
  XOR U4566 ( .A(n3962), .B(n3963), .Z(n3958) );
  ANDN U4567 ( .B(n3964), .A(n3965), .Z(n3962) );
  XNOR U4568 ( .A(b[1445]), .B(n3963), .Z(n3964) );
  XNOR U4569 ( .A(b[1445]), .B(n3965), .Z(c[1445]) );
  XNOR U4570 ( .A(a[1445]), .B(n3966), .Z(n3965) );
  IV U4571 ( .A(n3963), .Z(n3966) );
  XOR U4572 ( .A(n3967), .B(n3968), .Z(n3963) );
  ANDN U4573 ( .B(n3969), .A(n3970), .Z(n3967) );
  XNOR U4574 ( .A(b[1444]), .B(n3968), .Z(n3969) );
  XNOR U4575 ( .A(b[1444]), .B(n3970), .Z(c[1444]) );
  XNOR U4576 ( .A(a[1444]), .B(n3971), .Z(n3970) );
  IV U4577 ( .A(n3968), .Z(n3971) );
  XOR U4578 ( .A(n3972), .B(n3973), .Z(n3968) );
  ANDN U4579 ( .B(n3974), .A(n3975), .Z(n3972) );
  XNOR U4580 ( .A(b[1443]), .B(n3973), .Z(n3974) );
  XNOR U4581 ( .A(b[1443]), .B(n3975), .Z(c[1443]) );
  XNOR U4582 ( .A(a[1443]), .B(n3976), .Z(n3975) );
  IV U4583 ( .A(n3973), .Z(n3976) );
  XOR U4584 ( .A(n3977), .B(n3978), .Z(n3973) );
  ANDN U4585 ( .B(n3979), .A(n3980), .Z(n3977) );
  XNOR U4586 ( .A(b[1442]), .B(n3978), .Z(n3979) );
  XNOR U4587 ( .A(b[1442]), .B(n3980), .Z(c[1442]) );
  XNOR U4588 ( .A(a[1442]), .B(n3981), .Z(n3980) );
  IV U4589 ( .A(n3978), .Z(n3981) );
  XOR U4590 ( .A(n3982), .B(n3983), .Z(n3978) );
  ANDN U4591 ( .B(n3984), .A(n3985), .Z(n3982) );
  XNOR U4592 ( .A(b[1441]), .B(n3983), .Z(n3984) );
  XNOR U4593 ( .A(b[1441]), .B(n3985), .Z(c[1441]) );
  XNOR U4594 ( .A(a[1441]), .B(n3986), .Z(n3985) );
  IV U4595 ( .A(n3983), .Z(n3986) );
  XOR U4596 ( .A(n3987), .B(n3988), .Z(n3983) );
  ANDN U4597 ( .B(n3989), .A(n3990), .Z(n3987) );
  XNOR U4598 ( .A(b[1440]), .B(n3988), .Z(n3989) );
  XNOR U4599 ( .A(b[1440]), .B(n3990), .Z(c[1440]) );
  XNOR U4600 ( .A(a[1440]), .B(n3991), .Z(n3990) );
  IV U4601 ( .A(n3988), .Z(n3991) );
  XOR U4602 ( .A(n3992), .B(n3993), .Z(n3988) );
  ANDN U4603 ( .B(n3994), .A(n3995), .Z(n3992) );
  XNOR U4604 ( .A(b[1439]), .B(n3993), .Z(n3994) );
  XNOR U4605 ( .A(b[143]), .B(n3996), .Z(c[143]) );
  XNOR U4606 ( .A(b[1439]), .B(n3995), .Z(c[1439]) );
  XNOR U4607 ( .A(a[1439]), .B(n3997), .Z(n3995) );
  IV U4608 ( .A(n3993), .Z(n3997) );
  XOR U4609 ( .A(n3998), .B(n3999), .Z(n3993) );
  ANDN U4610 ( .B(n4000), .A(n4001), .Z(n3998) );
  XNOR U4611 ( .A(b[1438]), .B(n3999), .Z(n4000) );
  XNOR U4612 ( .A(b[1438]), .B(n4001), .Z(c[1438]) );
  XNOR U4613 ( .A(a[1438]), .B(n4002), .Z(n4001) );
  IV U4614 ( .A(n3999), .Z(n4002) );
  XOR U4615 ( .A(n4003), .B(n4004), .Z(n3999) );
  ANDN U4616 ( .B(n4005), .A(n4006), .Z(n4003) );
  XNOR U4617 ( .A(b[1437]), .B(n4004), .Z(n4005) );
  XNOR U4618 ( .A(b[1437]), .B(n4006), .Z(c[1437]) );
  XNOR U4619 ( .A(a[1437]), .B(n4007), .Z(n4006) );
  IV U4620 ( .A(n4004), .Z(n4007) );
  XOR U4621 ( .A(n4008), .B(n4009), .Z(n4004) );
  ANDN U4622 ( .B(n4010), .A(n4011), .Z(n4008) );
  XNOR U4623 ( .A(b[1436]), .B(n4009), .Z(n4010) );
  XNOR U4624 ( .A(b[1436]), .B(n4011), .Z(c[1436]) );
  XNOR U4625 ( .A(a[1436]), .B(n4012), .Z(n4011) );
  IV U4626 ( .A(n4009), .Z(n4012) );
  XOR U4627 ( .A(n4013), .B(n4014), .Z(n4009) );
  ANDN U4628 ( .B(n4015), .A(n4016), .Z(n4013) );
  XNOR U4629 ( .A(b[1435]), .B(n4014), .Z(n4015) );
  XNOR U4630 ( .A(b[1435]), .B(n4016), .Z(c[1435]) );
  XNOR U4631 ( .A(a[1435]), .B(n4017), .Z(n4016) );
  IV U4632 ( .A(n4014), .Z(n4017) );
  XOR U4633 ( .A(n4018), .B(n4019), .Z(n4014) );
  ANDN U4634 ( .B(n4020), .A(n4021), .Z(n4018) );
  XNOR U4635 ( .A(b[1434]), .B(n4019), .Z(n4020) );
  XNOR U4636 ( .A(b[1434]), .B(n4021), .Z(c[1434]) );
  XNOR U4637 ( .A(a[1434]), .B(n4022), .Z(n4021) );
  IV U4638 ( .A(n4019), .Z(n4022) );
  XOR U4639 ( .A(n4023), .B(n4024), .Z(n4019) );
  ANDN U4640 ( .B(n4025), .A(n4026), .Z(n4023) );
  XNOR U4641 ( .A(b[1433]), .B(n4024), .Z(n4025) );
  XNOR U4642 ( .A(b[1433]), .B(n4026), .Z(c[1433]) );
  XNOR U4643 ( .A(a[1433]), .B(n4027), .Z(n4026) );
  IV U4644 ( .A(n4024), .Z(n4027) );
  XOR U4645 ( .A(n4028), .B(n4029), .Z(n4024) );
  ANDN U4646 ( .B(n4030), .A(n4031), .Z(n4028) );
  XNOR U4647 ( .A(b[1432]), .B(n4029), .Z(n4030) );
  XNOR U4648 ( .A(b[1432]), .B(n4031), .Z(c[1432]) );
  XNOR U4649 ( .A(a[1432]), .B(n4032), .Z(n4031) );
  IV U4650 ( .A(n4029), .Z(n4032) );
  XOR U4651 ( .A(n4033), .B(n4034), .Z(n4029) );
  ANDN U4652 ( .B(n4035), .A(n4036), .Z(n4033) );
  XNOR U4653 ( .A(b[1431]), .B(n4034), .Z(n4035) );
  XNOR U4654 ( .A(b[1431]), .B(n4036), .Z(c[1431]) );
  XNOR U4655 ( .A(a[1431]), .B(n4037), .Z(n4036) );
  IV U4656 ( .A(n4034), .Z(n4037) );
  XOR U4657 ( .A(n4038), .B(n4039), .Z(n4034) );
  ANDN U4658 ( .B(n4040), .A(n4041), .Z(n4038) );
  XNOR U4659 ( .A(b[1430]), .B(n4039), .Z(n4040) );
  XNOR U4660 ( .A(b[1430]), .B(n4041), .Z(c[1430]) );
  XNOR U4661 ( .A(a[1430]), .B(n4042), .Z(n4041) );
  IV U4662 ( .A(n4039), .Z(n4042) );
  XOR U4663 ( .A(n4043), .B(n4044), .Z(n4039) );
  ANDN U4664 ( .B(n4045), .A(n4046), .Z(n4043) );
  XNOR U4665 ( .A(b[1429]), .B(n4044), .Z(n4045) );
  XNOR U4666 ( .A(b[142]), .B(n4047), .Z(c[142]) );
  XNOR U4667 ( .A(b[1429]), .B(n4046), .Z(c[1429]) );
  XNOR U4668 ( .A(a[1429]), .B(n4048), .Z(n4046) );
  IV U4669 ( .A(n4044), .Z(n4048) );
  XOR U4670 ( .A(n4049), .B(n4050), .Z(n4044) );
  ANDN U4671 ( .B(n4051), .A(n4052), .Z(n4049) );
  XNOR U4672 ( .A(b[1428]), .B(n4050), .Z(n4051) );
  XNOR U4673 ( .A(b[1428]), .B(n4052), .Z(c[1428]) );
  XNOR U4674 ( .A(a[1428]), .B(n4053), .Z(n4052) );
  IV U4675 ( .A(n4050), .Z(n4053) );
  XOR U4676 ( .A(n4054), .B(n4055), .Z(n4050) );
  ANDN U4677 ( .B(n4056), .A(n4057), .Z(n4054) );
  XNOR U4678 ( .A(b[1427]), .B(n4055), .Z(n4056) );
  XNOR U4679 ( .A(b[1427]), .B(n4057), .Z(c[1427]) );
  XNOR U4680 ( .A(a[1427]), .B(n4058), .Z(n4057) );
  IV U4681 ( .A(n4055), .Z(n4058) );
  XOR U4682 ( .A(n4059), .B(n4060), .Z(n4055) );
  ANDN U4683 ( .B(n4061), .A(n4062), .Z(n4059) );
  XNOR U4684 ( .A(b[1426]), .B(n4060), .Z(n4061) );
  XNOR U4685 ( .A(b[1426]), .B(n4062), .Z(c[1426]) );
  XNOR U4686 ( .A(a[1426]), .B(n4063), .Z(n4062) );
  IV U4687 ( .A(n4060), .Z(n4063) );
  XOR U4688 ( .A(n4064), .B(n4065), .Z(n4060) );
  ANDN U4689 ( .B(n4066), .A(n4067), .Z(n4064) );
  XNOR U4690 ( .A(b[1425]), .B(n4065), .Z(n4066) );
  XNOR U4691 ( .A(b[1425]), .B(n4067), .Z(c[1425]) );
  XNOR U4692 ( .A(a[1425]), .B(n4068), .Z(n4067) );
  IV U4693 ( .A(n4065), .Z(n4068) );
  XOR U4694 ( .A(n4069), .B(n4070), .Z(n4065) );
  ANDN U4695 ( .B(n4071), .A(n4072), .Z(n4069) );
  XNOR U4696 ( .A(b[1424]), .B(n4070), .Z(n4071) );
  XNOR U4697 ( .A(b[1424]), .B(n4072), .Z(c[1424]) );
  XNOR U4698 ( .A(a[1424]), .B(n4073), .Z(n4072) );
  IV U4699 ( .A(n4070), .Z(n4073) );
  XOR U4700 ( .A(n4074), .B(n4075), .Z(n4070) );
  ANDN U4701 ( .B(n4076), .A(n4077), .Z(n4074) );
  XNOR U4702 ( .A(b[1423]), .B(n4075), .Z(n4076) );
  XNOR U4703 ( .A(b[1423]), .B(n4077), .Z(c[1423]) );
  XNOR U4704 ( .A(a[1423]), .B(n4078), .Z(n4077) );
  IV U4705 ( .A(n4075), .Z(n4078) );
  XOR U4706 ( .A(n4079), .B(n4080), .Z(n4075) );
  ANDN U4707 ( .B(n4081), .A(n4082), .Z(n4079) );
  XNOR U4708 ( .A(b[1422]), .B(n4080), .Z(n4081) );
  XNOR U4709 ( .A(b[1422]), .B(n4082), .Z(c[1422]) );
  XNOR U4710 ( .A(a[1422]), .B(n4083), .Z(n4082) );
  IV U4711 ( .A(n4080), .Z(n4083) );
  XOR U4712 ( .A(n4084), .B(n4085), .Z(n4080) );
  ANDN U4713 ( .B(n4086), .A(n4087), .Z(n4084) );
  XNOR U4714 ( .A(b[1421]), .B(n4085), .Z(n4086) );
  XNOR U4715 ( .A(b[1421]), .B(n4087), .Z(c[1421]) );
  XNOR U4716 ( .A(a[1421]), .B(n4088), .Z(n4087) );
  IV U4717 ( .A(n4085), .Z(n4088) );
  XOR U4718 ( .A(n4089), .B(n4090), .Z(n4085) );
  ANDN U4719 ( .B(n4091), .A(n4092), .Z(n4089) );
  XNOR U4720 ( .A(b[1420]), .B(n4090), .Z(n4091) );
  XNOR U4721 ( .A(b[1420]), .B(n4092), .Z(c[1420]) );
  XNOR U4722 ( .A(a[1420]), .B(n4093), .Z(n4092) );
  IV U4723 ( .A(n4090), .Z(n4093) );
  XOR U4724 ( .A(n4094), .B(n4095), .Z(n4090) );
  ANDN U4725 ( .B(n4096), .A(n4097), .Z(n4094) );
  XNOR U4726 ( .A(b[1419]), .B(n4095), .Z(n4096) );
  XNOR U4727 ( .A(b[141]), .B(n4098), .Z(c[141]) );
  XNOR U4728 ( .A(b[1419]), .B(n4097), .Z(c[1419]) );
  XNOR U4729 ( .A(a[1419]), .B(n4099), .Z(n4097) );
  IV U4730 ( .A(n4095), .Z(n4099) );
  XOR U4731 ( .A(n4100), .B(n4101), .Z(n4095) );
  ANDN U4732 ( .B(n4102), .A(n4103), .Z(n4100) );
  XNOR U4733 ( .A(b[1418]), .B(n4101), .Z(n4102) );
  XNOR U4734 ( .A(b[1418]), .B(n4103), .Z(c[1418]) );
  XNOR U4735 ( .A(a[1418]), .B(n4104), .Z(n4103) );
  IV U4736 ( .A(n4101), .Z(n4104) );
  XOR U4737 ( .A(n4105), .B(n4106), .Z(n4101) );
  ANDN U4738 ( .B(n4107), .A(n4108), .Z(n4105) );
  XNOR U4739 ( .A(b[1417]), .B(n4106), .Z(n4107) );
  XNOR U4740 ( .A(b[1417]), .B(n4108), .Z(c[1417]) );
  XNOR U4741 ( .A(a[1417]), .B(n4109), .Z(n4108) );
  IV U4742 ( .A(n4106), .Z(n4109) );
  XOR U4743 ( .A(n4110), .B(n4111), .Z(n4106) );
  ANDN U4744 ( .B(n4112), .A(n4113), .Z(n4110) );
  XNOR U4745 ( .A(b[1416]), .B(n4111), .Z(n4112) );
  XNOR U4746 ( .A(b[1416]), .B(n4113), .Z(c[1416]) );
  XNOR U4747 ( .A(a[1416]), .B(n4114), .Z(n4113) );
  IV U4748 ( .A(n4111), .Z(n4114) );
  XOR U4749 ( .A(n4115), .B(n4116), .Z(n4111) );
  ANDN U4750 ( .B(n4117), .A(n4118), .Z(n4115) );
  XNOR U4751 ( .A(b[1415]), .B(n4116), .Z(n4117) );
  XNOR U4752 ( .A(b[1415]), .B(n4118), .Z(c[1415]) );
  XNOR U4753 ( .A(a[1415]), .B(n4119), .Z(n4118) );
  IV U4754 ( .A(n4116), .Z(n4119) );
  XOR U4755 ( .A(n4120), .B(n4121), .Z(n4116) );
  ANDN U4756 ( .B(n4122), .A(n4123), .Z(n4120) );
  XNOR U4757 ( .A(b[1414]), .B(n4121), .Z(n4122) );
  XNOR U4758 ( .A(b[1414]), .B(n4123), .Z(c[1414]) );
  XNOR U4759 ( .A(a[1414]), .B(n4124), .Z(n4123) );
  IV U4760 ( .A(n4121), .Z(n4124) );
  XOR U4761 ( .A(n4125), .B(n4126), .Z(n4121) );
  ANDN U4762 ( .B(n4127), .A(n4128), .Z(n4125) );
  XNOR U4763 ( .A(b[1413]), .B(n4126), .Z(n4127) );
  XNOR U4764 ( .A(b[1413]), .B(n4128), .Z(c[1413]) );
  XNOR U4765 ( .A(a[1413]), .B(n4129), .Z(n4128) );
  IV U4766 ( .A(n4126), .Z(n4129) );
  XOR U4767 ( .A(n4130), .B(n4131), .Z(n4126) );
  ANDN U4768 ( .B(n4132), .A(n4133), .Z(n4130) );
  XNOR U4769 ( .A(b[1412]), .B(n4131), .Z(n4132) );
  XNOR U4770 ( .A(b[1412]), .B(n4133), .Z(c[1412]) );
  XNOR U4771 ( .A(a[1412]), .B(n4134), .Z(n4133) );
  IV U4772 ( .A(n4131), .Z(n4134) );
  XOR U4773 ( .A(n4135), .B(n4136), .Z(n4131) );
  ANDN U4774 ( .B(n4137), .A(n4138), .Z(n4135) );
  XNOR U4775 ( .A(b[1411]), .B(n4136), .Z(n4137) );
  XNOR U4776 ( .A(b[1411]), .B(n4138), .Z(c[1411]) );
  XNOR U4777 ( .A(a[1411]), .B(n4139), .Z(n4138) );
  IV U4778 ( .A(n4136), .Z(n4139) );
  XOR U4779 ( .A(n4140), .B(n4141), .Z(n4136) );
  ANDN U4780 ( .B(n4142), .A(n4143), .Z(n4140) );
  XNOR U4781 ( .A(b[1410]), .B(n4141), .Z(n4142) );
  XNOR U4782 ( .A(b[1410]), .B(n4143), .Z(c[1410]) );
  XNOR U4783 ( .A(a[1410]), .B(n4144), .Z(n4143) );
  IV U4784 ( .A(n4141), .Z(n4144) );
  XOR U4785 ( .A(n4145), .B(n4146), .Z(n4141) );
  ANDN U4786 ( .B(n4147), .A(n4148), .Z(n4145) );
  XNOR U4787 ( .A(b[1409]), .B(n4146), .Z(n4147) );
  XNOR U4788 ( .A(b[140]), .B(n4149), .Z(c[140]) );
  XNOR U4789 ( .A(b[1409]), .B(n4148), .Z(c[1409]) );
  XNOR U4790 ( .A(a[1409]), .B(n4150), .Z(n4148) );
  IV U4791 ( .A(n4146), .Z(n4150) );
  XOR U4792 ( .A(n4151), .B(n4152), .Z(n4146) );
  ANDN U4793 ( .B(n4153), .A(n4154), .Z(n4151) );
  XNOR U4794 ( .A(b[1408]), .B(n4152), .Z(n4153) );
  XNOR U4795 ( .A(b[1408]), .B(n4154), .Z(c[1408]) );
  XNOR U4796 ( .A(a[1408]), .B(n4155), .Z(n4154) );
  IV U4797 ( .A(n4152), .Z(n4155) );
  XOR U4798 ( .A(n4156), .B(n4157), .Z(n4152) );
  ANDN U4799 ( .B(n4158), .A(n4159), .Z(n4156) );
  XNOR U4800 ( .A(b[1407]), .B(n4157), .Z(n4158) );
  XNOR U4801 ( .A(b[1407]), .B(n4159), .Z(c[1407]) );
  XNOR U4802 ( .A(a[1407]), .B(n4160), .Z(n4159) );
  IV U4803 ( .A(n4157), .Z(n4160) );
  XOR U4804 ( .A(n4161), .B(n4162), .Z(n4157) );
  ANDN U4805 ( .B(n4163), .A(n4164), .Z(n4161) );
  XNOR U4806 ( .A(b[1406]), .B(n4162), .Z(n4163) );
  XNOR U4807 ( .A(b[1406]), .B(n4164), .Z(c[1406]) );
  XNOR U4808 ( .A(a[1406]), .B(n4165), .Z(n4164) );
  IV U4809 ( .A(n4162), .Z(n4165) );
  XOR U4810 ( .A(n4166), .B(n4167), .Z(n4162) );
  ANDN U4811 ( .B(n4168), .A(n4169), .Z(n4166) );
  XNOR U4812 ( .A(b[1405]), .B(n4167), .Z(n4168) );
  XNOR U4813 ( .A(b[1405]), .B(n4169), .Z(c[1405]) );
  XNOR U4814 ( .A(a[1405]), .B(n4170), .Z(n4169) );
  IV U4815 ( .A(n4167), .Z(n4170) );
  XOR U4816 ( .A(n4171), .B(n4172), .Z(n4167) );
  ANDN U4817 ( .B(n4173), .A(n4174), .Z(n4171) );
  XNOR U4818 ( .A(b[1404]), .B(n4172), .Z(n4173) );
  XNOR U4819 ( .A(b[1404]), .B(n4174), .Z(c[1404]) );
  XNOR U4820 ( .A(a[1404]), .B(n4175), .Z(n4174) );
  IV U4821 ( .A(n4172), .Z(n4175) );
  XOR U4822 ( .A(n4176), .B(n4177), .Z(n4172) );
  ANDN U4823 ( .B(n4178), .A(n4179), .Z(n4176) );
  XNOR U4824 ( .A(b[1403]), .B(n4177), .Z(n4178) );
  XNOR U4825 ( .A(b[1403]), .B(n4179), .Z(c[1403]) );
  XNOR U4826 ( .A(a[1403]), .B(n4180), .Z(n4179) );
  IV U4827 ( .A(n4177), .Z(n4180) );
  XOR U4828 ( .A(n4181), .B(n4182), .Z(n4177) );
  ANDN U4829 ( .B(n4183), .A(n4184), .Z(n4181) );
  XNOR U4830 ( .A(b[1402]), .B(n4182), .Z(n4183) );
  XNOR U4831 ( .A(b[1402]), .B(n4184), .Z(c[1402]) );
  XNOR U4832 ( .A(a[1402]), .B(n4185), .Z(n4184) );
  IV U4833 ( .A(n4182), .Z(n4185) );
  XOR U4834 ( .A(n4186), .B(n4187), .Z(n4182) );
  ANDN U4835 ( .B(n4188), .A(n4189), .Z(n4186) );
  XNOR U4836 ( .A(b[1401]), .B(n4187), .Z(n4188) );
  XNOR U4837 ( .A(b[1401]), .B(n4189), .Z(c[1401]) );
  XNOR U4838 ( .A(a[1401]), .B(n4190), .Z(n4189) );
  IV U4839 ( .A(n4187), .Z(n4190) );
  XOR U4840 ( .A(n4191), .B(n4192), .Z(n4187) );
  ANDN U4841 ( .B(n4193), .A(n4194), .Z(n4191) );
  XNOR U4842 ( .A(b[1400]), .B(n4192), .Z(n4193) );
  XNOR U4843 ( .A(b[1400]), .B(n4194), .Z(c[1400]) );
  XNOR U4844 ( .A(a[1400]), .B(n4195), .Z(n4194) );
  IV U4845 ( .A(n4192), .Z(n4195) );
  XOR U4846 ( .A(n4196), .B(n4197), .Z(n4192) );
  ANDN U4847 ( .B(n4198), .A(n4199), .Z(n4196) );
  XNOR U4848 ( .A(b[1399]), .B(n4197), .Z(n4198) );
  XNOR U4849 ( .A(b[13]), .B(n4200), .Z(c[13]) );
  XNOR U4850 ( .A(b[139]), .B(n4201), .Z(c[139]) );
  XNOR U4851 ( .A(b[1399]), .B(n4199), .Z(c[1399]) );
  XNOR U4852 ( .A(a[1399]), .B(n4202), .Z(n4199) );
  IV U4853 ( .A(n4197), .Z(n4202) );
  XOR U4854 ( .A(n4203), .B(n4204), .Z(n4197) );
  ANDN U4855 ( .B(n4205), .A(n4206), .Z(n4203) );
  XNOR U4856 ( .A(b[1398]), .B(n4204), .Z(n4205) );
  XNOR U4857 ( .A(b[1398]), .B(n4206), .Z(c[1398]) );
  XNOR U4858 ( .A(a[1398]), .B(n4207), .Z(n4206) );
  IV U4859 ( .A(n4204), .Z(n4207) );
  XOR U4860 ( .A(n4208), .B(n4209), .Z(n4204) );
  ANDN U4861 ( .B(n4210), .A(n4211), .Z(n4208) );
  XNOR U4862 ( .A(b[1397]), .B(n4209), .Z(n4210) );
  XNOR U4863 ( .A(b[1397]), .B(n4211), .Z(c[1397]) );
  XNOR U4864 ( .A(a[1397]), .B(n4212), .Z(n4211) );
  IV U4865 ( .A(n4209), .Z(n4212) );
  XOR U4866 ( .A(n4213), .B(n4214), .Z(n4209) );
  ANDN U4867 ( .B(n4215), .A(n4216), .Z(n4213) );
  XNOR U4868 ( .A(b[1396]), .B(n4214), .Z(n4215) );
  XNOR U4869 ( .A(b[1396]), .B(n4216), .Z(c[1396]) );
  XNOR U4870 ( .A(a[1396]), .B(n4217), .Z(n4216) );
  IV U4871 ( .A(n4214), .Z(n4217) );
  XOR U4872 ( .A(n4218), .B(n4219), .Z(n4214) );
  ANDN U4873 ( .B(n4220), .A(n4221), .Z(n4218) );
  XNOR U4874 ( .A(b[1395]), .B(n4219), .Z(n4220) );
  XNOR U4875 ( .A(b[1395]), .B(n4221), .Z(c[1395]) );
  XNOR U4876 ( .A(a[1395]), .B(n4222), .Z(n4221) );
  IV U4877 ( .A(n4219), .Z(n4222) );
  XOR U4878 ( .A(n4223), .B(n4224), .Z(n4219) );
  ANDN U4879 ( .B(n4225), .A(n4226), .Z(n4223) );
  XNOR U4880 ( .A(b[1394]), .B(n4224), .Z(n4225) );
  XNOR U4881 ( .A(b[1394]), .B(n4226), .Z(c[1394]) );
  XNOR U4882 ( .A(a[1394]), .B(n4227), .Z(n4226) );
  IV U4883 ( .A(n4224), .Z(n4227) );
  XOR U4884 ( .A(n4228), .B(n4229), .Z(n4224) );
  ANDN U4885 ( .B(n4230), .A(n4231), .Z(n4228) );
  XNOR U4886 ( .A(b[1393]), .B(n4229), .Z(n4230) );
  XNOR U4887 ( .A(b[1393]), .B(n4231), .Z(c[1393]) );
  XNOR U4888 ( .A(a[1393]), .B(n4232), .Z(n4231) );
  IV U4889 ( .A(n4229), .Z(n4232) );
  XOR U4890 ( .A(n4233), .B(n4234), .Z(n4229) );
  ANDN U4891 ( .B(n4235), .A(n4236), .Z(n4233) );
  XNOR U4892 ( .A(b[1392]), .B(n4234), .Z(n4235) );
  XNOR U4893 ( .A(b[1392]), .B(n4236), .Z(c[1392]) );
  XNOR U4894 ( .A(a[1392]), .B(n4237), .Z(n4236) );
  IV U4895 ( .A(n4234), .Z(n4237) );
  XOR U4896 ( .A(n4238), .B(n4239), .Z(n4234) );
  ANDN U4897 ( .B(n4240), .A(n4241), .Z(n4238) );
  XNOR U4898 ( .A(b[1391]), .B(n4239), .Z(n4240) );
  XNOR U4899 ( .A(b[1391]), .B(n4241), .Z(c[1391]) );
  XNOR U4900 ( .A(a[1391]), .B(n4242), .Z(n4241) );
  IV U4901 ( .A(n4239), .Z(n4242) );
  XOR U4902 ( .A(n4243), .B(n4244), .Z(n4239) );
  ANDN U4903 ( .B(n4245), .A(n4246), .Z(n4243) );
  XNOR U4904 ( .A(b[1390]), .B(n4244), .Z(n4245) );
  XNOR U4905 ( .A(b[1390]), .B(n4246), .Z(c[1390]) );
  XNOR U4906 ( .A(a[1390]), .B(n4247), .Z(n4246) );
  IV U4907 ( .A(n4244), .Z(n4247) );
  XOR U4908 ( .A(n4248), .B(n4249), .Z(n4244) );
  ANDN U4909 ( .B(n4250), .A(n4251), .Z(n4248) );
  XNOR U4910 ( .A(b[1389]), .B(n4249), .Z(n4250) );
  XNOR U4911 ( .A(b[138]), .B(n4252), .Z(c[138]) );
  XNOR U4912 ( .A(b[1389]), .B(n4251), .Z(c[1389]) );
  XNOR U4913 ( .A(a[1389]), .B(n4253), .Z(n4251) );
  IV U4914 ( .A(n4249), .Z(n4253) );
  XOR U4915 ( .A(n4254), .B(n4255), .Z(n4249) );
  ANDN U4916 ( .B(n4256), .A(n4257), .Z(n4254) );
  XNOR U4917 ( .A(b[1388]), .B(n4255), .Z(n4256) );
  XNOR U4918 ( .A(b[1388]), .B(n4257), .Z(c[1388]) );
  XNOR U4919 ( .A(a[1388]), .B(n4258), .Z(n4257) );
  IV U4920 ( .A(n4255), .Z(n4258) );
  XOR U4921 ( .A(n4259), .B(n4260), .Z(n4255) );
  ANDN U4922 ( .B(n4261), .A(n4262), .Z(n4259) );
  XNOR U4923 ( .A(b[1387]), .B(n4260), .Z(n4261) );
  XNOR U4924 ( .A(b[1387]), .B(n4262), .Z(c[1387]) );
  XNOR U4925 ( .A(a[1387]), .B(n4263), .Z(n4262) );
  IV U4926 ( .A(n4260), .Z(n4263) );
  XOR U4927 ( .A(n4264), .B(n4265), .Z(n4260) );
  ANDN U4928 ( .B(n4266), .A(n4267), .Z(n4264) );
  XNOR U4929 ( .A(b[1386]), .B(n4265), .Z(n4266) );
  XNOR U4930 ( .A(b[1386]), .B(n4267), .Z(c[1386]) );
  XNOR U4931 ( .A(a[1386]), .B(n4268), .Z(n4267) );
  IV U4932 ( .A(n4265), .Z(n4268) );
  XOR U4933 ( .A(n4269), .B(n4270), .Z(n4265) );
  ANDN U4934 ( .B(n4271), .A(n4272), .Z(n4269) );
  XNOR U4935 ( .A(b[1385]), .B(n4270), .Z(n4271) );
  XNOR U4936 ( .A(b[1385]), .B(n4272), .Z(c[1385]) );
  XNOR U4937 ( .A(a[1385]), .B(n4273), .Z(n4272) );
  IV U4938 ( .A(n4270), .Z(n4273) );
  XOR U4939 ( .A(n4274), .B(n4275), .Z(n4270) );
  ANDN U4940 ( .B(n4276), .A(n4277), .Z(n4274) );
  XNOR U4941 ( .A(b[1384]), .B(n4275), .Z(n4276) );
  XNOR U4942 ( .A(b[1384]), .B(n4277), .Z(c[1384]) );
  XNOR U4943 ( .A(a[1384]), .B(n4278), .Z(n4277) );
  IV U4944 ( .A(n4275), .Z(n4278) );
  XOR U4945 ( .A(n4279), .B(n4280), .Z(n4275) );
  ANDN U4946 ( .B(n4281), .A(n4282), .Z(n4279) );
  XNOR U4947 ( .A(b[1383]), .B(n4280), .Z(n4281) );
  XNOR U4948 ( .A(b[1383]), .B(n4282), .Z(c[1383]) );
  XNOR U4949 ( .A(a[1383]), .B(n4283), .Z(n4282) );
  IV U4950 ( .A(n4280), .Z(n4283) );
  XOR U4951 ( .A(n4284), .B(n4285), .Z(n4280) );
  ANDN U4952 ( .B(n4286), .A(n4287), .Z(n4284) );
  XNOR U4953 ( .A(b[1382]), .B(n4285), .Z(n4286) );
  XNOR U4954 ( .A(b[1382]), .B(n4287), .Z(c[1382]) );
  XNOR U4955 ( .A(a[1382]), .B(n4288), .Z(n4287) );
  IV U4956 ( .A(n4285), .Z(n4288) );
  XOR U4957 ( .A(n4289), .B(n4290), .Z(n4285) );
  ANDN U4958 ( .B(n4291), .A(n4292), .Z(n4289) );
  XNOR U4959 ( .A(b[1381]), .B(n4290), .Z(n4291) );
  XNOR U4960 ( .A(b[1381]), .B(n4292), .Z(c[1381]) );
  XNOR U4961 ( .A(a[1381]), .B(n4293), .Z(n4292) );
  IV U4962 ( .A(n4290), .Z(n4293) );
  XOR U4963 ( .A(n4294), .B(n4295), .Z(n4290) );
  ANDN U4964 ( .B(n4296), .A(n4297), .Z(n4294) );
  XNOR U4965 ( .A(b[1380]), .B(n4295), .Z(n4296) );
  XNOR U4966 ( .A(b[1380]), .B(n4297), .Z(c[1380]) );
  XNOR U4967 ( .A(a[1380]), .B(n4298), .Z(n4297) );
  IV U4968 ( .A(n4295), .Z(n4298) );
  XOR U4969 ( .A(n4299), .B(n4300), .Z(n4295) );
  ANDN U4970 ( .B(n4301), .A(n4302), .Z(n4299) );
  XNOR U4971 ( .A(b[1379]), .B(n4300), .Z(n4301) );
  XNOR U4972 ( .A(b[137]), .B(n4303), .Z(c[137]) );
  XNOR U4973 ( .A(b[1379]), .B(n4302), .Z(c[1379]) );
  XNOR U4974 ( .A(a[1379]), .B(n4304), .Z(n4302) );
  IV U4975 ( .A(n4300), .Z(n4304) );
  XOR U4976 ( .A(n4305), .B(n4306), .Z(n4300) );
  ANDN U4977 ( .B(n4307), .A(n4308), .Z(n4305) );
  XNOR U4978 ( .A(b[1378]), .B(n4306), .Z(n4307) );
  XNOR U4979 ( .A(b[1378]), .B(n4308), .Z(c[1378]) );
  XNOR U4980 ( .A(a[1378]), .B(n4309), .Z(n4308) );
  IV U4981 ( .A(n4306), .Z(n4309) );
  XOR U4982 ( .A(n4310), .B(n4311), .Z(n4306) );
  ANDN U4983 ( .B(n4312), .A(n4313), .Z(n4310) );
  XNOR U4984 ( .A(b[1377]), .B(n4311), .Z(n4312) );
  XNOR U4985 ( .A(b[1377]), .B(n4313), .Z(c[1377]) );
  XNOR U4986 ( .A(a[1377]), .B(n4314), .Z(n4313) );
  IV U4987 ( .A(n4311), .Z(n4314) );
  XOR U4988 ( .A(n4315), .B(n4316), .Z(n4311) );
  ANDN U4989 ( .B(n4317), .A(n4318), .Z(n4315) );
  XNOR U4990 ( .A(b[1376]), .B(n4316), .Z(n4317) );
  XNOR U4991 ( .A(b[1376]), .B(n4318), .Z(c[1376]) );
  XNOR U4992 ( .A(a[1376]), .B(n4319), .Z(n4318) );
  IV U4993 ( .A(n4316), .Z(n4319) );
  XOR U4994 ( .A(n4320), .B(n4321), .Z(n4316) );
  ANDN U4995 ( .B(n4322), .A(n4323), .Z(n4320) );
  XNOR U4996 ( .A(b[1375]), .B(n4321), .Z(n4322) );
  XNOR U4997 ( .A(b[1375]), .B(n4323), .Z(c[1375]) );
  XNOR U4998 ( .A(a[1375]), .B(n4324), .Z(n4323) );
  IV U4999 ( .A(n4321), .Z(n4324) );
  XOR U5000 ( .A(n4325), .B(n4326), .Z(n4321) );
  ANDN U5001 ( .B(n4327), .A(n4328), .Z(n4325) );
  XNOR U5002 ( .A(b[1374]), .B(n4326), .Z(n4327) );
  XNOR U5003 ( .A(b[1374]), .B(n4328), .Z(c[1374]) );
  XNOR U5004 ( .A(a[1374]), .B(n4329), .Z(n4328) );
  IV U5005 ( .A(n4326), .Z(n4329) );
  XOR U5006 ( .A(n4330), .B(n4331), .Z(n4326) );
  ANDN U5007 ( .B(n4332), .A(n4333), .Z(n4330) );
  XNOR U5008 ( .A(b[1373]), .B(n4331), .Z(n4332) );
  XNOR U5009 ( .A(b[1373]), .B(n4333), .Z(c[1373]) );
  XNOR U5010 ( .A(a[1373]), .B(n4334), .Z(n4333) );
  IV U5011 ( .A(n4331), .Z(n4334) );
  XOR U5012 ( .A(n4335), .B(n4336), .Z(n4331) );
  ANDN U5013 ( .B(n4337), .A(n4338), .Z(n4335) );
  XNOR U5014 ( .A(b[1372]), .B(n4336), .Z(n4337) );
  XNOR U5015 ( .A(b[1372]), .B(n4338), .Z(c[1372]) );
  XNOR U5016 ( .A(a[1372]), .B(n4339), .Z(n4338) );
  IV U5017 ( .A(n4336), .Z(n4339) );
  XOR U5018 ( .A(n4340), .B(n4341), .Z(n4336) );
  ANDN U5019 ( .B(n4342), .A(n4343), .Z(n4340) );
  XNOR U5020 ( .A(b[1371]), .B(n4341), .Z(n4342) );
  XNOR U5021 ( .A(b[1371]), .B(n4343), .Z(c[1371]) );
  XNOR U5022 ( .A(a[1371]), .B(n4344), .Z(n4343) );
  IV U5023 ( .A(n4341), .Z(n4344) );
  XOR U5024 ( .A(n4345), .B(n4346), .Z(n4341) );
  ANDN U5025 ( .B(n4347), .A(n4348), .Z(n4345) );
  XNOR U5026 ( .A(b[1370]), .B(n4346), .Z(n4347) );
  XNOR U5027 ( .A(b[1370]), .B(n4348), .Z(c[1370]) );
  XNOR U5028 ( .A(a[1370]), .B(n4349), .Z(n4348) );
  IV U5029 ( .A(n4346), .Z(n4349) );
  XOR U5030 ( .A(n4350), .B(n4351), .Z(n4346) );
  ANDN U5031 ( .B(n4352), .A(n4353), .Z(n4350) );
  XNOR U5032 ( .A(b[1369]), .B(n4351), .Z(n4352) );
  XNOR U5033 ( .A(b[136]), .B(n4354), .Z(c[136]) );
  XNOR U5034 ( .A(b[1369]), .B(n4353), .Z(c[1369]) );
  XNOR U5035 ( .A(a[1369]), .B(n4355), .Z(n4353) );
  IV U5036 ( .A(n4351), .Z(n4355) );
  XOR U5037 ( .A(n4356), .B(n4357), .Z(n4351) );
  ANDN U5038 ( .B(n4358), .A(n4359), .Z(n4356) );
  XNOR U5039 ( .A(b[1368]), .B(n4357), .Z(n4358) );
  XNOR U5040 ( .A(b[1368]), .B(n4359), .Z(c[1368]) );
  XNOR U5041 ( .A(a[1368]), .B(n4360), .Z(n4359) );
  IV U5042 ( .A(n4357), .Z(n4360) );
  XOR U5043 ( .A(n4361), .B(n4362), .Z(n4357) );
  ANDN U5044 ( .B(n4363), .A(n4364), .Z(n4361) );
  XNOR U5045 ( .A(b[1367]), .B(n4362), .Z(n4363) );
  XNOR U5046 ( .A(b[1367]), .B(n4364), .Z(c[1367]) );
  XNOR U5047 ( .A(a[1367]), .B(n4365), .Z(n4364) );
  IV U5048 ( .A(n4362), .Z(n4365) );
  XOR U5049 ( .A(n4366), .B(n4367), .Z(n4362) );
  ANDN U5050 ( .B(n4368), .A(n4369), .Z(n4366) );
  XNOR U5051 ( .A(b[1366]), .B(n4367), .Z(n4368) );
  XNOR U5052 ( .A(b[1366]), .B(n4369), .Z(c[1366]) );
  XNOR U5053 ( .A(a[1366]), .B(n4370), .Z(n4369) );
  IV U5054 ( .A(n4367), .Z(n4370) );
  XOR U5055 ( .A(n4371), .B(n4372), .Z(n4367) );
  ANDN U5056 ( .B(n4373), .A(n4374), .Z(n4371) );
  XNOR U5057 ( .A(b[1365]), .B(n4372), .Z(n4373) );
  XNOR U5058 ( .A(b[1365]), .B(n4374), .Z(c[1365]) );
  XNOR U5059 ( .A(a[1365]), .B(n4375), .Z(n4374) );
  IV U5060 ( .A(n4372), .Z(n4375) );
  XOR U5061 ( .A(n4376), .B(n4377), .Z(n4372) );
  ANDN U5062 ( .B(n4378), .A(n4379), .Z(n4376) );
  XNOR U5063 ( .A(b[1364]), .B(n4377), .Z(n4378) );
  XNOR U5064 ( .A(b[1364]), .B(n4379), .Z(c[1364]) );
  XNOR U5065 ( .A(a[1364]), .B(n4380), .Z(n4379) );
  IV U5066 ( .A(n4377), .Z(n4380) );
  XOR U5067 ( .A(n4381), .B(n4382), .Z(n4377) );
  ANDN U5068 ( .B(n4383), .A(n4384), .Z(n4381) );
  XNOR U5069 ( .A(b[1363]), .B(n4382), .Z(n4383) );
  XNOR U5070 ( .A(b[1363]), .B(n4384), .Z(c[1363]) );
  XNOR U5071 ( .A(a[1363]), .B(n4385), .Z(n4384) );
  IV U5072 ( .A(n4382), .Z(n4385) );
  XOR U5073 ( .A(n4386), .B(n4387), .Z(n4382) );
  ANDN U5074 ( .B(n4388), .A(n4389), .Z(n4386) );
  XNOR U5075 ( .A(b[1362]), .B(n4387), .Z(n4388) );
  XNOR U5076 ( .A(b[1362]), .B(n4389), .Z(c[1362]) );
  XNOR U5077 ( .A(a[1362]), .B(n4390), .Z(n4389) );
  IV U5078 ( .A(n4387), .Z(n4390) );
  XOR U5079 ( .A(n4391), .B(n4392), .Z(n4387) );
  ANDN U5080 ( .B(n4393), .A(n4394), .Z(n4391) );
  XNOR U5081 ( .A(b[1361]), .B(n4392), .Z(n4393) );
  XNOR U5082 ( .A(b[1361]), .B(n4394), .Z(c[1361]) );
  XNOR U5083 ( .A(a[1361]), .B(n4395), .Z(n4394) );
  IV U5084 ( .A(n4392), .Z(n4395) );
  XOR U5085 ( .A(n4396), .B(n4397), .Z(n4392) );
  ANDN U5086 ( .B(n4398), .A(n4399), .Z(n4396) );
  XNOR U5087 ( .A(b[1360]), .B(n4397), .Z(n4398) );
  XNOR U5088 ( .A(b[1360]), .B(n4399), .Z(c[1360]) );
  XNOR U5089 ( .A(a[1360]), .B(n4400), .Z(n4399) );
  IV U5090 ( .A(n4397), .Z(n4400) );
  XOR U5091 ( .A(n4401), .B(n4402), .Z(n4397) );
  ANDN U5092 ( .B(n4403), .A(n4404), .Z(n4401) );
  XNOR U5093 ( .A(b[1359]), .B(n4402), .Z(n4403) );
  XNOR U5094 ( .A(b[135]), .B(n4405), .Z(c[135]) );
  XNOR U5095 ( .A(b[1359]), .B(n4404), .Z(c[1359]) );
  XNOR U5096 ( .A(a[1359]), .B(n4406), .Z(n4404) );
  IV U5097 ( .A(n4402), .Z(n4406) );
  XOR U5098 ( .A(n4407), .B(n4408), .Z(n4402) );
  ANDN U5099 ( .B(n4409), .A(n4410), .Z(n4407) );
  XNOR U5100 ( .A(b[1358]), .B(n4408), .Z(n4409) );
  XNOR U5101 ( .A(b[1358]), .B(n4410), .Z(c[1358]) );
  XNOR U5102 ( .A(a[1358]), .B(n4411), .Z(n4410) );
  IV U5103 ( .A(n4408), .Z(n4411) );
  XOR U5104 ( .A(n4412), .B(n4413), .Z(n4408) );
  ANDN U5105 ( .B(n4414), .A(n4415), .Z(n4412) );
  XNOR U5106 ( .A(b[1357]), .B(n4413), .Z(n4414) );
  XNOR U5107 ( .A(b[1357]), .B(n4415), .Z(c[1357]) );
  XNOR U5108 ( .A(a[1357]), .B(n4416), .Z(n4415) );
  IV U5109 ( .A(n4413), .Z(n4416) );
  XOR U5110 ( .A(n4417), .B(n4418), .Z(n4413) );
  ANDN U5111 ( .B(n4419), .A(n4420), .Z(n4417) );
  XNOR U5112 ( .A(b[1356]), .B(n4418), .Z(n4419) );
  XNOR U5113 ( .A(b[1356]), .B(n4420), .Z(c[1356]) );
  XNOR U5114 ( .A(a[1356]), .B(n4421), .Z(n4420) );
  IV U5115 ( .A(n4418), .Z(n4421) );
  XOR U5116 ( .A(n4422), .B(n4423), .Z(n4418) );
  ANDN U5117 ( .B(n4424), .A(n4425), .Z(n4422) );
  XNOR U5118 ( .A(b[1355]), .B(n4423), .Z(n4424) );
  XNOR U5119 ( .A(b[1355]), .B(n4425), .Z(c[1355]) );
  XNOR U5120 ( .A(a[1355]), .B(n4426), .Z(n4425) );
  IV U5121 ( .A(n4423), .Z(n4426) );
  XOR U5122 ( .A(n4427), .B(n4428), .Z(n4423) );
  ANDN U5123 ( .B(n4429), .A(n4430), .Z(n4427) );
  XNOR U5124 ( .A(b[1354]), .B(n4428), .Z(n4429) );
  XNOR U5125 ( .A(b[1354]), .B(n4430), .Z(c[1354]) );
  XNOR U5126 ( .A(a[1354]), .B(n4431), .Z(n4430) );
  IV U5127 ( .A(n4428), .Z(n4431) );
  XOR U5128 ( .A(n4432), .B(n4433), .Z(n4428) );
  ANDN U5129 ( .B(n4434), .A(n4435), .Z(n4432) );
  XNOR U5130 ( .A(b[1353]), .B(n4433), .Z(n4434) );
  XNOR U5131 ( .A(b[1353]), .B(n4435), .Z(c[1353]) );
  XNOR U5132 ( .A(a[1353]), .B(n4436), .Z(n4435) );
  IV U5133 ( .A(n4433), .Z(n4436) );
  XOR U5134 ( .A(n4437), .B(n4438), .Z(n4433) );
  ANDN U5135 ( .B(n4439), .A(n4440), .Z(n4437) );
  XNOR U5136 ( .A(b[1352]), .B(n4438), .Z(n4439) );
  XNOR U5137 ( .A(b[1352]), .B(n4440), .Z(c[1352]) );
  XNOR U5138 ( .A(a[1352]), .B(n4441), .Z(n4440) );
  IV U5139 ( .A(n4438), .Z(n4441) );
  XOR U5140 ( .A(n4442), .B(n4443), .Z(n4438) );
  ANDN U5141 ( .B(n4444), .A(n4445), .Z(n4442) );
  XNOR U5142 ( .A(b[1351]), .B(n4443), .Z(n4444) );
  XNOR U5143 ( .A(b[1351]), .B(n4445), .Z(c[1351]) );
  XNOR U5144 ( .A(a[1351]), .B(n4446), .Z(n4445) );
  IV U5145 ( .A(n4443), .Z(n4446) );
  XOR U5146 ( .A(n4447), .B(n4448), .Z(n4443) );
  ANDN U5147 ( .B(n4449), .A(n4450), .Z(n4447) );
  XNOR U5148 ( .A(b[1350]), .B(n4448), .Z(n4449) );
  XNOR U5149 ( .A(b[1350]), .B(n4450), .Z(c[1350]) );
  XNOR U5150 ( .A(a[1350]), .B(n4451), .Z(n4450) );
  IV U5151 ( .A(n4448), .Z(n4451) );
  XOR U5152 ( .A(n4452), .B(n4453), .Z(n4448) );
  ANDN U5153 ( .B(n4454), .A(n4455), .Z(n4452) );
  XNOR U5154 ( .A(b[1349]), .B(n4453), .Z(n4454) );
  XNOR U5155 ( .A(b[134]), .B(n4456), .Z(c[134]) );
  XNOR U5156 ( .A(b[1349]), .B(n4455), .Z(c[1349]) );
  XNOR U5157 ( .A(a[1349]), .B(n4457), .Z(n4455) );
  IV U5158 ( .A(n4453), .Z(n4457) );
  XOR U5159 ( .A(n4458), .B(n4459), .Z(n4453) );
  ANDN U5160 ( .B(n4460), .A(n4461), .Z(n4458) );
  XNOR U5161 ( .A(b[1348]), .B(n4459), .Z(n4460) );
  XNOR U5162 ( .A(b[1348]), .B(n4461), .Z(c[1348]) );
  XNOR U5163 ( .A(a[1348]), .B(n4462), .Z(n4461) );
  IV U5164 ( .A(n4459), .Z(n4462) );
  XOR U5165 ( .A(n4463), .B(n4464), .Z(n4459) );
  ANDN U5166 ( .B(n4465), .A(n4466), .Z(n4463) );
  XNOR U5167 ( .A(b[1347]), .B(n4464), .Z(n4465) );
  XNOR U5168 ( .A(b[1347]), .B(n4466), .Z(c[1347]) );
  XNOR U5169 ( .A(a[1347]), .B(n4467), .Z(n4466) );
  IV U5170 ( .A(n4464), .Z(n4467) );
  XOR U5171 ( .A(n4468), .B(n4469), .Z(n4464) );
  ANDN U5172 ( .B(n4470), .A(n4471), .Z(n4468) );
  XNOR U5173 ( .A(b[1346]), .B(n4469), .Z(n4470) );
  XNOR U5174 ( .A(b[1346]), .B(n4471), .Z(c[1346]) );
  XNOR U5175 ( .A(a[1346]), .B(n4472), .Z(n4471) );
  IV U5176 ( .A(n4469), .Z(n4472) );
  XOR U5177 ( .A(n4473), .B(n4474), .Z(n4469) );
  ANDN U5178 ( .B(n4475), .A(n4476), .Z(n4473) );
  XNOR U5179 ( .A(b[1345]), .B(n4474), .Z(n4475) );
  XNOR U5180 ( .A(b[1345]), .B(n4476), .Z(c[1345]) );
  XNOR U5181 ( .A(a[1345]), .B(n4477), .Z(n4476) );
  IV U5182 ( .A(n4474), .Z(n4477) );
  XOR U5183 ( .A(n4478), .B(n4479), .Z(n4474) );
  ANDN U5184 ( .B(n4480), .A(n4481), .Z(n4478) );
  XNOR U5185 ( .A(b[1344]), .B(n4479), .Z(n4480) );
  XNOR U5186 ( .A(b[1344]), .B(n4481), .Z(c[1344]) );
  XNOR U5187 ( .A(a[1344]), .B(n4482), .Z(n4481) );
  IV U5188 ( .A(n4479), .Z(n4482) );
  XOR U5189 ( .A(n4483), .B(n4484), .Z(n4479) );
  ANDN U5190 ( .B(n4485), .A(n4486), .Z(n4483) );
  XNOR U5191 ( .A(b[1343]), .B(n4484), .Z(n4485) );
  XNOR U5192 ( .A(b[1343]), .B(n4486), .Z(c[1343]) );
  XNOR U5193 ( .A(a[1343]), .B(n4487), .Z(n4486) );
  IV U5194 ( .A(n4484), .Z(n4487) );
  XOR U5195 ( .A(n4488), .B(n4489), .Z(n4484) );
  ANDN U5196 ( .B(n4490), .A(n4491), .Z(n4488) );
  XNOR U5197 ( .A(b[1342]), .B(n4489), .Z(n4490) );
  XNOR U5198 ( .A(b[1342]), .B(n4491), .Z(c[1342]) );
  XNOR U5199 ( .A(a[1342]), .B(n4492), .Z(n4491) );
  IV U5200 ( .A(n4489), .Z(n4492) );
  XOR U5201 ( .A(n4493), .B(n4494), .Z(n4489) );
  ANDN U5202 ( .B(n4495), .A(n4496), .Z(n4493) );
  XNOR U5203 ( .A(b[1341]), .B(n4494), .Z(n4495) );
  XNOR U5204 ( .A(b[1341]), .B(n4496), .Z(c[1341]) );
  XNOR U5205 ( .A(a[1341]), .B(n4497), .Z(n4496) );
  IV U5206 ( .A(n4494), .Z(n4497) );
  XOR U5207 ( .A(n4498), .B(n4499), .Z(n4494) );
  ANDN U5208 ( .B(n4500), .A(n4501), .Z(n4498) );
  XNOR U5209 ( .A(b[1340]), .B(n4499), .Z(n4500) );
  XNOR U5210 ( .A(b[1340]), .B(n4501), .Z(c[1340]) );
  XNOR U5211 ( .A(a[1340]), .B(n4502), .Z(n4501) );
  IV U5212 ( .A(n4499), .Z(n4502) );
  XOR U5213 ( .A(n4503), .B(n4504), .Z(n4499) );
  ANDN U5214 ( .B(n4505), .A(n4506), .Z(n4503) );
  XNOR U5215 ( .A(b[1339]), .B(n4504), .Z(n4505) );
  XNOR U5216 ( .A(b[133]), .B(n4507), .Z(c[133]) );
  XNOR U5217 ( .A(b[1339]), .B(n4506), .Z(c[1339]) );
  XNOR U5218 ( .A(a[1339]), .B(n4508), .Z(n4506) );
  IV U5219 ( .A(n4504), .Z(n4508) );
  XOR U5220 ( .A(n4509), .B(n4510), .Z(n4504) );
  ANDN U5221 ( .B(n4511), .A(n4512), .Z(n4509) );
  XNOR U5222 ( .A(b[1338]), .B(n4510), .Z(n4511) );
  XNOR U5223 ( .A(b[1338]), .B(n4512), .Z(c[1338]) );
  XNOR U5224 ( .A(a[1338]), .B(n4513), .Z(n4512) );
  IV U5225 ( .A(n4510), .Z(n4513) );
  XOR U5226 ( .A(n4514), .B(n4515), .Z(n4510) );
  ANDN U5227 ( .B(n4516), .A(n4517), .Z(n4514) );
  XNOR U5228 ( .A(b[1337]), .B(n4515), .Z(n4516) );
  XNOR U5229 ( .A(b[1337]), .B(n4517), .Z(c[1337]) );
  XNOR U5230 ( .A(a[1337]), .B(n4518), .Z(n4517) );
  IV U5231 ( .A(n4515), .Z(n4518) );
  XOR U5232 ( .A(n4519), .B(n4520), .Z(n4515) );
  ANDN U5233 ( .B(n4521), .A(n4522), .Z(n4519) );
  XNOR U5234 ( .A(b[1336]), .B(n4520), .Z(n4521) );
  XNOR U5235 ( .A(b[1336]), .B(n4522), .Z(c[1336]) );
  XNOR U5236 ( .A(a[1336]), .B(n4523), .Z(n4522) );
  IV U5237 ( .A(n4520), .Z(n4523) );
  XOR U5238 ( .A(n4524), .B(n4525), .Z(n4520) );
  ANDN U5239 ( .B(n4526), .A(n4527), .Z(n4524) );
  XNOR U5240 ( .A(b[1335]), .B(n4525), .Z(n4526) );
  XNOR U5241 ( .A(b[1335]), .B(n4527), .Z(c[1335]) );
  XNOR U5242 ( .A(a[1335]), .B(n4528), .Z(n4527) );
  IV U5243 ( .A(n4525), .Z(n4528) );
  XOR U5244 ( .A(n4529), .B(n4530), .Z(n4525) );
  ANDN U5245 ( .B(n4531), .A(n4532), .Z(n4529) );
  XNOR U5246 ( .A(b[1334]), .B(n4530), .Z(n4531) );
  XNOR U5247 ( .A(b[1334]), .B(n4532), .Z(c[1334]) );
  XNOR U5248 ( .A(a[1334]), .B(n4533), .Z(n4532) );
  IV U5249 ( .A(n4530), .Z(n4533) );
  XOR U5250 ( .A(n4534), .B(n4535), .Z(n4530) );
  ANDN U5251 ( .B(n4536), .A(n4537), .Z(n4534) );
  XNOR U5252 ( .A(b[1333]), .B(n4535), .Z(n4536) );
  XNOR U5253 ( .A(b[1333]), .B(n4537), .Z(c[1333]) );
  XNOR U5254 ( .A(a[1333]), .B(n4538), .Z(n4537) );
  IV U5255 ( .A(n4535), .Z(n4538) );
  XOR U5256 ( .A(n4539), .B(n4540), .Z(n4535) );
  ANDN U5257 ( .B(n4541), .A(n4542), .Z(n4539) );
  XNOR U5258 ( .A(b[1332]), .B(n4540), .Z(n4541) );
  XNOR U5259 ( .A(b[1332]), .B(n4542), .Z(c[1332]) );
  XNOR U5260 ( .A(a[1332]), .B(n4543), .Z(n4542) );
  IV U5261 ( .A(n4540), .Z(n4543) );
  XOR U5262 ( .A(n4544), .B(n4545), .Z(n4540) );
  ANDN U5263 ( .B(n4546), .A(n4547), .Z(n4544) );
  XNOR U5264 ( .A(b[1331]), .B(n4545), .Z(n4546) );
  XNOR U5265 ( .A(b[1331]), .B(n4547), .Z(c[1331]) );
  XNOR U5266 ( .A(a[1331]), .B(n4548), .Z(n4547) );
  IV U5267 ( .A(n4545), .Z(n4548) );
  XOR U5268 ( .A(n4549), .B(n4550), .Z(n4545) );
  ANDN U5269 ( .B(n4551), .A(n4552), .Z(n4549) );
  XNOR U5270 ( .A(b[1330]), .B(n4550), .Z(n4551) );
  XNOR U5271 ( .A(b[1330]), .B(n4552), .Z(c[1330]) );
  XNOR U5272 ( .A(a[1330]), .B(n4553), .Z(n4552) );
  IV U5273 ( .A(n4550), .Z(n4553) );
  XOR U5274 ( .A(n4554), .B(n4555), .Z(n4550) );
  ANDN U5275 ( .B(n4556), .A(n4557), .Z(n4554) );
  XNOR U5276 ( .A(b[1329]), .B(n4555), .Z(n4556) );
  XNOR U5277 ( .A(b[132]), .B(n4558), .Z(c[132]) );
  XNOR U5278 ( .A(b[1329]), .B(n4557), .Z(c[1329]) );
  XNOR U5279 ( .A(a[1329]), .B(n4559), .Z(n4557) );
  IV U5280 ( .A(n4555), .Z(n4559) );
  XOR U5281 ( .A(n4560), .B(n4561), .Z(n4555) );
  ANDN U5282 ( .B(n4562), .A(n4563), .Z(n4560) );
  XNOR U5283 ( .A(b[1328]), .B(n4561), .Z(n4562) );
  XNOR U5284 ( .A(b[1328]), .B(n4563), .Z(c[1328]) );
  XNOR U5285 ( .A(a[1328]), .B(n4564), .Z(n4563) );
  IV U5286 ( .A(n4561), .Z(n4564) );
  XOR U5287 ( .A(n4565), .B(n4566), .Z(n4561) );
  ANDN U5288 ( .B(n4567), .A(n4568), .Z(n4565) );
  XNOR U5289 ( .A(b[1327]), .B(n4566), .Z(n4567) );
  XNOR U5290 ( .A(b[1327]), .B(n4568), .Z(c[1327]) );
  XNOR U5291 ( .A(a[1327]), .B(n4569), .Z(n4568) );
  IV U5292 ( .A(n4566), .Z(n4569) );
  XOR U5293 ( .A(n4570), .B(n4571), .Z(n4566) );
  ANDN U5294 ( .B(n4572), .A(n4573), .Z(n4570) );
  XNOR U5295 ( .A(b[1326]), .B(n4571), .Z(n4572) );
  XNOR U5296 ( .A(b[1326]), .B(n4573), .Z(c[1326]) );
  XNOR U5297 ( .A(a[1326]), .B(n4574), .Z(n4573) );
  IV U5298 ( .A(n4571), .Z(n4574) );
  XOR U5299 ( .A(n4575), .B(n4576), .Z(n4571) );
  ANDN U5300 ( .B(n4577), .A(n4578), .Z(n4575) );
  XNOR U5301 ( .A(b[1325]), .B(n4576), .Z(n4577) );
  XNOR U5302 ( .A(b[1325]), .B(n4578), .Z(c[1325]) );
  XNOR U5303 ( .A(a[1325]), .B(n4579), .Z(n4578) );
  IV U5304 ( .A(n4576), .Z(n4579) );
  XOR U5305 ( .A(n4580), .B(n4581), .Z(n4576) );
  ANDN U5306 ( .B(n4582), .A(n4583), .Z(n4580) );
  XNOR U5307 ( .A(b[1324]), .B(n4581), .Z(n4582) );
  XNOR U5308 ( .A(b[1324]), .B(n4583), .Z(c[1324]) );
  XNOR U5309 ( .A(a[1324]), .B(n4584), .Z(n4583) );
  IV U5310 ( .A(n4581), .Z(n4584) );
  XOR U5311 ( .A(n4585), .B(n4586), .Z(n4581) );
  ANDN U5312 ( .B(n4587), .A(n4588), .Z(n4585) );
  XNOR U5313 ( .A(b[1323]), .B(n4586), .Z(n4587) );
  XNOR U5314 ( .A(b[1323]), .B(n4588), .Z(c[1323]) );
  XNOR U5315 ( .A(a[1323]), .B(n4589), .Z(n4588) );
  IV U5316 ( .A(n4586), .Z(n4589) );
  XOR U5317 ( .A(n4590), .B(n4591), .Z(n4586) );
  ANDN U5318 ( .B(n4592), .A(n4593), .Z(n4590) );
  XNOR U5319 ( .A(b[1322]), .B(n4591), .Z(n4592) );
  XNOR U5320 ( .A(b[1322]), .B(n4593), .Z(c[1322]) );
  XNOR U5321 ( .A(a[1322]), .B(n4594), .Z(n4593) );
  IV U5322 ( .A(n4591), .Z(n4594) );
  XOR U5323 ( .A(n4595), .B(n4596), .Z(n4591) );
  ANDN U5324 ( .B(n4597), .A(n4598), .Z(n4595) );
  XNOR U5325 ( .A(b[1321]), .B(n4596), .Z(n4597) );
  XNOR U5326 ( .A(b[1321]), .B(n4598), .Z(c[1321]) );
  XNOR U5327 ( .A(a[1321]), .B(n4599), .Z(n4598) );
  IV U5328 ( .A(n4596), .Z(n4599) );
  XOR U5329 ( .A(n4600), .B(n4601), .Z(n4596) );
  ANDN U5330 ( .B(n4602), .A(n4603), .Z(n4600) );
  XNOR U5331 ( .A(b[1320]), .B(n4601), .Z(n4602) );
  XNOR U5332 ( .A(b[1320]), .B(n4603), .Z(c[1320]) );
  XNOR U5333 ( .A(a[1320]), .B(n4604), .Z(n4603) );
  IV U5334 ( .A(n4601), .Z(n4604) );
  XOR U5335 ( .A(n4605), .B(n4606), .Z(n4601) );
  ANDN U5336 ( .B(n4607), .A(n4608), .Z(n4605) );
  XNOR U5337 ( .A(b[1319]), .B(n4606), .Z(n4607) );
  XNOR U5338 ( .A(b[131]), .B(n4609), .Z(c[131]) );
  XNOR U5339 ( .A(b[1319]), .B(n4608), .Z(c[1319]) );
  XNOR U5340 ( .A(a[1319]), .B(n4610), .Z(n4608) );
  IV U5341 ( .A(n4606), .Z(n4610) );
  XOR U5342 ( .A(n4611), .B(n4612), .Z(n4606) );
  ANDN U5343 ( .B(n4613), .A(n4614), .Z(n4611) );
  XNOR U5344 ( .A(b[1318]), .B(n4612), .Z(n4613) );
  XNOR U5345 ( .A(b[1318]), .B(n4614), .Z(c[1318]) );
  XNOR U5346 ( .A(a[1318]), .B(n4615), .Z(n4614) );
  IV U5347 ( .A(n4612), .Z(n4615) );
  XOR U5348 ( .A(n4616), .B(n4617), .Z(n4612) );
  ANDN U5349 ( .B(n4618), .A(n4619), .Z(n4616) );
  XNOR U5350 ( .A(b[1317]), .B(n4617), .Z(n4618) );
  XNOR U5351 ( .A(b[1317]), .B(n4619), .Z(c[1317]) );
  XNOR U5352 ( .A(a[1317]), .B(n4620), .Z(n4619) );
  IV U5353 ( .A(n4617), .Z(n4620) );
  XOR U5354 ( .A(n4621), .B(n4622), .Z(n4617) );
  ANDN U5355 ( .B(n4623), .A(n4624), .Z(n4621) );
  XNOR U5356 ( .A(b[1316]), .B(n4622), .Z(n4623) );
  XNOR U5357 ( .A(b[1316]), .B(n4624), .Z(c[1316]) );
  XNOR U5358 ( .A(a[1316]), .B(n4625), .Z(n4624) );
  IV U5359 ( .A(n4622), .Z(n4625) );
  XOR U5360 ( .A(n4626), .B(n4627), .Z(n4622) );
  ANDN U5361 ( .B(n4628), .A(n4629), .Z(n4626) );
  XNOR U5362 ( .A(b[1315]), .B(n4627), .Z(n4628) );
  XNOR U5363 ( .A(b[1315]), .B(n4629), .Z(c[1315]) );
  XNOR U5364 ( .A(a[1315]), .B(n4630), .Z(n4629) );
  IV U5365 ( .A(n4627), .Z(n4630) );
  XOR U5366 ( .A(n4631), .B(n4632), .Z(n4627) );
  ANDN U5367 ( .B(n4633), .A(n4634), .Z(n4631) );
  XNOR U5368 ( .A(b[1314]), .B(n4632), .Z(n4633) );
  XNOR U5369 ( .A(b[1314]), .B(n4634), .Z(c[1314]) );
  XNOR U5370 ( .A(a[1314]), .B(n4635), .Z(n4634) );
  IV U5371 ( .A(n4632), .Z(n4635) );
  XOR U5372 ( .A(n4636), .B(n4637), .Z(n4632) );
  ANDN U5373 ( .B(n4638), .A(n4639), .Z(n4636) );
  XNOR U5374 ( .A(b[1313]), .B(n4637), .Z(n4638) );
  XNOR U5375 ( .A(b[1313]), .B(n4639), .Z(c[1313]) );
  XNOR U5376 ( .A(a[1313]), .B(n4640), .Z(n4639) );
  IV U5377 ( .A(n4637), .Z(n4640) );
  XOR U5378 ( .A(n4641), .B(n4642), .Z(n4637) );
  ANDN U5379 ( .B(n4643), .A(n4644), .Z(n4641) );
  XNOR U5380 ( .A(b[1312]), .B(n4642), .Z(n4643) );
  XNOR U5381 ( .A(b[1312]), .B(n4644), .Z(c[1312]) );
  XNOR U5382 ( .A(a[1312]), .B(n4645), .Z(n4644) );
  IV U5383 ( .A(n4642), .Z(n4645) );
  XOR U5384 ( .A(n4646), .B(n4647), .Z(n4642) );
  ANDN U5385 ( .B(n4648), .A(n4649), .Z(n4646) );
  XNOR U5386 ( .A(b[1311]), .B(n4647), .Z(n4648) );
  XNOR U5387 ( .A(b[1311]), .B(n4649), .Z(c[1311]) );
  XNOR U5388 ( .A(a[1311]), .B(n4650), .Z(n4649) );
  IV U5389 ( .A(n4647), .Z(n4650) );
  XOR U5390 ( .A(n4651), .B(n4652), .Z(n4647) );
  ANDN U5391 ( .B(n4653), .A(n4654), .Z(n4651) );
  XNOR U5392 ( .A(b[1310]), .B(n4652), .Z(n4653) );
  XNOR U5393 ( .A(b[1310]), .B(n4654), .Z(c[1310]) );
  XNOR U5394 ( .A(a[1310]), .B(n4655), .Z(n4654) );
  IV U5395 ( .A(n4652), .Z(n4655) );
  XOR U5396 ( .A(n4656), .B(n4657), .Z(n4652) );
  ANDN U5397 ( .B(n4658), .A(n4659), .Z(n4656) );
  XNOR U5398 ( .A(b[1309]), .B(n4657), .Z(n4658) );
  XNOR U5399 ( .A(b[130]), .B(n4660), .Z(c[130]) );
  XNOR U5400 ( .A(b[1309]), .B(n4659), .Z(c[1309]) );
  XNOR U5401 ( .A(a[1309]), .B(n4661), .Z(n4659) );
  IV U5402 ( .A(n4657), .Z(n4661) );
  XOR U5403 ( .A(n4662), .B(n4663), .Z(n4657) );
  ANDN U5404 ( .B(n4664), .A(n4665), .Z(n4662) );
  XNOR U5405 ( .A(b[1308]), .B(n4663), .Z(n4664) );
  XNOR U5406 ( .A(b[1308]), .B(n4665), .Z(c[1308]) );
  XNOR U5407 ( .A(a[1308]), .B(n4666), .Z(n4665) );
  IV U5408 ( .A(n4663), .Z(n4666) );
  XOR U5409 ( .A(n4667), .B(n4668), .Z(n4663) );
  ANDN U5410 ( .B(n4669), .A(n4670), .Z(n4667) );
  XNOR U5411 ( .A(b[1307]), .B(n4668), .Z(n4669) );
  XNOR U5412 ( .A(b[1307]), .B(n4670), .Z(c[1307]) );
  XNOR U5413 ( .A(a[1307]), .B(n4671), .Z(n4670) );
  IV U5414 ( .A(n4668), .Z(n4671) );
  XOR U5415 ( .A(n4672), .B(n4673), .Z(n4668) );
  ANDN U5416 ( .B(n4674), .A(n4675), .Z(n4672) );
  XNOR U5417 ( .A(b[1306]), .B(n4673), .Z(n4674) );
  XNOR U5418 ( .A(b[1306]), .B(n4675), .Z(c[1306]) );
  XNOR U5419 ( .A(a[1306]), .B(n4676), .Z(n4675) );
  IV U5420 ( .A(n4673), .Z(n4676) );
  XOR U5421 ( .A(n4677), .B(n4678), .Z(n4673) );
  ANDN U5422 ( .B(n4679), .A(n4680), .Z(n4677) );
  XNOR U5423 ( .A(b[1305]), .B(n4678), .Z(n4679) );
  XNOR U5424 ( .A(b[1305]), .B(n4680), .Z(c[1305]) );
  XNOR U5425 ( .A(a[1305]), .B(n4681), .Z(n4680) );
  IV U5426 ( .A(n4678), .Z(n4681) );
  XOR U5427 ( .A(n4682), .B(n4683), .Z(n4678) );
  ANDN U5428 ( .B(n4684), .A(n4685), .Z(n4682) );
  XNOR U5429 ( .A(b[1304]), .B(n4683), .Z(n4684) );
  XNOR U5430 ( .A(b[1304]), .B(n4685), .Z(c[1304]) );
  XNOR U5431 ( .A(a[1304]), .B(n4686), .Z(n4685) );
  IV U5432 ( .A(n4683), .Z(n4686) );
  XOR U5433 ( .A(n4687), .B(n4688), .Z(n4683) );
  ANDN U5434 ( .B(n4689), .A(n4690), .Z(n4687) );
  XNOR U5435 ( .A(b[1303]), .B(n4688), .Z(n4689) );
  XNOR U5436 ( .A(b[1303]), .B(n4690), .Z(c[1303]) );
  XNOR U5437 ( .A(a[1303]), .B(n4691), .Z(n4690) );
  IV U5438 ( .A(n4688), .Z(n4691) );
  XOR U5439 ( .A(n4692), .B(n4693), .Z(n4688) );
  ANDN U5440 ( .B(n4694), .A(n4695), .Z(n4692) );
  XNOR U5441 ( .A(b[1302]), .B(n4693), .Z(n4694) );
  XNOR U5442 ( .A(b[1302]), .B(n4695), .Z(c[1302]) );
  XNOR U5443 ( .A(a[1302]), .B(n4696), .Z(n4695) );
  IV U5444 ( .A(n4693), .Z(n4696) );
  XOR U5445 ( .A(n4697), .B(n4698), .Z(n4693) );
  ANDN U5446 ( .B(n4699), .A(n4700), .Z(n4697) );
  XNOR U5447 ( .A(b[1301]), .B(n4698), .Z(n4699) );
  XNOR U5448 ( .A(b[1301]), .B(n4700), .Z(c[1301]) );
  XNOR U5449 ( .A(a[1301]), .B(n4701), .Z(n4700) );
  IV U5450 ( .A(n4698), .Z(n4701) );
  XOR U5451 ( .A(n4702), .B(n4703), .Z(n4698) );
  ANDN U5452 ( .B(n4704), .A(n4705), .Z(n4702) );
  XNOR U5453 ( .A(b[1300]), .B(n4703), .Z(n4704) );
  XNOR U5454 ( .A(b[1300]), .B(n4705), .Z(c[1300]) );
  XNOR U5455 ( .A(a[1300]), .B(n4706), .Z(n4705) );
  IV U5456 ( .A(n4703), .Z(n4706) );
  XOR U5457 ( .A(n4707), .B(n4708), .Z(n4703) );
  ANDN U5458 ( .B(n4709), .A(n4710), .Z(n4707) );
  XNOR U5459 ( .A(b[1299]), .B(n4708), .Z(n4709) );
  XNOR U5460 ( .A(b[12]), .B(n4711), .Z(c[12]) );
  XNOR U5461 ( .A(b[129]), .B(n4712), .Z(c[129]) );
  XNOR U5462 ( .A(b[1299]), .B(n4710), .Z(c[1299]) );
  XNOR U5463 ( .A(a[1299]), .B(n4713), .Z(n4710) );
  IV U5464 ( .A(n4708), .Z(n4713) );
  XOR U5465 ( .A(n4714), .B(n4715), .Z(n4708) );
  ANDN U5466 ( .B(n4716), .A(n4717), .Z(n4714) );
  XNOR U5467 ( .A(b[1298]), .B(n4715), .Z(n4716) );
  XNOR U5468 ( .A(b[1298]), .B(n4717), .Z(c[1298]) );
  XNOR U5469 ( .A(a[1298]), .B(n4718), .Z(n4717) );
  IV U5470 ( .A(n4715), .Z(n4718) );
  XOR U5471 ( .A(n4719), .B(n4720), .Z(n4715) );
  ANDN U5472 ( .B(n4721), .A(n4722), .Z(n4719) );
  XNOR U5473 ( .A(b[1297]), .B(n4720), .Z(n4721) );
  XNOR U5474 ( .A(b[1297]), .B(n4722), .Z(c[1297]) );
  XNOR U5475 ( .A(a[1297]), .B(n4723), .Z(n4722) );
  IV U5476 ( .A(n4720), .Z(n4723) );
  XOR U5477 ( .A(n4724), .B(n4725), .Z(n4720) );
  ANDN U5478 ( .B(n4726), .A(n4727), .Z(n4724) );
  XNOR U5479 ( .A(b[1296]), .B(n4725), .Z(n4726) );
  XNOR U5480 ( .A(b[1296]), .B(n4727), .Z(c[1296]) );
  XNOR U5481 ( .A(a[1296]), .B(n4728), .Z(n4727) );
  IV U5482 ( .A(n4725), .Z(n4728) );
  XOR U5483 ( .A(n4729), .B(n4730), .Z(n4725) );
  ANDN U5484 ( .B(n4731), .A(n4732), .Z(n4729) );
  XNOR U5485 ( .A(b[1295]), .B(n4730), .Z(n4731) );
  XNOR U5486 ( .A(b[1295]), .B(n4732), .Z(c[1295]) );
  XNOR U5487 ( .A(a[1295]), .B(n4733), .Z(n4732) );
  IV U5488 ( .A(n4730), .Z(n4733) );
  XOR U5489 ( .A(n4734), .B(n4735), .Z(n4730) );
  ANDN U5490 ( .B(n4736), .A(n4737), .Z(n4734) );
  XNOR U5491 ( .A(b[1294]), .B(n4735), .Z(n4736) );
  XNOR U5492 ( .A(b[1294]), .B(n4737), .Z(c[1294]) );
  XNOR U5493 ( .A(a[1294]), .B(n4738), .Z(n4737) );
  IV U5494 ( .A(n4735), .Z(n4738) );
  XOR U5495 ( .A(n4739), .B(n4740), .Z(n4735) );
  ANDN U5496 ( .B(n4741), .A(n4742), .Z(n4739) );
  XNOR U5497 ( .A(b[1293]), .B(n4740), .Z(n4741) );
  XNOR U5498 ( .A(b[1293]), .B(n4742), .Z(c[1293]) );
  XNOR U5499 ( .A(a[1293]), .B(n4743), .Z(n4742) );
  IV U5500 ( .A(n4740), .Z(n4743) );
  XOR U5501 ( .A(n4744), .B(n4745), .Z(n4740) );
  ANDN U5502 ( .B(n4746), .A(n4747), .Z(n4744) );
  XNOR U5503 ( .A(b[1292]), .B(n4745), .Z(n4746) );
  XNOR U5504 ( .A(b[1292]), .B(n4747), .Z(c[1292]) );
  XNOR U5505 ( .A(a[1292]), .B(n4748), .Z(n4747) );
  IV U5506 ( .A(n4745), .Z(n4748) );
  XOR U5507 ( .A(n4749), .B(n4750), .Z(n4745) );
  ANDN U5508 ( .B(n4751), .A(n4752), .Z(n4749) );
  XNOR U5509 ( .A(b[1291]), .B(n4750), .Z(n4751) );
  XNOR U5510 ( .A(b[1291]), .B(n4752), .Z(c[1291]) );
  XNOR U5511 ( .A(a[1291]), .B(n4753), .Z(n4752) );
  IV U5512 ( .A(n4750), .Z(n4753) );
  XOR U5513 ( .A(n4754), .B(n4755), .Z(n4750) );
  ANDN U5514 ( .B(n4756), .A(n4757), .Z(n4754) );
  XNOR U5515 ( .A(b[1290]), .B(n4755), .Z(n4756) );
  XNOR U5516 ( .A(b[1290]), .B(n4757), .Z(c[1290]) );
  XNOR U5517 ( .A(a[1290]), .B(n4758), .Z(n4757) );
  IV U5518 ( .A(n4755), .Z(n4758) );
  XOR U5519 ( .A(n4759), .B(n4760), .Z(n4755) );
  ANDN U5520 ( .B(n4761), .A(n4762), .Z(n4759) );
  XNOR U5521 ( .A(b[1289]), .B(n4760), .Z(n4761) );
  XNOR U5522 ( .A(b[128]), .B(n4763), .Z(c[128]) );
  XNOR U5523 ( .A(b[1289]), .B(n4762), .Z(c[1289]) );
  XNOR U5524 ( .A(a[1289]), .B(n4764), .Z(n4762) );
  IV U5525 ( .A(n4760), .Z(n4764) );
  XOR U5526 ( .A(n4765), .B(n4766), .Z(n4760) );
  ANDN U5527 ( .B(n4767), .A(n4768), .Z(n4765) );
  XNOR U5528 ( .A(b[1288]), .B(n4766), .Z(n4767) );
  XNOR U5529 ( .A(b[1288]), .B(n4768), .Z(c[1288]) );
  XNOR U5530 ( .A(a[1288]), .B(n4769), .Z(n4768) );
  IV U5531 ( .A(n4766), .Z(n4769) );
  XOR U5532 ( .A(n4770), .B(n4771), .Z(n4766) );
  ANDN U5533 ( .B(n4772), .A(n4773), .Z(n4770) );
  XNOR U5534 ( .A(b[1287]), .B(n4771), .Z(n4772) );
  XNOR U5535 ( .A(b[1287]), .B(n4773), .Z(c[1287]) );
  XNOR U5536 ( .A(a[1287]), .B(n4774), .Z(n4773) );
  IV U5537 ( .A(n4771), .Z(n4774) );
  XOR U5538 ( .A(n4775), .B(n4776), .Z(n4771) );
  ANDN U5539 ( .B(n4777), .A(n4778), .Z(n4775) );
  XNOR U5540 ( .A(b[1286]), .B(n4776), .Z(n4777) );
  XNOR U5541 ( .A(b[1286]), .B(n4778), .Z(c[1286]) );
  XNOR U5542 ( .A(a[1286]), .B(n4779), .Z(n4778) );
  IV U5543 ( .A(n4776), .Z(n4779) );
  XOR U5544 ( .A(n4780), .B(n4781), .Z(n4776) );
  ANDN U5545 ( .B(n4782), .A(n4783), .Z(n4780) );
  XNOR U5546 ( .A(b[1285]), .B(n4781), .Z(n4782) );
  XNOR U5547 ( .A(b[1285]), .B(n4783), .Z(c[1285]) );
  XNOR U5548 ( .A(a[1285]), .B(n4784), .Z(n4783) );
  IV U5549 ( .A(n4781), .Z(n4784) );
  XOR U5550 ( .A(n4785), .B(n4786), .Z(n4781) );
  ANDN U5551 ( .B(n4787), .A(n4788), .Z(n4785) );
  XNOR U5552 ( .A(b[1284]), .B(n4786), .Z(n4787) );
  XNOR U5553 ( .A(b[1284]), .B(n4788), .Z(c[1284]) );
  XNOR U5554 ( .A(a[1284]), .B(n4789), .Z(n4788) );
  IV U5555 ( .A(n4786), .Z(n4789) );
  XOR U5556 ( .A(n4790), .B(n4791), .Z(n4786) );
  ANDN U5557 ( .B(n4792), .A(n4793), .Z(n4790) );
  XNOR U5558 ( .A(b[1283]), .B(n4791), .Z(n4792) );
  XNOR U5559 ( .A(b[1283]), .B(n4793), .Z(c[1283]) );
  XNOR U5560 ( .A(a[1283]), .B(n4794), .Z(n4793) );
  IV U5561 ( .A(n4791), .Z(n4794) );
  XOR U5562 ( .A(n4795), .B(n4796), .Z(n4791) );
  ANDN U5563 ( .B(n4797), .A(n4798), .Z(n4795) );
  XNOR U5564 ( .A(b[1282]), .B(n4796), .Z(n4797) );
  XNOR U5565 ( .A(b[1282]), .B(n4798), .Z(c[1282]) );
  XNOR U5566 ( .A(a[1282]), .B(n4799), .Z(n4798) );
  IV U5567 ( .A(n4796), .Z(n4799) );
  XOR U5568 ( .A(n4800), .B(n4801), .Z(n4796) );
  ANDN U5569 ( .B(n4802), .A(n4803), .Z(n4800) );
  XNOR U5570 ( .A(b[1281]), .B(n4801), .Z(n4802) );
  XNOR U5571 ( .A(b[1281]), .B(n4803), .Z(c[1281]) );
  XNOR U5572 ( .A(a[1281]), .B(n4804), .Z(n4803) );
  IV U5573 ( .A(n4801), .Z(n4804) );
  XOR U5574 ( .A(n4805), .B(n4806), .Z(n4801) );
  ANDN U5575 ( .B(n4807), .A(n4808), .Z(n4805) );
  XNOR U5576 ( .A(b[1280]), .B(n4806), .Z(n4807) );
  XNOR U5577 ( .A(b[1280]), .B(n4808), .Z(c[1280]) );
  XNOR U5578 ( .A(a[1280]), .B(n4809), .Z(n4808) );
  IV U5579 ( .A(n4806), .Z(n4809) );
  XOR U5580 ( .A(n4810), .B(n4811), .Z(n4806) );
  ANDN U5581 ( .B(n4812), .A(n4813), .Z(n4810) );
  XNOR U5582 ( .A(b[1279]), .B(n4811), .Z(n4812) );
  XNOR U5583 ( .A(b[127]), .B(n4814), .Z(c[127]) );
  XNOR U5584 ( .A(b[1279]), .B(n4813), .Z(c[1279]) );
  XNOR U5585 ( .A(a[1279]), .B(n4815), .Z(n4813) );
  IV U5586 ( .A(n4811), .Z(n4815) );
  XOR U5587 ( .A(n4816), .B(n4817), .Z(n4811) );
  ANDN U5588 ( .B(n4818), .A(n4819), .Z(n4816) );
  XNOR U5589 ( .A(b[1278]), .B(n4817), .Z(n4818) );
  XNOR U5590 ( .A(b[1278]), .B(n4819), .Z(c[1278]) );
  XNOR U5591 ( .A(a[1278]), .B(n4820), .Z(n4819) );
  IV U5592 ( .A(n4817), .Z(n4820) );
  XOR U5593 ( .A(n4821), .B(n4822), .Z(n4817) );
  ANDN U5594 ( .B(n4823), .A(n4824), .Z(n4821) );
  XNOR U5595 ( .A(b[1277]), .B(n4822), .Z(n4823) );
  XNOR U5596 ( .A(b[1277]), .B(n4824), .Z(c[1277]) );
  XNOR U5597 ( .A(a[1277]), .B(n4825), .Z(n4824) );
  IV U5598 ( .A(n4822), .Z(n4825) );
  XOR U5599 ( .A(n4826), .B(n4827), .Z(n4822) );
  ANDN U5600 ( .B(n4828), .A(n4829), .Z(n4826) );
  XNOR U5601 ( .A(b[1276]), .B(n4827), .Z(n4828) );
  XNOR U5602 ( .A(b[1276]), .B(n4829), .Z(c[1276]) );
  XNOR U5603 ( .A(a[1276]), .B(n4830), .Z(n4829) );
  IV U5604 ( .A(n4827), .Z(n4830) );
  XOR U5605 ( .A(n4831), .B(n4832), .Z(n4827) );
  ANDN U5606 ( .B(n4833), .A(n4834), .Z(n4831) );
  XNOR U5607 ( .A(b[1275]), .B(n4832), .Z(n4833) );
  XNOR U5608 ( .A(b[1275]), .B(n4834), .Z(c[1275]) );
  XNOR U5609 ( .A(a[1275]), .B(n4835), .Z(n4834) );
  IV U5610 ( .A(n4832), .Z(n4835) );
  XOR U5611 ( .A(n4836), .B(n4837), .Z(n4832) );
  ANDN U5612 ( .B(n4838), .A(n4839), .Z(n4836) );
  XNOR U5613 ( .A(b[1274]), .B(n4837), .Z(n4838) );
  XNOR U5614 ( .A(b[1274]), .B(n4839), .Z(c[1274]) );
  XNOR U5615 ( .A(a[1274]), .B(n4840), .Z(n4839) );
  IV U5616 ( .A(n4837), .Z(n4840) );
  XOR U5617 ( .A(n4841), .B(n4842), .Z(n4837) );
  ANDN U5618 ( .B(n4843), .A(n4844), .Z(n4841) );
  XNOR U5619 ( .A(b[1273]), .B(n4842), .Z(n4843) );
  XNOR U5620 ( .A(b[1273]), .B(n4844), .Z(c[1273]) );
  XNOR U5621 ( .A(a[1273]), .B(n4845), .Z(n4844) );
  IV U5622 ( .A(n4842), .Z(n4845) );
  XOR U5623 ( .A(n4846), .B(n4847), .Z(n4842) );
  ANDN U5624 ( .B(n4848), .A(n4849), .Z(n4846) );
  XNOR U5625 ( .A(b[1272]), .B(n4847), .Z(n4848) );
  XNOR U5626 ( .A(b[1272]), .B(n4849), .Z(c[1272]) );
  XNOR U5627 ( .A(a[1272]), .B(n4850), .Z(n4849) );
  IV U5628 ( .A(n4847), .Z(n4850) );
  XOR U5629 ( .A(n4851), .B(n4852), .Z(n4847) );
  ANDN U5630 ( .B(n4853), .A(n4854), .Z(n4851) );
  XNOR U5631 ( .A(b[1271]), .B(n4852), .Z(n4853) );
  XNOR U5632 ( .A(b[1271]), .B(n4854), .Z(c[1271]) );
  XNOR U5633 ( .A(a[1271]), .B(n4855), .Z(n4854) );
  IV U5634 ( .A(n4852), .Z(n4855) );
  XOR U5635 ( .A(n4856), .B(n4857), .Z(n4852) );
  ANDN U5636 ( .B(n4858), .A(n4859), .Z(n4856) );
  XNOR U5637 ( .A(b[1270]), .B(n4857), .Z(n4858) );
  XNOR U5638 ( .A(b[1270]), .B(n4859), .Z(c[1270]) );
  XNOR U5639 ( .A(a[1270]), .B(n4860), .Z(n4859) );
  IV U5640 ( .A(n4857), .Z(n4860) );
  XOR U5641 ( .A(n4861), .B(n4862), .Z(n4857) );
  ANDN U5642 ( .B(n4863), .A(n4864), .Z(n4861) );
  XNOR U5643 ( .A(b[1269]), .B(n4862), .Z(n4863) );
  XNOR U5644 ( .A(b[126]), .B(n4865), .Z(c[126]) );
  XNOR U5645 ( .A(b[1269]), .B(n4864), .Z(c[1269]) );
  XNOR U5646 ( .A(a[1269]), .B(n4866), .Z(n4864) );
  IV U5647 ( .A(n4862), .Z(n4866) );
  XOR U5648 ( .A(n4867), .B(n4868), .Z(n4862) );
  ANDN U5649 ( .B(n4869), .A(n4870), .Z(n4867) );
  XNOR U5650 ( .A(b[1268]), .B(n4868), .Z(n4869) );
  XNOR U5651 ( .A(b[1268]), .B(n4870), .Z(c[1268]) );
  XNOR U5652 ( .A(a[1268]), .B(n4871), .Z(n4870) );
  IV U5653 ( .A(n4868), .Z(n4871) );
  XOR U5654 ( .A(n4872), .B(n4873), .Z(n4868) );
  ANDN U5655 ( .B(n4874), .A(n4875), .Z(n4872) );
  XNOR U5656 ( .A(b[1267]), .B(n4873), .Z(n4874) );
  XNOR U5657 ( .A(b[1267]), .B(n4875), .Z(c[1267]) );
  XNOR U5658 ( .A(a[1267]), .B(n4876), .Z(n4875) );
  IV U5659 ( .A(n4873), .Z(n4876) );
  XOR U5660 ( .A(n4877), .B(n4878), .Z(n4873) );
  ANDN U5661 ( .B(n4879), .A(n4880), .Z(n4877) );
  XNOR U5662 ( .A(b[1266]), .B(n4878), .Z(n4879) );
  XNOR U5663 ( .A(b[1266]), .B(n4880), .Z(c[1266]) );
  XNOR U5664 ( .A(a[1266]), .B(n4881), .Z(n4880) );
  IV U5665 ( .A(n4878), .Z(n4881) );
  XOR U5666 ( .A(n4882), .B(n4883), .Z(n4878) );
  ANDN U5667 ( .B(n4884), .A(n4885), .Z(n4882) );
  XNOR U5668 ( .A(b[1265]), .B(n4883), .Z(n4884) );
  XNOR U5669 ( .A(b[1265]), .B(n4885), .Z(c[1265]) );
  XNOR U5670 ( .A(a[1265]), .B(n4886), .Z(n4885) );
  IV U5671 ( .A(n4883), .Z(n4886) );
  XOR U5672 ( .A(n4887), .B(n4888), .Z(n4883) );
  ANDN U5673 ( .B(n4889), .A(n4890), .Z(n4887) );
  XNOR U5674 ( .A(b[1264]), .B(n4888), .Z(n4889) );
  XNOR U5675 ( .A(b[1264]), .B(n4890), .Z(c[1264]) );
  XNOR U5676 ( .A(a[1264]), .B(n4891), .Z(n4890) );
  IV U5677 ( .A(n4888), .Z(n4891) );
  XOR U5678 ( .A(n4892), .B(n4893), .Z(n4888) );
  ANDN U5679 ( .B(n4894), .A(n4895), .Z(n4892) );
  XNOR U5680 ( .A(b[1263]), .B(n4893), .Z(n4894) );
  XNOR U5681 ( .A(b[1263]), .B(n4895), .Z(c[1263]) );
  XNOR U5682 ( .A(a[1263]), .B(n4896), .Z(n4895) );
  IV U5683 ( .A(n4893), .Z(n4896) );
  XOR U5684 ( .A(n4897), .B(n4898), .Z(n4893) );
  ANDN U5685 ( .B(n4899), .A(n4900), .Z(n4897) );
  XNOR U5686 ( .A(b[1262]), .B(n4898), .Z(n4899) );
  XNOR U5687 ( .A(b[1262]), .B(n4900), .Z(c[1262]) );
  XNOR U5688 ( .A(a[1262]), .B(n4901), .Z(n4900) );
  IV U5689 ( .A(n4898), .Z(n4901) );
  XOR U5690 ( .A(n4902), .B(n4903), .Z(n4898) );
  ANDN U5691 ( .B(n4904), .A(n4905), .Z(n4902) );
  XNOR U5692 ( .A(b[1261]), .B(n4903), .Z(n4904) );
  XNOR U5693 ( .A(b[1261]), .B(n4905), .Z(c[1261]) );
  XNOR U5694 ( .A(a[1261]), .B(n4906), .Z(n4905) );
  IV U5695 ( .A(n4903), .Z(n4906) );
  XOR U5696 ( .A(n4907), .B(n4908), .Z(n4903) );
  ANDN U5697 ( .B(n4909), .A(n4910), .Z(n4907) );
  XNOR U5698 ( .A(b[1260]), .B(n4908), .Z(n4909) );
  XNOR U5699 ( .A(b[1260]), .B(n4910), .Z(c[1260]) );
  XNOR U5700 ( .A(a[1260]), .B(n4911), .Z(n4910) );
  IV U5701 ( .A(n4908), .Z(n4911) );
  XOR U5702 ( .A(n4912), .B(n4913), .Z(n4908) );
  ANDN U5703 ( .B(n4914), .A(n4915), .Z(n4912) );
  XNOR U5704 ( .A(b[1259]), .B(n4913), .Z(n4914) );
  XNOR U5705 ( .A(b[125]), .B(n4916), .Z(c[125]) );
  XNOR U5706 ( .A(b[1259]), .B(n4915), .Z(c[1259]) );
  XNOR U5707 ( .A(a[1259]), .B(n4917), .Z(n4915) );
  IV U5708 ( .A(n4913), .Z(n4917) );
  XOR U5709 ( .A(n4918), .B(n4919), .Z(n4913) );
  ANDN U5710 ( .B(n4920), .A(n4921), .Z(n4918) );
  XNOR U5711 ( .A(b[1258]), .B(n4919), .Z(n4920) );
  XNOR U5712 ( .A(b[1258]), .B(n4921), .Z(c[1258]) );
  XNOR U5713 ( .A(a[1258]), .B(n4922), .Z(n4921) );
  IV U5714 ( .A(n4919), .Z(n4922) );
  XOR U5715 ( .A(n4923), .B(n4924), .Z(n4919) );
  ANDN U5716 ( .B(n4925), .A(n4926), .Z(n4923) );
  XNOR U5717 ( .A(b[1257]), .B(n4924), .Z(n4925) );
  XNOR U5718 ( .A(b[1257]), .B(n4926), .Z(c[1257]) );
  XNOR U5719 ( .A(a[1257]), .B(n4927), .Z(n4926) );
  IV U5720 ( .A(n4924), .Z(n4927) );
  XOR U5721 ( .A(n4928), .B(n4929), .Z(n4924) );
  ANDN U5722 ( .B(n4930), .A(n4931), .Z(n4928) );
  XNOR U5723 ( .A(b[1256]), .B(n4929), .Z(n4930) );
  XNOR U5724 ( .A(b[1256]), .B(n4931), .Z(c[1256]) );
  XNOR U5725 ( .A(a[1256]), .B(n4932), .Z(n4931) );
  IV U5726 ( .A(n4929), .Z(n4932) );
  XOR U5727 ( .A(n4933), .B(n4934), .Z(n4929) );
  ANDN U5728 ( .B(n4935), .A(n4936), .Z(n4933) );
  XNOR U5729 ( .A(b[1255]), .B(n4934), .Z(n4935) );
  XNOR U5730 ( .A(b[1255]), .B(n4936), .Z(c[1255]) );
  XNOR U5731 ( .A(a[1255]), .B(n4937), .Z(n4936) );
  IV U5732 ( .A(n4934), .Z(n4937) );
  XOR U5733 ( .A(n4938), .B(n4939), .Z(n4934) );
  ANDN U5734 ( .B(n4940), .A(n4941), .Z(n4938) );
  XNOR U5735 ( .A(b[1254]), .B(n4939), .Z(n4940) );
  XNOR U5736 ( .A(b[1254]), .B(n4941), .Z(c[1254]) );
  XNOR U5737 ( .A(a[1254]), .B(n4942), .Z(n4941) );
  IV U5738 ( .A(n4939), .Z(n4942) );
  XOR U5739 ( .A(n4943), .B(n4944), .Z(n4939) );
  ANDN U5740 ( .B(n4945), .A(n4946), .Z(n4943) );
  XNOR U5741 ( .A(b[1253]), .B(n4944), .Z(n4945) );
  XNOR U5742 ( .A(b[1253]), .B(n4946), .Z(c[1253]) );
  XNOR U5743 ( .A(a[1253]), .B(n4947), .Z(n4946) );
  IV U5744 ( .A(n4944), .Z(n4947) );
  XOR U5745 ( .A(n4948), .B(n4949), .Z(n4944) );
  ANDN U5746 ( .B(n4950), .A(n4951), .Z(n4948) );
  XNOR U5747 ( .A(b[1252]), .B(n4949), .Z(n4950) );
  XNOR U5748 ( .A(b[1252]), .B(n4951), .Z(c[1252]) );
  XNOR U5749 ( .A(a[1252]), .B(n4952), .Z(n4951) );
  IV U5750 ( .A(n4949), .Z(n4952) );
  XOR U5751 ( .A(n4953), .B(n4954), .Z(n4949) );
  ANDN U5752 ( .B(n4955), .A(n4956), .Z(n4953) );
  XNOR U5753 ( .A(b[1251]), .B(n4954), .Z(n4955) );
  XNOR U5754 ( .A(b[1251]), .B(n4956), .Z(c[1251]) );
  XNOR U5755 ( .A(a[1251]), .B(n4957), .Z(n4956) );
  IV U5756 ( .A(n4954), .Z(n4957) );
  XOR U5757 ( .A(n4958), .B(n4959), .Z(n4954) );
  ANDN U5758 ( .B(n4960), .A(n4961), .Z(n4958) );
  XNOR U5759 ( .A(b[1250]), .B(n4959), .Z(n4960) );
  XNOR U5760 ( .A(b[1250]), .B(n4961), .Z(c[1250]) );
  XNOR U5761 ( .A(a[1250]), .B(n4962), .Z(n4961) );
  IV U5762 ( .A(n4959), .Z(n4962) );
  XOR U5763 ( .A(n4963), .B(n4964), .Z(n4959) );
  ANDN U5764 ( .B(n4965), .A(n4966), .Z(n4963) );
  XNOR U5765 ( .A(b[1249]), .B(n4964), .Z(n4965) );
  XNOR U5766 ( .A(b[124]), .B(n4967), .Z(c[124]) );
  XNOR U5767 ( .A(b[1249]), .B(n4966), .Z(c[1249]) );
  XNOR U5768 ( .A(a[1249]), .B(n4968), .Z(n4966) );
  IV U5769 ( .A(n4964), .Z(n4968) );
  XOR U5770 ( .A(n4969), .B(n4970), .Z(n4964) );
  ANDN U5771 ( .B(n4971), .A(n4972), .Z(n4969) );
  XNOR U5772 ( .A(b[1248]), .B(n4970), .Z(n4971) );
  XNOR U5773 ( .A(b[1248]), .B(n4972), .Z(c[1248]) );
  XNOR U5774 ( .A(a[1248]), .B(n4973), .Z(n4972) );
  IV U5775 ( .A(n4970), .Z(n4973) );
  XOR U5776 ( .A(n4974), .B(n4975), .Z(n4970) );
  ANDN U5777 ( .B(n4976), .A(n4977), .Z(n4974) );
  XNOR U5778 ( .A(b[1247]), .B(n4975), .Z(n4976) );
  XNOR U5779 ( .A(b[1247]), .B(n4977), .Z(c[1247]) );
  XNOR U5780 ( .A(a[1247]), .B(n4978), .Z(n4977) );
  IV U5781 ( .A(n4975), .Z(n4978) );
  XOR U5782 ( .A(n4979), .B(n4980), .Z(n4975) );
  ANDN U5783 ( .B(n4981), .A(n4982), .Z(n4979) );
  XNOR U5784 ( .A(b[1246]), .B(n4980), .Z(n4981) );
  XNOR U5785 ( .A(b[1246]), .B(n4982), .Z(c[1246]) );
  XNOR U5786 ( .A(a[1246]), .B(n4983), .Z(n4982) );
  IV U5787 ( .A(n4980), .Z(n4983) );
  XOR U5788 ( .A(n4984), .B(n4985), .Z(n4980) );
  ANDN U5789 ( .B(n4986), .A(n4987), .Z(n4984) );
  XNOR U5790 ( .A(b[1245]), .B(n4985), .Z(n4986) );
  XNOR U5791 ( .A(b[1245]), .B(n4987), .Z(c[1245]) );
  XNOR U5792 ( .A(a[1245]), .B(n4988), .Z(n4987) );
  IV U5793 ( .A(n4985), .Z(n4988) );
  XOR U5794 ( .A(n4989), .B(n4990), .Z(n4985) );
  ANDN U5795 ( .B(n4991), .A(n4992), .Z(n4989) );
  XNOR U5796 ( .A(b[1244]), .B(n4990), .Z(n4991) );
  XNOR U5797 ( .A(b[1244]), .B(n4992), .Z(c[1244]) );
  XNOR U5798 ( .A(a[1244]), .B(n4993), .Z(n4992) );
  IV U5799 ( .A(n4990), .Z(n4993) );
  XOR U5800 ( .A(n4994), .B(n4995), .Z(n4990) );
  ANDN U5801 ( .B(n4996), .A(n4997), .Z(n4994) );
  XNOR U5802 ( .A(b[1243]), .B(n4995), .Z(n4996) );
  XNOR U5803 ( .A(b[1243]), .B(n4997), .Z(c[1243]) );
  XNOR U5804 ( .A(a[1243]), .B(n4998), .Z(n4997) );
  IV U5805 ( .A(n4995), .Z(n4998) );
  XOR U5806 ( .A(n4999), .B(n5000), .Z(n4995) );
  ANDN U5807 ( .B(n5001), .A(n5002), .Z(n4999) );
  XNOR U5808 ( .A(b[1242]), .B(n5000), .Z(n5001) );
  XNOR U5809 ( .A(b[1242]), .B(n5002), .Z(c[1242]) );
  XNOR U5810 ( .A(a[1242]), .B(n5003), .Z(n5002) );
  IV U5811 ( .A(n5000), .Z(n5003) );
  XOR U5812 ( .A(n5004), .B(n5005), .Z(n5000) );
  ANDN U5813 ( .B(n5006), .A(n5007), .Z(n5004) );
  XNOR U5814 ( .A(b[1241]), .B(n5005), .Z(n5006) );
  XNOR U5815 ( .A(b[1241]), .B(n5007), .Z(c[1241]) );
  XNOR U5816 ( .A(a[1241]), .B(n5008), .Z(n5007) );
  IV U5817 ( .A(n5005), .Z(n5008) );
  XOR U5818 ( .A(n5009), .B(n5010), .Z(n5005) );
  ANDN U5819 ( .B(n5011), .A(n5012), .Z(n5009) );
  XNOR U5820 ( .A(b[1240]), .B(n5010), .Z(n5011) );
  XNOR U5821 ( .A(b[1240]), .B(n5012), .Z(c[1240]) );
  XNOR U5822 ( .A(a[1240]), .B(n5013), .Z(n5012) );
  IV U5823 ( .A(n5010), .Z(n5013) );
  XOR U5824 ( .A(n5014), .B(n5015), .Z(n5010) );
  ANDN U5825 ( .B(n5016), .A(n5017), .Z(n5014) );
  XNOR U5826 ( .A(b[1239]), .B(n5015), .Z(n5016) );
  XNOR U5827 ( .A(b[123]), .B(n5018), .Z(c[123]) );
  XNOR U5828 ( .A(b[1239]), .B(n5017), .Z(c[1239]) );
  XNOR U5829 ( .A(a[1239]), .B(n5019), .Z(n5017) );
  IV U5830 ( .A(n5015), .Z(n5019) );
  XOR U5831 ( .A(n5020), .B(n5021), .Z(n5015) );
  ANDN U5832 ( .B(n5022), .A(n5023), .Z(n5020) );
  XNOR U5833 ( .A(b[1238]), .B(n5021), .Z(n5022) );
  XNOR U5834 ( .A(b[1238]), .B(n5023), .Z(c[1238]) );
  XNOR U5835 ( .A(a[1238]), .B(n5024), .Z(n5023) );
  IV U5836 ( .A(n5021), .Z(n5024) );
  XOR U5837 ( .A(n5025), .B(n5026), .Z(n5021) );
  ANDN U5838 ( .B(n5027), .A(n5028), .Z(n5025) );
  XNOR U5839 ( .A(b[1237]), .B(n5026), .Z(n5027) );
  XNOR U5840 ( .A(b[1237]), .B(n5028), .Z(c[1237]) );
  XNOR U5841 ( .A(a[1237]), .B(n5029), .Z(n5028) );
  IV U5842 ( .A(n5026), .Z(n5029) );
  XOR U5843 ( .A(n5030), .B(n5031), .Z(n5026) );
  ANDN U5844 ( .B(n5032), .A(n5033), .Z(n5030) );
  XNOR U5845 ( .A(b[1236]), .B(n5031), .Z(n5032) );
  XNOR U5846 ( .A(b[1236]), .B(n5033), .Z(c[1236]) );
  XNOR U5847 ( .A(a[1236]), .B(n5034), .Z(n5033) );
  IV U5848 ( .A(n5031), .Z(n5034) );
  XOR U5849 ( .A(n5035), .B(n5036), .Z(n5031) );
  ANDN U5850 ( .B(n5037), .A(n5038), .Z(n5035) );
  XNOR U5851 ( .A(b[1235]), .B(n5036), .Z(n5037) );
  XNOR U5852 ( .A(b[1235]), .B(n5038), .Z(c[1235]) );
  XNOR U5853 ( .A(a[1235]), .B(n5039), .Z(n5038) );
  IV U5854 ( .A(n5036), .Z(n5039) );
  XOR U5855 ( .A(n5040), .B(n5041), .Z(n5036) );
  ANDN U5856 ( .B(n5042), .A(n5043), .Z(n5040) );
  XNOR U5857 ( .A(b[1234]), .B(n5041), .Z(n5042) );
  XNOR U5858 ( .A(b[1234]), .B(n5043), .Z(c[1234]) );
  XNOR U5859 ( .A(a[1234]), .B(n5044), .Z(n5043) );
  IV U5860 ( .A(n5041), .Z(n5044) );
  XOR U5861 ( .A(n5045), .B(n5046), .Z(n5041) );
  ANDN U5862 ( .B(n5047), .A(n5048), .Z(n5045) );
  XNOR U5863 ( .A(b[1233]), .B(n5046), .Z(n5047) );
  XNOR U5864 ( .A(b[1233]), .B(n5048), .Z(c[1233]) );
  XNOR U5865 ( .A(a[1233]), .B(n5049), .Z(n5048) );
  IV U5866 ( .A(n5046), .Z(n5049) );
  XOR U5867 ( .A(n5050), .B(n5051), .Z(n5046) );
  ANDN U5868 ( .B(n5052), .A(n5053), .Z(n5050) );
  XNOR U5869 ( .A(b[1232]), .B(n5051), .Z(n5052) );
  XNOR U5870 ( .A(b[1232]), .B(n5053), .Z(c[1232]) );
  XNOR U5871 ( .A(a[1232]), .B(n5054), .Z(n5053) );
  IV U5872 ( .A(n5051), .Z(n5054) );
  XOR U5873 ( .A(n5055), .B(n5056), .Z(n5051) );
  ANDN U5874 ( .B(n5057), .A(n5058), .Z(n5055) );
  XNOR U5875 ( .A(b[1231]), .B(n5056), .Z(n5057) );
  XNOR U5876 ( .A(b[1231]), .B(n5058), .Z(c[1231]) );
  XNOR U5877 ( .A(a[1231]), .B(n5059), .Z(n5058) );
  IV U5878 ( .A(n5056), .Z(n5059) );
  XOR U5879 ( .A(n5060), .B(n5061), .Z(n5056) );
  ANDN U5880 ( .B(n5062), .A(n5063), .Z(n5060) );
  XNOR U5881 ( .A(b[1230]), .B(n5061), .Z(n5062) );
  XNOR U5882 ( .A(b[1230]), .B(n5063), .Z(c[1230]) );
  XNOR U5883 ( .A(a[1230]), .B(n5064), .Z(n5063) );
  IV U5884 ( .A(n5061), .Z(n5064) );
  XOR U5885 ( .A(n5065), .B(n5066), .Z(n5061) );
  ANDN U5886 ( .B(n5067), .A(n5068), .Z(n5065) );
  XNOR U5887 ( .A(b[1229]), .B(n5066), .Z(n5067) );
  XNOR U5888 ( .A(b[122]), .B(n5069), .Z(c[122]) );
  XNOR U5889 ( .A(b[1229]), .B(n5068), .Z(c[1229]) );
  XNOR U5890 ( .A(a[1229]), .B(n5070), .Z(n5068) );
  IV U5891 ( .A(n5066), .Z(n5070) );
  XOR U5892 ( .A(n5071), .B(n5072), .Z(n5066) );
  ANDN U5893 ( .B(n5073), .A(n5074), .Z(n5071) );
  XNOR U5894 ( .A(b[1228]), .B(n5072), .Z(n5073) );
  XNOR U5895 ( .A(b[1228]), .B(n5074), .Z(c[1228]) );
  XNOR U5896 ( .A(a[1228]), .B(n5075), .Z(n5074) );
  IV U5897 ( .A(n5072), .Z(n5075) );
  XOR U5898 ( .A(n5076), .B(n5077), .Z(n5072) );
  ANDN U5899 ( .B(n5078), .A(n5079), .Z(n5076) );
  XNOR U5900 ( .A(b[1227]), .B(n5077), .Z(n5078) );
  XNOR U5901 ( .A(b[1227]), .B(n5079), .Z(c[1227]) );
  XNOR U5902 ( .A(a[1227]), .B(n5080), .Z(n5079) );
  IV U5903 ( .A(n5077), .Z(n5080) );
  XOR U5904 ( .A(n5081), .B(n5082), .Z(n5077) );
  ANDN U5905 ( .B(n5083), .A(n5084), .Z(n5081) );
  XNOR U5906 ( .A(b[1226]), .B(n5082), .Z(n5083) );
  XNOR U5907 ( .A(b[1226]), .B(n5084), .Z(c[1226]) );
  XNOR U5908 ( .A(a[1226]), .B(n5085), .Z(n5084) );
  IV U5909 ( .A(n5082), .Z(n5085) );
  XOR U5910 ( .A(n5086), .B(n5087), .Z(n5082) );
  ANDN U5911 ( .B(n5088), .A(n5089), .Z(n5086) );
  XNOR U5912 ( .A(b[1225]), .B(n5087), .Z(n5088) );
  XNOR U5913 ( .A(b[1225]), .B(n5089), .Z(c[1225]) );
  XNOR U5914 ( .A(a[1225]), .B(n5090), .Z(n5089) );
  IV U5915 ( .A(n5087), .Z(n5090) );
  XOR U5916 ( .A(n5091), .B(n5092), .Z(n5087) );
  ANDN U5917 ( .B(n5093), .A(n5094), .Z(n5091) );
  XNOR U5918 ( .A(b[1224]), .B(n5092), .Z(n5093) );
  XNOR U5919 ( .A(b[1224]), .B(n5094), .Z(c[1224]) );
  XNOR U5920 ( .A(a[1224]), .B(n5095), .Z(n5094) );
  IV U5921 ( .A(n5092), .Z(n5095) );
  XOR U5922 ( .A(n5096), .B(n5097), .Z(n5092) );
  ANDN U5923 ( .B(n5098), .A(n5099), .Z(n5096) );
  XNOR U5924 ( .A(b[1223]), .B(n5097), .Z(n5098) );
  XNOR U5925 ( .A(b[1223]), .B(n5099), .Z(c[1223]) );
  XNOR U5926 ( .A(a[1223]), .B(n5100), .Z(n5099) );
  IV U5927 ( .A(n5097), .Z(n5100) );
  XOR U5928 ( .A(n5101), .B(n5102), .Z(n5097) );
  ANDN U5929 ( .B(n5103), .A(n5104), .Z(n5101) );
  XNOR U5930 ( .A(b[1222]), .B(n5102), .Z(n5103) );
  XNOR U5931 ( .A(b[1222]), .B(n5104), .Z(c[1222]) );
  XNOR U5932 ( .A(a[1222]), .B(n5105), .Z(n5104) );
  IV U5933 ( .A(n5102), .Z(n5105) );
  XOR U5934 ( .A(n5106), .B(n5107), .Z(n5102) );
  ANDN U5935 ( .B(n5108), .A(n5109), .Z(n5106) );
  XNOR U5936 ( .A(b[1221]), .B(n5107), .Z(n5108) );
  XNOR U5937 ( .A(b[1221]), .B(n5109), .Z(c[1221]) );
  XNOR U5938 ( .A(a[1221]), .B(n5110), .Z(n5109) );
  IV U5939 ( .A(n5107), .Z(n5110) );
  XOR U5940 ( .A(n5111), .B(n5112), .Z(n5107) );
  ANDN U5941 ( .B(n5113), .A(n5114), .Z(n5111) );
  XNOR U5942 ( .A(b[1220]), .B(n5112), .Z(n5113) );
  XNOR U5943 ( .A(b[1220]), .B(n5114), .Z(c[1220]) );
  XNOR U5944 ( .A(a[1220]), .B(n5115), .Z(n5114) );
  IV U5945 ( .A(n5112), .Z(n5115) );
  XOR U5946 ( .A(n5116), .B(n5117), .Z(n5112) );
  ANDN U5947 ( .B(n5118), .A(n5119), .Z(n5116) );
  XNOR U5948 ( .A(b[1219]), .B(n5117), .Z(n5118) );
  XNOR U5949 ( .A(b[121]), .B(n5120), .Z(c[121]) );
  XNOR U5950 ( .A(b[1219]), .B(n5119), .Z(c[1219]) );
  XNOR U5951 ( .A(a[1219]), .B(n5121), .Z(n5119) );
  IV U5952 ( .A(n5117), .Z(n5121) );
  XOR U5953 ( .A(n5122), .B(n5123), .Z(n5117) );
  ANDN U5954 ( .B(n5124), .A(n5125), .Z(n5122) );
  XNOR U5955 ( .A(b[1218]), .B(n5123), .Z(n5124) );
  XNOR U5956 ( .A(b[1218]), .B(n5125), .Z(c[1218]) );
  XNOR U5957 ( .A(a[1218]), .B(n5126), .Z(n5125) );
  IV U5958 ( .A(n5123), .Z(n5126) );
  XOR U5959 ( .A(n5127), .B(n5128), .Z(n5123) );
  ANDN U5960 ( .B(n5129), .A(n5130), .Z(n5127) );
  XNOR U5961 ( .A(b[1217]), .B(n5128), .Z(n5129) );
  XNOR U5962 ( .A(b[1217]), .B(n5130), .Z(c[1217]) );
  XNOR U5963 ( .A(a[1217]), .B(n5131), .Z(n5130) );
  IV U5964 ( .A(n5128), .Z(n5131) );
  XOR U5965 ( .A(n5132), .B(n5133), .Z(n5128) );
  ANDN U5966 ( .B(n5134), .A(n5135), .Z(n5132) );
  XNOR U5967 ( .A(b[1216]), .B(n5133), .Z(n5134) );
  XNOR U5968 ( .A(b[1216]), .B(n5135), .Z(c[1216]) );
  XNOR U5969 ( .A(a[1216]), .B(n5136), .Z(n5135) );
  IV U5970 ( .A(n5133), .Z(n5136) );
  XOR U5971 ( .A(n5137), .B(n5138), .Z(n5133) );
  ANDN U5972 ( .B(n5139), .A(n5140), .Z(n5137) );
  XNOR U5973 ( .A(b[1215]), .B(n5138), .Z(n5139) );
  XNOR U5974 ( .A(b[1215]), .B(n5140), .Z(c[1215]) );
  XNOR U5975 ( .A(a[1215]), .B(n5141), .Z(n5140) );
  IV U5976 ( .A(n5138), .Z(n5141) );
  XOR U5977 ( .A(n5142), .B(n5143), .Z(n5138) );
  ANDN U5978 ( .B(n5144), .A(n5145), .Z(n5142) );
  XNOR U5979 ( .A(b[1214]), .B(n5143), .Z(n5144) );
  XNOR U5980 ( .A(b[1214]), .B(n5145), .Z(c[1214]) );
  XNOR U5981 ( .A(a[1214]), .B(n5146), .Z(n5145) );
  IV U5982 ( .A(n5143), .Z(n5146) );
  XOR U5983 ( .A(n5147), .B(n5148), .Z(n5143) );
  ANDN U5984 ( .B(n5149), .A(n5150), .Z(n5147) );
  XNOR U5985 ( .A(b[1213]), .B(n5148), .Z(n5149) );
  XNOR U5986 ( .A(b[1213]), .B(n5150), .Z(c[1213]) );
  XNOR U5987 ( .A(a[1213]), .B(n5151), .Z(n5150) );
  IV U5988 ( .A(n5148), .Z(n5151) );
  XOR U5989 ( .A(n5152), .B(n5153), .Z(n5148) );
  ANDN U5990 ( .B(n5154), .A(n5155), .Z(n5152) );
  XNOR U5991 ( .A(b[1212]), .B(n5153), .Z(n5154) );
  XNOR U5992 ( .A(b[1212]), .B(n5155), .Z(c[1212]) );
  XNOR U5993 ( .A(a[1212]), .B(n5156), .Z(n5155) );
  IV U5994 ( .A(n5153), .Z(n5156) );
  XOR U5995 ( .A(n5157), .B(n5158), .Z(n5153) );
  ANDN U5996 ( .B(n5159), .A(n5160), .Z(n5157) );
  XNOR U5997 ( .A(b[1211]), .B(n5158), .Z(n5159) );
  XNOR U5998 ( .A(b[1211]), .B(n5160), .Z(c[1211]) );
  XNOR U5999 ( .A(a[1211]), .B(n5161), .Z(n5160) );
  IV U6000 ( .A(n5158), .Z(n5161) );
  XOR U6001 ( .A(n5162), .B(n5163), .Z(n5158) );
  ANDN U6002 ( .B(n5164), .A(n5165), .Z(n5162) );
  XNOR U6003 ( .A(b[1210]), .B(n5163), .Z(n5164) );
  XNOR U6004 ( .A(b[1210]), .B(n5165), .Z(c[1210]) );
  XNOR U6005 ( .A(a[1210]), .B(n5166), .Z(n5165) );
  IV U6006 ( .A(n5163), .Z(n5166) );
  XOR U6007 ( .A(n5167), .B(n5168), .Z(n5163) );
  ANDN U6008 ( .B(n5169), .A(n5170), .Z(n5167) );
  XNOR U6009 ( .A(b[1209]), .B(n5168), .Z(n5169) );
  XNOR U6010 ( .A(b[120]), .B(n5171), .Z(c[120]) );
  XNOR U6011 ( .A(b[1209]), .B(n5170), .Z(c[1209]) );
  XNOR U6012 ( .A(a[1209]), .B(n5172), .Z(n5170) );
  IV U6013 ( .A(n5168), .Z(n5172) );
  XOR U6014 ( .A(n5173), .B(n5174), .Z(n5168) );
  ANDN U6015 ( .B(n5175), .A(n5176), .Z(n5173) );
  XNOR U6016 ( .A(b[1208]), .B(n5174), .Z(n5175) );
  XNOR U6017 ( .A(b[1208]), .B(n5176), .Z(c[1208]) );
  XNOR U6018 ( .A(a[1208]), .B(n5177), .Z(n5176) );
  IV U6019 ( .A(n5174), .Z(n5177) );
  XOR U6020 ( .A(n5178), .B(n5179), .Z(n5174) );
  ANDN U6021 ( .B(n5180), .A(n5181), .Z(n5178) );
  XNOR U6022 ( .A(b[1207]), .B(n5179), .Z(n5180) );
  XNOR U6023 ( .A(b[1207]), .B(n5181), .Z(c[1207]) );
  XNOR U6024 ( .A(a[1207]), .B(n5182), .Z(n5181) );
  IV U6025 ( .A(n5179), .Z(n5182) );
  XOR U6026 ( .A(n5183), .B(n5184), .Z(n5179) );
  ANDN U6027 ( .B(n5185), .A(n5186), .Z(n5183) );
  XNOR U6028 ( .A(b[1206]), .B(n5184), .Z(n5185) );
  XNOR U6029 ( .A(b[1206]), .B(n5186), .Z(c[1206]) );
  XNOR U6030 ( .A(a[1206]), .B(n5187), .Z(n5186) );
  IV U6031 ( .A(n5184), .Z(n5187) );
  XOR U6032 ( .A(n5188), .B(n5189), .Z(n5184) );
  ANDN U6033 ( .B(n5190), .A(n5191), .Z(n5188) );
  XNOR U6034 ( .A(b[1205]), .B(n5189), .Z(n5190) );
  XNOR U6035 ( .A(b[1205]), .B(n5191), .Z(c[1205]) );
  XNOR U6036 ( .A(a[1205]), .B(n5192), .Z(n5191) );
  IV U6037 ( .A(n5189), .Z(n5192) );
  XOR U6038 ( .A(n5193), .B(n5194), .Z(n5189) );
  ANDN U6039 ( .B(n5195), .A(n5196), .Z(n5193) );
  XNOR U6040 ( .A(b[1204]), .B(n5194), .Z(n5195) );
  XNOR U6041 ( .A(b[1204]), .B(n5196), .Z(c[1204]) );
  XNOR U6042 ( .A(a[1204]), .B(n5197), .Z(n5196) );
  IV U6043 ( .A(n5194), .Z(n5197) );
  XOR U6044 ( .A(n5198), .B(n5199), .Z(n5194) );
  ANDN U6045 ( .B(n5200), .A(n5201), .Z(n5198) );
  XNOR U6046 ( .A(b[1203]), .B(n5199), .Z(n5200) );
  XNOR U6047 ( .A(b[1203]), .B(n5201), .Z(c[1203]) );
  XNOR U6048 ( .A(a[1203]), .B(n5202), .Z(n5201) );
  IV U6049 ( .A(n5199), .Z(n5202) );
  XOR U6050 ( .A(n5203), .B(n5204), .Z(n5199) );
  ANDN U6051 ( .B(n5205), .A(n5206), .Z(n5203) );
  XNOR U6052 ( .A(b[1202]), .B(n5204), .Z(n5205) );
  XNOR U6053 ( .A(b[1202]), .B(n5206), .Z(c[1202]) );
  XNOR U6054 ( .A(a[1202]), .B(n5207), .Z(n5206) );
  IV U6055 ( .A(n5204), .Z(n5207) );
  XOR U6056 ( .A(n5208), .B(n5209), .Z(n5204) );
  ANDN U6057 ( .B(n5210), .A(n5211), .Z(n5208) );
  XNOR U6058 ( .A(b[1201]), .B(n5209), .Z(n5210) );
  XNOR U6059 ( .A(b[1201]), .B(n5211), .Z(c[1201]) );
  XNOR U6060 ( .A(a[1201]), .B(n5212), .Z(n5211) );
  IV U6061 ( .A(n5209), .Z(n5212) );
  XOR U6062 ( .A(n5213), .B(n5214), .Z(n5209) );
  ANDN U6063 ( .B(n5215), .A(n5216), .Z(n5213) );
  XNOR U6064 ( .A(b[1200]), .B(n5214), .Z(n5215) );
  XNOR U6065 ( .A(b[1200]), .B(n5216), .Z(c[1200]) );
  XNOR U6066 ( .A(a[1200]), .B(n5217), .Z(n5216) );
  IV U6067 ( .A(n5214), .Z(n5217) );
  XOR U6068 ( .A(n5218), .B(n5219), .Z(n5214) );
  ANDN U6069 ( .B(n5220), .A(n5221), .Z(n5218) );
  XNOR U6070 ( .A(b[1199]), .B(n5219), .Z(n5220) );
  XNOR U6071 ( .A(b[11]), .B(n5222), .Z(c[11]) );
  XNOR U6072 ( .A(b[119]), .B(n5223), .Z(c[119]) );
  XNOR U6073 ( .A(b[1199]), .B(n5221), .Z(c[1199]) );
  XNOR U6074 ( .A(a[1199]), .B(n5224), .Z(n5221) );
  IV U6075 ( .A(n5219), .Z(n5224) );
  XOR U6076 ( .A(n5225), .B(n5226), .Z(n5219) );
  ANDN U6077 ( .B(n5227), .A(n5228), .Z(n5225) );
  XNOR U6078 ( .A(b[1198]), .B(n5226), .Z(n5227) );
  XNOR U6079 ( .A(b[1198]), .B(n5228), .Z(c[1198]) );
  XNOR U6080 ( .A(a[1198]), .B(n5229), .Z(n5228) );
  IV U6081 ( .A(n5226), .Z(n5229) );
  XOR U6082 ( .A(n5230), .B(n5231), .Z(n5226) );
  ANDN U6083 ( .B(n5232), .A(n5233), .Z(n5230) );
  XNOR U6084 ( .A(b[1197]), .B(n5231), .Z(n5232) );
  XNOR U6085 ( .A(b[1197]), .B(n5233), .Z(c[1197]) );
  XNOR U6086 ( .A(a[1197]), .B(n5234), .Z(n5233) );
  IV U6087 ( .A(n5231), .Z(n5234) );
  XOR U6088 ( .A(n5235), .B(n5236), .Z(n5231) );
  ANDN U6089 ( .B(n5237), .A(n5238), .Z(n5235) );
  XNOR U6090 ( .A(b[1196]), .B(n5236), .Z(n5237) );
  XNOR U6091 ( .A(b[1196]), .B(n5238), .Z(c[1196]) );
  XNOR U6092 ( .A(a[1196]), .B(n5239), .Z(n5238) );
  IV U6093 ( .A(n5236), .Z(n5239) );
  XOR U6094 ( .A(n5240), .B(n5241), .Z(n5236) );
  ANDN U6095 ( .B(n5242), .A(n5243), .Z(n5240) );
  XNOR U6096 ( .A(b[1195]), .B(n5241), .Z(n5242) );
  XNOR U6097 ( .A(b[1195]), .B(n5243), .Z(c[1195]) );
  XNOR U6098 ( .A(a[1195]), .B(n5244), .Z(n5243) );
  IV U6099 ( .A(n5241), .Z(n5244) );
  XOR U6100 ( .A(n5245), .B(n5246), .Z(n5241) );
  ANDN U6101 ( .B(n5247), .A(n5248), .Z(n5245) );
  XNOR U6102 ( .A(b[1194]), .B(n5246), .Z(n5247) );
  XNOR U6103 ( .A(b[1194]), .B(n5248), .Z(c[1194]) );
  XNOR U6104 ( .A(a[1194]), .B(n5249), .Z(n5248) );
  IV U6105 ( .A(n5246), .Z(n5249) );
  XOR U6106 ( .A(n5250), .B(n5251), .Z(n5246) );
  ANDN U6107 ( .B(n5252), .A(n5253), .Z(n5250) );
  XNOR U6108 ( .A(b[1193]), .B(n5251), .Z(n5252) );
  XNOR U6109 ( .A(b[1193]), .B(n5253), .Z(c[1193]) );
  XNOR U6110 ( .A(a[1193]), .B(n5254), .Z(n5253) );
  IV U6111 ( .A(n5251), .Z(n5254) );
  XOR U6112 ( .A(n5255), .B(n5256), .Z(n5251) );
  ANDN U6113 ( .B(n5257), .A(n5258), .Z(n5255) );
  XNOR U6114 ( .A(b[1192]), .B(n5256), .Z(n5257) );
  XNOR U6115 ( .A(b[1192]), .B(n5258), .Z(c[1192]) );
  XNOR U6116 ( .A(a[1192]), .B(n5259), .Z(n5258) );
  IV U6117 ( .A(n5256), .Z(n5259) );
  XOR U6118 ( .A(n5260), .B(n5261), .Z(n5256) );
  ANDN U6119 ( .B(n5262), .A(n5263), .Z(n5260) );
  XNOR U6120 ( .A(b[1191]), .B(n5261), .Z(n5262) );
  XNOR U6121 ( .A(b[1191]), .B(n5263), .Z(c[1191]) );
  XNOR U6122 ( .A(a[1191]), .B(n5264), .Z(n5263) );
  IV U6123 ( .A(n5261), .Z(n5264) );
  XOR U6124 ( .A(n5265), .B(n5266), .Z(n5261) );
  ANDN U6125 ( .B(n5267), .A(n5268), .Z(n5265) );
  XNOR U6126 ( .A(b[1190]), .B(n5266), .Z(n5267) );
  XNOR U6127 ( .A(b[1190]), .B(n5268), .Z(c[1190]) );
  XNOR U6128 ( .A(a[1190]), .B(n5269), .Z(n5268) );
  IV U6129 ( .A(n5266), .Z(n5269) );
  XOR U6130 ( .A(n5270), .B(n5271), .Z(n5266) );
  ANDN U6131 ( .B(n5272), .A(n5273), .Z(n5270) );
  XNOR U6132 ( .A(b[1189]), .B(n5271), .Z(n5272) );
  XNOR U6133 ( .A(b[118]), .B(n5274), .Z(c[118]) );
  XNOR U6134 ( .A(b[1189]), .B(n5273), .Z(c[1189]) );
  XNOR U6135 ( .A(a[1189]), .B(n5275), .Z(n5273) );
  IV U6136 ( .A(n5271), .Z(n5275) );
  XOR U6137 ( .A(n5276), .B(n5277), .Z(n5271) );
  ANDN U6138 ( .B(n5278), .A(n5279), .Z(n5276) );
  XNOR U6139 ( .A(b[1188]), .B(n5277), .Z(n5278) );
  XNOR U6140 ( .A(b[1188]), .B(n5279), .Z(c[1188]) );
  XNOR U6141 ( .A(a[1188]), .B(n5280), .Z(n5279) );
  IV U6142 ( .A(n5277), .Z(n5280) );
  XOR U6143 ( .A(n5281), .B(n5282), .Z(n5277) );
  ANDN U6144 ( .B(n5283), .A(n5284), .Z(n5281) );
  XNOR U6145 ( .A(b[1187]), .B(n5282), .Z(n5283) );
  XNOR U6146 ( .A(b[1187]), .B(n5284), .Z(c[1187]) );
  XNOR U6147 ( .A(a[1187]), .B(n5285), .Z(n5284) );
  IV U6148 ( .A(n5282), .Z(n5285) );
  XOR U6149 ( .A(n5286), .B(n5287), .Z(n5282) );
  ANDN U6150 ( .B(n5288), .A(n5289), .Z(n5286) );
  XNOR U6151 ( .A(b[1186]), .B(n5287), .Z(n5288) );
  XNOR U6152 ( .A(b[1186]), .B(n5289), .Z(c[1186]) );
  XNOR U6153 ( .A(a[1186]), .B(n5290), .Z(n5289) );
  IV U6154 ( .A(n5287), .Z(n5290) );
  XOR U6155 ( .A(n5291), .B(n5292), .Z(n5287) );
  ANDN U6156 ( .B(n5293), .A(n5294), .Z(n5291) );
  XNOR U6157 ( .A(b[1185]), .B(n5292), .Z(n5293) );
  XNOR U6158 ( .A(b[1185]), .B(n5294), .Z(c[1185]) );
  XNOR U6159 ( .A(a[1185]), .B(n5295), .Z(n5294) );
  IV U6160 ( .A(n5292), .Z(n5295) );
  XOR U6161 ( .A(n5296), .B(n5297), .Z(n5292) );
  ANDN U6162 ( .B(n5298), .A(n5299), .Z(n5296) );
  XNOR U6163 ( .A(b[1184]), .B(n5297), .Z(n5298) );
  XNOR U6164 ( .A(b[1184]), .B(n5299), .Z(c[1184]) );
  XNOR U6165 ( .A(a[1184]), .B(n5300), .Z(n5299) );
  IV U6166 ( .A(n5297), .Z(n5300) );
  XOR U6167 ( .A(n5301), .B(n5302), .Z(n5297) );
  ANDN U6168 ( .B(n5303), .A(n5304), .Z(n5301) );
  XNOR U6169 ( .A(b[1183]), .B(n5302), .Z(n5303) );
  XNOR U6170 ( .A(b[1183]), .B(n5304), .Z(c[1183]) );
  XNOR U6171 ( .A(a[1183]), .B(n5305), .Z(n5304) );
  IV U6172 ( .A(n5302), .Z(n5305) );
  XOR U6173 ( .A(n5306), .B(n5307), .Z(n5302) );
  ANDN U6174 ( .B(n5308), .A(n5309), .Z(n5306) );
  XNOR U6175 ( .A(b[1182]), .B(n5307), .Z(n5308) );
  XNOR U6176 ( .A(b[1182]), .B(n5309), .Z(c[1182]) );
  XNOR U6177 ( .A(a[1182]), .B(n5310), .Z(n5309) );
  IV U6178 ( .A(n5307), .Z(n5310) );
  XOR U6179 ( .A(n5311), .B(n5312), .Z(n5307) );
  ANDN U6180 ( .B(n5313), .A(n5314), .Z(n5311) );
  XNOR U6181 ( .A(b[1181]), .B(n5312), .Z(n5313) );
  XNOR U6182 ( .A(b[1181]), .B(n5314), .Z(c[1181]) );
  XNOR U6183 ( .A(a[1181]), .B(n5315), .Z(n5314) );
  IV U6184 ( .A(n5312), .Z(n5315) );
  XOR U6185 ( .A(n5316), .B(n5317), .Z(n5312) );
  ANDN U6186 ( .B(n5318), .A(n5319), .Z(n5316) );
  XNOR U6187 ( .A(b[1180]), .B(n5317), .Z(n5318) );
  XNOR U6188 ( .A(b[1180]), .B(n5319), .Z(c[1180]) );
  XNOR U6189 ( .A(a[1180]), .B(n5320), .Z(n5319) );
  IV U6190 ( .A(n5317), .Z(n5320) );
  XOR U6191 ( .A(n5321), .B(n5322), .Z(n5317) );
  ANDN U6192 ( .B(n5323), .A(n5324), .Z(n5321) );
  XNOR U6193 ( .A(b[1179]), .B(n5322), .Z(n5323) );
  XNOR U6194 ( .A(b[117]), .B(n5325), .Z(c[117]) );
  XNOR U6195 ( .A(b[1179]), .B(n5324), .Z(c[1179]) );
  XNOR U6196 ( .A(a[1179]), .B(n5326), .Z(n5324) );
  IV U6197 ( .A(n5322), .Z(n5326) );
  XOR U6198 ( .A(n5327), .B(n5328), .Z(n5322) );
  ANDN U6199 ( .B(n5329), .A(n5330), .Z(n5327) );
  XNOR U6200 ( .A(b[1178]), .B(n5328), .Z(n5329) );
  XNOR U6201 ( .A(b[1178]), .B(n5330), .Z(c[1178]) );
  XNOR U6202 ( .A(a[1178]), .B(n5331), .Z(n5330) );
  IV U6203 ( .A(n5328), .Z(n5331) );
  XOR U6204 ( .A(n5332), .B(n5333), .Z(n5328) );
  ANDN U6205 ( .B(n5334), .A(n5335), .Z(n5332) );
  XNOR U6206 ( .A(b[1177]), .B(n5333), .Z(n5334) );
  XNOR U6207 ( .A(b[1177]), .B(n5335), .Z(c[1177]) );
  XNOR U6208 ( .A(a[1177]), .B(n5336), .Z(n5335) );
  IV U6209 ( .A(n5333), .Z(n5336) );
  XOR U6210 ( .A(n5337), .B(n5338), .Z(n5333) );
  ANDN U6211 ( .B(n5339), .A(n5340), .Z(n5337) );
  XNOR U6212 ( .A(b[1176]), .B(n5338), .Z(n5339) );
  XNOR U6213 ( .A(b[1176]), .B(n5340), .Z(c[1176]) );
  XNOR U6214 ( .A(a[1176]), .B(n5341), .Z(n5340) );
  IV U6215 ( .A(n5338), .Z(n5341) );
  XOR U6216 ( .A(n5342), .B(n5343), .Z(n5338) );
  ANDN U6217 ( .B(n5344), .A(n5345), .Z(n5342) );
  XNOR U6218 ( .A(b[1175]), .B(n5343), .Z(n5344) );
  XNOR U6219 ( .A(b[1175]), .B(n5345), .Z(c[1175]) );
  XNOR U6220 ( .A(a[1175]), .B(n5346), .Z(n5345) );
  IV U6221 ( .A(n5343), .Z(n5346) );
  XOR U6222 ( .A(n5347), .B(n5348), .Z(n5343) );
  ANDN U6223 ( .B(n5349), .A(n5350), .Z(n5347) );
  XNOR U6224 ( .A(b[1174]), .B(n5348), .Z(n5349) );
  XNOR U6225 ( .A(b[1174]), .B(n5350), .Z(c[1174]) );
  XNOR U6226 ( .A(a[1174]), .B(n5351), .Z(n5350) );
  IV U6227 ( .A(n5348), .Z(n5351) );
  XOR U6228 ( .A(n5352), .B(n5353), .Z(n5348) );
  ANDN U6229 ( .B(n5354), .A(n5355), .Z(n5352) );
  XNOR U6230 ( .A(b[1173]), .B(n5353), .Z(n5354) );
  XNOR U6231 ( .A(b[1173]), .B(n5355), .Z(c[1173]) );
  XNOR U6232 ( .A(a[1173]), .B(n5356), .Z(n5355) );
  IV U6233 ( .A(n5353), .Z(n5356) );
  XOR U6234 ( .A(n5357), .B(n5358), .Z(n5353) );
  ANDN U6235 ( .B(n5359), .A(n5360), .Z(n5357) );
  XNOR U6236 ( .A(b[1172]), .B(n5358), .Z(n5359) );
  XNOR U6237 ( .A(b[1172]), .B(n5360), .Z(c[1172]) );
  XNOR U6238 ( .A(a[1172]), .B(n5361), .Z(n5360) );
  IV U6239 ( .A(n5358), .Z(n5361) );
  XOR U6240 ( .A(n5362), .B(n5363), .Z(n5358) );
  ANDN U6241 ( .B(n5364), .A(n5365), .Z(n5362) );
  XNOR U6242 ( .A(b[1171]), .B(n5363), .Z(n5364) );
  XNOR U6243 ( .A(b[1171]), .B(n5365), .Z(c[1171]) );
  XNOR U6244 ( .A(a[1171]), .B(n5366), .Z(n5365) );
  IV U6245 ( .A(n5363), .Z(n5366) );
  XOR U6246 ( .A(n5367), .B(n5368), .Z(n5363) );
  ANDN U6247 ( .B(n5369), .A(n5370), .Z(n5367) );
  XNOR U6248 ( .A(b[1170]), .B(n5368), .Z(n5369) );
  XNOR U6249 ( .A(b[1170]), .B(n5370), .Z(c[1170]) );
  XNOR U6250 ( .A(a[1170]), .B(n5371), .Z(n5370) );
  IV U6251 ( .A(n5368), .Z(n5371) );
  XOR U6252 ( .A(n5372), .B(n5373), .Z(n5368) );
  ANDN U6253 ( .B(n5374), .A(n5375), .Z(n5372) );
  XNOR U6254 ( .A(b[1169]), .B(n5373), .Z(n5374) );
  XNOR U6255 ( .A(b[116]), .B(n5376), .Z(c[116]) );
  XNOR U6256 ( .A(b[1169]), .B(n5375), .Z(c[1169]) );
  XNOR U6257 ( .A(a[1169]), .B(n5377), .Z(n5375) );
  IV U6258 ( .A(n5373), .Z(n5377) );
  XOR U6259 ( .A(n5378), .B(n5379), .Z(n5373) );
  ANDN U6260 ( .B(n5380), .A(n5381), .Z(n5378) );
  XNOR U6261 ( .A(b[1168]), .B(n5379), .Z(n5380) );
  XNOR U6262 ( .A(b[1168]), .B(n5381), .Z(c[1168]) );
  XNOR U6263 ( .A(a[1168]), .B(n5382), .Z(n5381) );
  IV U6264 ( .A(n5379), .Z(n5382) );
  XOR U6265 ( .A(n5383), .B(n5384), .Z(n5379) );
  ANDN U6266 ( .B(n5385), .A(n5386), .Z(n5383) );
  XNOR U6267 ( .A(b[1167]), .B(n5384), .Z(n5385) );
  XNOR U6268 ( .A(b[1167]), .B(n5386), .Z(c[1167]) );
  XNOR U6269 ( .A(a[1167]), .B(n5387), .Z(n5386) );
  IV U6270 ( .A(n5384), .Z(n5387) );
  XOR U6271 ( .A(n5388), .B(n5389), .Z(n5384) );
  ANDN U6272 ( .B(n5390), .A(n5391), .Z(n5388) );
  XNOR U6273 ( .A(b[1166]), .B(n5389), .Z(n5390) );
  XNOR U6274 ( .A(b[1166]), .B(n5391), .Z(c[1166]) );
  XNOR U6275 ( .A(a[1166]), .B(n5392), .Z(n5391) );
  IV U6276 ( .A(n5389), .Z(n5392) );
  XOR U6277 ( .A(n5393), .B(n5394), .Z(n5389) );
  ANDN U6278 ( .B(n5395), .A(n5396), .Z(n5393) );
  XNOR U6279 ( .A(b[1165]), .B(n5394), .Z(n5395) );
  XNOR U6280 ( .A(b[1165]), .B(n5396), .Z(c[1165]) );
  XNOR U6281 ( .A(a[1165]), .B(n5397), .Z(n5396) );
  IV U6282 ( .A(n5394), .Z(n5397) );
  XOR U6283 ( .A(n5398), .B(n5399), .Z(n5394) );
  ANDN U6284 ( .B(n5400), .A(n5401), .Z(n5398) );
  XNOR U6285 ( .A(b[1164]), .B(n5399), .Z(n5400) );
  XNOR U6286 ( .A(b[1164]), .B(n5401), .Z(c[1164]) );
  XNOR U6287 ( .A(a[1164]), .B(n5402), .Z(n5401) );
  IV U6288 ( .A(n5399), .Z(n5402) );
  XOR U6289 ( .A(n5403), .B(n5404), .Z(n5399) );
  ANDN U6290 ( .B(n5405), .A(n5406), .Z(n5403) );
  XNOR U6291 ( .A(b[1163]), .B(n5404), .Z(n5405) );
  XNOR U6292 ( .A(b[1163]), .B(n5406), .Z(c[1163]) );
  XNOR U6293 ( .A(a[1163]), .B(n5407), .Z(n5406) );
  IV U6294 ( .A(n5404), .Z(n5407) );
  XOR U6295 ( .A(n5408), .B(n5409), .Z(n5404) );
  ANDN U6296 ( .B(n5410), .A(n5411), .Z(n5408) );
  XNOR U6297 ( .A(b[1162]), .B(n5409), .Z(n5410) );
  XNOR U6298 ( .A(b[1162]), .B(n5411), .Z(c[1162]) );
  XNOR U6299 ( .A(a[1162]), .B(n5412), .Z(n5411) );
  IV U6300 ( .A(n5409), .Z(n5412) );
  XOR U6301 ( .A(n5413), .B(n5414), .Z(n5409) );
  ANDN U6302 ( .B(n5415), .A(n5416), .Z(n5413) );
  XNOR U6303 ( .A(b[1161]), .B(n5414), .Z(n5415) );
  XNOR U6304 ( .A(b[1161]), .B(n5416), .Z(c[1161]) );
  XNOR U6305 ( .A(a[1161]), .B(n5417), .Z(n5416) );
  IV U6306 ( .A(n5414), .Z(n5417) );
  XOR U6307 ( .A(n5418), .B(n5419), .Z(n5414) );
  ANDN U6308 ( .B(n5420), .A(n5421), .Z(n5418) );
  XNOR U6309 ( .A(b[1160]), .B(n5419), .Z(n5420) );
  XNOR U6310 ( .A(b[1160]), .B(n5421), .Z(c[1160]) );
  XNOR U6311 ( .A(a[1160]), .B(n5422), .Z(n5421) );
  IV U6312 ( .A(n5419), .Z(n5422) );
  XOR U6313 ( .A(n5423), .B(n5424), .Z(n5419) );
  ANDN U6314 ( .B(n5425), .A(n5426), .Z(n5423) );
  XNOR U6315 ( .A(b[1159]), .B(n5424), .Z(n5425) );
  XNOR U6316 ( .A(b[115]), .B(n5427), .Z(c[115]) );
  XNOR U6317 ( .A(b[1159]), .B(n5426), .Z(c[1159]) );
  XNOR U6318 ( .A(a[1159]), .B(n5428), .Z(n5426) );
  IV U6319 ( .A(n5424), .Z(n5428) );
  XOR U6320 ( .A(n5429), .B(n5430), .Z(n5424) );
  ANDN U6321 ( .B(n5431), .A(n5432), .Z(n5429) );
  XNOR U6322 ( .A(b[1158]), .B(n5430), .Z(n5431) );
  XNOR U6323 ( .A(b[1158]), .B(n5432), .Z(c[1158]) );
  XNOR U6324 ( .A(a[1158]), .B(n5433), .Z(n5432) );
  IV U6325 ( .A(n5430), .Z(n5433) );
  XOR U6326 ( .A(n5434), .B(n5435), .Z(n5430) );
  ANDN U6327 ( .B(n5436), .A(n5437), .Z(n5434) );
  XNOR U6328 ( .A(b[1157]), .B(n5435), .Z(n5436) );
  XNOR U6329 ( .A(b[1157]), .B(n5437), .Z(c[1157]) );
  XNOR U6330 ( .A(a[1157]), .B(n5438), .Z(n5437) );
  IV U6331 ( .A(n5435), .Z(n5438) );
  XOR U6332 ( .A(n5439), .B(n5440), .Z(n5435) );
  ANDN U6333 ( .B(n5441), .A(n5442), .Z(n5439) );
  XNOR U6334 ( .A(b[1156]), .B(n5440), .Z(n5441) );
  XNOR U6335 ( .A(b[1156]), .B(n5442), .Z(c[1156]) );
  XNOR U6336 ( .A(a[1156]), .B(n5443), .Z(n5442) );
  IV U6337 ( .A(n5440), .Z(n5443) );
  XOR U6338 ( .A(n5444), .B(n5445), .Z(n5440) );
  ANDN U6339 ( .B(n5446), .A(n5447), .Z(n5444) );
  XNOR U6340 ( .A(b[1155]), .B(n5445), .Z(n5446) );
  XNOR U6341 ( .A(b[1155]), .B(n5447), .Z(c[1155]) );
  XNOR U6342 ( .A(a[1155]), .B(n5448), .Z(n5447) );
  IV U6343 ( .A(n5445), .Z(n5448) );
  XOR U6344 ( .A(n5449), .B(n5450), .Z(n5445) );
  ANDN U6345 ( .B(n5451), .A(n5452), .Z(n5449) );
  XNOR U6346 ( .A(b[1154]), .B(n5450), .Z(n5451) );
  XNOR U6347 ( .A(b[1154]), .B(n5452), .Z(c[1154]) );
  XNOR U6348 ( .A(a[1154]), .B(n5453), .Z(n5452) );
  IV U6349 ( .A(n5450), .Z(n5453) );
  XOR U6350 ( .A(n5454), .B(n5455), .Z(n5450) );
  ANDN U6351 ( .B(n5456), .A(n5457), .Z(n5454) );
  XNOR U6352 ( .A(b[1153]), .B(n5455), .Z(n5456) );
  XNOR U6353 ( .A(b[1153]), .B(n5457), .Z(c[1153]) );
  XNOR U6354 ( .A(a[1153]), .B(n5458), .Z(n5457) );
  IV U6355 ( .A(n5455), .Z(n5458) );
  XOR U6356 ( .A(n5459), .B(n5460), .Z(n5455) );
  ANDN U6357 ( .B(n5461), .A(n5462), .Z(n5459) );
  XNOR U6358 ( .A(b[1152]), .B(n5460), .Z(n5461) );
  XNOR U6359 ( .A(b[1152]), .B(n5462), .Z(c[1152]) );
  XNOR U6360 ( .A(a[1152]), .B(n5463), .Z(n5462) );
  IV U6361 ( .A(n5460), .Z(n5463) );
  XOR U6362 ( .A(n5464), .B(n5465), .Z(n5460) );
  ANDN U6363 ( .B(n5466), .A(n5467), .Z(n5464) );
  XNOR U6364 ( .A(b[1151]), .B(n5465), .Z(n5466) );
  XNOR U6365 ( .A(b[1151]), .B(n5467), .Z(c[1151]) );
  XNOR U6366 ( .A(a[1151]), .B(n5468), .Z(n5467) );
  IV U6367 ( .A(n5465), .Z(n5468) );
  XOR U6368 ( .A(n5469), .B(n5470), .Z(n5465) );
  ANDN U6369 ( .B(n5471), .A(n5472), .Z(n5469) );
  XNOR U6370 ( .A(b[1150]), .B(n5470), .Z(n5471) );
  XNOR U6371 ( .A(b[1150]), .B(n5472), .Z(c[1150]) );
  XNOR U6372 ( .A(a[1150]), .B(n5473), .Z(n5472) );
  IV U6373 ( .A(n5470), .Z(n5473) );
  XOR U6374 ( .A(n5474), .B(n5475), .Z(n5470) );
  ANDN U6375 ( .B(n5476), .A(n5477), .Z(n5474) );
  XNOR U6376 ( .A(b[1149]), .B(n5475), .Z(n5476) );
  XNOR U6377 ( .A(b[114]), .B(n5478), .Z(c[114]) );
  XNOR U6378 ( .A(b[1149]), .B(n5477), .Z(c[1149]) );
  XNOR U6379 ( .A(a[1149]), .B(n5479), .Z(n5477) );
  IV U6380 ( .A(n5475), .Z(n5479) );
  XOR U6381 ( .A(n5480), .B(n5481), .Z(n5475) );
  ANDN U6382 ( .B(n5482), .A(n5483), .Z(n5480) );
  XNOR U6383 ( .A(b[1148]), .B(n5481), .Z(n5482) );
  XNOR U6384 ( .A(b[1148]), .B(n5483), .Z(c[1148]) );
  XNOR U6385 ( .A(a[1148]), .B(n5484), .Z(n5483) );
  IV U6386 ( .A(n5481), .Z(n5484) );
  XOR U6387 ( .A(n5485), .B(n5486), .Z(n5481) );
  ANDN U6388 ( .B(n5487), .A(n5488), .Z(n5485) );
  XNOR U6389 ( .A(b[1147]), .B(n5486), .Z(n5487) );
  XNOR U6390 ( .A(b[1147]), .B(n5488), .Z(c[1147]) );
  XNOR U6391 ( .A(a[1147]), .B(n5489), .Z(n5488) );
  IV U6392 ( .A(n5486), .Z(n5489) );
  XOR U6393 ( .A(n5490), .B(n5491), .Z(n5486) );
  ANDN U6394 ( .B(n5492), .A(n5493), .Z(n5490) );
  XNOR U6395 ( .A(b[1146]), .B(n5491), .Z(n5492) );
  XNOR U6396 ( .A(b[1146]), .B(n5493), .Z(c[1146]) );
  XNOR U6397 ( .A(a[1146]), .B(n5494), .Z(n5493) );
  IV U6398 ( .A(n5491), .Z(n5494) );
  XOR U6399 ( .A(n5495), .B(n5496), .Z(n5491) );
  ANDN U6400 ( .B(n5497), .A(n5498), .Z(n5495) );
  XNOR U6401 ( .A(b[1145]), .B(n5496), .Z(n5497) );
  XNOR U6402 ( .A(b[1145]), .B(n5498), .Z(c[1145]) );
  XNOR U6403 ( .A(a[1145]), .B(n5499), .Z(n5498) );
  IV U6404 ( .A(n5496), .Z(n5499) );
  XOR U6405 ( .A(n5500), .B(n5501), .Z(n5496) );
  ANDN U6406 ( .B(n5502), .A(n5503), .Z(n5500) );
  XNOR U6407 ( .A(b[1144]), .B(n5501), .Z(n5502) );
  XNOR U6408 ( .A(b[1144]), .B(n5503), .Z(c[1144]) );
  XNOR U6409 ( .A(a[1144]), .B(n5504), .Z(n5503) );
  IV U6410 ( .A(n5501), .Z(n5504) );
  XOR U6411 ( .A(n5505), .B(n5506), .Z(n5501) );
  ANDN U6412 ( .B(n5507), .A(n5508), .Z(n5505) );
  XNOR U6413 ( .A(b[1143]), .B(n5506), .Z(n5507) );
  XNOR U6414 ( .A(b[1143]), .B(n5508), .Z(c[1143]) );
  XNOR U6415 ( .A(a[1143]), .B(n5509), .Z(n5508) );
  IV U6416 ( .A(n5506), .Z(n5509) );
  XOR U6417 ( .A(n5510), .B(n5511), .Z(n5506) );
  ANDN U6418 ( .B(n5512), .A(n5513), .Z(n5510) );
  XNOR U6419 ( .A(b[1142]), .B(n5511), .Z(n5512) );
  XNOR U6420 ( .A(b[1142]), .B(n5513), .Z(c[1142]) );
  XNOR U6421 ( .A(a[1142]), .B(n5514), .Z(n5513) );
  IV U6422 ( .A(n5511), .Z(n5514) );
  XOR U6423 ( .A(n5515), .B(n5516), .Z(n5511) );
  ANDN U6424 ( .B(n5517), .A(n5518), .Z(n5515) );
  XNOR U6425 ( .A(b[1141]), .B(n5516), .Z(n5517) );
  XNOR U6426 ( .A(b[1141]), .B(n5518), .Z(c[1141]) );
  XNOR U6427 ( .A(a[1141]), .B(n5519), .Z(n5518) );
  IV U6428 ( .A(n5516), .Z(n5519) );
  XOR U6429 ( .A(n5520), .B(n5521), .Z(n5516) );
  ANDN U6430 ( .B(n5522), .A(n5523), .Z(n5520) );
  XNOR U6431 ( .A(b[1140]), .B(n5521), .Z(n5522) );
  XNOR U6432 ( .A(b[1140]), .B(n5523), .Z(c[1140]) );
  XNOR U6433 ( .A(a[1140]), .B(n5524), .Z(n5523) );
  IV U6434 ( .A(n5521), .Z(n5524) );
  XOR U6435 ( .A(n5525), .B(n5526), .Z(n5521) );
  ANDN U6436 ( .B(n5527), .A(n5528), .Z(n5525) );
  XNOR U6437 ( .A(b[1139]), .B(n5526), .Z(n5527) );
  XNOR U6438 ( .A(b[113]), .B(n5529), .Z(c[113]) );
  XNOR U6439 ( .A(b[1139]), .B(n5528), .Z(c[1139]) );
  XNOR U6440 ( .A(a[1139]), .B(n5530), .Z(n5528) );
  IV U6441 ( .A(n5526), .Z(n5530) );
  XOR U6442 ( .A(n5531), .B(n5532), .Z(n5526) );
  ANDN U6443 ( .B(n5533), .A(n5534), .Z(n5531) );
  XNOR U6444 ( .A(b[1138]), .B(n5532), .Z(n5533) );
  XNOR U6445 ( .A(b[1138]), .B(n5534), .Z(c[1138]) );
  XNOR U6446 ( .A(a[1138]), .B(n5535), .Z(n5534) );
  IV U6447 ( .A(n5532), .Z(n5535) );
  XOR U6448 ( .A(n5536), .B(n5537), .Z(n5532) );
  ANDN U6449 ( .B(n5538), .A(n5539), .Z(n5536) );
  XNOR U6450 ( .A(b[1137]), .B(n5537), .Z(n5538) );
  XNOR U6451 ( .A(b[1137]), .B(n5539), .Z(c[1137]) );
  XNOR U6452 ( .A(a[1137]), .B(n5540), .Z(n5539) );
  IV U6453 ( .A(n5537), .Z(n5540) );
  XOR U6454 ( .A(n5541), .B(n5542), .Z(n5537) );
  ANDN U6455 ( .B(n5543), .A(n5544), .Z(n5541) );
  XNOR U6456 ( .A(b[1136]), .B(n5542), .Z(n5543) );
  XNOR U6457 ( .A(b[1136]), .B(n5544), .Z(c[1136]) );
  XNOR U6458 ( .A(a[1136]), .B(n5545), .Z(n5544) );
  IV U6459 ( .A(n5542), .Z(n5545) );
  XOR U6460 ( .A(n5546), .B(n5547), .Z(n5542) );
  ANDN U6461 ( .B(n5548), .A(n5549), .Z(n5546) );
  XNOR U6462 ( .A(b[1135]), .B(n5547), .Z(n5548) );
  XNOR U6463 ( .A(b[1135]), .B(n5549), .Z(c[1135]) );
  XNOR U6464 ( .A(a[1135]), .B(n5550), .Z(n5549) );
  IV U6465 ( .A(n5547), .Z(n5550) );
  XOR U6466 ( .A(n5551), .B(n5552), .Z(n5547) );
  ANDN U6467 ( .B(n5553), .A(n5554), .Z(n5551) );
  XNOR U6468 ( .A(b[1134]), .B(n5552), .Z(n5553) );
  XNOR U6469 ( .A(b[1134]), .B(n5554), .Z(c[1134]) );
  XNOR U6470 ( .A(a[1134]), .B(n5555), .Z(n5554) );
  IV U6471 ( .A(n5552), .Z(n5555) );
  XOR U6472 ( .A(n5556), .B(n5557), .Z(n5552) );
  ANDN U6473 ( .B(n5558), .A(n5559), .Z(n5556) );
  XNOR U6474 ( .A(b[1133]), .B(n5557), .Z(n5558) );
  XNOR U6475 ( .A(b[1133]), .B(n5559), .Z(c[1133]) );
  XNOR U6476 ( .A(a[1133]), .B(n5560), .Z(n5559) );
  IV U6477 ( .A(n5557), .Z(n5560) );
  XOR U6478 ( .A(n5561), .B(n5562), .Z(n5557) );
  ANDN U6479 ( .B(n5563), .A(n5564), .Z(n5561) );
  XNOR U6480 ( .A(b[1132]), .B(n5562), .Z(n5563) );
  XNOR U6481 ( .A(b[1132]), .B(n5564), .Z(c[1132]) );
  XNOR U6482 ( .A(a[1132]), .B(n5565), .Z(n5564) );
  IV U6483 ( .A(n5562), .Z(n5565) );
  XOR U6484 ( .A(n5566), .B(n5567), .Z(n5562) );
  ANDN U6485 ( .B(n5568), .A(n5569), .Z(n5566) );
  XNOR U6486 ( .A(b[1131]), .B(n5567), .Z(n5568) );
  XNOR U6487 ( .A(b[1131]), .B(n5569), .Z(c[1131]) );
  XNOR U6488 ( .A(a[1131]), .B(n5570), .Z(n5569) );
  IV U6489 ( .A(n5567), .Z(n5570) );
  XOR U6490 ( .A(n5571), .B(n5572), .Z(n5567) );
  ANDN U6491 ( .B(n5573), .A(n5574), .Z(n5571) );
  XNOR U6492 ( .A(b[1130]), .B(n5572), .Z(n5573) );
  XNOR U6493 ( .A(b[1130]), .B(n5574), .Z(c[1130]) );
  XNOR U6494 ( .A(a[1130]), .B(n5575), .Z(n5574) );
  IV U6495 ( .A(n5572), .Z(n5575) );
  XOR U6496 ( .A(n5576), .B(n5577), .Z(n5572) );
  ANDN U6497 ( .B(n5578), .A(n5579), .Z(n5576) );
  XNOR U6498 ( .A(b[1129]), .B(n5577), .Z(n5578) );
  XNOR U6499 ( .A(b[112]), .B(n5580), .Z(c[112]) );
  XNOR U6500 ( .A(b[1129]), .B(n5579), .Z(c[1129]) );
  XNOR U6501 ( .A(a[1129]), .B(n5581), .Z(n5579) );
  IV U6502 ( .A(n5577), .Z(n5581) );
  XOR U6503 ( .A(n5582), .B(n5583), .Z(n5577) );
  ANDN U6504 ( .B(n5584), .A(n5585), .Z(n5582) );
  XNOR U6505 ( .A(b[1128]), .B(n5583), .Z(n5584) );
  XNOR U6506 ( .A(b[1128]), .B(n5585), .Z(c[1128]) );
  XNOR U6507 ( .A(a[1128]), .B(n5586), .Z(n5585) );
  IV U6508 ( .A(n5583), .Z(n5586) );
  XOR U6509 ( .A(n5587), .B(n5588), .Z(n5583) );
  ANDN U6510 ( .B(n5589), .A(n5590), .Z(n5587) );
  XNOR U6511 ( .A(b[1127]), .B(n5588), .Z(n5589) );
  XNOR U6512 ( .A(b[1127]), .B(n5590), .Z(c[1127]) );
  XNOR U6513 ( .A(a[1127]), .B(n5591), .Z(n5590) );
  IV U6514 ( .A(n5588), .Z(n5591) );
  XOR U6515 ( .A(n5592), .B(n5593), .Z(n5588) );
  ANDN U6516 ( .B(n5594), .A(n5595), .Z(n5592) );
  XNOR U6517 ( .A(b[1126]), .B(n5593), .Z(n5594) );
  XNOR U6518 ( .A(b[1126]), .B(n5595), .Z(c[1126]) );
  XNOR U6519 ( .A(a[1126]), .B(n5596), .Z(n5595) );
  IV U6520 ( .A(n5593), .Z(n5596) );
  XOR U6521 ( .A(n5597), .B(n5598), .Z(n5593) );
  ANDN U6522 ( .B(n5599), .A(n5600), .Z(n5597) );
  XNOR U6523 ( .A(b[1125]), .B(n5598), .Z(n5599) );
  XNOR U6524 ( .A(b[1125]), .B(n5600), .Z(c[1125]) );
  XNOR U6525 ( .A(a[1125]), .B(n5601), .Z(n5600) );
  IV U6526 ( .A(n5598), .Z(n5601) );
  XOR U6527 ( .A(n5602), .B(n5603), .Z(n5598) );
  ANDN U6528 ( .B(n5604), .A(n5605), .Z(n5602) );
  XNOR U6529 ( .A(b[1124]), .B(n5603), .Z(n5604) );
  XNOR U6530 ( .A(b[1124]), .B(n5605), .Z(c[1124]) );
  XNOR U6531 ( .A(a[1124]), .B(n5606), .Z(n5605) );
  IV U6532 ( .A(n5603), .Z(n5606) );
  XOR U6533 ( .A(n5607), .B(n5608), .Z(n5603) );
  ANDN U6534 ( .B(n5609), .A(n5610), .Z(n5607) );
  XNOR U6535 ( .A(b[1123]), .B(n5608), .Z(n5609) );
  XNOR U6536 ( .A(b[1123]), .B(n5610), .Z(c[1123]) );
  XNOR U6537 ( .A(a[1123]), .B(n5611), .Z(n5610) );
  IV U6538 ( .A(n5608), .Z(n5611) );
  XOR U6539 ( .A(n5612), .B(n5613), .Z(n5608) );
  ANDN U6540 ( .B(n5614), .A(n5615), .Z(n5612) );
  XNOR U6541 ( .A(b[1122]), .B(n5613), .Z(n5614) );
  XNOR U6542 ( .A(b[1122]), .B(n5615), .Z(c[1122]) );
  XNOR U6543 ( .A(a[1122]), .B(n5616), .Z(n5615) );
  IV U6544 ( .A(n5613), .Z(n5616) );
  XOR U6545 ( .A(n5617), .B(n5618), .Z(n5613) );
  ANDN U6546 ( .B(n5619), .A(n5620), .Z(n5617) );
  XNOR U6547 ( .A(b[1121]), .B(n5618), .Z(n5619) );
  XNOR U6548 ( .A(b[1121]), .B(n5620), .Z(c[1121]) );
  XNOR U6549 ( .A(a[1121]), .B(n5621), .Z(n5620) );
  IV U6550 ( .A(n5618), .Z(n5621) );
  XOR U6551 ( .A(n5622), .B(n5623), .Z(n5618) );
  ANDN U6552 ( .B(n5624), .A(n5625), .Z(n5622) );
  XNOR U6553 ( .A(b[1120]), .B(n5623), .Z(n5624) );
  XNOR U6554 ( .A(b[1120]), .B(n5625), .Z(c[1120]) );
  XNOR U6555 ( .A(a[1120]), .B(n5626), .Z(n5625) );
  IV U6556 ( .A(n5623), .Z(n5626) );
  XOR U6557 ( .A(n5627), .B(n5628), .Z(n5623) );
  ANDN U6558 ( .B(n5629), .A(n5630), .Z(n5627) );
  XNOR U6559 ( .A(b[1119]), .B(n5628), .Z(n5629) );
  XNOR U6560 ( .A(b[111]), .B(n5631), .Z(c[111]) );
  XNOR U6561 ( .A(b[1119]), .B(n5630), .Z(c[1119]) );
  XNOR U6562 ( .A(a[1119]), .B(n5632), .Z(n5630) );
  IV U6563 ( .A(n5628), .Z(n5632) );
  XOR U6564 ( .A(n5633), .B(n5634), .Z(n5628) );
  ANDN U6565 ( .B(n5635), .A(n5636), .Z(n5633) );
  XNOR U6566 ( .A(b[1118]), .B(n5634), .Z(n5635) );
  XNOR U6567 ( .A(b[1118]), .B(n5636), .Z(c[1118]) );
  XNOR U6568 ( .A(a[1118]), .B(n5637), .Z(n5636) );
  IV U6569 ( .A(n5634), .Z(n5637) );
  XOR U6570 ( .A(n5638), .B(n5639), .Z(n5634) );
  ANDN U6571 ( .B(n5640), .A(n5641), .Z(n5638) );
  XNOR U6572 ( .A(b[1117]), .B(n5639), .Z(n5640) );
  XNOR U6573 ( .A(b[1117]), .B(n5641), .Z(c[1117]) );
  XNOR U6574 ( .A(a[1117]), .B(n5642), .Z(n5641) );
  IV U6575 ( .A(n5639), .Z(n5642) );
  XOR U6576 ( .A(n5643), .B(n5644), .Z(n5639) );
  ANDN U6577 ( .B(n5645), .A(n5646), .Z(n5643) );
  XNOR U6578 ( .A(b[1116]), .B(n5644), .Z(n5645) );
  XNOR U6579 ( .A(b[1116]), .B(n5646), .Z(c[1116]) );
  XNOR U6580 ( .A(a[1116]), .B(n5647), .Z(n5646) );
  IV U6581 ( .A(n5644), .Z(n5647) );
  XOR U6582 ( .A(n5648), .B(n5649), .Z(n5644) );
  ANDN U6583 ( .B(n5650), .A(n5651), .Z(n5648) );
  XNOR U6584 ( .A(b[1115]), .B(n5649), .Z(n5650) );
  XNOR U6585 ( .A(b[1115]), .B(n5651), .Z(c[1115]) );
  XNOR U6586 ( .A(a[1115]), .B(n5652), .Z(n5651) );
  IV U6587 ( .A(n5649), .Z(n5652) );
  XOR U6588 ( .A(n5653), .B(n5654), .Z(n5649) );
  ANDN U6589 ( .B(n5655), .A(n5656), .Z(n5653) );
  XNOR U6590 ( .A(b[1114]), .B(n5654), .Z(n5655) );
  XNOR U6591 ( .A(b[1114]), .B(n5656), .Z(c[1114]) );
  XNOR U6592 ( .A(a[1114]), .B(n5657), .Z(n5656) );
  IV U6593 ( .A(n5654), .Z(n5657) );
  XOR U6594 ( .A(n5658), .B(n5659), .Z(n5654) );
  ANDN U6595 ( .B(n5660), .A(n5661), .Z(n5658) );
  XNOR U6596 ( .A(b[1113]), .B(n5659), .Z(n5660) );
  XNOR U6597 ( .A(b[1113]), .B(n5661), .Z(c[1113]) );
  XNOR U6598 ( .A(a[1113]), .B(n5662), .Z(n5661) );
  IV U6599 ( .A(n5659), .Z(n5662) );
  XOR U6600 ( .A(n5663), .B(n5664), .Z(n5659) );
  ANDN U6601 ( .B(n5665), .A(n5666), .Z(n5663) );
  XNOR U6602 ( .A(b[1112]), .B(n5664), .Z(n5665) );
  XNOR U6603 ( .A(b[1112]), .B(n5666), .Z(c[1112]) );
  XNOR U6604 ( .A(a[1112]), .B(n5667), .Z(n5666) );
  IV U6605 ( .A(n5664), .Z(n5667) );
  XOR U6606 ( .A(n5668), .B(n5669), .Z(n5664) );
  ANDN U6607 ( .B(n5670), .A(n5671), .Z(n5668) );
  XNOR U6608 ( .A(b[1111]), .B(n5669), .Z(n5670) );
  XNOR U6609 ( .A(b[1111]), .B(n5671), .Z(c[1111]) );
  XNOR U6610 ( .A(a[1111]), .B(n5672), .Z(n5671) );
  IV U6611 ( .A(n5669), .Z(n5672) );
  XOR U6612 ( .A(n5673), .B(n5674), .Z(n5669) );
  ANDN U6613 ( .B(n5675), .A(n5676), .Z(n5673) );
  XNOR U6614 ( .A(b[1110]), .B(n5674), .Z(n5675) );
  XNOR U6615 ( .A(b[1110]), .B(n5676), .Z(c[1110]) );
  XNOR U6616 ( .A(a[1110]), .B(n5677), .Z(n5676) );
  IV U6617 ( .A(n5674), .Z(n5677) );
  XOR U6618 ( .A(n5678), .B(n5679), .Z(n5674) );
  ANDN U6619 ( .B(n5680), .A(n5681), .Z(n5678) );
  XNOR U6620 ( .A(b[1109]), .B(n5679), .Z(n5680) );
  XNOR U6621 ( .A(b[110]), .B(n5682), .Z(c[110]) );
  XNOR U6622 ( .A(b[1109]), .B(n5681), .Z(c[1109]) );
  XNOR U6623 ( .A(a[1109]), .B(n5683), .Z(n5681) );
  IV U6624 ( .A(n5679), .Z(n5683) );
  XOR U6625 ( .A(n5684), .B(n5685), .Z(n5679) );
  ANDN U6626 ( .B(n5686), .A(n5687), .Z(n5684) );
  XNOR U6627 ( .A(b[1108]), .B(n5685), .Z(n5686) );
  XNOR U6628 ( .A(b[1108]), .B(n5687), .Z(c[1108]) );
  XNOR U6629 ( .A(a[1108]), .B(n5688), .Z(n5687) );
  IV U6630 ( .A(n5685), .Z(n5688) );
  XOR U6631 ( .A(n5689), .B(n5690), .Z(n5685) );
  ANDN U6632 ( .B(n5691), .A(n5692), .Z(n5689) );
  XNOR U6633 ( .A(b[1107]), .B(n5690), .Z(n5691) );
  XNOR U6634 ( .A(b[1107]), .B(n5692), .Z(c[1107]) );
  XNOR U6635 ( .A(a[1107]), .B(n5693), .Z(n5692) );
  IV U6636 ( .A(n5690), .Z(n5693) );
  XOR U6637 ( .A(n5694), .B(n5695), .Z(n5690) );
  ANDN U6638 ( .B(n5696), .A(n5697), .Z(n5694) );
  XNOR U6639 ( .A(b[1106]), .B(n5695), .Z(n5696) );
  XNOR U6640 ( .A(b[1106]), .B(n5697), .Z(c[1106]) );
  XNOR U6641 ( .A(a[1106]), .B(n5698), .Z(n5697) );
  IV U6642 ( .A(n5695), .Z(n5698) );
  XOR U6643 ( .A(n5699), .B(n5700), .Z(n5695) );
  ANDN U6644 ( .B(n5701), .A(n5702), .Z(n5699) );
  XNOR U6645 ( .A(b[1105]), .B(n5700), .Z(n5701) );
  XNOR U6646 ( .A(b[1105]), .B(n5702), .Z(c[1105]) );
  XNOR U6647 ( .A(a[1105]), .B(n5703), .Z(n5702) );
  IV U6648 ( .A(n5700), .Z(n5703) );
  XOR U6649 ( .A(n5704), .B(n5705), .Z(n5700) );
  ANDN U6650 ( .B(n5706), .A(n5707), .Z(n5704) );
  XNOR U6651 ( .A(b[1104]), .B(n5705), .Z(n5706) );
  XNOR U6652 ( .A(b[1104]), .B(n5707), .Z(c[1104]) );
  XNOR U6653 ( .A(a[1104]), .B(n5708), .Z(n5707) );
  IV U6654 ( .A(n5705), .Z(n5708) );
  XOR U6655 ( .A(n5709), .B(n5710), .Z(n5705) );
  ANDN U6656 ( .B(n5711), .A(n5712), .Z(n5709) );
  XNOR U6657 ( .A(b[1103]), .B(n5710), .Z(n5711) );
  XNOR U6658 ( .A(b[1103]), .B(n5712), .Z(c[1103]) );
  XNOR U6659 ( .A(a[1103]), .B(n5713), .Z(n5712) );
  IV U6660 ( .A(n5710), .Z(n5713) );
  XOR U6661 ( .A(n5714), .B(n5715), .Z(n5710) );
  ANDN U6662 ( .B(n5716), .A(n5717), .Z(n5714) );
  XNOR U6663 ( .A(b[1102]), .B(n5715), .Z(n5716) );
  XNOR U6664 ( .A(b[1102]), .B(n5717), .Z(c[1102]) );
  XNOR U6665 ( .A(a[1102]), .B(n5718), .Z(n5717) );
  IV U6666 ( .A(n5715), .Z(n5718) );
  XOR U6667 ( .A(n5719), .B(n5720), .Z(n5715) );
  ANDN U6668 ( .B(n5721), .A(n5722), .Z(n5719) );
  XNOR U6669 ( .A(b[1101]), .B(n5720), .Z(n5721) );
  XNOR U6670 ( .A(b[1101]), .B(n5722), .Z(c[1101]) );
  XNOR U6671 ( .A(a[1101]), .B(n5723), .Z(n5722) );
  IV U6672 ( .A(n5720), .Z(n5723) );
  XOR U6673 ( .A(n5724), .B(n5725), .Z(n5720) );
  ANDN U6674 ( .B(n5726), .A(n5727), .Z(n5724) );
  XNOR U6675 ( .A(b[1100]), .B(n5725), .Z(n5726) );
  XNOR U6676 ( .A(b[1100]), .B(n5727), .Z(c[1100]) );
  XNOR U6677 ( .A(a[1100]), .B(n5728), .Z(n5727) );
  IV U6678 ( .A(n5725), .Z(n5728) );
  XOR U6679 ( .A(n5729), .B(n5730), .Z(n5725) );
  ANDN U6680 ( .B(n5731), .A(n5732), .Z(n5729) );
  XNOR U6681 ( .A(b[1099]), .B(n5730), .Z(n5731) );
  XNOR U6682 ( .A(b[10]), .B(n5733), .Z(c[10]) );
  XNOR U6683 ( .A(b[109]), .B(n5734), .Z(c[109]) );
  XNOR U6684 ( .A(b[1099]), .B(n5732), .Z(c[1099]) );
  XNOR U6685 ( .A(a[1099]), .B(n5735), .Z(n5732) );
  IV U6686 ( .A(n5730), .Z(n5735) );
  XOR U6687 ( .A(n5736), .B(n5737), .Z(n5730) );
  ANDN U6688 ( .B(n5738), .A(n5739), .Z(n5736) );
  XNOR U6689 ( .A(b[1098]), .B(n5737), .Z(n5738) );
  XNOR U6690 ( .A(b[1098]), .B(n5739), .Z(c[1098]) );
  XNOR U6691 ( .A(a[1098]), .B(n5740), .Z(n5739) );
  IV U6692 ( .A(n5737), .Z(n5740) );
  XOR U6693 ( .A(n5741), .B(n5742), .Z(n5737) );
  ANDN U6694 ( .B(n5743), .A(n5744), .Z(n5741) );
  XNOR U6695 ( .A(b[1097]), .B(n5742), .Z(n5743) );
  XNOR U6696 ( .A(b[1097]), .B(n5744), .Z(c[1097]) );
  XNOR U6697 ( .A(a[1097]), .B(n5745), .Z(n5744) );
  IV U6698 ( .A(n5742), .Z(n5745) );
  XOR U6699 ( .A(n5746), .B(n5747), .Z(n5742) );
  ANDN U6700 ( .B(n5748), .A(n5749), .Z(n5746) );
  XNOR U6701 ( .A(b[1096]), .B(n5747), .Z(n5748) );
  XNOR U6702 ( .A(b[1096]), .B(n5749), .Z(c[1096]) );
  XNOR U6703 ( .A(a[1096]), .B(n5750), .Z(n5749) );
  IV U6704 ( .A(n5747), .Z(n5750) );
  XOR U6705 ( .A(n5751), .B(n5752), .Z(n5747) );
  ANDN U6706 ( .B(n5753), .A(n5754), .Z(n5751) );
  XNOR U6707 ( .A(b[1095]), .B(n5752), .Z(n5753) );
  XNOR U6708 ( .A(b[1095]), .B(n5754), .Z(c[1095]) );
  XNOR U6709 ( .A(a[1095]), .B(n5755), .Z(n5754) );
  IV U6710 ( .A(n5752), .Z(n5755) );
  XOR U6711 ( .A(n5756), .B(n5757), .Z(n5752) );
  ANDN U6712 ( .B(n5758), .A(n5759), .Z(n5756) );
  XNOR U6713 ( .A(b[1094]), .B(n5757), .Z(n5758) );
  XNOR U6714 ( .A(b[1094]), .B(n5759), .Z(c[1094]) );
  XNOR U6715 ( .A(a[1094]), .B(n5760), .Z(n5759) );
  IV U6716 ( .A(n5757), .Z(n5760) );
  XOR U6717 ( .A(n5761), .B(n5762), .Z(n5757) );
  ANDN U6718 ( .B(n5763), .A(n5764), .Z(n5761) );
  XNOR U6719 ( .A(b[1093]), .B(n5762), .Z(n5763) );
  XNOR U6720 ( .A(b[1093]), .B(n5764), .Z(c[1093]) );
  XNOR U6721 ( .A(a[1093]), .B(n5765), .Z(n5764) );
  IV U6722 ( .A(n5762), .Z(n5765) );
  XOR U6723 ( .A(n5766), .B(n5767), .Z(n5762) );
  ANDN U6724 ( .B(n5768), .A(n5769), .Z(n5766) );
  XNOR U6725 ( .A(b[1092]), .B(n5767), .Z(n5768) );
  XNOR U6726 ( .A(b[1092]), .B(n5769), .Z(c[1092]) );
  XNOR U6727 ( .A(a[1092]), .B(n5770), .Z(n5769) );
  IV U6728 ( .A(n5767), .Z(n5770) );
  XOR U6729 ( .A(n5771), .B(n5772), .Z(n5767) );
  ANDN U6730 ( .B(n5773), .A(n5774), .Z(n5771) );
  XNOR U6731 ( .A(b[1091]), .B(n5772), .Z(n5773) );
  XNOR U6732 ( .A(b[1091]), .B(n5774), .Z(c[1091]) );
  XNOR U6733 ( .A(a[1091]), .B(n5775), .Z(n5774) );
  IV U6734 ( .A(n5772), .Z(n5775) );
  XOR U6735 ( .A(n5776), .B(n5777), .Z(n5772) );
  ANDN U6736 ( .B(n5778), .A(n5779), .Z(n5776) );
  XNOR U6737 ( .A(b[1090]), .B(n5777), .Z(n5778) );
  XNOR U6738 ( .A(b[1090]), .B(n5779), .Z(c[1090]) );
  XNOR U6739 ( .A(a[1090]), .B(n5780), .Z(n5779) );
  IV U6740 ( .A(n5777), .Z(n5780) );
  XOR U6741 ( .A(n5781), .B(n5782), .Z(n5777) );
  ANDN U6742 ( .B(n5783), .A(n5784), .Z(n5781) );
  XNOR U6743 ( .A(b[1089]), .B(n5782), .Z(n5783) );
  XNOR U6744 ( .A(b[108]), .B(n5785), .Z(c[108]) );
  XNOR U6745 ( .A(b[1089]), .B(n5784), .Z(c[1089]) );
  XNOR U6746 ( .A(a[1089]), .B(n5786), .Z(n5784) );
  IV U6747 ( .A(n5782), .Z(n5786) );
  XOR U6748 ( .A(n5787), .B(n5788), .Z(n5782) );
  ANDN U6749 ( .B(n5789), .A(n5790), .Z(n5787) );
  XNOR U6750 ( .A(b[1088]), .B(n5788), .Z(n5789) );
  XNOR U6751 ( .A(b[1088]), .B(n5790), .Z(c[1088]) );
  XNOR U6752 ( .A(a[1088]), .B(n5791), .Z(n5790) );
  IV U6753 ( .A(n5788), .Z(n5791) );
  XOR U6754 ( .A(n5792), .B(n5793), .Z(n5788) );
  ANDN U6755 ( .B(n5794), .A(n5795), .Z(n5792) );
  XNOR U6756 ( .A(b[1087]), .B(n5793), .Z(n5794) );
  XNOR U6757 ( .A(b[1087]), .B(n5795), .Z(c[1087]) );
  XNOR U6758 ( .A(a[1087]), .B(n5796), .Z(n5795) );
  IV U6759 ( .A(n5793), .Z(n5796) );
  XOR U6760 ( .A(n5797), .B(n5798), .Z(n5793) );
  ANDN U6761 ( .B(n5799), .A(n5800), .Z(n5797) );
  XNOR U6762 ( .A(b[1086]), .B(n5798), .Z(n5799) );
  XNOR U6763 ( .A(b[1086]), .B(n5800), .Z(c[1086]) );
  XNOR U6764 ( .A(a[1086]), .B(n5801), .Z(n5800) );
  IV U6765 ( .A(n5798), .Z(n5801) );
  XOR U6766 ( .A(n5802), .B(n5803), .Z(n5798) );
  ANDN U6767 ( .B(n5804), .A(n5805), .Z(n5802) );
  XNOR U6768 ( .A(b[1085]), .B(n5803), .Z(n5804) );
  XNOR U6769 ( .A(b[1085]), .B(n5805), .Z(c[1085]) );
  XNOR U6770 ( .A(a[1085]), .B(n5806), .Z(n5805) );
  IV U6771 ( .A(n5803), .Z(n5806) );
  XOR U6772 ( .A(n5807), .B(n5808), .Z(n5803) );
  ANDN U6773 ( .B(n5809), .A(n5810), .Z(n5807) );
  XNOR U6774 ( .A(b[1084]), .B(n5808), .Z(n5809) );
  XNOR U6775 ( .A(b[1084]), .B(n5810), .Z(c[1084]) );
  XNOR U6776 ( .A(a[1084]), .B(n5811), .Z(n5810) );
  IV U6777 ( .A(n5808), .Z(n5811) );
  XOR U6778 ( .A(n5812), .B(n5813), .Z(n5808) );
  ANDN U6779 ( .B(n5814), .A(n5815), .Z(n5812) );
  XNOR U6780 ( .A(b[1083]), .B(n5813), .Z(n5814) );
  XNOR U6781 ( .A(b[1083]), .B(n5815), .Z(c[1083]) );
  XNOR U6782 ( .A(a[1083]), .B(n5816), .Z(n5815) );
  IV U6783 ( .A(n5813), .Z(n5816) );
  XOR U6784 ( .A(n5817), .B(n5818), .Z(n5813) );
  ANDN U6785 ( .B(n5819), .A(n5820), .Z(n5817) );
  XNOR U6786 ( .A(b[1082]), .B(n5818), .Z(n5819) );
  XNOR U6787 ( .A(b[1082]), .B(n5820), .Z(c[1082]) );
  XNOR U6788 ( .A(a[1082]), .B(n5821), .Z(n5820) );
  IV U6789 ( .A(n5818), .Z(n5821) );
  XOR U6790 ( .A(n5822), .B(n5823), .Z(n5818) );
  ANDN U6791 ( .B(n5824), .A(n5825), .Z(n5822) );
  XNOR U6792 ( .A(b[1081]), .B(n5823), .Z(n5824) );
  XNOR U6793 ( .A(b[1081]), .B(n5825), .Z(c[1081]) );
  XNOR U6794 ( .A(a[1081]), .B(n5826), .Z(n5825) );
  IV U6795 ( .A(n5823), .Z(n5826) );
  XOR U6796 ( .A(n5827), .B(n5828), .Z(n5823) );
  ANDN U6797 ( .B(n5829), .A(n5830), .Z(n5827) );
  XNOR U6798 ( .A(b[1080]), .B(n5828), .Z(n5829) );
  XNOR U6799 ( .A(b[1080]), .B(n5830), .Z(c[1080]) );
  XNOR U6800 ( .A(a[1080]), .B(n5831), .Z(n5830) );
  IV U6801 ( .A(n5828), .Z(n5831) );
  XOR U6802 ( .A(n5832), .B(n5833), .Z(n5828) );
  ANDN U6803 ( .B(n5834), .A(n5835), .Z(n5832) );
  XNOR U6804 ( .A(b[1079]), .B(n5833), .Z(n5834) );
  XNOR U6805 ( .A(b[107]), .B(n5836), .Z(c[107]) );
  XNOR U6806 ( .A(b[1079]), .B(n5835), .Z(c[1079]) );
  XNOR U6807 ( .A(a[1079]), .B(n5837), .Z(n5835) );
  IV U6808 ( .A(n5833), .Z(n5837) );
  XOR U6809 ( .A(n5838), .B(n5839), .Z(n5833) );
  ANDN U6810 ( .B(n5840), .A(n5841), .Z(n5838) );
  XNOR U6811 ( .A(b[1078]), .B(n5839), .Z(n5840) );
  XNOR U6812 ( .A(b[1078]), .B(n5841), .Z(c[1078]) );
  XNOR U6813 ( .A(a[1078]), .B(n5842), .Z(n5841) );
  IV U6814 ( .A(n5839), .Z(n5842) );
  XOR U6815 ( .A(n5843), .B(n5844), .Z(n5839) );
  ANDN U6816 ( .B(n5845), .A(n5846), .Z(n5843) );
  XNOR U6817 ( .A(b[1077]), .B(n5844), .Z(n5845) );
  XNOR U6818 ( .A(b[1077]), .B(n5846), .Z(c[1077]) );
  XNOR U6819 ( .A(a[1077]), .B(n5847), .Z(n5846) );
  IV U6820 ( .A(n5844), .Z(n5847) );
  XOR U6821 ( .A(n5848), .B(n5849), .Z(n5844) );
  ANDN U6822 ( .B(n5850), .A(n5851), .Z(n5848) );
  XNOR U6823 ( .A(b[1076]), .B(n5849), .Z(n5850) );
  XNOR U6824 ( .A(b[1076]), .B(n5851), .Z(c[1076]) );
  XNOR U6825 ( .A(a[1076]), .B(n5852), .Z(n5851) );
  IV U6826 ( .A(n5849), .Z(n5852) );
  XOR U6827 ( .A(n5853), .B(n5854), .Z(n5849) );
  ANDN U6828 ( .B(n5855), .A(n5856), .Z(n5853) );
  XNOR U6829 ( .A(b[1075]), .B(n5854), .Z(n5855) );
  XNOR U6830 ( .A(b[1075]), .B(n5856), .Z(c[1075]) );
  XNOR U6831 ( .A(a[1075]), .B(n5857), .Z(n5856) );
  IV U6832 ( .A(n5854), .Z(n5857) );
  XOR U6833 ( .A(n5858), .B(n5859), .Z(n5854) );
  ANDN U6834 ( .B(n5860), .A(n5861), .Z(n5858) );
  XNOR U6835 ( .A(b[1074]), .B(n5859), .Z(n5860) );
  XNOR U6836 ( .A(b[1074]), .B(n5861), .Z(c[1074]) );
  XNOR U6837 ( .A(a[1074]), .B(n5862), .Z(n5861) );
  IV U6838 ( .A(n5859), .Z(n5862) );
  XOR U6839 ( .A(n5863), .B(n5864), .Z(n5859) );
  ANDN U6840 ( .B(n5865), .A(n5866), .Z(n5863) );
  XNOR U6841 ( .A(b[1073]), .B(n5864), .Z(n5865) );
  XNOR U6842 ( .A(b[1073]), .B(n5866), .Z(c[1073]) );
  XNOR U6843 ( .A(a[1073]), .B(n5867), .Z(n5866) );
  IV U6844 ( .A(n5864), .Z(n5867) );
  XOR U6845 ( .A(n5868), .B(n5869), .Z(n5864) );
  ANDN U6846 ( .B(n5870), .A(n5871), .Z(n5868) );
  XNOR U6847 ( .A(b[1072]), .B(n5869), .Z(n5870) );
  XNOR U6848 ( .A(b[1072]), .B(n5871), .Z(c[1072]) );
  XNOR U6849 ( .A(a[1072]), .B(n5872), .Z(n5871) );
  IV U6850 ( .A(n5869), .Z(n5872) );
  XOR U6851 ( .A(n5873), .B(n5874), .Z(n5869) );
  ANDN U6852 ( .B(n5875), .A(n5876), .Z(n5873) );
  XNOR U6853 ( .A(b[1071]), .B(n5874), .Z(n5875) );
  XNOR U6854 ( .A(b[1071]), .B(n5876), .Z(c[1071]) );
  XNOR U6855 ( .A(a[1071]), .B(n5877), .Z(n5876) );
  IV U6856 ( .A(n5874), .Z(n5877) );
  XOR U6857 ( .A(n5878), .B(n5879), .Z(n5874) );
  ANDN U6858 ( .B(n5880), .A(n5881), .Z(n5878) );
  XNOR U6859 ( .A(b[1070]), .B(n5879), .Z(n5880) );
  XNOR U6860 ( .A(b[1070]), .B(n5881), .Z(c[1070]) );
  XNOR U6861 ( .A(a[1070]), .B(n5882), .Z(n5881) );
  IV U6862 ( .A(n5879), .Z(n5882) );
  XOR U6863 ( .A(n5883), .B(n5884), .Z(n5879) );
  ANDN U6864 ( .B(n5885), .A(n5886), .Z(n5883) );
  XNOR U6865 ( .A(b[1069]), .B(n5884), .Z(n5885) );
  XNOR U6866 ( .A(b[106]), .B(n5887), .Z(c[106]) );
  XNOR U6867 ( .A(b[1069]), .B(n5886), .Z(c[1069]) );
  XNOR U6868 ( .A(a[1069]), .B(n5888), .Z(n5886) );
  IV U6869 ( .A(n5884), .Z(n5888) );
  XOR U6870 ( .A(n5889), .B(n5890), .Z(n5884) );
  ANDN U6871 ( .B(n5891), .A(n5892), .Z(n5889) );
  XNOR U6872 ( .A(b[1068]), .B(n5890), .Z(n5891) );
  XNOR U6873 ( .A(b[1068]), .B(n5892), .Z(c[1068]) );
  XNOR U6874 ( .A(a[1068]), .B(n5893), .Z(n5892) );
  IV U6875 ( .A(n5890), .Z(n5893) );
  XOR U6876 ( .A(n5894), .B(n5895), .Z(n5890) );
  ANDN U6877 ( .B(n5896), .A(n5897), .Z(n5894) );
  XNOR U6878 ( .A(b[1067]), .B(n5895), .Z(n5896) );
  XNOR U6879 ( .A(b[1067]), .B(n5897), .Z(c[1067]) );
  XNOR U6880 ( .A(a[1067]), .B(n5898), .Z(n5897) );
  IV U6881 ( .A(n5895), .Z(n5898) );
  XOR U6882 ( .A(n5899), .B(n5900), .Z(n5895) );
  ANDN U6883 ( .B(n5901), .A(n5902), .Z(n5899) );
  XNOR U6884 ( .A(b[1066]), .B(n5900), .Z(n5901) );
  XNOR U6885 ( .A(b[1066]), .B(n5902), .Z(c[1066]) );
  XNOR U6886 ( .A(a[1066]), .B(n5903), .Z(n5902) );
  IV U6887 ( .A(n5900), .Z(n5903) );
  XOR U6888 ( .A(n5904), .B(n5905), .Z(n5900) );
  ANDN U6889 ( .B(n5906), .A(n5907), .Z(n5904) );
  XNOR U6890 ( .A(b[1065]), .B(n5905), .Z(n5906) );
  XNOR U6891 ( .A(b[1065]), .B(n5907), .Z(c[1065]) );
  XNOR U6892 ( .A(a[1065]), .B(n5908), .Z(n5907) );
  IV U6893 ( .A(n5905), .Z(n5908) );
  XOR U6894 ( .A(n5909), .B(n5910), .Z(n5905) );
  ANDN U6895 ( .B(n5911), .A(n5912), .Z(n5909) );
  XNOR U6896 ( .A(b[1064]), .B(n5910), .Z(n5911) );
  XNOR U6897 ( .A(b[1064]), .B(n5912), .Z(c[1064]) );
  XNOR U6898 ( .A(a[1064]), .B(n5913), .Z(n5912) );
  IV U6899 ( .A(n5910), .Z(n5913) );
  XOR U6900 ( .A(n5914), .B(n5915), .Z(n5910) );
  ANDN U6901 ( .B(n5916), .A(n5917), .Z(n5914) );
  XNOR U6902 ( .A(b[1063]), .B(n5915), .Z(n5916) );
  XNOR U6903 ( .A(b[1063]), .B(n5917), .Z(c[1063]) );
  XNOR U6904 ( .A(a[1063]), .B(n5918), .Z(n5917) );
  IV U6905 ( .A(n5915), .Z(n5918) );
  XOR U6906 ( .A(n5919), .B(n5920), .Z(n5915) );
  ANDN U6907 ( .B(n5921), .A(n5922), .Z(n5919) );
  XNOR U6908 ( .A(b[1062]), .B(n5920), .Z(n5921) );
  XNOR U6909 ( .A(b[1062]), .B(n5922), .Z(c[1062]) );
  XNOR U6910 ( .A(a[1062]), .B(n5923), .Z(n5922) );
  IV U6911 ( .A(n5920), .Z(n5923) );
  XOR U6912 ( .A(n5924), .B(n5925), .Z(n5920) );
  ANDN U6913 ( .B(n5926), .A(n5927), .Z(n5924) );
  XNOR U6914 ( .A(b[1061]), .B(n5925), .Z(n5926) );
  XNOR U6915 ( .A(b[1061]), .B(n5927), .Z(c[1061]) );
  XNOR U6916 ( .A(a[1061]), .B(n5928), .Z(n5927) );
  IV U6917 ( .A(n5925), .Z(n5928) );
  XOR U6918 ( .A(n5929), .B(n5930), .Z(n5925) );
  ANDN U6919 ( .B(n5931), .A(n5932), .Z(n5929) );
  XNOR U6920 ( .A(b[1060]), .B(n5930), .Z(n5931) );
  XNOR U6921 ( .A(b[1060]), .B(n5932), .Z(c[1060]) );
  XNOR U6922 ( .A(a[1060]), .B(n5933), .Z(n5932) );
  IV U6923 ( .A(n5930), .Z(n5933) );
  XOR U6924 ( .A(n5934), .B(n5935), .Z(n5930) );
  ANDN U6925 ( .B(n5936), .A(n5937), .Z(n5934) );
  XNOR U6926 ( .A(b[1059]), .B(n5935), .Z(n5936) );
  XNOR U6927 ( .A(b[105]), .B(n5938), .Z(c[105]) );
  XNOR U6928 ( .A(b[1059]), .B(n5937), .Z(c[1059]) );
  XNOR U6929 ( .A(a[1059]), .B(n5939), .Z(n5937) );
  IV U6930 ( .A(n5935), .Z(n5939) );
  XOR U6931 ( .A(n5940), .B(n5941), .Z(n5935) );
  ANDN U6932 ( .B(n5942), .A(n5943), .Z(n5940) );
  XNOR U6933 ( .A(b[1058]), .B(n5941), .Z(n5942) );
  XNOR U6934 ( .A(b[1058]), .B(n5943), .Z(c[1058]) );
  XNOR U6935 ( .A(a[1058]), .B(n5944), .Z(n5943) );
  IV U6936 ( .A(n5941), .Z(n5944) );
  XOR U6937 ( .A(n5945), .B(n5946), .Z(n5941) );
  ANDN U6938 ( .B(n5947), .A(n5948), .Z(n5945) );
  XNOR U6939 ( .A(b[1057]), .B(n5946), .Z(n5947) );
  XNOR U6940 ( .A(b[1057]), .B(n5948), .Z(c[1057]) );
  XNOR U6941 ( .A(a[1057]), .B(n5949), .Z(n5948) );
  IV U6942 ( .A(n5946), .Z(n5949) );
  XOR U6943 ( .A(n5950), .B(n5951), .Z(n5946) );
  ANDN U6944 ( .B(n5952), .A(n5953), .Z(n5950) );
  XNOR U6945 ( .A(b[1056]), .B(n5951), .Z(n5952) );
  XNOR U6946 ( .A(b[1056]), .B(n5953), .Z(c[1056]) );
  XNOR U6947 ( .A(a[1056]), .B(n5954), .Z(n5953) );
  IV U6948 ( .A(n5951), .Z(n5954) );
  XOR U6949 ( .A(n5955), .B(n5956), .Z(n5951) );
  ANDN U6950 ( .B(n5957), .A(n5958), .Z(n5955) );
  XNOR U6951 ( .A(b[1055]), .B(n5956), .Z(n5957) );
  XNOR U6952 ( .A(b[1055]), .B(n5958), .Z(c[1055]) );
  XNOR U6953 ( .A(a[1055]), .B(n5959), .Z(n5958) );
  IV U6954 ( .A(n5956), .Z(n5959) );
  XOR U6955 ( .A(n5960), .B(n5961), .Z(n5956) );
  ANDN U6956 ( .B(n5962), .A(n5963), .Z(n5960) );
  XNOR U6957 ( .A(b[1054]), .B(n5961), .Z(n5962) );
  XNOR U6958 ( .A(b[1054]), .B(n5963), .Z(c[1054]) );
  XNOR U6959 ( .A(a[1054]), .B(n5964), .Z(n5963) );
  IV U6960 ( .A(n5961), .Z(n5964) );
  XOR U6961 ( .A(n5965), .B(n5966), .Z(n5961) );
  ANDN U6962 ( .B(n5967), .A(n5968), .Z(n5965) );
  XNOR U6963 ( .A(b[1053]), .B(n5966), .Z(n5967) );
  XNOR U6964 ( .A(b[1053]), .B(n5968), .Z(c[1053]) );
  XNOR U6965 ( .A(a[1053]), .B(n5969), .Z(n5968) );
  IV U6966 ( .A(n5966), .Z(n5969) );
  XOR U6967 ( .A(n5970), .B(n5971), .Z(n5966) );
  ANDN U6968 ( .B(n5972), .A(n5973), .Z(n5970) );
  XNOR U6969 ( .A(b[1052]), .B(n5971), .Z(n5972) );
  XNOR U6970 ( .A(b[1052]), .B(n5973), .Z(c[1052]) );
  XNOR U6971 ( .A(a[1052]), .B(n5974), .Z(n5973) );
  IV U6972 ( .A(n5971), .Z(n5974) );
  XOR U6973 ( .A(n5975), .B(n5976), .Z(n5971) );
  ANDN U6974 ( .B(n5977), .A(n5978), .Z(n5975) );
  XNOR U6975 ( .A(b[1051]), .B(n5976), .Z(n5977) );
  XNOR U6976 ( .A(b[1051]), .B(n5978), .Z(c[1051]) );
  XNOR U6977 ( .A(a[1051]), .B(n5979), .Z(n5978) );
  IV U6978 ( .A(n5976), .Z(n5979) );
  XOR U6979 ( .A(n5980), .B(n5981), .Z(n5976) );
  ANDN U6980 ( .B(n5982), .A(n5983), .Z(n5980) );
  XNOR U6981 ( .A(b[1050]), .B(n5981), .Z(n5982) );
  XNOR U6982 ( .A(b[1050]), .B(n5983), .Z(c[1050]) );
  XNOR U6983 ( .A(a[1050]), .B(n5984), .Z(n5983) );
  IV U6984 ( .A(n5981), .Z(n5984) );
  XOR U6985 ( .A(n5985), .B(n5986), .Z(n5981) );
  ANDN U6986 ( .B(n5987), .A(n5988), .Z(n5985) );
  XNOR U6987 ( .A(b[1049]), .B(n5986), .Z(n5987) );
  XNOR U6988 ( .A(b[104]), .B(n5989), .Z(c[104]) );
  XNOR U6989 ( .A(b[1049]), .B(n5988), .Z(c[1049]) );
  XNOR U6990 ( .A(a[1049]), .B(n5990), .Z(n5988) );
  IV U6991 ( .A(n5986), .Z(n5990) );
  XOR U6992 ( .A(n5991), .B(n5992), .Z(n5986) );
  ANDN U6993 ( .B(n5993), .A(n5994), .Z(n5991) );
  XNOR U6994 ( .A(b[1048]), .B(n5992), .Z(n5993) );
  XNOR U6995 ( .A(b[1048]), .B(n5994), .Z(c[1048]) );
  XNOR U6996 ( .A(a[1048]), .B(n5995), .Z(n5994) );
  IV U6997 ( .A(n5992), .Z(n5995) );
  XOR U6998 ( .A(n5996), .B(n5997), .Z(n5992) );
  ANDN U6999 ( .B(n5998), .A(n5999), .Z(n5996) );
  XNOR U7000 ( .A(b[1047]), .B(n5997), .Z(n5998) );
  XNOR U7001 ( .A(b[1047]), .B(n5999), .Z(c[1047]) );
  XNOR U7002 ( .A(a[1047]), .B(n6000), .Z(n5999) );
  IV U7003 ( .A(n5997), .Z(n6000) );
  XOR U7004 ( .A(n6001), .B(n6002), .Z(n5997) );
  ANDN U7005 ( .B(n6003), .A(n6004), .Z(n6001) );
  XNOR U7006 ( .A(b[1046]), .B(n6002), .Z(n6003) );
  XNOR U7007 ( .A(b[1046]), .B(n6004), .Z(c[1046]) );
  XNOR U7008 ( .A(a[1046]), .B(n6005), .Z(n6004) );
  IV U7009 ( .A(n6002), .Z(n6005) );
  XOR U7010 ( .A(n6006), .B(n6007), .Z(n6002) );
  ANDN U7011 ( .B(n6008), .A(n6009), .Z(n6006) );
  XNOR U7012 ( .A(b[1045]), .B(n6007), .Z(n6008) );
  XNOR U7013 ( .A(b[1045]), .B(n6009), .Z(c[1045]) );
  XNOR U7014 ( .A(a[1045]), .B(n6010), .Z(n6009) );
  IV U7015 ( .A(n6007), .Z(n6010) );
  XOR U7016 ( .A(n6011), .B(n6012), .Z(n6007) );
  ANDN U7017 ( .B(n6013), .A(n6014), .Z(n6011) );
  XNOR U7018 ( .A(b[1044]), .B(n6012), .Z(n6013) );
  XNOR U7019 ( .A(b[1044]), .B(n6014), .Z(c[1044]) );
  XNOR U7020 ( .A(a[1044]), .B(n6015), .Z(n6014) );
  IV U7021 ( .A(n6012), .Z(n6015) );
  XOR U7022 ( .A(n6016), .B(n6017), .Z(n6012) );
  ANDN U7023 ( .B(n6018), .A(n6019), .Z(n6016) );
  XNOR U7024 ( .A(b[1043]), .B(n6017), .Z(n6018) );
  XNOR U7025 ( .A(b[1043]), .B(n6019), .Z(c[1043]) );
  XNOR U7026 ( .A(a[1043]), .B(n6020), .Z(n6019) );
  IV U7027 ( .A(n6017), .Z(n6020) );
  XOR U7028 ( .A(n6021), .B(n6022), .Z(n6017) );
  ANDN U7029 ( .B(n6023), .A(n6024), .Z(n6021) );
  XNOR U7030 ( .A(b[1042]), .B(n6022), .Z(n6023) );
  XNOR U7031 ( .A(b[1042]), .B(n6024), .Z(c[1042]) );
  XNOR U7032 ( .A(a[1042]), .B(n6025), .Z(n6024) );
  IV U7033 ( .A(n6022), .Z(n6025) );
  XOR U7034 ( .A(n6026), .B(n6027), .Z(n6022) );
  ANDN U7035 ( .B(n6028), .A(n6029), .Z(n6026) );
  XNOR U7036 ( .A(b[1041]), .B(n6027), .Z(n6028) );
  XNOR U7037 ( .A(b[1041]), .B(n6029), .Z(c[1041]) );
  XNOR U7038 ( .A(a[1041]), .B(n6030), .Z(n6029) );
  IV U7039 ( .A(n6027), .Z(n6030) );
  XOR U7040 ( .A(n6031), .B(n6032), .Z(n6027) );
  ANDN U7041 ( .B(n6033), .A(n6034), .Z(n6031) );
  XNOR U7042 ( .A(b[1040]), .B(n6032), .Z(n6033) );
  XNOR U7043 ( .A(b[1040]), .B(n6034), .Z(c[1040]) );
  XNOR U7044 ( .A(a[1040]), .B(n6035), .Z(n6034) );
  IV U7045 ( .A(n6032), .Z(n6035) );
  XOR U7046 ( .A(n6036), .B(n6037), .Z(n6032) );
  ANDN U7047 ( .B(n6038), .A(n6039), .Z(n6036) );
  XNOR U7048 ( .A(b[1039]), .B(n6037), .Z(n6038) );
  XNOR U7049 ( .A(b[103]), .B(n6040), .Z(c[103]) );
  XNOR U7050 ( .A(b[1039]), .B(n6039), .Z(c[1039]) );
  XNOR U7051 ( .A(a[1039]), .B(n6041), .Z(n6039) );
  IV U7052 ( .A(n6037), .Z(n6041) );
  XOR U7053 ( .A(n6042), .B(n6043), .Z(n6037) );
  ANDN U7054 ( .B(n6044), .A(n6045), .Z(n6042) );
  XNOR U7055 ( .A(b[1038]), .B(n6043), .Z(n6044) );
  XNOR U7056 ( .A(b[1038]), .B(n6045), .Z(c[1038]) );
  XNOR U7057 ( .A(a[1038]), .B(n6046), .Z(n6045) );
  IV U7058 ( .A(n6043), .Z(n6046) );
  XOR U7059 ( .A(n6047), .B(n6048), .Z(n6043) );
  ANDN U7060 ( .B(n6049), .A(n6050), .Z(n6047) );
  XNOR U7061 ( .A(b[1037]), .B(n6048), .Z(n6049) );
  XNOR U7062 ( .A(b[1037]), .B(n6050), .Z(c[1037]) );
  XNOR U7063 ( .A(a[1037]), .B(n6051), .Z(n6050) );
  IV U7064 ( .A(n6048), .Z(n6051) );
  XOR U7065 ( .A(n6052), .B(n6053), .Z(n6048) );
  ANDN U7066 ( .B(n6054), .A(n6055), .Z(n6052) );
  XNOR U7067 ( .A(b[1036]), .B(n6053), .Z(n6054) );
  XNOR U7068 ( .A(b[1036]), .B(n6055), .Z(c[1036]) );
  XNOR U7069 ( .A(a[1036]), .B(n6056), .Z(n6055) );
  IV U7070 ( .A(n6053), .Z(n6056) );
  XOR U7071 ( .A(n6057), .B(n6058), .Z(n6053) );
  ANDN U7072 ( .B(n6059), .A(n6060), .Z(n6057) );
  XNOR U7073 ( .A(b[1035]), .B(n6058), .Z(n6059) );
  XNOR U7074 ( .A(b[1035]), .B(n6060), .Z(c[1035]) );
  XNOR U7075 ( .A(a[1035]), .B(n6061), .Z(n6060) );
  IV U7076 ( .A(n6058), .Z(n6061) );
  XOR U7077 ( .A(n6062), .B(n6063), .Z(n6058) );
  ANDN U7078 ( .B(n6064), .A(n6065), .Z(n6062) );
  XNOR U7079 ( .A(b[1034]), .B(n6063), .Z(n6064) );
  XNOR U7080 ( .A(b[1034]), .B(n6065), .Z(c[1034]) );
  XNOR U7081 ( .A(a[1034]), .B(n6066), .Z(n6065) );
  IV U7082 ( .A(n6063), .Z(n6066) );
  XOR U7083 ( .A(n6067), .B(n6068), .Z(n6063) );
  ANDN U7084 ( .B(n6069), .A(n6070), .Z(n6067) );
  XNOR U7085 ( .A(b[1033]), .B(n6068), .Z(n6069) );
  XNOR U7086 ( .A(b[1033]), .B(n6070), .Z(c[1033]) );
  XNOR U7087 ( .A(a[1033]), .B(n6071), .Z(n6070) );
  IV U7088 ( .A(n6068), .Z(n6071) );
  XOR U7089 ( .A(n6072), .B(n6073), .Z(n6068) );
  ANDN U7090 ( .B(n6074), .A(n6075), .Z(n6072) );
  XNOR U7091 ( .A(b[1032]), .B(n6073), .Z(n6074) );
  XNOR U7092 ( .A(b[1032]), .B(n6075), .Z(c[1032]) );
  XNOR U7093 ( .A(a[1032]), .B(n6076), .Z(n6075) );
  IV U7094 ( .A(n6073), .Z(n6076) );
  XOR U7095 ( .A(n6077), .B(n6078), .Z(n6073) );
  ANDN U7096 ( .B(n6079), .A(n6080), .Z(n6077) );
  XNOR U7097 ( .A(b[1031]), .B(n6078), .Z(n6079) );
  XNOR U7098 ( .A(b[1031]), .B(n6080), .Z(c[1031]) );
  XNOR U7099 ( .A(a[1031]), .B(n6081), .Z(n6080) );
  IV U7100 ( .A(n6078), .Z(n6081) );
  XOR U7101 ( .A(n6082), .B(n6083), .Z(n6078) );
  ANDN U7102 ( .B(n6084), .A(n6085), .Z(n6082) );
  XNOR U7103 ( .A(b[1030]), .B(n6083), .Z(n6084) );
  XNOR U7104 ( .A(b[1030]), .B(n6085), .Z(c[1030]) );
  XNOR U7105 ( .A(a[1030]), .B(n6086), .Z(n6085) );
  IV U7106 ( .A(n6083), .Z(n6086) );
  XOR U7107 ( .A(n6087), .B(n6088), .Z(n6083) );
  ANDN U7108 ( .B(n6089), .A(n6090), .Z(n6087) );
  XNOR U7109 ( .A(b[1029]), .B(n6088), .Z(n6089) );
  XNOR U7110 ( .A(b[102]), .B(n6091), .Z(c[102]) );
  XNOR U7111 ( .A(b[1029]), .B(n6090), .Z(c[1029]) );
  XNOR U7112 ( .A(a[1029]), .B(n6092), .Z(n6090) );
  IV U7113 ( .A(n6088), .Z(n6092) );
  XOR U7114 ( .A(n6093), .B(n6094), .Z(n6088) );
  ANDN U7115 ( .B(n6095), .A(n6096), .Z(n6093) );
  XNOR U7116 ( .A(b[1028]), .B(n6094), .Z(n6095) );
  XNOR U7117 ( .A(b[1028]), .B(n6096), .Z(c[1028]) );
  XNOR U7118 ( .A(a[1028]), .B(n6097), .Z(n6096) );
  IV U7119 ( .A(n6094), .Z(n6097) );
  XOR U7120 ( .A(n6098), .B(n6099), .Z(n6094) );
  ANDN U7121 ( .B(n6100), .A(n6101), .Z(n6098) );
  XNOR U7122 ( .A(b[1027]), .B(n6099), .Z(n6100) );
  XNOR U7123 ( .A(b[1027]), .B(n6101), .Z(c[1027]) );
  XNOR U7124 ( .A(a[1027]), .B(n6102), .Z(n6101) );
  IV U7125 ( .A(n6099), .Z(n6102) );
  XOR U7126 ( .A(n6103), .B(n6104), .Z(n6099) );
  ANDN U7127 ( .B(n6105), .A(n6106), .Z(n6103) );
  XNOR U7128 ( .A(b[1026]), .B(n6104), .Z(n6105) );
  XNOR U7129 ( .A(b[1026]), .B(n6106), .Z(c[1026]) );
  XNOR U7130 ( .A(a[1026]), .B(n6107), .Z(n6106) );
  IV U7131 ( .A(n6104), .Z(n6107) );
  XOR U7132 ( .A(n6108), .B(n6109), .Z(n6104) );
  ANDN U7133 ( .B(n6110), .A(n6111), .Z(n6108) );
  XNOR U7134 ( .A(b[1025]), .B(n6109), .Z(n6110) );
  XNOR U7135 ( .A(b[1025]), .B(n6111), .Z(c[1025]) );
  XNOR U7136 ( .A(a[1025]), .B(n6112), .Z(n6111) );
  IV U7137 ( .A(n6109), .Z(n6112) );
  XOR U7138 ( .A(n6113), .B(n6114), .Z(n6109) );
  ANDN U7139 ( .B(n6115), .A(n6116), .Z(n6113) );
  XNOR U7140 ( .A(b[1024]), .B(n6114), .Z(n6115) );
  XNOR U7141 ( .A(b[1024]), .B(n6116), .Z(c[1024]) );
  XNOR U7142 ( .A(a[1024]), .B(n6117), .Z(n6116) );
  IV U7143 ( .A(n6114), .Z(n6117) );
  XOR U7144 ( .A(n6118), .B(n6119), .Z(n6114) );
  ANDN U7145 ( .B(n6120), .A(n6121), .Z(n6118) );
  XNOR U7146 ( .A(b[1023]), .B(n6119), .Z(n6120) );
  XNOR U7147 ( .A(b[1023]), .B(n6121), .Z(c[1023]) );
  XNOR U7148 ( .A(a[1023]), .B(n6122), .Z(n6121) );
  IV U7149 ( .A(n6119), .Z(n6122) );
  XOR U7150 ( .A(n6123), .B(n6124), .Z(n6119) );
  ANDN U7151 ( .B(n6125), .A(n6126), .Z(n6123) );
  XNOR U7152 ( .A(b[1022]), .B(n6124), .Z(n6125) );
  XNOR U7153 ( .A(b[1022]), .B(n6126), .Z(c[1022]) );
  XNOR U7154 ( .A(a[1022]), .B(n6127), .Z(n6126) );
  IV U7155 ( .A(n6124), .Z(n6127) );
  XOR U7156 ( .A(n6128), .B(n6129), .Z(n6124) );
  ANDN U7157 ( .B(n6130), .A(n6131), .Z(n6128) );
  XNOR U7158 ( .A(b[1021]), .B(n6129), .Z(n6130) );
  XNOR U7159 ( .A(b[1021]), .B(n6131), .Z(c[1021]) );
  XNOR U7160 ( .A(a[1021]), .B(n6132), .Z(n6131) );
  IV U7161 ( .A(n6129), .Z(n6132) );
  XOR U7162 ( .A(n6133), .B(n6134), .Z(n6129) );
  ANDN U7163 ( .B(n6135), .A(n6136), .Z(n6133) );
  XNOR U7164 ( .A(b[1020]), .B(n6134), .Z(n6135) );
  XNOR U7165 ( .A(b[1020]), .B(n6136), .Z(c[1020]) );
  XNOR U7166 ( .A(a[1020]), .B(n6137), .Z(n6136) );
  IV U7167 ( .A(n6134), .Z(n6137) );
  XOR U7168 ( .A(n6138), .B(n6139), .Z(n6134) );
  ANDN U7169 ( .B(n6140), .A(n6141), .Z(n6138) );
  XNOR U7170 ( .A(b[1019]), .B(n6139), .Z(n6140) );
  XNOR U7171 ( .A(b[101]), .B(n6142), .Z(c[101]) );
  XNOR U7172 ( .A(b[1019]), .B(n6141), .Z(c[1019]) );
  XNOR U7173 ( .A(a[1019]), .B(n6143), .Z(n6141) );
  IV U7174 ( .A(n6139), .Z(n6143) );
  XOR U7175 ( .A(n6144), .B(n6145), .Z(n6139) );
  ANDN U7176 ( .B(n6146), .A(n6147), .Z(n6144) );
  XNOR U7177 ( .A(b[1018]), .B(n6145), .Z(n6146) );
  XNOR U7178 ( .A(b[1018]), .B(n6147), .Z(c[1018]) );
  XNOR U7179 ( .A(a[1018]), .B(n6148), .Z(n6147) );
  IV U7180 ( .A(n6145), .Z(n6148) );
  XOR U7181 ( .A(n6149), .B(n6150), .Z(n6145) );
  ANDN U7182 ( .B(n6151), .A(n6152), .Z(n6149) );
  XNOR U7183 ( .A(b[1017]), .B(n6150), .Z(n6151) );
  XNOR U7184 ( .A(b[1017]), .B(n6152), .Z(c[1017]) );
  XNOR U7185 ( .A(a[1017]), .B(n6153), .Z(n6152) );
  IV U7186 ( .A(n6150), .Z(n6153) );
  XOR U7187 ( .A(n6154), .B(n6155), .Z(n6150) );
  ANDN U7188 ( .B(n6156), .A(n6157), .Z(n6154) );
  XNOR U7189 ( .A(b[1016]), .B(n6155), .Z(n6156) );
  XNOR U7190 ( .A(b[1016]), .B(n6157), .Z(c[1016]) );
  XNOR U7191 ( .A(a[1016]), .B(n6158), .Z(n6157) );
  IV U7192 ( .A(n6155), .Z(n6158) );
  XOR U7193 ( .A(n6159), .B(n6160), .Z(n6155) );
  ANDN U7194 ( .B(n6161), .A(n6162), .Z(n6159) );
  XNOR U7195 ( .A(b[1015]), .B(n6160), .Z(n6161) );
  XNOR U7196 ( .A(b[1015]), .B(n6162), .Z(c[1015]) );
  XNOR U7197 ( .A(a[1015]), .B(n6163), .Z(n6162) );
  IV U7198 ( .A(n6160), .Z(n6163) );
  XOR U7199 ( .A(n6164), .B(n6165), .Z(n6160) );
  ANDN U7200 ( .B(n6166), .A(n6167), .Z(n6164) );
  XNOR U7201 ( .A(b[1014]), .B(n6165), .Z(n6166) );
  XNOR U7202 ( .A(b[1014]), .B(n6167), .Z(c[1014]) );
  XNOR U7203 ( .A(a[1014]), .B(n6168), .Z(n6167) );
  IV U7204 ( .A(n6165), .Z(n6168) );
  XOR U7205 ( .A(n6169), .B(n6170), .Z(n6165) );
  ANDN U7206 ( .B(n6171), .A(n6172), .Z(n6169) );
  XNOR U7207 ( .A(b[1013]), .B(n6170), .Z(n6171) );
  XNOR U7208 ( .A(b[1013]), .B(n6172), .Z(c[1013]) );
  XNOR U7209 ( .A(a[1013]), .B(n6173), .Z(n6172) );
  IV U7210 ( .A(n6170), .Z(n6173) );
  XOR U7211 ( .A(n6174), .B(n6175), .Z(n6170) );
  ANDN U7212 ( .B(n6176), .A(n6177), .Z(n6174) );
  XNOR U7213 ( .A(b[1012]), .B(n6175), .Z(n6176) );
  XNOR U7214 ( .A(b[1012]), .B(n6177), .Z(c[1012]) );
  XNOR U7215 ( .A(a[1012]), .B(n6178), .Z(n6177) );
  IV U7216 ( .A(n6175), .Z(n6178) );
  XOR U7217 ( .A(n6179), .B(n6180), .Z(n6175) );
  ANDN U7218 ( .B(n6181), .A(n6182), .Z(n6179) );
  XNOR U7219 ( .A(b[1011]), .B(n6180), .Z(n6181) );
  XNOR U7220 ( .A(b[1011]), .B(n6182), .Z(c[1011]) );
  XNOR U7221 ( .A(a[1011]), .B(n6183), .Z(n6182) );
  IV U7222 ( .A(n6180), .Z(n6183) );
  XOR U7223 ( .A(n6184), .B(n6185), .Z(n6180) );
  ANDN U7224 ( .B(n6186), .A(n6187), .Z(n6184) );
  XNOR U7225 ( .A(b[1010]), .B(n6185), .Z(n6186) );
  XNOR U7226 ( .A(b[1010]), .B(n6187), .Z(c[1010]) );
  XNOR U7227 ( .A(a[1010]), .B(n6188), .Z(n6187) );
  IV U7228 ( .A(n6185), .Z(n6188) );
  XOR U7229 ( .A(n6189), .B(n6190), .Z(n6185) );
  ANDN U7230 ( .B(n6191), .A(n6192), .Z(n6189) );
  XNOR U7231 ( .A(b[1009]), .B(n6190), .Z(n6191) );
  XNOR U7232 ( .A(b[100]), .B(n6193), .Z(c[100]) );
  XNOR U7233 ( .A(b[1009]), .B(n6192), .Z(c[1009]) );
  XNOR U7234 ( .A(a[1009]), .B(n6194), .Z(n6192) );
  IV U7235 ( .A(n6190), .Z(n6194) );
  XOR U7236 ( .A(n6195), .B(n6196), .Z(n6190) );
  ANDN U7237 ( .B(n6197), .A(n6198), .Z(n6195) );
  XNOR U7238 ( .A(b[1008]), .B(n6196), .Z(n6197) );
  XNOR U7239 ( .A(b[1008]), .B(n6198), .Z(c[1008]) );
  XNOR U7240 ( .A(a[1008]), .B(n6199), .Z(n6198) );
  IV U7241 ( .A(n6196), .Z(n6199) );
  XOR U7242 ( .A(n6200), .B(n6201), .Z(n6196) );
  ANDN U7243 ( .B(n6202), .A(n6203), .Z(n6200) );
  XNOR U7244 ( .A(b[1007]), .B(n6201), .Z(n6202) );
  XNOR U7245 ( .A(b[1007]), .B(n6203), .Z(c[1007]) );
  XNOR U7246 ( .A(a[1007]), .B(n6204), .Z(n6203) );
  IV U7247 ( .A(n6201), .Z(n6204) );
  XOR U7248 ( .A(n6205), .B(n6206), .Z(n6201) );
  ANDN U7249 ( .B(n6207), .A(n6208), .Z(n6205) );
  XNOR U7250 ( .A(b[1006]), .B(n6206), .Z(n6207) );
  XNOR U7251 ( .A(b[1006]), .B(n6208), .Z(c[1006]) );
  XNOR U7252 ( .A(a[1006]), .B(n6209), .Z(n6208) );
  IV U7253 ( .A(n6206), .Z(n6209) );
  XOR U7254 ( .A(n6210), .B(n6211), .Z(n6206) );
  ANDN U7255 ( .B(n6212), .A(n6213), .Z(n6210) );
  XNOR U7256 ( .A(b[1005]), .B(n6211), .Z(n6212) );
  XNOR U7257 ( .A(b[1005]), .B(n6213), .Z(c[1005]) );
  XNOR U7258 ( .A(a[1005]), .B(n6214), .Z(n6213) );
  IV U7259 ( .A(n6211), .Z(n6214) );
  XOR U7260 ( .A(n6215), .B(n6216), .Z(n6211) );
  ANDN U7261 ( .B(n6217), .A(n6218), .Z(n6215) );
  XNOR U7262 ( .A(b[1004]), .B(n6216), .Z(n6217) );
  XNOR U7263 ( .A(b[1004]), .B(n6218), .Z(c[1004]) );
  XNOR U7264 ( .A(a[1004]), .B(n6219), .Z(n6218) );
  IV U7265 ( .A(n6216), .Z(n6219) );
  XOR U7266 ( .A(n6220), .B(n6221), .Z(n6216) );
  ANDN U7267 ( .B(n6222), .A(n6223), .Z(n6220) );
  XNOR U7268 ( .A(b[1003]), .B(n6221), .Z(n6222) );
  XNOR U7269 ( .A(b[1003]), .B(n6223), .Z(c[1003]) );
  XNOR U7270 ( .A(a[1003]), .B(n6224), .Z(n6223) );
  IV U7271 ( .A(n6221), .Z(n6224) );
  XOR U7272 ( .A(n6225), .B(n6226), .Z(n6221) );
  ANDN U7273 ( .B(n6227), .A(n6228), .Z(n6225) );
  XNOR U7274 ( .A(b[1002]), .B(n6226), .Z(n6227) );
  XNOR U7275 ( .A(b[1002]), .B(n6228), .Z(c[1002]) );
  XNOR U7276 ( .A(a[1002]), .B(n6229), .Z(n6228) );
  IV U7277 ( .A(n6226), .Z(n6229) );
  XOR U7278 ( .A(n6230), .B(n6231), .Z(n6226) );
  ANDN U7279 ( .B(n6232), .A(n6233), .Z(n6230) );
  XNOR U7280 ( .A(b[1001]), .B(n6231), .Z(n6232) );
  XNOR U7281 ( .A(b[1001]), .B(n6233), .Z(c[1001]) );
  XNOR U7282 ( .A(a[1001]), .B(n6234), .Z(n6233) );
  IV U7283 ( .A(n6231), .Z(n6234) );
  XOR U7284 ( .A(n6235), .B(n6236), .Z(n6231) );
  ANDN U7285 ( .B(n6237), .A(n6238), .Z(n6235) );
  XNOR U7286 ( .A(b[1000]), .B(n6236), .Z(n6237) );
  XNOR U7287 ( .A(b[1000]), .B(n6238), .Z(c[1000]) );
  XNOR U7288 ( .A(a[1000]), .B(n6239), .Z(n6238) );
  IV U7289 ( .A(n6236), .Z(n6239) );
  XOR U7290 ( .A(n6240), .B(n6241), .Z(n6236) );
  ANDN U7291 ( .B(n6242), .A(n8), .Z(n6240) );
  XNOR U7292 ( .A(a[999]), .B(n6243), .Z(n8) );
  IV U7293 ( .A(n6241), .Z(n6243) );
  XNOR U7294 ( .A(b[999]), .B(n6241), .Z(n6242) );
  XOR U7295 ( .A(n6244), .B(n6245), .Z(n6241) );
  ANDN U7296 ( .B(n6246), .A(n9), .Z(n6244) );
  XNOR U7297 ( .A(a[998]), .B(n6247), .Z(n9) );
  IV U7298 ( .A(n6245), .Z(n6247) );
  XNOR U7299 ( .A(b[998]), .B(n6245), .Z(n6246) );
  XOR U7300 ( .A(n6248), .B(n6249), .Z(n6245) );
  ANDN U7301 ( .B(n6250), .A(n10), .Z(n6248) );
  XNOR U7302 ( .A(a[997]), .B(n6251), .Z(n10) );
  IV U7303 ( .A(n6249), .Z(n6251) );
  XNOR U7304 ( .A(b[997]), .B(n6249), .Z(n6250) );
  XOR U7305 ( .A(n6252), .B(n6253), .Z(n6249) );
  ANDN U7306 ( .B(n6254), .A(n11), .Z(n6252) );
  XNOR U7307 ( .A(a[996]), .B(n6255), .Z(n11) );
  IV U7308 ( .A(n6253), .Z(n6255) );
  XNOR U7309 ( .A(b[996]), .B(n6253), .Z(n6254) );
  XOR U7310 ( .A(n6256), .B(n6257), .Z(n6253) );
  ANDN U7311 ( .B(n6258), .A(n12), .Z(n6256) );
  XNOR U7312 ( .A(a[995]), .B(n6259), .Z(n12) );
  IV U7313 ( .A(n6257), .Z(n6259) );
  XNOR U7314 ( .A(b[995]), .B(n6257), .Z(n6258) );
  XOR U7315 ( .A(n6260), .B(n6261), .Z(n6257) );
  ANDN U7316 ( .B(n6262), .A(n13), .Z(n6260) );
  XNOR U7317 ( .A(a[994]), .B(n6263), .Z(n13) );
  IV U7318 ( .A(n6261), .Z(n6263) );
  XNOR U7319 ( .A(b[994]), .B(n6261), .Z(n6262) );
  XOR U7320 ( .A(n6264), .B(n6265), .Z(n6261) );
  ANDN U7321 ( .B(n6266), .A(n14), .Z(n6264) );
  XNOR U7322 ( .A(a[993]), .B(n6267), .Z(n14) );
  IV U7323 ( .A(n6265), .Z(n6267) );
  XNOR U7324 ( .A(b[993]), .B(n6265), .Z(n6266) );
  XOR U7325 ( .A(n6268), .B(n6269), .Z(n6265) );
  ANDN U7326 ( .B(n6270), .A(n15), .Z(n6268) );
  XNOR U7327 ( .A(a[992]), .B(n6271), .Z(n15) );
  IV U7328 ( .A(n6269), .Z(n6271) );
  XNOR U7329 ( .A(b[992]), .B(n6269), .Z(n6270) );
  XOR U7330 ( .A(n6272), .B(n6273), .Z(n6269) );
  ANDN U7331 ( .B(n6274), .A(n16), .Z(n6272) );
  XNOR U7332 ( .A(a[991]), .B(n6275), .Z(n16) );
  IV U7333 ( .A(n6273), .Z(n6275) );
  XNOR U7334 ( .A(b[991]), .B(n6273), .Z(n6274) );
  XOR U7335 ( .A(n6276), .B(n6277), .Z(n6273) );
  ANDN U7336 ( .B(n6278), .A(n17), .Z(n6276) );
  XNOR U7337 ( .A(a[990]), .B(n6279), .Z(n17) );
  IV U7338 ( .A(n6277), .Z(n6279) );
  XNOR U7339 ( .A(b[990]), .B(n6277), .Z(n6278) );
  XOR U7340 ( .A(n6280), .B(n6281), .Z(n6277) );
  ANDN U7341 ( .B(n6282), .A(n19), .Z(n6280) );
  XNOR U7342 ( .A(a[989]), .B(n6283), .Z(n19) );
  IV U7343 ( .A(n6281), .Z(n6283) );
  XNOR U7344 ( .A(b[989]), .B(n6281), .Z(n6282) );
  XOR U7345 ( .A(n6284), .B(n6285), .Z(n6281) );
  ANDN U7346 ( .B(n6286), .A(n20), .Z(n6284) );
  XNOR U7347 ( .A(a[988]), .B(n6287), .Z(n20) );
  IV U7348 ( .A(n6285), .Z(n6287) );
  XNOR U7349 ( .A(b[988]), .B(n6285), .Z(n6286) );
  XOR U7350 ( .A(n6288), .B(n6289), .Z(n6285) );
  ANDN U7351 ( .B(n6290), .A(n21), .Z(n6288) );
  XNOR U7352 ( .A(a[987]), .B(n6291), .Z(n21) );
  IV U7353 ( .A(n6289), .Z(n6291) );
  XNOR U7354 ( .A(b[987]), .B(n6289), .Z(n6290) );
  XOR U7355 ( .A(n6292), .B(n6293), .Z(n6289) );
  ANDN U7356 ( .B(n6294), .A(n22), .Z(n6292) );
  XNOR U7357 ( .A(a[986]), .B(n6295), .Z(n22) );
  IV U7358 ( .A(n6293), .Z(n6295) );
  XNOR U7359 ( .A(b[986]), .B(n6293), .Z(n6294) );
  XOR U7360 ( .A(n6296), .B(n6297), .Z(n6293) );
  ANDN U7361 ( .B(n6298), .A(n23), .Z(n6296) );
  XNOR U7362 ( .A(a[985]), .B(n6299), .Z(n23) );
  IV U7363 ( .A(n6297), .Z(n6299) );
  XNOR U7364 ( .A(b[985]), .B(n6297), .Z(n6298) );
  XOR U7365 ( .A(n6300), .B(n6301), .Z(n6297) );
  ANDN U7366 ( .B(n6302), .A(n24), .Z(n6300) );
  XNOR U7367 ( .A(a[984]), .B(n6303), .Z(n24) );
  IV U7368 ( .A(n6301), .Z(n6303) );
  XNOR U7369 ( .A(b[984]), .B(n6301), .Z(n6302) );
  XOR U7370 ( .A(n6304), .B(n6305), .Z(n6301) );
  ANDN U7371 ( .B(n6306), .A(n25), .Z(n6304) );
  XNOR U7372 ( .A(a[983]), .B(n6307), .Z(n25) );
  IV U7373 ( .A(n6305), .Z(n6307) );
  XNOR U7374 ( .A(b[983]), .B(n6305), .Z(n6306) );
  XOR U7375 ( .A(n6308), .B(n6309), .Z(n6305) );
  ANDN U7376 ( .B(n6310), .A(n26), .Z(n6308) );
  XNOR U7377 ( .A(a[982]), .B(n6311), .Z(n26) );
  IV U7378 ( .A(n6309), .Z(n6311) );
  XNOR U7379 ( .A(b[982]), .B(n6309), .Z(n6310) );
  XOR U7380 ( .A(n6312), .B(n6313), .Z(n6309) );
  ANDN U7381 ( .B(n6314), .A(n27), .Z(n6312) );
  XNOR U7382 ( .A(a[981]), .B(n6315), .Z(n27) );
  IV U7383 ( .A(n6313), .Z(n6315) );
  XNOR U7384 ( .A(b[981]), .B(n6313), .Z(n6314) );
  XOR U7385 ( .A(n6316), .B(n6317), .Z(n6313) );
  ANDN U7386 ( .B(n6318), .A(n28), .Z(n6316) );
  XNOR U7387 ( .A(a[980]), .B(n6319), .Z(n28) );
  IV U7388 ( .A(n6317), .Z(n6319) );
  XNOR U7389 ( .A(b[980]), .B(n6317), .Z(n6318) );
  XOR U7390 ( .A(n6320), .B(n6321), .Z(n6317) );
  ANDN U7391 ( .B(n6322), .A(n30), .Z(n6320) );
  XNOR U7392 ( .A(a[979]), .B(n6323), .Z(n30) );
  IV U7393 ( .A(n6321), .Z(n6323) );
  XNOR U7394 ( .A(b[979]), .B(n6321), .Z(n6322) );
  XOR U7395 ( .A(n6324), .B(n6325), .Z(n6321) );
  ANDN U7396 ( .B(n6326), .A(n31), .Z(n6324) );
  XNOR U7397 ( .A(a[978]), .B(n6327), .Z(n31) );
  IV U7398 ( .A(n6325), .Z(n6327) );
  XNOR U7399 ( .A(b[978]), .B(n6325), .Z(n6326) );
  XOR U7400 ( .A(n6328), .B(n6329), .Z(n6325) );
  ANDN U7401 ( .B(n6330), .A(n32), .Z(n6328) );
  XNOR U7402 ( .A(a[977]), .B(n6331), .Z(n32) );
  IV U7403 ( .A(n6329), .Z(n6331) );
  XNOR U7404 ( .A(b[977]), .B(n6329), .Z(n6330) );
  XOR U7405 ( .A(n6332), .B(n6333), .Z(n6329) );
  ANDN U7406 ( .B(n6334), .A(n33), .Z(n6332) );
  XNOR U7407 ( .A(a[976]), .B(n6335), .Z(n33) );
  IV U7408 ( .A(n6333), .Z(n6335) );
  XNOR U7409 ( .A(b[976]), .B(n6333), .Z(n6334) );
  XOR U7410 ( .A(n6336), .B(n6337), .Z(n6333) );
  ANDN U7411 ( .B(n6338), .A(n34), .Z(n6336) );
  XNOR U7412 ( .A(a[975]), .B(n6339), .Z(n34) );
  IV U7413 ( .A(n6337), .Z(n6339) );
  XNOR U7414 ( .A(b[975]), .B(n6337), .Z(n6338) );
  XOR U7415 ( .A(n6340), .B(n6341), .Z(n6337) );
  ANDN U7416 ( .B(n6342), .A(n35), .Z(n6340) );
  XNOR U7417 ( .A(a[974]), .B(n6343), .Z(n35) );
  IV U7418 ( .A(n6341), .Z(n6343) );
  XNOR U7419 ( .A(b[974]), .B(n6341), .Z(n6342) );
  XOR U7420 ( .A(n6344), .B(n6345), .Z(n6341) );
  ANDN U7421 ( .B(n6346), .A(n36), .Z(n6344) );
  XNOR U7422 ( .A(a[973]), .B(n6347), .Z(n36) );
  IV U7423 ( .A(n6345), .Z(n6347) );
  XNOR U7424 ( .A(b[973]), .B(n6345), .Z(n6346) );
  XOR U7425 ( .A(n6348), .B(n6349), .Z(n6345) );
  ANDN U7426 ( .B(n6350), .A(n37), .Z(n6348) );
  XNOR U7427 ( .A(a[972]), .B(n6351), .Z(n37) );
  IV U7428 ( .A(n6349), .Z(n6351) );
  XNOR U7429 ( .A(b[972]), .B(n6349), .Z(n6350) );
  XOR U7430 ( .A(n6352), .B(n6353), .Z(n6349) );
  ANDN U7431 ( .B(n6354), .A(n38), .Z(n6352) );
  XNOR U7432 ( .A(a[971]), .B(n6355), .Z(n38) );
  IV U7433 ( .A(n6353), .Z(n6355) );
  XNOR U7434 ( .A(b[971]), .B(n6353), .Z(n6354) );
  XOR U7435 ( .A(n6356), .B(n6357), .Z(n6353) );
  ANDN U7436 ( .B(n6358), .A(n39), .Z(n6356) );
  XNOR U7437 ( .A(a[970]), .B(n6359), .Z(n39) );
  IV U7438 ( .A(n6357), .Z(n6359) );
  XNOR U7439 ( .A(b[970]), .B(n6357), .Z(n6358) );
  XOR U7440 ( .A(n6360), .B(n6361), .Z(n6357) );
  ANDN U7441 ( .B(n6362), .A(n41), .Z(n6360) );
  XNOR U7442 ( .A(a[969]), .B(n6363), .Z(n41) );
  IV U7443 ( .A(n6361), .Z(n6363) );
  XNOR U7444 ( .A(b[969]), .B(n6361), .Z(n6362) );
  XOR U7445 ( .A(n6364), .B(n6365), .Z(n6361) );
  ANDN U7446 ( .B(n6366), .A(n42), .Z(n6364) );
  XNOR U7447 ( .A(a[968]), .B(n6367), .Z(n42) );
  IV U7448 ( .A(n6365), .Z(n6367) );
  XNOR U7449 ( .A(b[968]), .B(n6365), .Z(n6366) );
  XOR U7450 ( .A(n6368), .B(n6369), .Z(n6365) );
  ANDN U7451 ( .B(n6370), .A(n43), .Z(n6368) );
  XNOR U7452 ( .A(a[967]), .B(n6371), .Z(n43) );
  IV U7453 ( .A(n6369), .Z(n6371) );
  XNOR U7454 ( .A(b[967]), .B(n6369), .Z(n6370) );
  XOR U7455 ( .A(n6372), .B(n6373), .Z(n6369) );
  ANDN U7456 ( .B(n6374), .A(n44), .Z(n6372) );
  XNOR U7457 ( .A(a[966]), .B(n6375), .Z(n44) );
  IV U7458 ( .A(n6373), .Z(n6375) );
  XNOR U7459 ( .A(b[966]), .B(n6373), .Z(n6374) );
  XOR U7460 ( .A(n6376), .B(n6377), .Z(n6373) );
  ANDN U7461 ( .B(n6378), .A(n45), .Z(n6376) );
  XNOR U7462 ( .A(a[965]), .B(n6379), .Z(n45) );
  IV U7463 ( .A(n6377), .Z(n6379) );
  XNOR U7464 ( .A(b[965]), .B(n6377), .Z(n6378) );
  XOR U7465 ( .A(n6380), .B(n6381), .Z(n6377) );
  ANDN U7466 ( .B(n6382), .A(n46), .Z(n6380) );
  XNOR U7467 ( .A(a[964]), .B(n6383), .Z(n46) );
  IV U7468 ( .A(n6381), .Z(n6383) );
  XNOR U7469 ( .A(b[964]), .B(n6381), .Z(n6382) );
  XOR U7470 ( .A(n6384), .B(n6385), .Z(n6381) );
  ANDN U7471 ( .B(n6386), .A(n47), .Z(n6384) );
  XNOR U7472 ( .A(a[963]), .B(n6387), .Z(n47) );
  IV U7473 ( .A(n6385), .Z(n6387) );
  XNOR U7474 ( .A(b[963]), .B(n6385), .Z(n6386) );
  XOR U7475 ( .A(n6388), .B(n6389), .Z(n6385) );
  ANDN U7476 ( .B(n6390), .A(n48), .Z(n6388) );
  XNOR U7477 ( .A(a[962]), .B(n6391), .Z(n48) );
  IV U7478 ( .A(n6389), .Z(n6391) );
  XNOR U7479 ( .A(b[962]), .B(n6389), .Z(n6390) );
  XOR U7480 ( .A(n6392), .B(n6393), .Z(n6389) );
  ANDN U7481 ( .B(n6394), .A(n49), .Z(n6392) );
  XNOR U7482 ( .A(a[961]), .B(n6395), .Z(n49) );
  IV U7483 ( .A(n6393), .Z(n6395) );
  XNOR U7484 ( .A(b[961]), .B(n6393), .Z(n6394) );
  XOR U7485 ( .A(n6396), .B(n6397), .Z(n6393) );
  ANDN U7486 ( .B(n6398), .A(n50), .Z(n6396) );
  XNOR U7487 ( .A(a[960]), .B(n6399), .Z(n50) );
  IV U7488 ( .A(n6397), .Z(n6399) );
  XNOR U7489 ( .A(b[960]), .B(n6397), .Z(n6398) );
  XOR U7490 ( .A(n6400), .B(n6401), .Z(n6397) );
  ANDN U7491 ( .B(n6402), .A(n52), .Z(n6400) );
  XNOR U7492 ( .A(a[959]), .B(n6403), .Z(n52) );
  IV U7493 ( .A(n6401), .Z(n6403) );
  XNOR U7494 ( .A(b[959]), .B(n6401), .Z(n6402) );
  XOR U7495 ( .A(n6404), .B(n6405), .Z(n6401) );
  ANDN U7496 ( .B(n6406), .A(n53), .Z(n6404) );
  XNOR U7497 ( .A(a[958]), .B(n6407), .Z(n53) );
  IV U7498 ( .A(n6405), .Z(n6407) );
  XNOR U7499 ( .A(b[958]), .B(n6405), .Z(n6406) );
  XOR U7500 ( .A(n6408), .B(n6409), .Z(n6405) );
  ANDN U7501 ( .B(n6410), .A(n54), .Z(n6408) );
  XNOR U7502 ( .A(a[957]), .B(n6411), .Z(n54) );
  IV U7503 ( .A(n6409), .Z(n6411) );
  XNOR U7504 ( .A(b[957]), .B(n6409), .Z(n6410) );
  XOR U7505 ( .A(n6412), .B(n6413), .Z(n6409) );
  ANDN U7506 ( .B(n6414), .A(n55), .Z(n6412) );
  XNOR U7507 ( .A(a[956]), .B(n6415), .Z(n55) );
  IV U7508 ( .A(n6413), .Z(n6415) );
  XNOR U7509 ( .A(b[956]), .B(n6413), .Z(n6414) );
  XOR U7510 ( .A(n6416), .B(n6417), .Z(n6413) );
  ANDN U7511 ( .B(n6418), .A(n56), .Z(n6416) );
  XNOR U7512 ( .A(a[955]), .B(n6419), .Z(n56) );
  IV U7513 ( .A(n6417), .Z(n6419) );
  XNOR U7514 ( .A(b[955]), .B(n6417), .Z(n6418) );
  XOR U7515 ( .A(n6420), .B(n6421), .Z(n6417) );
  ANDN U7516 ( .B(n6422), .A(n57), .Z(n6420) );
  XNOR U7517 ( .A(a[954]), .B(n6423), .Z(n57) );
  IV U7518 ( .A(n6421), .Z(n6423) );
  XNOR U7519 ( .A(b[954]), .B(n6421), .Z(n6422) );
  XOR U7520 ( .A(n6424), .B(n6425), .Z(n6421) );
  ANDN U7521 ( .B(n6426), .A(n58), .Z(n6424) );
  XNOR U7522 ( .A(a[953]), .B(n6427), .Z(n58) );
  IV U7523 ( .A(n6425), .Z(n6427) );
  XNOR U7524 ( .A(b[953]), .B(n6425), .Z(n6426) );
  XOR U7525 ( .A(n6428), .B(n6429), .Z(n6425) );
  ANDN U7526 ( .B(n6430), .A(n59), .Z(n6428) );
  XNOR U7527 ( .A(a[952]), .B(n6431), .Z(n59) );
  IV U7528 ( .A(n6429), .Z(n6431) );
  XNOR U7529 ( .A(b[952]), .B(n6429), .Z(n6430) );
  XOR U7530 ( .A(n6432), .B(n6433), .Z(n6429) );
  ANDN U7531 ( .B(n6434), .A(n60), .Z(n6432) );
  XNOR U7532 ( .A(a[951]), .B(n6435), .Z(n60) );
  IV U7533 ( .A(n6433), .Z(n6435) );
  XNOR U7534 ( .A(b[951]), .B(n6433), .Z(n6434) );
  XOR U7535 ( .A(n6436), .B(n6437), .Z(n6433) );
  ANDN U7536 ( .B(n6438), .A(n61), .Z(n6436) );
  XNOR U7537 ( .A(a[950]), .B(n6439), .Z(n61) );
  IV U7538 ( .A(n6437), .Z(n6439) );
  XNOR U7539 ( .A(b[950]), .B(n6437), .Z(n6438) );
  XOR U7540 ( .A(n6440), .B(n6441), .Z(n6437) );
  ANDN U7541 ( .B(n6442), .A(n63), .Z(n6440) );
  XNOR U7542 ( .A(a[949]), .B(n6443), .Z(n63) );
  IV U7543 ( .A(n6441), .Z(n6443) );
  XNOR U7544 ( .A(b[949]), .B(n6441), .Z(n6442) );
  XOR U7545 ( .A(n6444), .B(n6445), .Z(n6441) );
  ANDN U7546 ( .B(n6446), .A(n64), .Z(n6444) );
  XNOR U7547 ( .A(a[948]), .B(n6447), .Z(n64) );
  IV U7548 ( .A(n6445), .Z(n6447) );
  XNOR U7549 ( .A(b[948]), .B(n6445), .Z(n6446) );
  XOR U7550 ( .A(n6448), .B(n6449), .Z(n6445) );
  ANDN U7551 ( .B(n6450), .A(n65), .Z(n6448) );
  XNOR U7552 ( .A(a[947]), .B(n6451), .Z(n65) );
  IV U7553 ( .A(n6449), .Z(n6451) );
  XNOR U7554 ( .A(b[947]), .B(n6449), .Z(n6450) );
  XOR U7555 ( .A(n6452), .B(n6453), .Z(n6449) );
  ANDN U7556 ( .B(n6454), .A(n66), .Z(n6452) );
  XNOR U7557 ( .A(a[946]), .B(n6455), .Z(n66) );
  IV U7558 ( .A(n6453), .Z(n6455) );
  XNOR U7559 ( .A(b[946]), .B(n6453), .Z(n6454) );
  XOR U7560 ( .A(n6456), .B(n6457), .Z(n6453) );
  ANDN U7561 ( .B(n6458), .A(n67), .Z(n6456) );
  XNOR U7562 ( .A(a[945]), .B(n6459), .Z(n67) );
  IV U7563 ( .A(n6457), .Z(n6459) );
  XNOR U7564 ( .A(b[945]), .B(n6457), .Z(n6458) );
  XOR U7565 ( .A(n6460), .B(n6461), .Z(n6457) );
  ANDN U7566 ( .B(n6462), .A(n68), .Z(n6460) );
  XNOR U7567 ( .A(a[944]), .B(n6463), .Z(n68) );
  IV U7568 ( .A(n6461), .Z(n6463) );
  XNOR U7569 ( .A(b[944]), .B(n6461), .Z(n6462) );
  XOR U7570 ( .A(n6464), .B(n6465), .Z(n6461) );
  ANDN U7571 ( .B(n6466), .A(n69), .Z(n6464) );
  XNOR U7572 ( .A(a[943]), .B(n6467), .Z(n69) );
  IV U7573 ( .A(n6465), .Z(n6467) );
  XNOR U7574 ( .A(b[943]), .B(n6465), .Z(n6466) );
  XOR U7575 ( .A(n6468), .B(n6469), .Z(n6465) );
  ANDN U7576 ( .B(n6470), .A(n70), .Z(n6468) );
  XNOR U7577 ( .A(a[942]), .B(n6471), .Z(n70) );
  IV U7578 ( .A(n6469), .Z(n6471) );
  XNOR U7579 ( .A(b[942]), .B(n6469), .Z(n6470) );
  XOR U7580 ( .A(n6472), .B(n6473), .Z(n6469) );
  ANDN U7581 ( .B(n6474), .A(n71), .Z(n6472) );
  XNOR U7582 ( .A(a[941]), .B(n6475), .Z(n71) );
  IV U7583 ( .A(n6473), .Z(n6475) );
  XNOR U7584 ( .A(b[941]), .B(n6473), .Z(n6474) );
  XOR U7585 ( .A(n6476), .B(n6477), .Z(n6473) );
  ANDN U7586 ( .B(n6478), .A(n72), .Z(n6476) );
  XNOR U7587 ( .A(a[940]), .B(n6479), .Z(n72) );
  IV U7588 ( .A(n6477), .Z(n6479) );
  XNOR U7589 ( .A(b[940]), .B(n6477), .Z(n6478) );
  XOR U7590 ( .A(n6480), .B(n6481), .Z(n6477) );
  ANDN U7591 ( .B(n6482), .A(n74), .Z(n6480) );
  XNOR U7592 ( .A(a[939]), .B(n6483), .Z(n74) );
  IV U7593 ( .A(n6481), .Z(n6483) );
  XNOR U7594 ( .A(b[939]), .B(n6481), .Z(n6482) );
  XOR U7595 ( .A(n6484), .B(n6485), .Z(n6481) );
  ANDN U7596 ( .B(n6486), .A(n75), .Z(n6484) );
  XNOR U7597 ( .A(a[938]), .B(n6487), .Z(n75) );
  IV U7598 ( .A(n6485), .Z(n6487) );
  XNOR U7599 ( .A(b[938]), .B(n6485), .Z(n6486) );
  XOR U7600 ( .A(n6488), .B(n6489), .Z(n6485) );
  ANDN U7601 ( .B(n6490), .A(n76), .Z(n6488) );
  XNOR U7602 ( .A(a[937]), .B(n6491), .Z(n76) );
  IV U7603 ( .A(n6489), .Z(n6491) );
  XNOR U7604 ( .A(b[937]), .B(n6489), .Z(n6490) );
  XOR U7605 ( .A(n6492), .B(n6493), .Z(n6489) );
  ANDN U7606 ( .B(n6494), .A(n77), .Z(n6492) );
  XNOR U7607 ( .A(a[936]), .B(n6495), .Z(n77) );
  IV U7608 ( .A(n6493), .Z(n6495) );
  XNOR U7609 ( .A(b[936]), .B(n6493), .Z(n6494) );
  XOR U7610 ( .A(n6496), .B(n6497), .Z(n6493) );
  ANDN U7611 ( .B(n6498), .A(n78), .Z(n6496) );
  XNOR U7612 ( .A(a[935]), .B(n6499), .Z(n78) );
  IV U7613 ( .A(n6497), .Z(n6499) );
  XNOR U7614 ( .A(b[935]), .B(n6497), .Z(n6498) );
  XOR U7615 ( .A(n6500), .B(n6501), .Z(n6497) );
  ANDN U7616 ( .B(n6502), .A(n79), .Z(n6500) );
  XNOR U7617 ( .A(a[934]), .B(n6503), .Z(n79) );
  IV U7618 ( .A(n6501), .Z(n6503) );
  XNOR U7619 ( .A(b[934]), .B(n6501), .Z(n6502) );
  XOR U7620 ( .A(n6504), .B(n6505), .Z(n6501) );
  ANDN U7621 ( .B(n6506), .A(n80), .Z(n6504) );
  XNOR U7622 ( .A(a[933]), .B(n6507), .Z(n80) );
  IV U7623 ( .A(n6505), .Z(n6507) );
  XNOR U7624 ( .A(b[933]), .B(n6505), .Z(n6506) );
  XOR U7625 ( .A(n6508), .B(n6509), .Z(n6505) );
  ANDN U7626 ( .B(n6510), .A(n81), .Z(n6508) );
  XNOR U7627 ( .A(a[932]), .B(n6511), .Z(n81) );
  IV U7628 ( .A(n6509), .Z(n6511) );
  XNOR U7629 ( .A(b[932]), .B(n6509), .Z(n6510) );
  XOR U7630 ( .A(n6512), .B(n6513), .Z(n6509) );
  ANDN U7631 ( .B(n6514), .A(n82), .Z(n6512) );
  XNOR U7632 ( .A(a[931]), .B(n6515), .Z(n82) );
  IV U7633 ( .A(n6513), .Z(n6515) );
  XNOR U7634 ( .A(b[931]), .B(n6513), .Z(n6514) );
  XOR U7635 ( .A(n6516), .B(n6517), .Z(n6513) );
  ANDN U7636 ( .B(n6518), .A(n83), .Z(n6516) );
  XNOR U7637 ( .A(a[930]), .B(n6519), .Z(n83) );
  IV U7638 ( .A(n6517), .Z(n6519) );
  XNOR U7639 ( .A(b[930]), .B(n6517), .Z(n6518) );
  XOR U7640 ( .A(n6520), .B(n6521), .Z(n6517) );
  ANDN U7641 ( .B(n6522), .A(n85), .Z(n6520) );
  XNOR U7642 ( .A(a[929]), .B(n6523), .Z(n85) );
  IV U7643 ( .A(n6521), .Z(n6523) );
  XNOR U7644 ( .A(b[929]), .B(n6521), .Z(n6522) );
  XOR U7645 ( .A(n6524), .B(n6525), .Z(n6521) );
  ANDN U7646 ( .B(n6526), .A(n86), .Z(n6524) );
  XNOR U7647 ( .A(a[928]), .B(n6527), .Z(n86) );
  IV U7648 ( .A(n6525), .Z(n6527) );
  XNOR U7649 ( .A(b[928]), .B(n6525), .Z(n6526) );
  XOR U7650 ( .A(n6528), .B(n6529), .Z(n6525) );
  ANDN U7651 ( .B(n6530), .A(n87), .Z(n6528) );
  XNOR U7652 ( .A(a[927]), .B(n6531), .Z(n87) );
  IV U7653 ( .A(n6529), .Z(n6531) );
  XNOR U7654 ( .A(b[927]), .B(n6529), .Z(n6530) );
  XOR U7655 ( .A(n6532), .B(n6533), .Z(n6529) );
  ANDN U7656 ( .B(n6534), .A(n88), .Z(n6532) );
  XNOR U7657 ( .A(a[926]), .B(n6535), .Z(n88) );
  IV U7658 ( .A(n6533), .Z(n6535) );
  XNOR U7659 ( .A(b[926]), .B(n6533), .Z(n6534) );
  XOR U7660 ( .A(n6536), .B(n6537), .Z(n6533) );
  ANDN U7661 ( .B(n6538), .A(n89), .Z(n6536) );
  XNOR U7662 ( .A(a[925]), .B(n6539), .Z(n89) );
  IV U7663 ( .A(n6537), .Z(n6539) );
  XNOR U7664 ( .A(b[925]), .B(n6537), .Z(n6538) );
  XOR U7665 ( .A(n6540), .B(n6541), .Z(n6537) );
  ANDN U7666 ( .B(n6542), .A(n90), .Z(n6540) );
  XNOR U7667 ( .A(a[924]), .B(n6543), .Z(n90) );
  IV U7668 ( .A(n6541), .Z(n6543) );
  XNOR U7669 ( .A(b[924]), .B(n6541), .Z(n6542) );
  XOR U7670 ( .A(n6544), .B(n6545), .Z(n6541) );
  ANDN U7671 ( .B(n6546), .A(n91), .Z(n6544) );
  XNOR U7672 ( .A(a[923]), .B(n6547), .Z(n91) );
  IV U7673 ( .A(n6545), .Z(n6547) );
  XNOR U7674 ( .A(b[923]), .B(n6545), .Z(n6546) );
  XOR U7675 ( .A(n6548), .B(n6549), .Z(n6545) );
  ANDN U7676 ( .B(n6550), .A(n92), .Z(n6548) );
  XNOR U7677 ( .A(a[922]), .B(n6551), .Z(n92) );
  IV U7678 ( .A(n6549), .Z(n6551) );
  XNOR U7679 ( .A(b[922]), .B(n6549), .Z(n6550) );
  XOR U7680 ( .A(n6552), .B(n6553), .Z(n6549) );
  ANDN U7681 ( .B(n6554), .A(n93), .Z(n6552) );
  XNOR U7682 ( .A(a[921]), .B(n6555), .Z(n93) );
  IV U7683 ( .A(n6553), .Z(n6555) );
  XNOR U7684 ( .A(b[921]), .B(n6553), .Z(n6554) );
  XOR U7685 ( .A(n6556), .B(n6557), .Z(n6553) );
  ANDN U7686 ( .B(n6558), .A(n94), .Z(n6556) );
  XNOR U7687 ( .A(a[920]), .B(n6559), .Z(n94) );
  IV U7688 ( .A(n6557), .Z(n6559) );
  XNOR U7689 ( .A(b[920]), .B(n6557), .Z(n6558) );
  XOR U7690 ( .A(n6560), .B(n6561), .Z(n6557) );
  ANDN U7691 ( .B(n6562), .A(n96), .Z(n6560) );
  XNOR U7692 ( .A(a[919]), .B(n6563), .Z(n96) );
  IV U7693 ( .A(n6561), .Z(n6563) );
  XNOR U7694 ( .A(b[919]), .B(n6561), .Z(n6562) );
  XOR U7695 ( .A(n6564), .B(n6565), .Z(n6561) );
  ANDN U7696 ( .B(n6566), .A(n97), .Z(n6564) );
  XNOR U7697 ( .A(a[918]), .B(n6567), .Z(n97) );
  IV U7698 ( .A(n6565), .Z(n6567) );
  XNOR U7699 ( .A(b[918]), .B(n6565), .Z(n6566) );
  XOR U7700 ( .A(n6568), .B(n6569), .Z(n6565) );
  ANDN U7701 ( .B(n6570), .A(n98), .Z(n6568) );
  XNOR U7702 ( .A(a[917]), .B(n6571), .Z(n98) );
  IV U7703 ( .A(n6569), .Z(n6571) );
  XNOR U7704 ( .A(b[917]), .B(n6569), .Z(n6570) );
  XOR U7705 ( .A(n6572), .B(n6573), .Z(n6569) );
  ANDN U7706 ( .B(n6574), .A(n99), .Z(n6572) );
  XNOR U7707 ( .A(a[916]), .B(n6575), .Z(n99) );
  IV U7708 ( .A(n6573), .Z(n6575) );
  XNOR U7709 ( .A(b[916]), .B(n6573), .Z(n6574) );
  XOR U7710 ( .A(n6576), .B(n6577), .Z(n6573) );
  ANDN U7711 ( .B(n6578), .A(n100), .Z(n6576) );
  XNOR U7712 ( .A(a[915]), .B(n6579), .Z(n100) );
  IV U7713 ( .A(n6577), .Z(n6579) );
  XNOR U7714 ( .A(b[915]), .B(n6577), .Z(n6578) );
  XOR U7715 ( .A(n6580), .B(n6581), .Z(n6577) );
  ANDN U7716 ( .B(n6582), .A(n101), .Z(n6580) );
  XNOR U7717 ( .A(a[914]), .B(n6583), .Z(n101) );
  IV U7718 ( .A(n6581), .Z(n6583) );
  XNOR U7719 ( .A(b[914]), .B(n6581), .Z(n6582) );
  XOR U7720 ( .A(n6584), .B(n6585), .Z(n6581) );
  ANDN U7721 ( .B(n6586), .A(n102), .Z(n6584) );
  XNOR U7722 ( .A(a[913]), .B(n6587), .Z(n102) );
  IV U7723 ( .A(n6585), .Z(n6587) );
  XNOR U7724 ( .A(b[913]), .B(n6585), .Z(n6586) );
  XOR U7725 ( .A(n6588), .B(n6589), .Z(n6585) );
  ANDN U7726 ( .B(n6590), .A(n103), .Z(n6588) );
  XNOR U7727 ( .A(a[912]), .B(n6591), .Z(n103) );
  IV U7728 ( .A(n6589), .Z(n6591) );
  XNOR U7729 ( .A(b[912]), .B(n6589), .Z(n6590) );
  XOR U7730 ( .A(n6592), .B(n6593), .Z(n6589) );
  ANDN U7731 ( .B(n6594), .A(n104), .Z(n6592) );
  XNOR U7732 ( .A(a[911]), .B(n6595), .Z(n104) );
  IV U7733 ( .A(n6593), .Z(n6595) );
  XNOR U7734 ( .A(b[911]), .B(n6593), .Z(n6594) );
  XOR U7735 ( .A(n6596), .B(n6597), .Z(n6593) );
  ANDN U7736 ( .B(n6598), .A(n105), .Z(n6596) );
  XNOR U7737 ( .A(a[910]), .B(n6599), .Z(n105) );
  IV U7738 ( .A(n6597), .Z(n6599) );
  XNOR U7739 ( .A(b[910]), .B(n6597), .Z(n6598) );
  XOR U7740 ( .A(n6600), .B(n6601), .Z(n6597) );
  ANDN U7741 ( .B(n6602), .A(n107), .Z(n6600) );
  XNOR U7742 ( .A(a[909]), .B(n6603), .Z(n107) );
  IV U7743 ( .A(n6601), .Z(n6603) );
  XNOR U7744 ( .A(b[909]), .B(n6601), .Z(n6602) );
  XOR U7745 ( .A(n6604), .B(n6605), .Z(n6601) );
  ANDN U7746 ( .B(n6606), .A(n108), .Z(n6604) );
  XNOR U7747 ( .A(a[908]), .B(n6607), .Z(n108) );
  IV U7748 ( .A(n6605), .Z(n6607) );
  XNOR U7749 ( .A(b[908]), .B(n6605), .Z(n6606) );
  XOR U7750 ( .A(n6608), .B(n6609), .Z(n6605) );
  ANDN U7751 ( .B(n6610), .A(n109), .Z(n6608) );
  XNOR U7752 ( .A(a[907]), .B(n6611), .Z(n109) );
  IV U7753 ( .A(n6609), .Z(n6611) );
  XNOR U7754 ( .A(b[907]), .B(n6609), .Z(n6610) );
  XOR U7755 ( .A(n6612), .B(n6613), .Z(n6609) );
  ANDN U7756 ( .B(n6614), .A(n110), .Z(n6612) );
  XNOR U7757 ( .A(a[906]), .B(n6615), .Z(n110) );
  IV U7758 ( .A(n6613), .Z(n6615) );
  XNOR U7759 ( .A(b[906]), .B(n6613), .Z(n6614) );
  XOR U7760 ( .A(n6616), .B(n6617), .Z(n6613) );
  ANDN U7761 ( .B(n6618), .A(n111), .Z(n6616) );
  XNOR U7762 ( .A(a[905]), .B(n6619), .Z(n111) );
  IV U7763 ( .A(n6617), .Z(n6619) );
  XNOR U7764 ( .A(b[905]), .B(n6617), .Z(n6618) );
  XOR U7765 ( .A(n6620), .B(n6621), .Z(n6617) );
  ANDN U7766 ( .B(n6622), .A(n112), .Z(n6620) );
  XNOR U7767 ( .A(a[904]), .B(n6623), .Z(n112) );
  IV U7768 ( .A(n6621), .Z(n6623) );
  XNOR U7769 ( .A(b[904]), .B(n6621), .Z(n6622) );
  XOR U7770 ( .A(n6624), .B(n6625), .Z(n6621) );
  ANDN U7771 ( .B(n6626), .A(n113), .Z(n6624) );
  XNOR U7772 ( .A(a[903]), .B(n6627), .Z(n113) );
  IV U7773 ( .A(n6625), .Z(n6627) );
  XNOR U7774 ( .A(b[903]), .B(n6625), .Z(n6626) );
  XOR U7775 ( .A(n6628), .B(n6629), .Z(n6625) );
  ANDN U7776 ( .B(n6630), .A(n114), .Z(n6628) );
  XNOR U7777 ( .A(a[902]), .B(n6631), .Z(n114) );
  IV U7778 ( .A(n6629), .Z(n6631) );
  XNOR U7779 ( .A(b[902]), .B(n6629), .Z(n6630) );
  XOR U7780 ( .A(n6632), .B(n6633), .Z(n6629) );
  ANDN U7781 ( .B(n6634), .A(n115), .Z(n6632) );
  XNOR U7782 ( .A(a[901]), .B(n6635), .Z(n115) );
  IV U7783 ( .A(n6633), .Z(n6635) );
  XNOR U7784 ( .A(b[901]), .B(n6633), .Z(n6634) );
  XOR U7785 ( .A(n6636), .B(n6637), .Z(n6633) );
  ANDN U7786 ( .B(n6638), .A(n116), .Z(n6636) );
  XNOR U7787 ( .A(a[900]), .B(n6639), .Z(n116) );
  IV U7788 ( .A(n6637), .Z(n6639) );
  XNOR U7789 ( .A(b[900]), .B(n6637), .Z(n6638) );
  XOR U7790 ( .A(n6640), .B(n6641), .Z(n6637) );
  ANDN U7791 ( .B(n6642), .A(n119), .Z(n6640) );
  XNOR U7792 ( .A(a[899]), .B(n6643), .Z(n119) );
  IV U7793 ( .A(n6641), .Z(n6643) );
  XNOR U7794 ( .A(b[899]), .B(n6641), .Z(n6642) );
  XOR U7795 ( .A(n6644), .B(n6645), .Z(n6641) );
  ANDN U7796 ( .B(n6646), .A(n120), .Z(n6644) );
  XNOR U7797 ( .A(a[898]), .B(n6647), .Z(n120) );
  IV U7798 ( .A(n6645), .Z(n6647) );
  XNOR U7799 ( .A(b[898]), .B(n6645), .Z(n6646) );
  XOR U7800 ( .A(n6648), .B(n6649), .Z(n6645) );
  ANDN U7801 ( .B(n6650), .A(n121), .Z(n6648) );
  XNOR U7802 ( .A(a[897]), .B(n6651), .Z(n121) );
  IV U7803 ( .A(n6649), .Z(n6651) );
  XNOR U7804 ( .A(b[897]), .B(n6649), .Z(n6650) );
  XOR U7805 ( .A(n6652), .B(n6653), .Z(n6649) );
  ANDN U7806 ( .B(n6654), .A(n122), .Z(n6652) );
  XNOR U7807 ( .A(a[896]), .B(n6655), .Z(n122) );
  IV U7808 ( .A(n6653), .Z(n6655) );
  XNOR U7809 ( .A(b[896]), .B(n6653), .Z(n6654) );
  XOR U7810 ( .A(n6656), .B(n6657), .Z(n6653) );
  ANDN U7811 ( .B(n6658), .A(n123), .Z(n6656) );
  XNOR U7812 ( .A(a[895]), .B(n6659), .Z(n123) );
  IV U7813 ( .A(n6657), .Z(n6659) );
  XNOR U7814 ( .A(b[895]), .B(n6657), .Z(n6658) );
  XOR U7815 ( .A(n6660), .B(n6661), .Z(n6657) );
  ANDN U7816 ( .B(n6662), .A(n124), .Z(n6660) );
  XNOR U7817 ( .A(a[894]), .B(n6663), .Z(n124) );
  IV U7818 ( .A(n6661), .Z(n6663) );
  XNOR U7819 ( .A(b[894]), .B(n6661), .Z(n6662) );
  XOR U7820 ( .A(n6664), .B(n6665), .Z(n6661) );
  ANDN U7821 ( .B(n6666), .A(n125), .Z(n6664) );
  XNOR U7822 ( .A(a[893]), .B(n6667), .Z(n125) );
  IV U7823 ( .A(n6665), .Z(n6667) );
  XNOR U7824 ( .A(b[893]), .B(n6665), .Z(n6666) );
  XOR U7825 ( .A(n6668), .B(n6669), .Z(n6665) );
  ANDN U7826 ( .B(n6670), .A(n126), .Z(n6668) );
  XNOR U7827 ( .A(a[892]), .B(n6671), .Z(n126) );
  IV U7828 ( .A(n6669), .Z(n6671) );
  XNOR U7829 ( .A(b[892]), .B(n6669), .Z(n6670) );
  XOR U7830 ( .A(n6672), .B(n6673), .Z(n6669) );
  ANDN U7831 ( .B(n6674), .A(n127), .Z(n6672) );
  XNOR U7832 ( .A(a[891]), .B(n6675), .Z(n127) );
  IV U7833 ( .A(n6673), .Z(n6675) );
  XNOR U7834 ( .A(b[891]), .B(n6673), .Z(n6674) );
  XOR U7835 ( .A(n6676), .B(n6677), .Z(n6673) );
  ANDN U7836 ( .B(n6678), .A(n128), .Z(n6676) );
  XNOR U7837 ( .A(a[890]), .B(n6679), .Z(n128) );
  IV U7838 ( .A(n6677), .Z(n6679) );
  XNOR U7839 ( .A(b[890]), .B(n6677), .Z(n6678) );
  XOR U7840 ( .A(n6680), .B(n6681), .Z(n6677) );
  ANDN U7841 ( .B(n6682), .A(n130), .Z(n6680) );
  XNOR U7842 ( .A(a[889]), .B(n6683), .Z(n130) );
  IV U7843 ( .A(n6681), .Z(n6683) );
  XNOR U7844 ( .A(b[889]), .B(n6681), .Z(n6682) );
  XOR U7845 ( .A(n6684), .B(n6685), .Z(n6681) );
  ANDN U7846 ( .B(n6686), .A(n131), .Z(n6684) );
  XNOR U7847 ( .A(a[888]), .B(n6687), .Z(n131) );
  IV U7848 ( .A(n6685), .Z(n6687) );
  XNOR U7849 ( .A(b[888]), .B(n6685), .Z(n6686) );
  XOR U7850 ( .A(n6688), .B(n6689), .Z(n6685) );
  ANDN U7851 ( .B(n6690), .A(n132), .Z(n6688) );
  XNOR U7852 ( .A(a[887]), .B(n6691), .Z(n132) );
  IV U7853 ( .A(n6689), .Z(n6691) );
  XNOR U7854 ( .A(b[887]), .B(n6689), .Z(n6690) );
  XOR U7855 ( .A(n6692), .B(n6693), .Z(n6689) );
  ANDN U7856 ( .B(n6694), .A(n133), .Z(n6692) );
  XNOR U7857 ( .A(a[886]), .B(n6695), .Z(n133) );
  IV U7858 ( .A(n6693), .Z(n6695) );
  XNOR U7859 ( .A(b[886]), .B(n6693), .Z(n6694) );
  XOR U7860 ( .A(n6696), .B(n6697), .Z(n6693) );
  ANDN U7861 ( .B(n6698), .A(n134), .Z(n6696) );
  XNOR U7862 ( .A(a[885]), .B(n6699), .Z(n134) );
  IV U7863 ( .A(n6697), .Z(n6699) );
  XNOR U7864 ( .A(b[885]), .B(n6697), .Z(n6698) );
  XOR U7865 ( .A(n6700), .B(n6701), .Z(n6697) );
  ANDN U7866 ( .B(n6702), .A(n135), .Z(n6700) );
  XNOR U7867 ( .A(a[884]), .B(n6703), .Z(n135) );
  IV U7868 ( .A(n6701), .Z(n6703) );
  XNOR U7869 ( .A(b[884]), .B(n6701), .Z(n6702) );
  XOR U7870 ( .A(n6704), .B(n6705), .Z(n6701) );
  ANDN U7871 ( .B(n6706), .A(n136), .Z(n6704) );
  XNOR U7872 ( .A(a[883]), .B(n6707), .Z(n136) );
  IV U7873 ( .A(n6705), .Z(n6707) );
  XNOR U7874 ( .A(b[883]), .B(n6705), .Z(n6706) );
  XOR U7875 ( .A(n6708), .B(n6709), .Z(n6705) );
  ANDN U7876 ( .B(n6710), .A(n137), .Z(n6708) );
  XNOR U7877 ( .A(a[882]), .B(n6711), .Z(n137) );
  IV U7878 ( .A(n6709), .Z(n6711) );
  XNOR U7879 ( .A(b[882]), .B(n6709), .Z(n6710) );
  XOR U7880 ( .A(n6712), .B(n6713), .Z(n6709) );
  ANDN U7881 ( .B(n6714), .A(n138), .Z(n6712) );
  XNOR U7882 ( .A(a[881]), .B(n6715), .Z(n138) );
  IV U7883 ( .A(n6713), .Z(n6715) );
  XNOR U7884 ( .A(b[881]), .B(n6713), .Z(n6714) );
  XOR U7885 ( .A(n6716), .B(n6717), .Z(n6713) );
  ANDN U7886 ( .B(n6718), .A(n139), .Z(n6716) );
  XNOR U7887 ( .A(a[880]), .B(n6719), .Z(n139) );
  IV U7888 ( .A(n6717), .Z(n6719) );
  XNOR U7889 ( .A(b[880]), .B(n6717), .Z(n6718) );
  XOR U7890 ( .A(n6720), .B(n6721), .Z(n6717) );
  ANDN U7891 ( .B(n6722), .A(n141), .Z(n6720) );
  XNOR U7892 ( .A(a[879]), .B(n6723), .Z(n141) );
  IV U7893 ( .A(n6721), .Z(n6723) );
  XNOR U7894 ( .A(b[879]), .B(n6721), .Z(n6722) );
  XOR U7895 ( .A(n6724), .B(n6725), .Z(n6721) );
  ANDN U7896 ( .B(n6726), .A(n142), .Z(n6724) );
  XNOR U7897 ( .A(a[878]), .B(n6727), .Z(n142) );
  IV U7898 ( .A(n6725), .Z(n6727) );
  XNOR U7899 ( .A(b[878]), .B(n6725), .Z(n6726) );
  XOR U7900 ( .A(n6728), .B(n6729), .Z(n6725) );
  ANDN U7901 ( .B(n6730), .A(n143), .Z(n6728) );
  XNOR U7902 ( .A(a[877]), .B(n6731), .Z(n143) );
  IV U7903 ( .A(n6729), .Z(n6731) );
  XNOR U7904 ( .A(b[877]), .B(n6729), .Z(n6730) );
  XOR U7905 ( .A(n6732), .B(n6733), .Z(n6729) );
  ANDN U7906 ( .B(n6734), .A(n144), .Z(n6732) );
  XNOR U7907 ( .A(a[876]), .B(n6735), .Z(n144) );
  IV U7908 ( .A(n6733), .Z(n6735) );
  XNOR U7909 ( .A(b[876]), .B(n6733), .Z(n6734) );
  XOR U7910 ( .A(n6736), .B(n6737), .Z(n6733) );
  ANDN U7911 ( .B(n6738), .A(n145), .Z(n6736) );
  XNOR U7912 ( .A(a[875]), .B(n6739), .Z(n145) );
  IV U7913 ( .A(n6737), .Z(n6739) );
  XNOR U7914 ( .A(b[875]), .B(n6737), .Z(n6738) );
  XOR U7915 ( .A(n6740), .B(n6741), .Z(n6737) );
  ANDN U7916 ( .B(n6742), .A(n146), .Z(n6740) );
  XNOR U7917 ( .A(a[874]), .B(n6743), .Z(n146) );
  IV U7918 ( .A(n6741), .Z(n6743) );
  XNOR U7919 ( .A(b[874]), .B(n6741), .Z(n6742) );
  XOR U7920 ( .A(n6744), .B(n6745), .Z(n6741) );
  ANDN U7921 ( .B(n6746), .A(n147), .Z(n6744) );
  XNOR U7922 ( .A(a[873]), .B(n6747), .Z(n147) );
  IV U7923 ( .A(n6745), .Z(n6747) );
  XNOR U7924 ( .A(b[873]), .B(n6745), .Z(n6746) );
  XOR U7925 ( .A(n6748), .B(n6749), .Z(n6745) );
  ANDN U7926 ( .B(n6750), .A(n148), .Z(n6748) );
  XNOR U7927 ( .A(a[872]), .B(n6751), .Z(n148) );
  IV U7928 ( .A(n6749), .Z(n6751) );
  XNOR U7929 ( .A(b[872]), .B(n6749), .Z(n6750) );
  XOR U7930 ( .A(n6752), .B(n6753), .Z(n6749) );
  ANDN U7931 ( .B(n6754), .A(n149), .Z(n6752) );
  XNOR U7932 ( .A(a[871]), .B(n6755), .Z(n149) );
  IV U7933 ( .A(n6753), .Z(n6755) );
  XNOR U7934 ( .A(b[871]), .B(n6753), .Z(n6754) );
  XOR U7935 ( .A(n6756), .B(n6757), .Z(n6753) );
  ANDN U7936 ( .B(n6758), .A(n150), .Z(n6756) );
  XNOR U7937 ( .A(a[870]), .B(n6759), .Z(n150) );
  IV U7938 ( .A(n6757), .Z(n6759) );
  XNOR U7939 ( .A(b[870]), .B(n6757), .Z(n6758) );
  XOR U7940 ( .A(n6760), .B(n6761), .Z(n6757) );
  ANDN U7941 ( .B(n6762), .A(n152), .Z(n6760) );
  XNOR U7942 ( .A(a[869]), .B(n6763), .Z(n152) );
  IV U7943 ( .A(n6761), .Z(n6763) );
  XNOR U7944 ( .A(b[869]), .B(n6761), .Z(n6762) );
  XOR U7945 ( .A(n6764), .B(n6765), .Z(n6761) );
  ANDN U7946 ( .B(n6766), .A(n153), .Z(n6764) );
  XNOR U7947 ( .A(a[868]), .B(n6767), .Z(n153) );
  IV U7948 ( .A(n6765), .Z(n6767) );
  XNOR U7949 ( .A(b[868]), .B(n6765), .Z(n6766) );
  XOR U7950 ( .A(n6768), .B(n6769), .Z(n6765) );
  ANDN U7951 ( .B(n6770), .A(n154), .Z(n6768) );
  XNOR U7952 ( .A(a[867]), .B(n6771), .Z(n154) );
  IV U7953 ( .A(n6769), .Z(n6771) );
  XNOR U7954 ( .A(b[867]), .B(n6769), .Z(n6770) );
  XOR U7955 ( .A(n6772), .B(n6773), .Z(n6769) );
  ANDN U7956 ( .B(n6774), .A(n155), .Z(n6772) );
  XNOR U7957 ( .A(a[866]), .B(n6775), .Z(n155) );
  IV U7958 ( .A(n6773), .Z(n6775) );
  XNOR U7959 ( .A(b[866]), .B(n6773), .Z(n6774) );
  XOR U7960 ( .A(n6776), .B(n6777), .Z(n6773) );
  ANDN U7961 ( .B(n6778), .A(n156), .Z(n6776) );
  XNOR U7962 ( .A(a[865]), .B(n6779), .Z(n156) );
  IV U7963 ( .A(n6777), .Z(n6779) );
  XNOR U7964 ( .A(b[865]), .B(n6777), .Z(n6778) );
  XOR U7965 ( .A(n6780), .B(n6781), .Z(n6777) );
  ANDN U7966 ( .B(n6782), .A(n157), .Z(n6780) );
  XNOR U7967 ( .A(a[864]), .B(n6783), .Z(n157) );
  IV U7968 ( .A(n6781), .Z(n6783) );
  XNOR U7969 ( .A(b[864]), .B(n6781), .Z(n6782) );
  XOR U7970 ( .A(n6784), .B(n6785), .Z(n6781) );
  ANDN U7971 ( .B(n6786), .A(n158), .Z(n6784) );
  XNOR U7972 ( .A(a[863]), .B(n6787), .Z(n158) );
  IV U7973 ( .A(n6785), .Z(n6787) );
  XNOR U7974 ( .A(b[863]), .B(n6785), .Z(n6786) );
  XOR U7975 ( .A(n6788), .B(n6789), .Z(n6785) );
  ANDN U7976 ( .B(n6790), .A(n159), .Z(n6788) );
  XNOR U7977 ( .A(a[862]), .B(n6791), .Z(n159) );
  IV U7978 ( .A(n6789), .Z(n6791) );
  XNOR U7979 ( .A(b[862]), .B(n6789), .Z(n6790) );
  XOR U7980 ( .A(n6792), .B(n6793), .Z(n6789) );
  ANDN U7981 ( .B(n6794), .A(n160), .Z(n6792) );
  XNOR U7982 ( .A(a[861]), .B(n6795), .Z(n160) );
  IV U7983 ( .A(n6793), .Z(n6795) );
  XNOR U7984 ( .A(b[861]), .B(n6793), .Z(n6794) );
  XOR U7985 ( .A(n6796), .B(n6797), .Z(n6793) );
  ANDN U7986 ( .B(n6798), .A(n161), .Z(n6796) );
  XNOR U7987 ( .A(a[860]), .B(n6799), .Z(n161) );
  IV U7988 ( .A(n6797), .Z(n6799) );
  XNOR U7989 ( .A(b[860]), .B(n6797), .Z(n6798) );
  XOR U7990 ( .A(n6800), .B(n6801), .Z(n6797) );
  ANDN U7991 ( .B(n6802), .A(n163), .Z(n6800) );
  XNOR U7992 ( .A(a[859]), .B(n6803), .Z(n163) );
  IV U7993 ( .A(n6801), .Z(n6803) );
  XNOR U7994 ( .A(b[859]), .B(n6801), .Z(n6802) );
  XOR U7995 ( .A(n6804), .B(n6805), .Z(n6801) );
  ANDN U7996 ( .B(n6806), .A(n164), .Z(n6804) );
  XNOR U7997 ( .A(a[858]), .B(n6807), .Z(n164) );
  IV U7998 ( .A(n6805), .Z(n6807) );
  XNOR U7999 ( .A(b[858]), .B(n6805), .Z(n6806) );
  XOR U8000 ( .A(n6808), .B(n6809), .Z(n6805) );
  ANDN U8001 ( .B(n6810), .A(n165), .Z(n6808) );
  XNOR U8002 ( .A(a[857]), .B(n6811), .Z(n165) );
  IV U8003 ( .A(n6809), .Z(n6811) );
  XNOR U8004 ( .A(b[857]), .B(n6809), .Z(n6810) );
  XOR U8005 ( .A(n6812), .B(n6813), .Z(n6809) );
  ANDN U8006 ( .B(n6814), .A(n166), .Z(n6812) );
  XNOR U8007 ( .A(a[856]), .B(n6815), .Z(n166) );
  IV U8008 ( .A(n6813), .Z(n6815) );
  XNOR U8009 ( .A(b[856]), .B(n6813), .Z(n6814) );
  XOR U8010 ( .A(n6816), .B(n6817), .Z(n6813) );
  ANDN U8011 ( .B(n6818), .A(n167), .Z(n6816) );
  XNOR U8012 ( .A(a[855]), .B(n6819), .Z(n167) );
  IV U8013 ( .A(n6817), .Z(n6819) );
  XNOR U8014 ( .A(b[855]), .B(n6817), .Z(n6818) );
  XOR U8015 ( .A(n6820), .B(n6821), .Z(n6817) );
  ANDN U8016 ( .B(n6822), .A(n168), .Z(n6820) );
  XNOR U8017 ( .A(a[854]), .B(n6823), .Z(n168) );
  IV U8018 ( .A(n6821), .Z(n6823) );
  XNOR U8019 ( .A(b[854]), .B(n6821), .Z(n6822) );
  XOR U8020 ( .A(n6824), .B(n6825), .Z(n6821) );
  ANDN U8021 ( .B(n6826), .A(n169), .Z(n6824) );
  XNOR U8022 ( .A(a[853]), .B(n6827), .Z(n169) );
  IV U8023 ( .A(n6825), .Z(n6827) );
  XNOR U8024 ( .A(b[853]), .B(n6825), .Z(n6826) );
  XOR U8025 ( .A(n6828), .B(n6829), .Z(n6825) );
  ANDN U8026 ( .B(n6830), .A(n170), .Z(n6828) );
  XNOR U8027 ( .A(a[852]), .B(n6831), .Z(n170) );
  IV U8028 ( .A(n6829), .Z(n6831) );
  XNOR U8029 ( .A(b[852]), .B(n6829), .Z(n6830) );
  XOR U8030 ( .A(n6832), .B(n6833), .Z(n6829) );
  ANDN U8031 ( .B(n6834), .A(n171), .Z(n6832) );
  XNOR U8032 ( .A(a[851]), .B(n6835), .Z(n171) );
  IV U8033 ( .A(n6833), .Z(n6835) );
  XNOR U8034 ( .A(b[851]), .B(n6833), .Z(n6834) );
  XOR U8035 ( .A(n6836), .B(n6837), .Z(n6833) );
  ANDN U8036 ( .B(n6838), .A(n172), .Z(n6836) );
  XNOR U8037 ( .A(a[850]), .B(n6839), .Z(n172) );
  IV U8038 ( .A(n6837), .Z(n6839) );
  XNOR U8039 ( .A(b[850]), .B(n6837), .Z(n6838) );
  XOR U8040 ( .A(n6840), .B(n6841), .Z(n6837) );
  ANDN U8041 ( .B(n6842), .A(n174), .Z(n6840) );
  XNOR U8042 ( .A(a[849]), .B(n6843), .Z(n174) );
  IV U8043 ( .A(n6841), .Z(n6843) );
  XNOR U8044 ( .A(b[849]), .B(n6841), .Z(n6842) );
  XOR U8045 ( .A(n6844), .B(n6845), .Z(n6841) );
  ANDN U8046 ( .B(n6846), .A(n175), .Z(n6844) );
  XNOR U8047 ( .A(a[848]), .B(n6847), .Z(n175) );
  IV U8048 ( .A(n6845), .Z(n6847) );
  XNOR U8049 ( .A(b[848]), .B(n6845), .Z(n6846) );
  XOR U8050 ( .A(n6848), .B(n6849), .Z(n6845) );
  ANDN U8051 ( .B(n6850), .A(n176), .Z(n6848) );
  XNOR U8052 ( .A(a[847]), .B(n6851), .Z(n176) );
  IV U8053 ( .A(n6849), .Z(n6851) );
  XNOR U8054 ( .A(b[847]), .B(n6849), .Z(n6850) );
  XOR U8055 ( .A(n6852), .B(n6853), .Z(n6849) );
  ANDN U8056 ( .B(n6854), .A(n177), .Z(n6852) );
  XNOR U8057 ( .A(a[846]), .B(n6855), .Z(n177) );
  IV U8058 ( .A(n6853), .Z(n6855) );
  XNOR U8059 ( .A(b[846]), .B(n6853), .Z(n6854) );
  XOR U8060 ( .A(n6856), .B(n6857), .Z(n6853) );
  ANDN U8061 ( .B(n6858), .A(n178), .Z(n6856) );
  XNOR U8062 ( .A(a[845]), .B(n6859), .Z(n178) );
  IV U8063 ( .A(n6857), .Z(n6859) );
  XNOR U8064 ( .A(b[845]), .B(n6857), .Z(n6858) );
  XOR U8065 ( .A(n6860), .B(n6861), .Z(n6857) );
  ANDN U8066 ( .B(n6862), .A(n179), .Z(n6860) );
  XNOR U8067 ( .A(a[844]), .B(n6863), .Z(n179) );
  IV U8068 ( .A(n6861), .Z(n6863) );
  XNOR U8069 ( .A(b[844]), .B(n6861), .Z(n6862) );
  XOR U8070 ( .A(n6864), .B(n6865), .Z(n6861) );
  ANDN U8071 ( .B(n6866), .A(n180), .Z(n6864) );
  XNOR U8072 ( .A(a[843]), .B(n6867), .Z(n180) );
  IV U8073 ( .A(n6865), .Z(n6867) );
  XNOR U8074 ( .A(b[843]), .B(n6865), .Z(n6866) );
  XOR U8075 ( .A(n6868), .B(n6869), .Z(n6865) );
  ANDN U8076 ( .B(n6870), .A(n181), .Z(n6868) );
  XNOR U8077 ( .A(a[842]), .B(n6871), .Z(n181) );
  IV U8078 ( .A(n6869), .Z(n6871) );
  XNOR U8079 ( .A(b[842]), .B(n6869), .Z(n6870) );
  XOR U8080 ( .A(n6872), .B(n6873), .Z(n6869) );
  ANDN U8081 ( .B(n6874), .A(n182), .Z(n6872) );
  XNOR U8082 ( .A(a[841]), .B(n6875), .Z(n182) );
  IV U8083 ( .A(n6873), .Z(n6875) );
  XNOR U8084 ( .A(b[841]), .B(n6873), .Z(n6874) );
  XOR U8085 ( .A(n6876), .B(n6877), .Z(n6873) );
  ANDN U8086 ( .B(n6878), .A(n183), .Z(n6876) );
  XNOR U8087 ( .A(a[840]), .B(n6879), .Z(n183) );
  IV U8088 ( .A(n6877), .Z(n6879) );
  XNOR U8089 ( .A(b[840]), .B(n6877), .Z(n6878) );
  XOR U8090 ( .A(n6880), .B(n6881), .Z(n6877) );
  ANDN U8091 ( .B(n6882), .A(n185), .Z(n6880) );
  XNOR U8092 ( .A(a[839]), .B(n6883), .Z(n185) );
  IV U8093 ( .A(n6881), .Z(n6883) );
  XNOR U8094 ( .A(b[839]), .B(n6881), .Z(n6882) );
  XOR U8095 ( .A(n6884), .B(n6885), .Z(n6881) );
  ANDN U8096 ( .B(n6886), .A(n186), .Z(n6884) );
  XNOR U8097 ( .A(a[838]), .B(n6887), .Z(n186) );
  IV U8098 ( .A(n6885), .Z(n6887) );
  XNOR U8099 ( .A(b[838]), .B(n6885), .Z(n6886) );
  XOR U8100 ( .A(n6888), .B(n6889), .Z(n6885) );
  ANDN U8101 ( .B(n6890), .A(n187), .Z(n6888) );
  XNOR U8102 ( .A(a[837]), .B(n6891), .Z(n187) );
  IV U8103 ( .A(n6889), .Z(n6891) );
  XNOR U8104 ( .A(b[837]), .B(n6889), .Z(n6890) );
  XOR U8105 ( .A(n6892), .B(n6893), .Z(n6889) );
  ANDN U8106 ( .B(n6894), .A(n188), .Z(n6892) );
  XNOR U8107 ( .A(a[836]), .B(n6895), .Z(n188) );
  IV U8108 ( .A(n6893), .Z(n6895) );
  XNOR U8109 ( .A(b[836]), .B(n6893), .Z(n6894) );
  XOR U8110 ( .A(n6896), .B(n6897), .Z(n6893) );
  ANDN U8111 ( .B(n6898), .A(n189), .Z(n6896) );
  XNOR U8112 ( .A(a[835]), .B(n6899), .Z(n189) );
  IV U8113 ( .A(n6897), .Z(n6899) );
  XNOR U8114 ( .A(b[835]), .B(n6897), .Z(n6898) );
  XOR U8115 ( .A(n6900), .B(n6901), .Z(n6897) );
  ANDN U8116 ( .B(n6902), .A(n190), .Z(n6900) );
  XNOR U8117 ( .A(a[834]), .B(n6903), .Z(n190) );
  IV U8118 ( .A(n6901), .Z(n6903) );
  XNOR U8119 ( .A(b[834]), .B(n6901), .Z(n6902) );
  XOR U8120 ( .A(n6904), .B(n6905), .Z(n6901) );
  ANDN U8121 ( .B(n6906), .A(n191), .Z(n6904) );
  XNOR U8122 ( .A(a[833]), .B(n6907), .Z(n191) );
  IV U8123 ( .A(n6905), .Z(n6907) );
  XNOR U8124 ( .A(b[833]), .B(n6905), .Z(n6906) );
  XOR U8125 ( .A(n6908), .B(n6909), .Z(n6905) );
  ANDN U8126 ( .B(n6910), .A(n192), .Z(n6908) );
  XNOR U8127 ( .A(a[832]), .B(n6911), .Z(n192) );
  IV U8128 ( .A(n6909), .Z(n6911) );
  XNOR U8129 ( .A(b[832]), .B(n6909), .Z(n6910) );
  XOR U8130 ( .A(n6912), .B(n6913), .Z(n6909) );
  ANDN U8131 ( .B(n6914), .A(n193), .Z(n6912) );
  XNOR U8132 ( .A(a[831]), .B(n6915), .Z(n193) );
  IV U8133 ( .A(n6913), .Z(n6915) );
  XNOR U8134 ( .A(b[831]), .B(n6913), .Z(n6914) );
  XOR U8135 ( .A(n6916), .B(n6917), .Z(n6913) );
  ANDN U8136 ( .B(n6918), .A(n194), .Z(n6916) );
  XNOR U8137 ( .A(a[830]), .B(n6919), .Z(n194) );
  IV U8138 ( .A(n6917), .Z(n6919) );
  XNOR U8139 ( .A(b[830]), .B(n6917), .Z(n6918) );
  XOR U8140 ( .A(n6920), .B(n6921), .Z(n6917) );
  ANDN U8141 ( .B(n6922), .A(n196), .Z(n6920) );
  XNOR U8142 ( .A(a[829]), .B(n6923), .Z(n196) );
  IV U8143 ( .A(n6921), .Z(n6923) );
  XNOR U8144 ( .A(b[829]), .B(n6921), .Z(n6922) );
  XOR U8145 ( .A(n6924), .B(n6925), .Z(n6921) );
  ANDN U8146 ( .B(n6926), .A(n197), .Z(n6924) );
  XNOR U8147 ( .A(a[828]), .B(n6927), .Z(n197) );
  IV U8148 ( .A(n6925), .Z(n6927) );
  XNOR U8149 ( .A(b[828]), .B(n6925), .Z(n6926) );
  XOR U8150 ( .A(n6928), .B(n6929), .Z(n6925) );
  ANDN U8151 ( .B(n6930), .A(n198), .Z(n6928) );
  XNOR U8152 ( .A(a[827]), .B(n6931), .Z(n198) );
  IV U8153 ( .A(n6929), .Z(n6931) );
  XNOR U8154 ( .A(b[827]), .B(n6929), .Z(n6930) );
  XOR U8155 ( .A(n6932), .B(n6933), .Z(n6929) );
  ANDN U8156 ( .B(n6934), .A(n199), .Z(n6932) );
  XNOR U8157 ( .A(a[826]), .B(n6935), .Z(n199) );
  IV U8158 ( .A(n6933), .Z(n6935) );
  XNOR U8159 ( .A(b[826]), .B(n6933), .Z(n6934) );
  XOR U8160 ( .A(n6936), .B(n6937), .Z(n6933) );
  ANDN U8161 ( .B(n6938), .A(n200), .Z(n6936) );
  XNOR U8162 ( .A(a[825]), .B(n6939), .Z(n200) );
  IV U8163 ( .A(n6937), .Z(n6939) );
  XNOR U8164 ( .A(b[825]), .B(n6937), .Z(n6938) );
  XOR U8165 ( .A(n6940), .B(n6941), .Z(n6937) );
  ANDN U8166 ( .B(n6942), .A(n201), .Z(n6940) );
  XNOR U8167 ( .A(a[824]), .B(n6943), .Z(n201) );
  IV U8168 ( .A(n6941), .Z(n6943) );
  XNOR U8169 ( .A(b[824]), .B(n6941), .Z(n6942) );
  XOR U8170 ( .A(n6944), .B(n6945), .Z(n6941) );
  ANDN U8171 ( .B(n6946), .A(n202), .Z(n6944) );
  XNOR U8172 ( .A(a[823]), .B(n6947), .Z(n202) );
  IV U8173 ( .A(n6945), .Z(n6947) );
  XNOR U8174 ( .A(b[823]), .B(n6945), .Z(n6946) );
  XOR U8175 ( .A(n6948), .B(n6949), .Z(n6945) );
  ANDN U8176 ( .B(n6950), .A(n203), .Z(n6948) );
  XNOR U8177 ( .A(a[822]), .B(n6951), .Z(n203) );
  IV U8178 ( .A(n6949), .Z(n6951) );
  XNOR U8179 ( .A(b[822]), .B(n6949), .Z(n6950) );
  XOR U8180 ( .A(n6952), .B(n6953), .Z(n6949) );
  ANDN U8181 ( .B(n6954), .A(n204), .Z(n6952) );
  XNOR U8182 ( .A(a[821]), .B(n6955), .Z(n204) );
  IV U8183 ( .A(n6953), .Z(n6955) );
  XNOR U8184 ( .A(b[821]), .B(n6953), .Z(n6954) );
  XOR U8185 ( .A(n6956), .B(n6957), .Z(n6953) );
  ANDN U8186 ( .B(n6958), .A(n205), .Z(n6956) );
  XNOR U8187 ( .A(a[820]), .B(n6959), .Z(n205) );
  IV U8188 ( .A(n6957), .Z(n6959) );
  XNOR U8189 ( .A(b[820]), .B(n6957), .Z(n6958) );
  XOR U8190 ( .A(n6960), .B(n6961), .Z(n6957) );
  ANDN U8191 ( .B(n6962), .A(n207), .Z(n6960) );
  XNOR U8192 ( .A(a[819]), .B(n6963), .Z(n207) );
  IV U8193 ( .A(n6961), .Z(n6963) );
  XNOR U8194 ( .A(b[819]), .B(n6961), .Z(n6962) );
  XOR U8195 ( .A(n6964), .B(n6965), .Z(n6961) );
  ANDN U8196 ( .B(n6966), .A(n208), .Z(n6964) );
  XNOR U8197 ( .A(a[818]), .B(n6967), .Z(n208) );
  IV U8198 ( .A(n6965), .Z(n6967) );
  XNOR U8199 ( .A(b[818]), .B(n6965), .Z(n6966) );
  XOR U8200 ( .A(n6968), .B(n6969), .Z(n6965) );
  ANDN U8201 ( .B(n6970), .A(n209), .Z(n6968) );
  XNOR U8202 ( .A(a[817]), .B(n6971), .Z(n209) );
  IV U8203 ( .A(n6969), .Z(n6971) );
  XNOR U8204 ( .A(b[817]), .B(n6969), .Z(n6970) );
  XOR U8205 ( .A(n6972), .B(n6973), .Z(n6969) );
  ANDN U8206 ( .B(n6974), .A(n210), .Z(n6972) );
  XNOR U8207 ( .A(a[816]), .B(n6975), .Z(n210) );
  IV U8208 ( .A(n6973), .Z(n6975) );
  XNOR U8209 ( .A(b[816]), .B(n6973), .Z(n6974) );
  XOR U8210 ( .A(n6976), .B(n6977), .Z(n6973) );
  ANDN U8211 ( .B(n6978), .A(n211), .Z(n6976) );
  XNOR U8212 ( .A(a[815]), .B(n6979), .Z(n211) );
  IV U8213 ( .A(n6977), .Z(n6979) );
  XNOR U8214 ( .A(b[815]), .B(n6977), .Z(n6978) );
  XOR U8215 ( .A(n6980), .B(n6981), .Z(n6977) );
  ANDN U8216 ( .B(n6982), .A(n212), .Z(n6980) );
  XNOR U8217 ( .A(a[814]), .B(n6983), .Z(n212) );
  IV U8218 ( .A(n6981), .Z(n6983) );
  XNOR U8219 ( .A(b[814]), .B(n6981), .Z(n6982) );
  XOR U8220 ( .A(n6984), .B(n6985), .Z(n6981) );
  ANDN U8221 ( .B(n6986), .A(n213), .Z(n6984) );
  XNOR U8222 ( .A(a[813]), .B(n6987), .Z(n213) );
  IV U8223 ( .A(n6985), .Z(n6987) );
  XNOR U8224 ( .A(b[813]), .B(n6985), .Z(n6986) );
  XOR U8225 ( .A(n6988), .B(n6989), .Z(n6985) );
  ANDN U8226 ( .B(n6990), .A(n214), .Z(n6988) );
  XNOR U8227 ( .A(a[812]), .B(n6991), .Z(n214) );
  IV U8228 ( .A(n6989), .Z(n6991) );
  XNOR U8229 ( .A(b[812]), .B(n6989), .Z(n6990) );
  XOR U8230 ( .A(n6992), .B(n6993), .Z(n6989) );
  ANDN U8231 ( .B(n6994), .A(n215), .Z(n6992) );
  XNOR U8232 ( .A(a[811]), .B(n6995), .Z(n215) );
  IV U8233 ( .A(n6993), .Z(n6995) );
  XNOR U8234 ( .A(b[811]), .B(n6993), .Z(n6994) );
  XOR U8235 ( .A(n6996), .B(n6997), .Z(n6993) );
  ANDN U8236 ( .B(n6998), .A(n216), .Z(n6996) );
  XNOR U8237 ( .A(a[810]), .B(n6999), .Z(n216) );
  IV U8238 ( .A(n6997), .Z(n6999) );
  XNOR U8239 ( .A(b[810]), .B(n6997), .Z(n6998) );
  XOR U8240 ( .A(n7000), .B(n7001), .Z(n6997) );
  ANDN U8241 ( .B(n7002), .A(n218), .Z(n7000) );
  XNOR U8242 ( .A(a[809]), .B(n7003), .Z(n218) );
  IV U8243 ( .A(n7001), .Z(n7003) );
  XNOR U8244 ( .A(b[809]), .B(n7001), .Z(n7002) );
  XOR U8245 ( .A(n7004), .B(n7005), .Z(n7001) );
  ANDN U8246 ( .B(n7006), .A(n219), .Z(n7004) );
  XNOR U8247 ( .A(a[808]), .B(n7007), .Z(n219) );
  IV U8248 ( .A(n7005), .Z(n7007) );
  XNOR U8249 ( .A(b[808]), .B(n7005), .Z(n7006) );
  XOR U8250 ( .A(n7008), .B(n7009), .Z(n7005) );
  ANDN U8251 ( .B(n7010), .A(n220), .Z(n7008) );
  XNOR U8252 ( .A(a[807]), .B(n7011), .Z(n220) );
  IV U8253 ( .A(n7009), .Z(n7011) );
  XNOR U8254 ( .A(b[807]), .B(n7009), .Z(n7010) );
  XOR U8255 ( .A(n7012), .B(n7013), .Z(n7009) );
  ANDN U8256 ( .B(n7014), .A(n221), .Z(n7012) );
  XNOR U8257 ( .A(a[806]), .B(n7015), .Z(n221) );
  IV U8258 ( .A(n7013), .Z(n7015) );
  XNOR U8259 ( .A(b[806]), .B(n7013), .Z(n7014) );
  XOR U8260 ( .A(n7016), .B(n7017), .Z(n7013) );
  ANDN U8261 ( .B(n7018), .A(n222), .Z(n7016) );
  XNOR U8262 ( .A(a[805]), .B(n7019), .Z(n222) );
  IV U8263 ( .A(n7017), .Z(n7019) );
  XNOR U8264 ( .A(b[805]), .B(n7017), .Z(n7018) );
  XOR U8265 ( .A(n7020), .B(n7021), .Z(n7017) );
  ANDN U8266 ( .B(n7022), .A(n223), .Z(n7020) );
  XNOR U8267 ( .A(a[804]), .B(n7023), .Z(n223) );
  IV U8268 ( .A(n7021), .Z(n7023) );
  XNOR U8269 ( .A(b[804]), .B(n7021), .Z(n7022) );
  XOR U8270 ( .A(n7024), .B(n7025), .Z(n7021) );
  ANDN U8271 ( .B(n7026), .A(n224), .Z(n7024) );
  XNOR U8272 ( .A(a[803]), .B(n7027), .Z(n224) );
  IV U8273 ( .A(n7025), .Z(n7027) );
  XNOR U8274 ( .A(b[803]), .B(n7025), .Z(n7026) );
  XOR U8275 ( .A(n7028), .B(n7029), .Z(n7025) );
  ANDN U8276 ( .B(n7030), .A(n225), .Z(n7028) );
  XNOR U8277 ( .A(a[802]), .B(n7031), .Z(n225) );
  IV U8278 ( .A(n7029), .Z(n7031) );
  XNOR U8279 ( .A(b[802]), .B(n7029), .Z(n7030) );
  XOR U8280 ( .A(n7032), .B(n7033), .Z(n7029) );
  ANDN U8281 ( .B(n7034), .A(n226), .Z(n7032) );
  XNOR U8282 ( .A(a[801]), .B(n7035), .Z(n226) );
  IV U8283 ( .A(n7033), .Z(n7035) );
  XNOR U8284 ( .A(b[801]), .B(n7033), .Z(n7034) );
  XOR U8285 ( .A(n7036), .B(n7037), .Z(n7033) );
  ANDN U8286 ( .B(n7038), .A(n227), .Z(n7036) );
  XNOR U8287 ( .A(a[800]), .B(n7039), .Z(n227) );
  IV U8288 ( .A(n7037), .Z(n7039) );
  XNOR U8289 ( .A(b[800]), .B(n7037), .Z(n7038) );
  XOR U8290 ( .A(n7040), .B(n7041), .Z(n7037) );
  ANDN U8291 ( .B(n7042), .A(n230), .Z(n7040) );
  XNOR U8292 ( .A(a[799]), .B(n7043), .Z(n230) );
  IV U8293 ( .A(n7041), .Z(n7043) );
  XNOR U8294 ( .A(b[799]), .B(n7041), .Z(n7042) );
  XOR U8295 ( .A(n7044), .B(n7045), .Z(n7041) );
  ANDN U8296 ( .B(n7046), .A(n231), .Z(n7044) );
  XNOR U8297 ( .A(a[798]), .B(n7047), .Z(n231) );
  IV U8298 ( .A(n7045), .Z(n7047) );
  XNOR U8299 ( .A(b[798]), .B(n7045), .Z(n7046) );
  XOR U8300 ( .A(n7048), .B(n7049), .Z(n7045) );
  ANDN U8301 ( .B(n7050), .A(n232), .Z(n7048) );
  XNOR U8302 ( .A(a[797]), .B(n7051), .Z(n232) );
  IV U8303 ( .A(n7049), .Z(n7051) );
  XNOR U8304 ( .A(b[797]), .B(n7049), .Z(n7050) );
  XOR U8305 ( .A(n7052), .B(n7053), .Z(n7049) );
  ANDN U8306 ( .B(n7054), .A(n233), .Z(n7052) );
  XNOR U8307 ( .A(a[796]), .B(n7055), .Z(n233) );
  IV U8308 ( .A(n7053), .Z(n7055) );
  XNOR U8309 ( .A(b[796]), .B(n7053), .Z(n7054) );
  XOR U8310 ( .A(n7056), .B(n7057), .Z(n7053) );
  ANDN U8311 ( .B(n7058), .A(n234), .Z(n7056) );
  XNOR U8312 ( .A(a[795]), .B(n7059), .Z(n234) );
  IV U8313 ( .A(n7057), .Z(n7059) );
  XNOR U8314 ( .A(b[795]), .B(n7057), .Z(n7058) );
  XOR U8315 ( .A(n7060), .B(n7061), .Z(n7057) );
  ANDN U8316 ( .B(n7062), .A(n235), .Z(n7060) );
  XNOR U8317 ( .A(a[794]), .B(n7063), .Z(n235) );
  IV U8318 ( .A(n7061), .Z(n7063) );
  XNOR U8319 ( .A(b[794]), .B(n7061), .Z(n7062) );
  XOR U8320 ( .A(n7064), .B(n7065), .Z(n7061) );
  ANDN U8321 ( .B(n7066), .A(n236), .Z(n7064) );
  XNOR U8322 ( .A(a[793]), .B(n7067), .Z(n236) );
  IV U8323 ( .A(n7065), .Z(n7067) );
  XNOR U8324 ( .A(b[793]), .B(n7065), .Z(n7066) );
  XOR U8325 ( .A(n7068), .B(n7069), .Z(n7065) );
  ANDN U8326 ( .B(n7070), .A(n237), .Z(n7068) );
  XNOR U8327 ( .A(a[792]), .B(n7071), .Z(n237) );
  IV U8328 ( .A(n7069), .Z(n7071) );
  XNOR U8329 ( .A(b[792]), .B(n7069), .Z(n7070) );
  XOR U8330 ( .A(n7072), .B(n7073), .Z(n7069) );
  ANDN U8331 ( .B(n7074), .A(n238), .Z(n7072) );
  XNOR U8332 ( .A(a[791]), .B(n7075), .Z(n238) );
  IV U8333 ( .A(n7073), .Z(n7075) );
  XNOR U8334 ( .A(b[791]), .B(n7073), .Z(n7074) );
  XOR U8335 ( .A(n7076), .B(n7077), .Z(n7073) );
  ANDN U8336 ( .B(n7078), .A(n239), .Z(n7076) );
  XNOR U8337 ( .A(a[790]), .B(n7079), .Z(n239) );
  IV U8338 ( .A(n7077), .Z(n7079) );
  XNOR U8339 ( .A(b[790]), .B(n7077), .Z(n7078) );
  XOR U8340 ( .A(n7080), .B(n7081), .Z(n7077) );
  ANDN U8341 ( .B(n7082), .A(n241), .Z(n7080) );
  XNOR U8342 ( .A(a[789]), .B(n7083), .Z(n241) );
  IV U8343 ( .A(n7081), .Z(n7083) );
  XNOR U8344 ( .A(b[789]), .B(n7081), .Z(n7082) );
  XOR U8345 ( .A(n7084), .B(n7085), .Z(n7081) );
  ANDN U8346 ( .B(n7086), .A(n242), .Z(n7084) );
  XNOR U8347 ( .A(a[788]), .B(n7087), .Z(n242) );
  IV U8348 ( .A(n7085), .Z(n7087) );
  XNOR U8349 ( .A(b[788]), .B(n7085), .Z(n7086) );
  XOR U8350 ( .A(n7088), .B(n7089), .Z(n7085) );
  ANDN U8351 ( .B(n7090), .A(n243), .Z(n7088) );
  XNOR U8352 ( .A(a[787]), .B(n7091), .Z(n243) );
  IV U8353 ( .A(n7089), .Z(n7091) );
  XNOR U8354 ( .A(b[787]), .B(n7089), .Z(n7090) );
  XOR U8355 ( .A(n7092), .B(n7093), .Z(n7089) );
  ANDN U8356 ( .B(n7094), .A(n244), .Z(n7092) );
  XNOR U8357 ( .A(a[786]), .B(n7095), .Z(n244) );
  IV U8358 ( .A(n7093), .Z(n7095) );
  XNOR U8359 ( .A(b[786]), .B(n7093), .Z(n7094) );
  XOR U8360 ( .A(n7096), .B(n7097), .Z(n7093) );
  ANDN U8361 ( .B(n7098), .A(n245), .Z(n7096) );
  XNOR U8362 ( .A(a[785]), .B(n7099), .Z(n245) );
  IV U8363 ( .A(n7097), .Z(n7099) );
  XNOR U8364 ( .A(b[785]), .B(n7097), .Z(n7098) );
  XOR U8365 ( .A(n7100), .B(n7101), .Z(n7097) );
  ANDN U8366 ( .B(n7102), .A(n246), .Z(n7100) );
  XNOR U8367 ( .A(a[784]), .B(n7103), .Z(n246) );
  IV U8368 ( .A(n7101), .Z(n7103) );
  XNOR U8369 ( .A(b[784]), .B(n7101), .Z(n7102) );
  XOR U8370 ( .A(n7104), .B(n7105), .Z(n7101) );
  ANDN U8371 ( .B(n7106), .A(n247), .Z(n7104) );
  XNOR U8372 ( .A(a[783]), .B(n7107), .Z(n247) );
  IV U8373 ( .A(n7105), .Z(n7107) );
  XNOR U8374 ( .A(b[783]), .B(n7105), .Z(n7106) );
  XOR U8375 ( .A(n7108), .B(n7109), .Z(n7105) );
  ANDN U8376 ( .B(n7110), .A(n248), .Z(n7108) );
  XNOR U8377 ( .A(a[782]), .B(n7111), .Z(n248) );
  IV U8378 ( .A(n7109), .Z(n7111) );
  XNOR U8379 ( .A(b[782]), .B(n7109), .Z(n7110) );
  XOR U8380 ( .A(n7112), .B(n7113), .Z(n7109) );
  ANDN U8381 ( .B(n7114), .A(n249), .Z(n7112) );
  XNOR U8382 ( .A(a[781]), .B(n7115), .Z(n249) );
  IV U8383 ( .A(n7113), .Z(n7115) );
  XNOR U8384 ( .A(b[781]), .B(n7113), .Z(n7114) );
  XOR U8385 ( .A(n7116), .B(n7117), .Z(n7113) );
  ANDN U8386 ( .B(n7118), .A(n250), .Z(n7116) );
  XNOR U8387 ( .A(a[780]), .B(n7119), .Z(n250) );
  IV U8388 ( .A(n7117), .Z(n7119) );
  XNOR U8389 ( .A(b[780]), .B(n7117), .Z(n7118) );
  XOR U8390 ( .A(n7120), .B(n7121), .Z(n7117) );
  ANDN U8391 ( .B(n7122), .A(n252), .Z(n7120) );
  XNOR U8392 ( .A(a[779]), .B(n7123), .Z(n252) );
  IV U8393 ( .A(n7121), .Z(n7123) );
  XNOR U8394 ( .A(b[779]), .B(n7121), .Z(n7122) );
  XOR U8395 ( .A(n7124), .B(n7125), .Z(n7121) );
  ANDN U8396 ( .B(n7126), .A(n253), .Z(n7124) );
  XNOR U8397 ( .A(a[778]), .B(n7127), .Z(n253) );
  IV U8398 ( .A(n7125), .Z(n7127) );
  XNOR U8399 ( .A(b[778]), .B(n7125), .Z(n7126) );
  XOR U8400 ( .A(n7128), .B(n7129), .Z(n7125) );
  ANDN U8401 ( .B(n7130), .A(n254), .Z(n7128) );
  XNOR U8402 ( .A(a[777]), .B(n7131), .Z(n254) );
  IV U8403 ( .A(n7129), .Z(n7131) );
  XNOR U8404 ( .A(b[777]), .B(n7129), .Z(n7130) );
  XOR U8405 ( .A(n7132), .B(n7133), .Z(n7129) );
  ANDN U8406 ( .B(n7134), .A(n255), .Z(n7132) );
  XNOR U8407 ( .A(a[776]), .B(n7135), .Z(n255) );
  IV U8408 ( .A(n7133), .Z(n7135) );
  XNOR U8409 ( .A(b[776]), .B(n7133), .Z(n7134) );
  XOR U8410 ( .A(n7136), .B(n7137), .Z(n7133) );
  ANDN U8411 ( .B(n7138), .A(n256), .Z(n7136) );
  XNOR U8412 ( .A(a[775]), .B(n7139), .Z(n256) );
  IV U8413 ( .A(n7137), .Z(n7139) );
  XNOR U8414 ( .A(b[775]), .B(n7137), .Z(n7138) );
  XOR U8415 ( .A(n7140), .B(n7141), .Z(n7137) );
  ANDN U8416 ( .B(n7142), .A(n257), .Z(n7140) );
  XNOR U8417 ( .A(a[774]), .B(n7143), .Z(n257) );
  IV U8418 ( .A(n7141), .Z(n7143) );
  XNOR U8419 ( .A(b[774]), .B(n7141), .Z(n7142) );
  XOR U8420 ( .A(n7144), .B(n7145), .Z(n7141) );
  ANDN U8421 ( .B(n7146), .A(n258), .Z(n7144) );
  XNOR U8422 ( .A(a[773]), .B(n7147), .Z(n258) );
  IV U8423 ( .A(n7145), .Z(n7147) );
  XNOR U8424 ( .A(b[773]), .B(n7145), .Z(n7146) );
  XOR U8425 ( .A(n7148), .B(n7149), .Z(n7145) );
  ANDN U8426 ( .B(n7150), .A(n259), .Z(n7148) );
  XNOR U8427 ( .A(a[772]), .B(n7151), .Z(n259) );
  IV U8428 ( .A(n7149), .Z(n7151) );
  XNOR U8429 ( .A(b[772]), .B(n7149), .Z(n7150) );
  XOR U8430 ( .A(n7152), .B(n7153), .Z(n7149) );
  ANDN U8431 ( .B(n7154), .A(n260), .Z(n7152) );
  XNOR U8432 ( .A(a[771]), .B(n7155), .Z(n260) );
  IV U8433 ( .A(n7153), .Z(n7155) );
  XNOR U8434 ( .A(b[771]), .B(n7153), .Z(n7154) );
  XOR U8435 ( .A(n7156), .B(n7157), .Z(n7153) );
  ANDN U8436 ( .B(n7158), .A(n261), .Z(n7156) );
  XNOR U8437 ( .A(a[770]), .B(n7159), .Z(n261) );
  IV U8438 ( .A(n7157), .Z(n7159) );
  XNOR U8439 ( .A(b[770]), .B(n7157), .Z(n7158) );
  XOR U8440 ( .A(n7160), .B(n7161), .Z(n7157) );
  ANDN U8441 ( .B(n7162), .A(n263), .Z(n7160) );
  XNOR U8442 ( .A(a[769]), .B(n7163), .Z(n263) );
  IV U8443 ( .A(n7161), .Z(n7163) );
  XNOR U8444 ( .A(b[769]), .B(n7161), .Z(n7162) );
  XOR U8445 ( .A(n7164), .B(n7165), .Z(n7161) );
  ANDN U8446 ( .B(n7166), .A(n264), .Z(n7164) );
  XNOR U8447 ( .A(a[768]), .B(n7167), .Z(n264) );
  IV U8448 ( .A(n7165), .Z(n7167) );
  XNOR U8449 ( .A(b[768]), .B(n7165), .Z(n7166) );
  XOR U8450 ( .A(n7168), .B(n7169), .Z(n7165) );
  ANDN U8451 ( .B(n7170), .A(n265), .Z(n7168) );
  XNOR U8452 ( .A(a[767]), .B(n7171), .Z(n265) );
  IV U8453 ( .A(n7169), .Z(n7171) );
  XNOR U8454 ( .A(b[767]), .B(n7169), .Z(n7170) );
  XOR U8455 ( .A(n7172), .B(n7173), .Z(n7169) );
  ANDN U8456 ( .B(n7174), .A(n266), .Z(n7172) );
  XNOR U8457 ( .A(a[766]), .B(n7175), .Z(n266) );
  IV U8458 ( .A(n7173), .Z(n7175) );
  XNOR U8459 ( .A(b[766]), .B(n7173), .Z(n7174) );
  XOR U8460 ( .A(n7176), .B(n7177), .Z(n7173) );
  ANDN U8461 ( .B(n7178), .A(n267), .Z(n7176) );
  XNOR U8462 ( .A(a[765]), .B(n7179), .Z(n267) );
  IV U8463 ( .A(n7177), .Z(n7179) );
  XNOR U8464 ( .A(b[765]), .B(n7177), .Z(n7178) );
  XOR U8465 ( .A(n7180), .B(n7181), .Z(n7177) );
  ANDN U8466 ( .B(n7182), .A(n268), .Z(n7180) );
  XNOR U8467 ( .A(a[764]), .B(n7183), .Z(n268) );
  IV U8468 ( .A(n7181), .Z(n7183) );
  XNOR U8469 ( .A(b[764]), .B(n7181), .Z(n7182) );
  XOR U8470 ( .A(n7184), .B(n7185), .Z(n7181) );
  ANDN U8471 ( .B(n7186), .A(n269), .Z(n7184) );
  XNOR U8472 ( .A(a[763]), .B(n7187), .Z(n269) );
  IV U8473 ( .A(n7185), .Z(n7187) );
  XNOR U8474 ( .A(b[763]), .B(n7185), .Z(n7186) );
  XOR U8475 ( .A(n7188), .B(n7189), .Z(n7185) );
  ANDN U8476 ( .B(n7190), .A(n270), .Z(n7188) );
  XNOR U8477 ( .A(a[762]), .B(n7191), .Z(n270) );
  IV U8478 ( .A(n7189), .Z(n7191) );
  XNOR U8479 ( .A(b[762]), .B(n7189), .Z(n7190) );
  XOR U8480 ( .A(n7192), .B(n7193), .Z(n7189) );
  ANDN U8481 ( .B(n7194), .A(n271), .Z(n7192) );
  XNOR U8482 ( .A(a[761]), .B(n7195), .Z(n271) );
  IV U8483 ( .A(n7193), .Z(n7195) );
  XNOR U8484 ( .A(b[761]), .B(n7193), .Z(n7194) );
  XOR U8485 ( .A(n7196), .B(n7197), .Z(n7193) );
  ANDN U8486 ( .B(n7198), .A(n272), .Z(n7196) );
  XNOR U8487 ( .A(a[760]), .B(n7199), .Z(n272) );
  IV U8488 ( .A(n7197), .Z(n7199) );
  XNOR U8489 ( .A(b[760]), .B(n7197), .Z(n7198) );
  XOR U8490 ( .A(n7200), .B(n7201), .Z(n7197) );
  ANDN U8491 ( .B(n7202), .A(n274), .Z(n7200) );
  XNOR U8492 ( .A(a[759]), .B(n7203), .Z(n274) );
  IV U8493 ( .A(n7201), .Z(n7203) );
  XNOR U8494 ( .A(b[759]), .B(n7201), .Z(n7202) );
  XOR U8495 ( .A(n7204), .B(n7205), .Z(n7201) );
  ANDN U8496 ( .B(n7206), .A(n275), .Z(n7204) );
  XNOR U8497 ( .A(a[758]), .B(n7207), .Z(n275) );
  IV U8498 ( .A(n7205), .Z(n7207) );
  XNOR U8499 ( .A(b[758]), .B(n7205), .Z(n7206) );
  XOR U8500 ( .A(n7208), .B(n7209), .Z(n7205) );
  ANDN U8501 ( .B(n7210), .A(n276), .Z(n7208) );
  XNOR U8502 ( .A(a[757]), .B(n7211), .Z(n276) );
  IV U8503 ( .A(n7209), .Z(n7211) );
  XNOR U8504 ( .A(b[757]), .B(n7209), .Z(n7210) );
  XOR U8505 ( .A(n7212), .B(n7213), .Z(n7209) );
  ANDN U8506 ( .B(n7214), .A(n277), .Z(n7212) );
  XNOR U8507 ( .A(a[756]), .B(n7215), .Z(n277) );
  IV U8508 ( .A(n7213), .Z(n7215) );
  XNOR U8509 ( .A(b[756]), .B(n7213), .Z(n7214) );
  XOR U8510 ( .A(n7216), .B(n7217), .Z(n7213) );
  ANDN U8511 ( .B(n7218), .A(n278), .Z(n7216) );
  XNOR U8512 ( .A(a[755]), .B(n7219), .Z(n278) );
  IV U8513 ( .A(n7217), .Z(n7219) );
  XNOR U8514 ( .A(b[755]), .B(n7217), .Z(n7218) );
  XOR U8515 ( .A(n7220), .B(n7221), .Z(n7217) );
  ANDN U8516 ( .B(n7222), .A(n279), .Z(n7220) );
  XNOR U8517 ( .A(a[754]), .B(n7223), .Z(n279) );
  IV U8518 ( .A(n7221), .Z(n7223) );
  XNOR U8519 ( .A(b[754]), .B(n7221), .Z(n7222) );
  XOR U8520 ( .A(n7224), .B(n7225), .Z(n7221) );
  ANDN U8521 ( .B(n7226), .A(n280), .Z(n7224) );
  XNOR U8522 ( .A(a[753]), .B(n7227), .Z(n280) );
  IV U8523 ( .A(n7225), .Z(n7227) );
  XNOR U8524 ( .A(b[753]), .B(n7225), .Z(n7226) );
  XOR U8525 ( .A(n7228), .B(n7229), .Z(n7225) );
  ANDN U8526 ( .B(n7230), .A(n281), .Z(n7228) );
  XNOR U8527 ( .A(a[752]), .B(n7231), .Z(n281) );
  IV U8528 ( .A(n7229), .Z(n7231) );
  XNOR U8529 ( .A(b[752]), .B(n7229), .Z(n7230) );
  XOR U8530 ( .A(n7232), .B(n7233), .Z(n7229) );
  ANDN U8531 ( .B(n7234), .A(n282), .Z(n7232) );
  XNOR U8532 ( .A(a[751]), .B(n7235), .Z(n282) );
  IV U8533 ( .A(n7233), .Z(n7235) );
  XNOR U8534 ( .A(b[751]), .B(n7233), .Z(n7234) );
  XOR U8535 ( .A(n7236), .B(n7237), .Z(n7233) );
  ANDN U8536 ( .B(n7238), .A(n283), .Z(n7236) );
  XNOR U8537 ( .A(a[750]), .B(n7239), .Z(n283) );
  IV U8538 ( .A(n7237), .Z(n7239) );
  XNOR U8539 ( .A(b[750]), .B(n7237), .Z(n7238) );
  XOR U8540 ( .A(n7240), .B(n7241), .Z(n7237) );
  ANDN U8541 ( .B(n7242), .A(n285), .Z(n7240) );
  XNOR U8542 ( .A(a[749]), .B(n7243), .Z(n285) );
  IV U8543 ( .A(n7241), .Z(n7243) );
  XNOR U8544 ( .A(b[749]), .B(n7241), .Z(n7242) );
  XOR U8545 ( .A(n7244), .B(n7245), .Z(n7241) );
  ANDN U8546 ( .B(n7246), .A(n286), .Z(n7244) );
  XNOR U8547 ( .A(a[748]), .B(n7247), .Z(n286) );
  IV U8548 ( .A(n7245), .Z(n7247) );
  XNOR U8549 ( .A(b[748]), .B(n7245), .Z(n7246) );
  XOR U8550 ( .A(n7248), .B(n7249), .Z(n7245) );
  ANDN U8551 ( .B(n7250), .A(n287), .Z(n7248) );
  XNOR U8552 ( .A(a[747]), .B(n7251), .Z(n287) );
  IV U8553 ( .A(n7249), .Z(n7251) );
  XNOR U8554 ( .A(b[747]), .B(n7249), .Z(n7250) );
  XOR U8555 ( .A(n7252), .B(n7253), .Z(n7249) );
  ANDN U8556 ( .B(n7254), .A(n288), .Z(n7252) );
  XNOR U8557 ( .A(a[746]), .B(n7255), .Z(n288) );
  IV U8558 ( .A(n7253), .Z(n7255) );
  XNOR U8559 ( .A(b[746]), .B(n7253), .Z(n7254) );
  XOR U8560 ( .A(n7256), .B(n7257), .Z(n7253) );
  ANDN U8561 ( .B(n7258), .A(n289), .Z(n7256) );
  XNOR U8562 ( .A(a[745]), .B(n7259), .Z(n289) );
  IV U8563 ( .A(n7257), .Z(n7259) );
  XNOR U8564 ( .A(b[745]), .B(n7257), .Z(n7258) );
  XOR U8565 ( .A(n7260), .B(n7261), .Z(n7257) );
  ANDN U8566 ( .B(n7262), .A(n290), .Z(n7260) );
  XNOR U8567 ( .A(a[744]), .B(n7263), .Z(n290) );
  IV U8568 ( .A(n7261), .Z(n7263) );
  XNOR U8569 ( .A(b[744]), .B(n7261), .Z(n7262) );
  XOR U8570 ( .A(n7264), .B(n7265), .Z(n7261) );
  ANDN U8571 ( .B(n7266), .A(n291), .Z(n7264) );
  XNOR U8572 ( .A(a[743]), .B(n7267), .Z(n291) );
  IV U8573 ( .A(n7265), .Z(n7267) );
  XNOR U8574 ( .A(b[743]), .B(n7265), .Z(n7266) );
  XOR U8575 ( .A(n7268), .B(n7269), .Z(n7265) );
  ANDN U8576 ( .B(n7270), .A(n292), .Z(n7268) );
  XNOR U8577 ( .A(a[742]), .B(n7271), .Z(n292) );
  IV U8578 ( .A(n7269), .Z(n7271) );
  XNOR U8579 ( .A(b[742]), .B(n7269), .Z(n7270) );
  XOR U8580 ( .A(n7272), .B(n7273), .Z(n7269) );
  ANDN U8581 ( .B(n7274), .A(n293), .Z(n7272) );
  XNOR U8582 ( .A(a[741]), .B(n7275), .Z(n293) );
  IV U8583 ( .A(n7273), .Z(n7275) );
  XNOR U8584 ( .A(b[741]), .B(n7273), .Z(n7274) );
  XOR U8585 ( .A(n7276), .B(n7277), .Z(n7273) );
  ANDN U8586 ( .B(n7278), .A(n294), .Z(n7276) );
  XNOR U8587 ( .A(a[740]), .B(n7279), .Z(n294) );
  IV U8588 ( .A(n7277), .Z(n7279) );
  XNOR U8589 ( .A(b[740]), .B(n7277), .Z(n7278) );
  XOR U8590 ( .A(n7280), .B(n7281), .Z(n7277) );
  ANDN U8591 ( .B(n7282), .A(n296), .Z(n7280) );
  XNOR U8592 ( .A(a[739]), .B(n7283), .Z(n296) );
  IV U8593 ( .A(n7281), .Z(n7283) );
  XNOR U8594 ( .A(b[739]), .B(n7281), .Z(n7282) );
  XOR U8595 ( .A(n7284), .B(n7285), .Z(n7281) );
  ANDN U8596 ( .B(n7286), .A(n297), .Z(n7284) );
  XNOR U8597 ( .A(a[738]), .B(n7287), .Z(n297) );
  IV U8598 ( .A(n7285), .Z(n7287) );
  XNOR U8599 ( .A(b[738]), .B(n7285), .Z(n7286) );
  XOR U8600 ( .A(n7288), .B(n7289), .Z(n7285) );
  ANDN U8601 ( .B(n7290), .A(n298), .Z(n7288) );
  XNOR U8602 ( .A(a[737]), .B(n7291), .Z(n298) );
  IV U8603 ( .A(n7289), .Z(n7291) );
  XNOR U8604 ( .A(b[737]), .B(n7289), .Z(n7290) );
  XOR U8605 ( .A(n7292), .B(n7293), .Z(n7289) );
  ANDN U8606 ( .B(n7294), .A(n299), .Z(n7292) );
  XNOR U8607 ( .A(a[736]), .B(n7295), .Z(n299) );
  IV U8608 ( .A(n7293), .Z(n7295) );
  XNOR U8609 ( .A(b[736]), .B(n7293), .Z(n7294) );
  XOR U8610 ( .A(n7296), .B(n7297), .Z(n7293) );
  ANDN U8611 ( .B(n7298), .A(n300), .Z(n7296) );
  XNOR U8612 ( .A(a[735]), .B(n7299), .Z(n300) );
  IV U8613 ( .A(n7297), .Z(n7299) );
  XNOR U8614 ( .A(b[735]), .B(n7297), .Z(n7298) );
  XOR U8615 ( .A(n7300), .B(n7301), .Z(n7297) );
  ANDN U8616 ( .B(n7302), .A(n301), .Z(n7300) );
  XNOR U8617 ( .A(a[734]), .B(n7303), .Z(n301) );
  IV U8618 ( .A(n7301), .Z(n7303) );
  XNOR U8619 ( .A(b[734]), .B(n7301), .Z(n7302) );
  XOR U8620 ( .A(n7304), .B(n7305), .Z(n7301) );
  ANDN U8621 ( .B(n7306), .A(n302), .Z(n7304) );
  XNOR U8622 ( .A(a[733]), .B(n7307), .Z(n302) );
  IV U8623 ( .A(n7305), .Z(n7307) );
  XNOR U8624 ( .A(b[733]), .B(n7305), .Z(n7306) );
  XOR U8625 ( .A(n7308), .B(n7309), .Z(n7305) );
  ANDN U8626 ( .B(n7310), .A(n303), .Z(n7308) );
  XNOR U8627 ( .A(a[732]), .B(n7311), .Z(n303) );
  IV U8628 ( .A(n7309), .Z(n7311) );
  XNOR U8629 ( .A(b[732]), .B(n7309), .Z(n7310) );
  XOR U8630 ( .A(n7312), .B(n7313), .Z(n7309) );
  ANDN U8631 ( .B(n7314), .A(n304), .Z(n7312) );
  XNOR U8632 ( .A(a[731]), .B(n7315), .Z(n304) );
  IV U8633 ( .A(n7313), .Z(n7315) );
  XNOR U8634 ( .A(b[731]), .B(n7313), .Z(n7314) );
  XOR U8635 ( .A(n7316), .B(n7317), .Z(n7313) );
  ANDN U8636 ( .B(n7318), .A(n305), .Z(n7316) );
  XNOR U8637 ( .A(a[730]), .B(n7319), .Z(n305) );
  IV U8638 ( .A(n7317), .Z(n7319) );
  XNOR U8639 ( .A(b[730]), .B(n7317), .Z(n7318) );
  XOR U8640 ( .A(n7320), .B(n7321), .Z(n7317) );
  ANDN U8641 ( .B(n7322), .A(n307), .Z(n7320) );
  XNOR U8642 ( .A(a[729]), .B(n7323), .Z(n307) );
  IV U8643 ( .A(n7321), .Z(n7323) );
  XNOR U8644 ( .A(b[729]), .B(n7321), .Z(n7322) );
  XOR U8645 ( .A(n7324), .B(n7325), .Z(n7321) );
  ANDN U8646 ( .B(n7326), .A(n308), .Z(n7324) );
  XNOR U8647 ( .A(a[728]), .B(n7327), .Z(n308) );
  IV U8648 ( .A(n7325), .Z(n7327) );
  XNOR U8649 ( .A(b[728]), .B(n7325), .Z(n7326) );
  XOR U8650 ( .A(n7328), .B(n7329), .Z(n7325) );
  ANDN U8651 ( .B(n7330), .A(n309), .Z(n7328) );
  XNOR U8652 ( .A(a[727]), .B(n7331), .Z(n309) );
  IV U8653 ( .A(n7329), .Z(n7331) );
  XNOR U8654 ( .A(b[727]), .B(n7329), .Z(n7330) );
  XOR U8655 ( .A(n7332), .B(n7333), .Z(n7329) );
  ANDN U8656 ( .B(n7334), .A(n310), .Z(n7332) );
  XNOR U8657 ( .A(a[726]), .B(n7335), .Z(n310) );
  IV U8658 ( .A(n7333), .Z(n7335) );
  XNOR U8659 ( .A(b[726]), .B(n7333), .Z(n7334) );
  XOR U8660 ( .A(n7336), .B(n7337), .Z(n7333) );
  ANDN U8661 ( .B(n7338), .A(n311), .Z(n7336) );
  XNOR U8662 ( .A(a[725]), .B(n7339), .Z(n311) );
  IV U8663 ( .A(n7337), .Z(n7339) );
  XNOR U8664 ( .A(b[725]), .B(n7337), .Z(n7338) );
  XOR U8665 ( .A(n7340), .B(n7341), .Z(n7337) );
  ANDN U8666 ( .B(n7342), .A(n312), .Z(n7340) );
  XNOR U8667 ( .A(a[724]), .B(n7343), .Z(n312) );
  IV U8668 ( .A(n7341), .Z(n7343) );
  XNOR U8669 ( .A(b[724]), .B(n7341), .Z(n7342) );
  XOR U8670 ( .A(n7344), .B(n7345), .Z(n7341) );
  ANDN U8671 ( .B(n7346), .A(n313), .Z(n7344) );
  XNOR U8672 ( .A(a[723]), .B(n7347), .Z(n313) );
  IV U8673 ( .A(n7345), .Z(n7347) );
  XNOR U8674 ( .A(b[723]), .B(n7345), .Z(n7346) );
  XOR U8675 ( .A(n7348), .B(n7349), .Z(n7345) );
  ANDN U8676 ( .B(n7350), .A(n314), .Z(n7348) );
  XNOR U8677 ( .A(a[722]), .B(n7351), .Z(n314) );
  IV U8678 ( .A(n7349), .Z(n7351) );
  XNOR U8679 ( .A(b[722]), .B(n7349), .Z(n7350) );
  XOR U8680 ( .A(n7352), .B(n7353), .Z(n7349) );
  ANDN U8681 ( .B(n7354), .A(n315), .Z(n7352) );
  XNOR U8682 ( .A(a[721]), .B(n7355), .Z(n315) );
  IV U8683 ( .A(n7353), .Z(n7355) );
  XNOR U8684 ( .A(b[721]), .B(n7353), .Z(n7354) );
  XOR U8685 ( .A(n7356), .B(n7357), .Z(n7353) );
  ANDN U8686 ( .B(n7358), .A(n316), .Z(n7356) );
  XNOR U8687 ( .A(a[720]), .B(n7359), .Z(n316) );
  IV U8688 ( .A(n7357), .Z(n7359) );
  XNOR U8689 ( .A(b[720]), .B(n7357), .Z(n7358) );
  XOR U8690 ( .A(n7360), .B(n7361), .Z(n7357) );
  ANDN U8691 ( .B(n7362), .A(n318), .Z(n7360) );
  XNOR U8692 ( .A(a[719]), .B(n7363), .Z(n318) );
  IV U8693 ( .A(n7361), .Z(n7363) );
  XNOR U8694 ( .A(b[719]), .B(n7361), .Z(n7362) );
  XOR U8695 ( .A(n7364), .B(n7365), .Z(n7361) );
  ANDN U8696 ( .B(n7366), .A(n319), .Z(n7364) );
  XNOR U8697 ( .A(a[718]), .B(n7367), .Z(n319) );
  IV U8698 ( .A(n7365), .Z(n7367) );
  XNOR U8699 ( .A(b[718]), .B(n7365), .Z(n7366) );
  XOR U8700 ( .A(n7368), .B(n7369), .Z(n7365) );
  ANDN U8701 ( .B(n7370), .A(n320), .Z(n7368) );
  XNOR U8702 ( .A(a[717]), .B(n7371), .Z(n320) );
  IV U8703 ( .A(n7369), .Z(n7371) );
  XNOR U8704 ( .A(b[717]), .B(n7369), .Z(n7370) );
  XOR U8705 ( .A(n7372), .B(n7373), .Z(n7369) );
  ANDN U8706 ( .B(n7374), .A(n321), .Z(n7372) );
  XNOR U8707 ( .A(a[716]), .B(n7375), .Z(n321) );
  IV U8708 ( .A(n7373), .Z(n7375) );
  XNOR U8709 ( .A(b[716]), .B(n7373), .Z(n7374) );
  XOR U8710 ( .A(n7376), .B(n7377), .Z(n7373) );
  ANDN U8711 ( .B(n7378), .A(n322), .Z(n7376) );
  XNOR U8712 ( .A(a[715]), .B(n7379), .Z(n322) );
  IV U8713 ( .A(n7377), .Z(n7379) );
  XNOR U8714 ( .A(b[715]), .B(n7377), .Z(n7378) );
  XOR U8715 ( .A(n7380), .B(n7381), .Z(n7377) );
  ANDN U8716 ( .B(n7382), .A(n323), .Z(n7380) );
  XNOR U8717 ( .A(a[714]), .B(n7383), .Z(n323) );
  IV U8718 ( .A(n7381), .Z(n7383) );
  XNOR U8719 ( .A(b[714]), .B(n7381), .Z(n7382) );
  XOR U8720 ( .A(n7384), .B(n7385), .Z(n7381) );
  ANDN U8721 ( .B(n7386), .A(n324), .Z(n7384) );
  XNOR U8722 ( .A(a[713]), .B(n7387), .Z(n324) );
  IV U8723 ( .A(n7385), .Z(n7387) );
  XNOR U8724 ( .A(b[713]), .B(n7385), .Z(n7386) );
  XOR U8725 ( .A(n7388), .B(n7389), .Z(n7385) );
  ANDN U8726 ( .B(n7390), .A(n325), .Z(n7388) );
  XNOR U8727 ( .A(a[712]), .B(n7391), .Z(n325) );
  IV U8728 ( .A(n7389), .Z(n7391) );
  XNOR U8729 ( .A(b[712]), .B(n7389), .Z(n7390) );
  XOR U8730 ( .A(n7392), .B(n7393), .Z(n7389) );
  ANDN U8731 ( .B(n7394), .A(n326), .Z(n7392) );
  XNOR U8732 ( .A(a[711]), .B(n7395), .Z(n326) );
  IV U8733 ( .A(n7393), .Z(n7395) );
  XNOR U8734 ( .A(b[711]), .B(n7393), .Z(n7394) );
  XOR U8735 ( .A(n7396), .B(n7397), .Z(n7393) );
  ANDN U8736 ( .B(n7398), .A(n327), .Z(n7396) );
  XNOR U8737 ( .A(a[710]), .B(n7399), .Z(n327) );
  IV U8738 ( .A(n7397), .Z(n7399) );
  XNOR U8739 ( .A(b[710]), .B(n7397), .Z(n7398) );
  XOR U8740 ( .A(n7400), .B(n7401), .Z(n7397) );
  ANDN U8741 ( .B(n7402), .A(n329), .Z(n7400) );
  XNOR U8742 ( .A(a[709]), .B(n7403), .Z(n329) );
  IV U8743 ( .A(n7401), .Z(n7403) );
  XNOR U8744 ( .A(b[709]), .B(n7401), .Z(n7402) );
  XOR U8745 ( .A(n7404), .B(n7405), .Z(n7401) );
  ANDN U8746 ( .B(n7406), .A(n330), .Z(n7404) );
  XNOR U8747 ( .A(a[708]), .B(n7407), .Z(n330) );
  IV U8748 ( .A(n7405), .Z(n7407) );
  XNOR U8749 ( .A(b[708]), .B(n7405), .Z(n7406) );
  XOR U8750 ( .A(n7408), .B(n7409), .Z(n7405) );
  ANDN U8751 ( .B(n7410), .A(n331), .Z(n7408) );
  XNOR U8752 ( .A(a[707]), .B(n7411), .Z(n331) );
  IV U8753 ( .A(n7409), .Z(n7411) );
  XNOR U8754 ( .A(b[707]), .B(n7409), .Z(n7410) );
  XOR U8755 ( .A(n7412), .B(n7413), .Z(n7409) );
  ANDN U8756 ( .B(n7414), .A(n332), .Z(n7412) );
  XNOR U8757 ( .A(a[706]), .B(n7415), .Z(n332) );
  IV U8758 ( .A(n7413), .Z(n7415) );
  XNOR U8759 ( .A(b[706]), .B(n7413), .Z(n7414) );
  XOR U8760 ( .A(n7416), .B(n7417), .Z(n7413) );
  ANDN U8761 ( .B(n7418), .A(n333), .Z(n7416) );
  XNOR U8762 ( .A(a[705]), .B(n7419), .Z(n333) );
  IV U8763 ( .A(n7417), .Z(n7419) );
  XNOR U8764 ( .A(b[705]), .B(n7417), .Z(n7418) );
  XOR U8765 ( .A(n7420), .B(n7421), .Z(n7417) );
  ANDN U8766 ( .B(n7422), .A(n334), .Z(n7420) );
  XNOR U8767 ( .A(a[704]), .B(n7423), .Z(n334) );
  IV U8768 ( .A(n7421), .Z(n7423) );
  XNOR U8769 ( .A(b[704]), .B(n7421), .Z(n7422) );
  XOR U8770 ( .A(n7424), .B(n7425), .Z(n7421) );
  ANDN U8771 ( .B(n7426), .A(n335), .Z(n7424) );
  XNOR U8772 ( .A(a[703]), .B(n7427), .Z(n335) );
  IV U8773 ( .A(n7425), .Z(n7427) );
  XNOR U8774 ( .A(b[703]), .B(n7425), .Z(n7426) );
  XOR U8775 ( .A(n7428), .B(n7429), .Z(n7425) );
  ANDN U8776 ( .B(n7430), .A(n336), .Z(n7428) );
  XNOR U8777 ( .A(a[702]), .B(n7431), .Z(n336) );
  IV U8778 ( .A(n7429), .Z(n7431) );
  XNOR U8779 ( .A(b[702]), .B(n7429), .Z(n7430) );
  XOR U8780 ( .A(n7432), .B(n7433), .Z(n7429) );
  ANDN U8781 ( .B(n7434), .A(n337), .Z(n7432) );
  XNOR U8782 ( .A(a[701]), .B(n7435), .Z(n337) );
  IV U8783 ( .A(n7433), .Z(n7435) );
  XNOR U8784 ( .A(b[701]), .B(n7433), .Z(n7434) );
  XOR U8785 ( .A(n7436), .B(n7437), .Z(n7433) );
  ANDN U8786 ( .B(n7438), .A(n338), .Z(n7436) );
  XNOR U8787 ( .A(a[700]), .B(n7439), .Z(n338) );
  IV U8788 ( .A(n7437), .Z(n7439) );
  XNOR U8789 ( .A(b[700]), .B(n7437), .Z(n7438) );
  XOR U8790 ( .A(n7440), .B(n7441), .Z(n7437) );
  ANDN U8791 ( .B(n7442), .A(n341), .Z(n7440) );
  XNOR U8792 ( .A(a[699]), .B(n7443), .Z(n341) );
  IV U8793 ( .A(n7441), .Z(n7443) );
  XNOR U8794 ( .A(b[699]), .B(n7441), .Z(n7442) );
  XOR U8795 ( .A(n7444), .B(n7445), .Z(n7441) );
  ANDN U8796 ( .B(n7446), .A(n342), .Z(n7444) );
  XNOR U8797 ( .A(a[698]), .B(n7447), .Z(n342) );
  IV U8798 ( .A(n7445), .Z(n7447) );
  XNOR U8799 ( .A(b[698]), .B(n7445), .Z(n7446) );
  XOR U8800 ( .A(n7448), .B(n7449), .Z(n7445) );
  ANDN U8801 ( .B(n7450), .A(n343), .Z(n7448) );
  XNOR U8802 ( .A(a[697]), .B(n7451), .Z(n343) );
  IV U8803 ( .A(n7449), .Z(n7451) );
  XNOR U8804 ( .A(b[697]), .B(n7449), .Z(n7450) );
  XOR U8805 ( .A(n7452), .B(n7453), .Z(n7449) );
  ANDN U8806 ( .B(n7454), .A(n344), .Z(n7452) );
  XNOR U8807 ( .A(a[696]), .B(n7455), .Z(n344) );
  IV U8808 ( .A(n7453), .Z(n7455) );
  XNOR U8809 ( .A(b[696]), .B(n7453), .Z(n7454) );
  XOR U8810 ( .A(n7456), .B(n7457), .Z(n7453) );
  ANDN U8811 ( .B(n7458), .A(n345), .Z(n7456) );
  XNOR U8812 ( .A(a[695]), .B(n7459), .Z(n345) );
  IV U8813 ( .A(n7457), .Z(n7459) );
  XNOR U8814 ( .A(b[695]), .B(n7457), .Z(n7458) );
  XOR U8815 ( .A(n7460), .B(n7461), .Z(n7457) );
  ANDN U8816 ( .B(n7462), .A(n346), .Z(n7460) );
  XNOR U8817 ( .A(a[694]), .B(n7463), .Z(n346) );
  IV U8818 ( .A(n7461), .Z(n7463) );
  XNOR U8819 ( .A(b[694]), .B(n7461), .Z(n7462) );
  XOR U8820 ( .A(n7464), .B(n7465), .Z(n7461) );
  ANDN U8821 ( .B(n7466), .A(n347), .Z(n7464) );
  XNOR U8822 ( .A(a[693]), .B(n7467), .Z(n347) );
  IV U8823 ( .A(n7465), .Z(n7467) );
  XNOR U8824 ( .A(b[693]), .B(n7465), .Z(n7466) );
  XOR U8825 ( .A(n7468), .B(n7469), .Z(n7465) );
  ANDN U8826 ( .B(n7470), .A(n348), .Z(n7468) );
  XNOR U8827 ( .A(a[692]), .B(n7471), .Z(n348) );
  IV U8828 ( .A(n7469), .Z(n7471) );
  XNOR U8829 ( .A(b[692]), .B(n7469), .Z(n7470) );
  XOR U8830 ( .A(n7472), .B(n7473), .Z(n7469) );
  ANDN U8831 ( .B(n7474), .A(n349), .Z(n7472) );
  XNOR U8832 ( .A(a[691]), .B(n7475), .Z(n349) );
  IV U8833 ( .A(n7473), .Z(n7475) );
  XNOR U8834 ( .A(b[691]), .B(n7473), .Z(n7474) );
  XOR U8835 ( .A(n7476), .B(n7477), .Z(n7473) );
  ANDN U8836 ( .B(n7478), .A(n350), .Z(n7476) );
  XNOR U8837 ( .A(a[690]), .B(n7479), .Z(n350) );
  IV U8838 ( .A(n7477), .Z(n7479) );
  XNOR U8839 ( .A(b[690]), .B(n7477), .Z(n7478) );
  XOR U8840 ( .A(n7480), .B(n7481), .Z(n7477) );
  ANDN U8841 ( .B(n7482), .A(n352), .Z(n7480) );
  XNOR U8842 ( .A(a[689]), .B(n7483), .Z(n352) );
  IV U8843 ( .A(n7481), .Z(n7483) );
  XNOR U8844 ( .A(b[689]), .B(n7481), .Z(n7482) );
  XOR U8845 ( .A(n7484), .B(n7485), .Z(n7481) );
  ANDN U8846 ( .B(n7486), .A(n353), .Z(n7484) );
  XNOR U8847 ( .A(a[688]), .B(n7487), .Z(n353) );
  IV U8848 ( .A(n7485), .Z(n7487) );
  XNOR U8849 ( .A(b[688]), .B(n7485), .Z(n7486) );
  XOR U8850 ( .A(n7488), .B(n7489), .Z(n7485) );
  ANDN U8851 ( .B(n7490), .A(n354), .Z(n7488) );
  XNOR U8852 ( .A(a[687]), .B(n7491), .Z(n354) );
  IV U8853 ( .A(n7489), .Z(n7491) );
  XNOR U8854 ( .A(b[687]), .B(n7489), .Z(n7490) );
  XOR U8855 ( .A(n7492), .B(n7493), .Z(n7489) );
  ANDN U8856 ( .B(n7494), .A(n355), .Z(n7492) );
  XNOR U8857 ( .A(a[686]), .B(n7495), .Z(n355) );
  IV U8858 ( .A(n7493), .Z(n7495) );
  XNOR U8859 ( .A(b[686]), .B(n7493), .Z(n7494) );
  XOR U8860 ( .A(n7496), .B(n7497), .Z(n7493) );
  ANDN U8861 ( .B(n7498), .A(n356), .Z(n7496) );
  XNOR U8862 ( .A(a[685]), .B(n7499), .Z(n356) );
  IV U8863 ( .A(n7497), .Z(n7499) );
  XNOR U8864 ( .A(b[685]), .B(n7497), .Z(n7498) );
  XOR U8865 ( .A(n7500), .B(n7501), .Z(n7497) );
  ANDN U8866 ( .B(n7502), .A(n357), .Z(n7500) );
  XNOR U8867 ( .A(a[684]), .B(n7503), .Z(n357) );
  IV U8868 ( .A(n7501), .Z(n7503) );
  XNOR U8869 ( .A(b[684]), .B(n7501), .Z(n7502) );
  XOR U8870 ( .A(n7504), .B(n7505), .Z(n7501) );
  ANDN U8871 ( .B(n7506), .A(n358), .Z(n7504) );
  XNOR U8872 ( .A(a[683]), .B(n7507), .Z(n358) );
  IV U8873 ( .A(n7505), .Z(n7507) );
  XNOR U8874 ( .A(b[683]), .B(n7505), .Z(n7506) );
  XOR U8875 ( .A(n7508), .B(n7509), .Z(n7505) );
  ANDN U8876 ( .B(n7510), .A(n359), .Z(n7508) );
  XNOR U8877 ( .A(a[682]), .B(n7511), .Z(n359) );
  IV U8878 ( .A(n7509), .Z(n7511) );
  XNOR U8879 ( .A(b[682]), .B(n7509), .Z(n7510) );
  XOR U8880 ( .A(n7512), .B(n7513), .Z(n7509) );
  ANDN U8881 ( .B(n7514), .A(n360), .Z(n7512) );
  XNOR U8882 ( .A(a[681]), .B(n7515), .Z(n360) );
  IV U8883 ( .A(n7513), .Z(n7515) );
  XNOR U8884 ( .A(b[681]), .B(n7513), .Z(n7514) );
  XOR U8885 ( .A(n7516), .B(n7517), .Z(n7513) );
  ANDN U8886 ( .B(n7518), .A(n361), .Z(n7516) );
  XNOR U8887 ( .A(a[680]), .B(n7519), .Z(n361) );
  IV U8888 ( .A(n7517), .Z(n7519) );
  XNOR U8889 ( .A(b[680]), .B(n7517), .Z(n7518) );
  XOR U8890 ( .A(n7520), .B(n7521), .Z(n7517) );
  ANDN U8891 ( .B(n7522), .A(n363), .Z(n7520) );
  XNOR U8892 ( .A(a[679]), .B(n7523), .Z(n363) );
  IV U8893 ( .A(n7521), .Z(n7523) );
  XNOR U8894 ( .A(b[679]), .B(n7521), .Z(n7522) );
  XOR U8895 ( .A(n7524), .B(n7525), .Z(n7521) );
  ANDN U8896 ( .B(n7526), .A(n364), .Z(n7524) );
  XNOR U8897 ( .A(a[678]), .B(n7527), .Z(n364) );
  IV U8898 ( .A(n7525), .Z(n7527) );
  XNOR U8899 ( .A(b[678]), .B(n7525), .Z(n7526) );
  XOR U8900 ( .A(n7528), .B(n7529), .Z(n7525) );
  ANDN U8901 ( .B(n7530), .A(n365), .Z(n7528) );
  XNOR U8902 ( .A(a[677]), .B(n7531), .Z(n365) );
  IV U8903 ( .A(n7529), .Z(n7531) );
  XNOR U8904 ( .A(b[677]), .B(n7529), .Z(n7530) );
  XOR U8905 ( .A(n7532), .B(n7533), .Z(n7529) );
  ANDN U8906 ( .B(n7534), .A(n366), .Z(n7532) );
  XNOR U8907 ( .A(a[676]), .B(n7535), .Z(n366) );
  IV U8908 ( .A(n7533), .Z(n7535) );
  XNOR U8909 ( .A(b[676]), .B(n7533), .Z(n7534) );
  XOR U8910 ( .A(n7536), .B(n7537), .Z(n7533) );
  ANDN U8911 ( .B(n7538), .A(n367), .Z(n7536) );
  XNOR U8912 ( .A(a[675]), .B(n7539), .Z(n367) );
  IV U8913 ( .A(n7537), .Z(n7539) );
  XNOR U8914 ( .A(b[675]), .B(n7537), .Z(n7538) );
  XOR U8915 ( .A(n7540), .B(n7541), .Z(n7537) );
  ANDN U8916 ( .B(n7542), .A(n368), .Z(n7540) );
  XNOR U8917 ( .A(a[674]), .B(n7543), .Z(n368) );
  IV U8918 ( .A(n7541), .Z(n7543) );
  XNOR U8919 ( .A(b[674]), .B(n7541), .Z(n7542) );
  XOR U8920 ( .A(n7544), .B(n7545), .Z(n7541) );
  ANDN U8921 ( .B(n7546), .A(n369), .Z(n7544) );
  XNOR U8922 ( .A(a[673]), .B(n7547), .Z(n369) );
  IV U8923 ( .A(n7545), .Z(n7547) );
  XNOR U8924 ( .A(b[673]), .B(n7545), .Z(n7546) );
  XOR U8925 ( .A(n7548), .B(n7549), .Z(n7545) );
  ANDN U8926 ( .B(n7550), .A(n370), .Z(n7548) );
  XNOR U8927 ( .A(a[672]), .B(n7551), .Z(n370) );
  IV U8928 ( .A(n7549), .Z(n7551) );
  XNOR U8929 ( .A(b[672]), .B(n7549), .Z(n7550) );
  XOR U8930 ( .A(n7552), .B(n7553), .Z(n7549) );
  ANDN U8931 ( .B(n7554), .A(n371), .Z(n7552) );
  XNOR U8932 ( .A(a[671]), .B(n7555), .Z(n371) );
  IV U8933 ( .A(n7553), .Z(n7555) );
  XNOR U8934 ( .A(b[671]), .B(n7553), .Z(n7554) );
  XOR U8935 ( .A(n7556), .B(n7557), .Z(n7553) );
  ANDN U8936 ( .B(n7558), .A(n372), .Z(n7556) );
  XNOR U8937 ( .A(a[670]), .B(n7559), .Z(n372) );
  IV U8938 ( .A(n7557), .Z(n7559) );
  XNOR U8939 ( .A(b[670]), .B(n7557), .Z(n7558) );
  XOR U8940 ( .A(n7560), .B(n7561), .Z(n7557) );
  ANDN U8941 ( .B(n7562), .A(n374), .Z(n7560) );
  XNOR U8942 ( .A(a[669]), .B(n7563), .Z(n374) );
  IV U8943 ( .A(n7561), .Z(n7563) );
  XNOR U8944 ( .A(b[669]), .B(n7561), .Z(n7562) );
  XOR U8945 ( .A(n7564), .B(n7565), .Z(n7561) );
  ANDN U8946 ( .B(n7566), .A(n375), .Z(n7564) );
  XNOR U8947 ( .A(a[668]), .B(n7567), .Z(n375) );
  IV U8948 ( .A(n7565), .Z(n7567) );
  XNOR U8949 ( .A(b[668]), .B(n7565), .Z(n7566) );
  XOR U8950 ( .A(n7568), .B(n7569), .Z(n7565) );
  ANDN U8951 ( .B(n7570), .A(n376), .Z(n7568) );
  XNOR U8952 ( .A(a[667]), .B(n7571), .Z(n376) );
  IV U8953 ( .A(n7569), .Z(n7571) );
  XNOR U8954 ( .A(b[667]), .B(n7569), .Z(n7570) );
  XOR U8955 ( .A(n7572), .B(n7573), .Z(n7569) );
  ANDN U8956 ( .B(n7574), .A(n377), .Z(n7572) );
  XNOR U8957 ( .A(a[666]), .B(n7575), .Z(n377) );
  IV U8958 ( .A(n7573), .Z(n7575) );
  XNOR U8959 ( .A(b[666]), .B(n7573), .Z(n7574) );
  XOR U8960 ( .A(n7576), .B(n7577), .Z(n7573) );
  ANDN U8961 ( .B(n7578), .A(n378), .Z(n7576) );
  XNOR U8962 ( .A(a[665]), .B(n7579), .Z(n378) );
  IV U8963 ( .A(n7577), .Z(n7579) );
  XNOR U8964 ( .A(b[665]), .B(n7577), .Z(n7578) );
  XOR U8965 ( .A(n7580), .B(n7581), .Z(n7577) );
  ANDN U8966 ( .B(n7582), .A(n379), .Z(n7580) );
  XNOR U8967 ( .A(a[664]), .B(n7583), .Z(n379) );
  IV U8968 ( .A(n7581), .Z(n7583) );
  XNOR U8969 ( .A(b[664]), .B(n7581), .Z(n7582) );
  XOR U8970 ( .A(n7584), .B(n7585), .Z(n7581) );
  ANDN U8971 ( .B(n7586), .A(n380), .Z(n7584) );
  XNOR U8972 ( .A(a[663]), .B(n7587), .Z(n380) );
  IV U8973 ( .A(n7585), .Z(n7587) );
  XNOR U8974 ( .A(b[663]), .B(n7585), .Z(n7586) );
  XOR U8975 ( .A(n7588), .B(n7589), .Z(n7585) );
  ANDN U8976 ( .B(n7590), .A(n381), .Z(n7588) );
  XNOR U8977 ( .A(a[662]), .B(n7591), .Z(n381) );
  IV U8978 ( .A(n7589), .Z(n7591) );
  XNOR U8979 ( .A(b[662]), .B(n7589), .Z(n7590) );
  XOR U8980 ( .A(n7592), .B(n7593), .Z(n7589) );
  ANDN U8981 ( .B(n7594), .A(n382), .Z(n7592) );
  XNOR U8982 ( .A(a[661]), .B(n7595), .Z(n382) );
  IV U8983 ( .A(n7593), .Z(n7595) );
  XNOR U8984 ( .A(b[661]), .B(n7593), .Z(n7594) );
  XOR U8985 ( .A(n7596), .B(n7597), .Z(n7593) );
  ANDN U8986 ( .B(n7598), .A(n383), .Z(n7596) );
  XNOR U8987 ( .A(a[660]), .B(n7599), .Z(n383) );
  IV U8988 ( .A(n7597), .Z(n7599) );
  XNOR U8989 ( .A(b[660]), .B(n7597), .Z(n7598) );
  XOR U8990 ( .A(n7600), .B(n7601), .Z(n7597) );
  ANDN U8991 ( .B(n7602), .A(n385), .Z(n7600) );
  XNOR U8992 ( .A(a[659]), .B(n7603), .Z(n385) );
  IV U8993 ( .A(n7601), .Z(n7603) );
  XNOR U8994 ( .A(b[659]), .B(n7601), .Z(n7602) );
  XOR U8995 ( .A(n7604), .B(n7605), .Z(n7601) );
  ANDN U8996 ( .B(n7606), .A(n386), .Z(n7604) );
  XNOR U8997 ( .A(a[658]), .B(n7607), .Z(n386) );
  IV U8998 ( .A(n7605), .Z(n7607) );
  XNOR U8999 ( .A(b[658]), .B(n7605), .Z(n7606) );
  XOR U9000 ( .A(n7608), .B(n7609), .Z(n7605) );
  ANDN U9001 ( .B(n7610), .A(n387), .Z(n7608) );
  XNOR U9002 ( .A(a[657]), .B(n7611), .Z(n387) );
  IV U9003 ( .A(n7609), .Z(n7611) );
  XNOR U9004 ( .A(b[657]), .B(n7609), .Z(n7610) );
  XOR U9005 ( .A(n7612), .B(n7613), .Z(n7609) );
  ANDN U9006 ( .B(n7614), .A(n388), .Z(n7612) );
  XNOR U9007 ( .A(a[656]), .B(n7615), .Z(n388) );
  IV U9008 ( .A(n7613), .Z(n7615) );
  XNOR U9009 ( .A(b[656]), .B(n7613), .Z(n7614) );
  XOR U9010 ( .A(n7616), .B(n7617), .Z(n7613) );
  ANDN U9011 ( .B(n7618), .A(n389), .Z(n7616) );
  XNOR U9012 ( .A(a[655]), .B(n7619), .Z(n389) );
  IV U9013 ( .A(n7617), .Z(n7619) );
  XNOR U9014 ( .A(b[655]), .B(n7617), .Z(n7618) );
  XOR U9015 ( .A(n7620), .B(n7621), .Z(n7617) );
  ANDN U9016 ( .B(n7622), .A(n390), .Z(n7620) );
  XNOR U9017 ( .A(a[654]), .B(n7623), .Z(n390) );
  IV U9018 ( .A(n7621), .Z(n7623) );
  XNOR U9019 ( .A(b[654]), .B(n7621), .Z(n7622) );
  XOR U9020 ( .A(n7624), .B(n7625), .Z(n7621) );
  ANDN U9021 ( .B(n7626), .A(n391), .Z(n7624) );
  XNOR U9022 ( .A(a[653]), .B(n7627), .Z(n391) );
  IV U9023 ( .A(n7625), .Z(n7627) );
  XNOR U9024 ( .A(b[653]), .B(n7625), .Z(n7626) );
  XOR U9025 ( .A(n7628), .B(n7629), .Z(n7625) );
  ANDN U9026 ( .B(n7630), .A(n392), .Z(n7628) );
  XNOR U9027 ( .A(a[652]), .B(n7631), .Z(n392) );
  IV U9028 ( .A(n7629), .Z(n7631) );
  XNOR U9029 ( .A(b[652]), .B(n7629), .Z(n7630) );
  XOR U9030 ( .A(n7632), .B(n7633), .Z(n7629) );
  ANDN U9031 ( .B(n7634), .A(n393), .Z(n7632) );
  XNOR U9032 ( .A(a[651]), .B(n7635), .Z(n393) );
  IV U9033 ( .A(n7633), .Z(n7635) );
  XNOR U9034 ( .A(b[651]), .B(n7633), .Z(n7634) );
  XOR U9035 ( .A(n7636), .B(n7637), .Z(n7633) );
  ANDN U9036 ( .B(n7638), .A(n394), .Z(n7636) );
  XNOR U9037 ( .A(a[650]), .B(n7639), .Z(n394) );
  IV U9038 ( .A(n7637), .Z(n7639) );
  XNOR U9039 ( .A(b[650]), .B(n7637), .Z(n7638) );
  XOR U9040 ( .A(n7640), .B(n7641), .Z(n7637) );
  ANDN U9041 ( .B(n7642), .A(n396), .Z(n7640) );
  XNOR U9042 ( .A(a[649]), .B(n7643), .Z(n396) );
  IV U9043 ( .A(n7641), .Z(n7643) );
  XNOR U9044 ( .A(b[649]), .B(n7641), .Z(n7642) );
  XOR U9045 ( .A(n7644), .B(n7645), .Z(n7641) );
  ANDN U9046 ( .B(n7646), .A(n397), .Z(n7644) );
  XNOR U9047 ( .A(a[648]), .B(n7647), .Z(n397) );
  IV U9048 ( .A(n7645), .Z(n7647) );
  XNOR U9049 ( .A(b[648]), .B(n7645), .Z(n7646) );
  XOR U9050 ( .A(n7648), .B(n7649), .Z(n7645) );
  ANDN U9051 ( .B(n7650), .A(n398), .Z(n7648) );
  XNOR U9052 ( .A(a[647]), .B(n7651), .Z(n398) );
  IV U9053 ( .A(n7649), .Z(n7651) );
  XNOR U9054 ( .A(b[647]), .B(n7649), .Z(n7650) );
  XOR U9055 ( .A(n7652), .B(n7653), .Z(n7649) );
  ANDN U9056 ( .B(n7654), .A(n399), .Z(n7652) );
  XNOR U9057 ( .A(a[646]), .B(n7655), .Z(n399) );
  IV U9058 ( .A(n7653), .Z(n7655) );
  XNOR U9059 ( .A(b[646]), .B(n7653), .Z(n7654) );
  XOR U9060 ( .A(n7656), .B(n7657), .Z(n7653) );
  ANDN U9061 ( .B(n7658), .A(n400), .Z(n7656) );
  XNOR U9062 ( .A(a[645]), .B(n7659), .Z(n400) );
  IV U9063 ( .A(n7657), .Z(n7659) );
  XNOR U9064 ( .A(b[645]), .B(n7657), .Z(n7658) );
  XOR U9065 ( .A(n7660), .B(n7661), .Z(n7657) );
  ANDN U9066 ( .B(n7662), .A(n401), .Z(n7660) );
  XNOR U9067 ( .A(a[644]), .B(n7663), .Z(n401) );
  IV U9068 ( .A(n7661), .Z(n7663) );
  XNOR U9069 ( .A(b[644]), .B(n7661), .Z(n7662) );
  XOR U9070 ( .A(n7664), .B(n7665), .Z(n7661) );
  ANDN U9071 ( .B(n7666), .A(n402), .Z(n7664) );
  XNOR U9072 ( .A(a[643]), .B(n7667), .Z(n402) );
  IV U9073 ( .A(n7665), .Z(n7667) );
  XNOR U9074 ( .A(b[643]), .B(n7665), .Z(n7666) );
  XOR U9075 ( .A(n7668), .B(n7669), .Z(n7665) );
  ANDN U9076 ( .B(n7670), .A(n403), .Z(n7668) );
  XNOR U9077 ( .A(a[642]), .B(n7671), .Z(n403) );
  IV U9078 ( .A(n7669), .Z(n7671) );
  XNOR U9079 ( .A(b[642]), .B(n7669), .Z(n7670) );
  XOR U9080 ( .A(n7672), .B(n7673), .Z(n7669) );
  ANDN U9081 ( .B(n7674), .A(n404), .Z(n7672) );
  XNOR U9082 ( .A(a[641]), .B(n7675), .Z(n404) );
  IV U9083 ( .A(n7673), .Z(n7675) );
  XNOR U9084 ( .A(b[641]), .B(n7673), .Z(n7674) );
  XOR U9085 ( .A(n7676), .B(n7677), .Z(n7673) );
  ANDN U9086 ( .B(n7678), .A(n405), .Z(n7676) );
  XNOR U9087 ( .A(a[640]), .B(n7679), .Z(n405) );
  IV U9088 ( .A(n7677), .Z(n7679) );
  XNOR U9089 ( .A(b[640]), .B(n7677), .Z(n7678) );
  XOR U9090 ( .A(n7680), .B(n7681), .Z(n7677) );
  ANDN U9091 ( .B(n7682), .A(n407), .Z(n7680) );
  XNOR U9092 ( .A(a[639]), .B(n7683), .Z(n407) );
  IV U9093 ( .A(n7681), .Z(n7683) );
  XNOR U9094 ( .A(b[639]), .B(n7681), .Z(n7682) );
  XOR U9095 ( .A(n7684), .B(n7685), .Z(n7681) );
  ANDN U9096 ( .B(n7686), .A(n408), .Z(n7684) );
  XNOR U9097 ( .A(a[638]), .B(n7687), .Z(n408) );
  IV U9098 ( .A(n7685), .Z(n7687) );
  XNOR U9099 ( .A(b[638]), .B(n7685), .Z(n7686) );
  XOR U9100 ( .A(n7688), .B(n7689), .Z(n7685) );
  ANDN U9101 ( .B(n7690), .A(n409), .Z(n7688) );
  XNOR U9102 ( .A(a[637]), .B(n7691), .Z(n409) );
  IV U9103 ( .A(n7689), .Z(n7691) );
  XNOR U9104 ( .A(b[637]), .B(n7689), .Z(n7690) );
  XOR U9105 ( .A(n7692), .B(n7693), .Z(n7689) );
  ANDN U9106 ( .B(n7694), .A(n410), .Z(n7692) );
  XNOR U9107 ( .A(a[636]), .B(n7695), .Z(n410) );
  IV U9108 ( .A(n7693), .Z(n7695) );
  XNOR U9109 ( .A(b[636]), .B(n7693), .Z(n7694) );
  XOR U9110 ( .A(n7696), .B(n7697), .Z(n7693) );
  ANDN U9111 ( .B(n7698), .A(n411), .Z(n7696) );
  XNOR U9112 ( .A(a[635]), .B(n7699), .Z(n411) );
  IV U9113 ( .A(n7697), .Z(n7699) );
  XNOR U9114 ( .A(b[635]), .B(n7697), .Z(n7698) );
  XOR U9115 ( .A(n7700), .B(n7701), .Z(n7697) );
  ANDN U9116 ( .B(n7702), .A(n412), .Z(n7700) );
  XNOR U9117 ( .A(a[634]), .B(n7703), .Z(n412) );
  IV U9118 ( .A(n7701), .Z(n7703) );
  XNOR U9119 ( .A(b[634]), .B(n7701), .Z(n7702) );
  XOR U9120 ( .A(n7704), .B(n7705), .Z(n7701) );
  ANDN U9121 ( .B(n7706), .A(n413), .Z(n7704) );
  XNOR U9122 ( .A(a[633]), .B(n7707), .Z(n413) );
  IV U9123 ( .A(n7705), .Z(n7707) );
  XNOR U9124 ( .A(b[633]), .B(n7705), .Z(n7706) );
  XOR U9125 ( .A(n7708), .B(n7709), .Z(n7705) );
  ANDN U9126 ( .B(n7710), .A(n414), .Z(n7708) );
  XNOR U9127 ( .A(a[632]), .B(n7711), .Z(n414) );
  IV U9128 ( .A(n7709), .Z(n7711) );
  XNOR U9129 ( .A(b[632]), .B(n7709), .Z(n7710) );
  XOR U9130 ( .A(n7712), .B(n7713), .Z(n7709) );
  ANDN U9131 ( .B(n7714), .A(n415), .Z(n7712) );
  XNOR U9132 ( .A(a[631]), .B(n7715), .Z(n415) );
  IV U9133 ( .A(n7713), .Z(n7715) );
  XNOR U9134 ( .A(b[631]), .B(n7713), .Z(n7714) );
  XOR U9135 ( .A(n7716), .B(n7717), .Z(n7713) );
  ANDN U9136 ( .B(n7718), .A(n416), .Z(n7716) );
  XNOR U9137 ( .A(a[630]), .B(n7719), .Z(n416) );
  IV U9138 ( .A(n7717), .Z(n7719) );
  XNOR U9139 ( .A(b[630]), .B(n7717), .Z(n7718) );
  XOR U9140 ( .A(n7720), .B(n7721), .Z(n7717) );
  ANDN U9141 ( .B(n7722), .A(n418), .Z(n7720) );
  XNOR U9142 ( .A(a[629]), .B(n7723), .Z(n418) );
  IV U9143 ( .A(n7721), .Z(n7723) );
  XNOR U9144 ( .A(b[629]), .B(n7721), .Z(n7722) );
  XOR U9145 ( .A(n7724), .B(n7725), .Z(n7721) );
  ANDN U9146 ( .B(n7726), .A(n419), .Z(n7724) );
  XNOR U9147 ( .A(a[628]), .B(n7727), .Z(n419) );
  IV U9148 ( .A(n7725), .Z(n7727) );
  XNOR U9149 ( .A(b[628]), .B(n7725), .Z(n7726) );
  XOR U9150 ( .A(n7728), .B(n7729), .Z(n7725) );
  ANDN U9151 ( .B(n7730), .A(n420), .Z(n7728) );
  XNOR U9152 ( .A(a[627]), .B(n7731), .Z(n420) );
  IV U9153 ( .A(n7729), .Z(n7731) );
  XNOR U9154 ( .A(b[627]), .B(n7729), .Z(n7730) );
  XOR U9155 ( .A(n7732), .B(n7733), .Z(n7729) );
  ANDN U9156 ( .B(n7734), .A(n421), .Z(n7732) );
  XNOR U9157 ( .A(a[626]), .B(n7735), .Z(n421) );
  IV U9158 ( .A(n7733), .Z(n7735) );
  XNOR U9159 ( .A(b[626]), .B(n7733), .Z(n7734) );
  XOR U9160 ( .A(n7736), .B(n7737), .Z(n7733) );
  ANDN U9161 ( .B(n7738), .A(n422), .Z(n7736) );
  XNOR U9162 ( .A(a[625]), .B(n7739), .Z(n422) );
  IV U9163 ( .A(n7737), .Z(n7739) );
  XNOR U9164 ( .A(b[625]), .B(n7737), .Z(n7738) );
  XOR U9165 ( .A(n7740), .B(n7741), .Z(n7737) );
  ANDN U9166 ( .B(n7742), .A(n423), .Z(n7740) );
  XNOR U9167 ( .A(a[624]), .B(n7743), .Z(n423) );
  IV U9168 ( .A(n7741), .Z(n7743) );
  XNOR U9169 ( .A(b[624]), .B(n7741), .Z(n7742) );
  XOR U9170 ( .A(n7744), .B(n7745), .Z(n7741) );
  ANDN U9171 ( .B(n7746), .A(n424), .Z(n7744) );
  XNOR U9172 ( .A(a[623]), .B(n7747), .Z(n424) );
  IV U9173 ( .A(n7745), .Z(n7747) );
  XNOR U9174 ( .A(b[623]), .B(n7745), .Z(n7746) );
  XOR U9175 ( .A(n7748), .B(n7749), .Z(n7745) );
  ANDN U9176 ( .B(n7750), .A(n425), .Z(n7748) );
  XNOR U9177 ( .A(a[622]), .B(n7751), .Z(n425) );
  IV U9178 ( .A(n7749), .Z(n7751) );
  XNOR U9179 ( .A(b[622]), .B(n7749), .Z(n7750) );
  XOR U9180 ( .A(n7752), .B(n7753), .Z(n7749) );
  ANDN U9181 ( .B(n7754), .A(n426), .Z(n7752) );
  XNOR U9182 ( .A(a[621]), .B(n7755), .Z(n426) );
  IV U9183 ( .A(n7753), .Z(n7755) );
  XNOR U9184 ( .A(b[621]), .B(n7753), .Z(n7754) );
  XOR U9185 ( .A(n7756), .B(n7757), .Z(n7753) );
  ANDN U9186 ( .B(n7758), .A(n427), .Z(n7756) );
  XNOR U9187 ( .A(a[620]), .B(n7759), .Z(n427) );
  IV U9188 ( .A(n7757), .Z(n7759) );
  XNOR U9189 ( .A(b[620]), .B(n7757), .Z(n7758) );
  XOR U9190 ( .A(n7760), .B(n7761), .Z(n7757) );
  ANDN U9191 ( .B(n7762), .A(n429), .Z(n7760) );
  XNOR U9192 ( .A(a[619]), .B(n7763), .Z(n429) );
  IV U9193 ( .A(n7761), .Z(n7763) );
  XNOR U9194 ( .A(b[619]), .B(n7761), .Z(n7762) );
  XOR U9195 ( .A(n7764), .B(n7765), .Z(n7761) );
  ANDN U9196 ( .B(n7766), .A(n430), .Z(n7764) );
  XNOR U9197 ( .A(a[618]), .B(n7767), .Z(n430) );
  IV U9198 ( .A(n7765), .Z(n7767) );
  XNOR U9199 ( .A(b[618]), .B(n7765), .Z(n7766) );
  XOR U9200 ( .A(n7768), .B(n7769), .Z(n7765) );
  ANDN U9201 ( .B(n7770), .A(n431), .Z(n7768) );
  XNOR U9202 ( .A(a[617]), .B(n7771), .Z(n431) );
  IV U9203 ( .A(n7769), .Z(n7771) );
  XNOR U9204 ( .A(b[617]), .B(n7769), .Z(n7770) );
  XOR U9205 ( .A(n7772), .B(n7773), .Z(n7769) );
  ANDN U9206 ( .B(n7774), .A(n432), .Z(n7772) );
  XNOR U9207 ( .A(a[616]), .B(n7775), .Z(n432) );
  IV U9208 ( .A(n7773), .Z(n7775) );
  XNOR U9209 ( .A(b[616]), .B(n7773), .Z(n7774) );
  XOR U9210 ( .A(n7776), .B(n7777), .Z(n7773) );
  ANDN U9211 ( .B(n7778), .A(n433), .Z(n7776) );
  XNOR U9212 ( .A(a[615]), .B(n7779), .Z(n433) );
  IV U9213 ( .A(n7777), .Z(n7779) );
  XNOR U9214 ( .A(b[615]), .B(n7777), .Z(n7778) );
  XOR U9215 ( .A(n7780), .B(n7781), .Z(n7777) );
  ANDN U9216 ( .B(n7782), .A(n434), .Z(n7780) );
  XNOR U9217 ( .A(a[614]), .B(n7783), .Z(n434) );
  IV U9218 ( .A(n7781), .Z(n7783) );
  XNOR U9219 ( .A(b[614]), .B(n7781), .Z(n7782) );
  XOR U9220 ( .A(n7784), .B(n7785), .Z(n7781) );
  ANDN U9221 ( .B(n7786), .A(n435), .Z(n7784) );
  XNOR U9222 ( .A(a[613]), .B(n7787), .Z(n435) );
  IV U9223 ( .A(n7785), .Z(n7787) );
  XNOR U9224 ( .A(b[613]), .B(n7785), .Z(n7786) );
  XOR U9225 ( .A(n7788), .B(n7789), .Z(n7785) );
  ANDN U9226 ( .B(n7790), .A(n436), .Z(n7788) );
  XNOR U9227 ( .A(a[612]), .B(n7791), .Z(n436) );
  IV U9228 ( .A(n7789), .Z(n7791) );
  XNOR U9229 ( .A(b[612]), .B(n7789), .Z(n7790) );
  XOR U9230 ( .A(n7792), .B(n7793), .Z(n7789) );
  ANDN U9231 ( .B(n7794), .A(n437), .Z(n7792) );
  XNOR U9232 ( .A(a[611]), .B(n7795), .Z(n437) );
  IV U9233 ( .A(n7793), .Z(n7795) );
  XNOR U9234 ( .A(b[611]), .B(n7793), .Z(n7794) );
  XOR U9235 ( .A(n7796), .B(n7797), .Z(n7793) );
  ANDN U9236 ( .B(n7798), .A(n438), .Z(n7796) );
  XNOR U9237 ( .A(a[610]), .B(n7799), .Z(n438) );
  IV U9238 ( .A(n7797), .Z(n7799) );
  XNOR U9239 ( .A(b[610]), .B(n7797), .Z(n7798) );
  XOR U9240 ( .A(n7800), .B(n7801), .Z(n7797) );
  ANDN U9241 ( .B(n7802), .A(n440), .Z(n7800) );
  XNOR U9242 ( .A(a[609]), .B(n7803), .Z(n440) );
  IV U9243 ( .A(n7801), .Z(n7803) );
  XNOR U9244 ( .A(b[609]), .B(n7801), .Z(n7802) );
  XOR U9245 ( .A(n7804), .B(n7805), .Z(n7801) );
  ANDN U9246 ( .B(n7806), .A(n441), .Z(n7804) );
  XNOR U9247 ( .A(a[608]), .B(n7807), .Z(n441) );
  IV U9248 ( .A(n7805), .Z(n7807) );
  XNOR U9249 ( .A(b[608]), .B(n7805), .Z(n7806) );
  XOR U9250 ( .A(n7808), .B(n7809), .Z(n7805) );
  ANDN U9251 ( .B(n7810), .A(n442), .Z(n7808) );
  XNOR U9252 ( .A(a[607]), .B(n7811), .Z(n442) );
  IV U9253 ( .A(n7809), .Z(n7811) );
  XNOR U9254 ( .A(b[607]), .B(n7809), .Z(n7810) );
  XOR U9255 ( .A(n7812), .B(n7813), .Z(n7809) );
  ANDN U9256 ( .B(n7814), .A(n443), .Z(n7812) );
  XNOR U9257 ( .A(a[606]), .B(n7815), .Z(n443) );
  IV U9258 ( .A(n7813), .Z(n7815) );
  XNOR U9259 ( .A(b[606]), .B(n7813), .Z(n7814) );
  XOR U9260 ( .A(n7816), .B(n7817), .Z(n7813) );
  ANDN U9261 ( .B(n7818), .A(n444), .Z(n7816) );
  XNOR U9262 ( .A(a[605]), .B(n7819), .Z(n444) );
  IV U9263 ( .A(n7817), .Z(n7819) );
  XNOR U9264 ( .A(b[605]), .B(n7817), .Z(n7818) );
  XOR U9265 ( .A(n7820), .B(n7821), .Z(n7817) );
  ANDN U9266 ( .B(n7822), .A(n445), .Z(n7820) );
  XNOR U9267 ( .A(a[604]), .B(n7823), .Z(n445) );
  IV U9268 ( .A(n7821), .Z(n7823) );
  XNOR U9269 ( .A(b[604]), .B(n7821), .Z(n7822) );
  XOR U9270 ( .A(n7824), .B(n7825), .Z(n7821) );
  ANDN U9271 ( .B(n7826), .A(n446), .Z(n7824) );
  XNOR U9272 ( .A(a[603]), .B(n7827), .Z(n446) );
  IV U9273 ( .A(n7825), .Z(n7827) );
  XNOR U9274 ( .A(b[603]), .B(n7825), .Z(n7826) );
  XOR U9275 ( .A(n7828), .B(n7829), .Z(n7825) );
  ANDN U9276 ( .B(n7830), .A(n447), .Z(n7828) );
  XNOR U9277 ( .A(a[602]), .B(n7831), .Z(n447) );
  IV U9278 ( .A(n7829), .Z(n7831) );
  XNOR U9279 ( .A(b[602]), .B(n7829), .Z(n7830) );
  XOR U9280 ( .A(n7832), .B(n7833), .Z(n7829) );
  ANDN U9281 ( .B(n7834), .A(n448), .Z(n7832) );
  XNOR U9282 ( .A(a[601]), .B(n7835), .Z(n448) );
  IV U9283 ( .A(n7833), .Z(n7835) );
  XNOR U9284 ( .A(b[601]), .B(n7833), .Z(n7834) );
  XOR U9285 ( .A(n7836), .B(n7837), .Z(n7833) );
  ANDN U9286 ( .B(n7838), .A(n449), .Z(n7836) );
  XNOR U9287 ( .A(a[600]), .B(n7839), .Z(n449) );
  IV U9288 ( .A(n7837), .Z(n7839) );
  XNOR U9289 ( .A(b[600]), .B(n7837), .Z(n7838) );
  XOR U9290 ( .A(n7840), .B(n7841), .Z(n7837) );
  ANDN U9291 ( .B(n7842), .A(n452), .Z(n7840) );
  XNOR U9292 ( .A(a[599]), .B(n7843), .Z(n452) );
  IV U9293 ( .A(n7841), .Z(n7843) );
  XNOR U9294 ( .A(b[599]), .B(n7841), .Z(n7842) );
  XOR U9295 ( .A(n7844), .B(n7845), .Z(n7841) );
  ANDN U9296 ( .B(n7846), .A(n453), .Z(n7844) );
  XNOR U9297 ( .A(a[598]), .B(n7847), .Z(n453) );
  IV U9298 ( .A(n7845), .Z(n7847) );
  XNOR U9299 ( .A(b[598]), .B(n7845), .Z(n7846) );
  XOR U9300 ( .A(n7848), .B(n7849), .Z(n7845) );
  ANDN U9301 ( .B(n7850), .A(n454), .Z(n7848) );
  XNOR U9302 ( .A(a[597]), .B(n7851), .Z(n454) );
  IV U9303 ( .A(n7849), .Z(n7851) );
  XNOR U9304 ( .A(b[597]), .B(n7849), .Z(n7850) );
  XOR U9305 ( .A(n7852), .B(n7853), .Z(n7849) );
  ANDN U9306 ( .B(n7854), .A(n455), .Z(n7852) );
  XNOR U9307 ( .A(a[596]), .B(n7855), .Z(n455) );
  IV U9308 ( .A(n7853), .Z(n7855) );
  XNOR U9309 ( .A(b[596]), .B(n7853), .Z(n7854) );
  XOR U9310 ( .A(n7856), .B(n7857), .Z(n7853) );
  ANDN U9311 ( .B(n7858), .A(n456), .Z(n7856) );
  XNOR U9312 ( .A(a[595]), .B(n7859), .Z(n456) );
  IV U9313 ( .A(n7857), .Z(n7859) );
  XNOR U9314 ( .A(b[595]), .B(n7857), .Z(n7858) );
  XOR U9315 ( .A(n7860), .B(n7861), .Z(n7857) );
  ANDN U9316 ( .B(n7862), .A(n457), .Z(n7860) );
  XNOR U9317 ( .A(a[594]), .B(n7863), .Z(n457) );
  IV U9318 ( .A(n7861), .Z(n7863) );
  XNOR U9319 ( .A(b[594]), .B(n7861), .Z(n7862) );
  XOR U9320 ( .A(n7864), .B(n7865), .Z(n7861) );
  ANDN U9321 ( .B(n7866), .A(n458), .Z(n7864) );
  XNOR U9322 ( .A(a[593]), .B(n7867), .Z(n458) );
  IV U9323 ( .A(n7865), .Z(n7867) );
  XNOR U9324 ( .A(b[593]), .B(n7865), .Z(n7866) );
  XOR U9325 ( .A(n7868), .B(n7869), .Z(n7865) );
  ANDN U9326 ( .B(n7870), .A(n459), .Z(n7868) );
  XNOR U9327 ( .A(a[592]), .B(n7871), .Z(n459) );
  IV U9328 ( .A(n7869), .Z(n7871) );
  XNOR U9329 ( .A(b[592]), .B(n7869), .Z(n7870) );
  XOR U9330 ( .A(n7872), .B(n7873), .Z(n7869) );
  ANDN U9331 ( .B(n7874), .A(n460), .Z(n7872) );
  XNOR U9332 ( .A(a[591]), .B(n7875), .Z(n460) );
  IV U9333 ( .A(n7873), .Z(n7875) );
  XNOR U9334 ( .A(b[591]), .B(n7873), .Z(n7874) );
  XOR U9335 ( .A(n7876), .B(n7877), .Z(n7873) );
  ANDN U9336 ( .B(n7878), .A(n461), .Z(n7876) );
  XNOR U9337 ( .A(a[590]), .B(n7879), .Z(n461) );
  IV U9338 ( .A(n7877), .Z(n7879) );
  XNOR U9339 ( .A(b[590]), .B(n7877), .Z(n7878) );
  XOR U9340 ( .A(n7880), .B(n7881), .Z(n7877) );
  ANDN U9341 ( .B(n7882), .A(n463), .Z(n7880) );
  XNOR U9342 ( .A(a[589]), .B(n7883), .Z(n463) );
  IV U9343 ( .A(n7881), .Z(n7883) );
  XNOR U9344 ( .A(b[589]), .B(n7881), .Z(n7882) );
  XOR U9345 ( .A(n7884), .B(n7885), .Z(n7881) );
  ANDN U9346 ( .B(n7886), .A(n464), .Z(n7884) );
  XNOR U9347 ( .A(a[588]), .B(n7887), .Z(n464) );
  IV U9348 ( .A(n7885), .Z(n7887) );
  XNOR U9349 ( .A(b[588]), .B(n7885), .Z(n7886) );
  XOR U9350 ( .A(n7888), .B(n7889), .Z(n7885) );
  ANDN U9351 ( .B(n7890), .A(n465), .Z(n7888) );
  XNOR U9352 ( .A(a[587]), .B(n7891), .Z(n465) );
  IV U9353 ( .A(n7889), .Z(n7891) );
  XNOR U9354 ( .A(b[587]), .B(n7889), .Z(n7890) );
  XOR U9355 ( .A(n7892), .B(n7893), .Z(n7889) );
  ANDN U9356 ( .B(n7894), .A(n466), .Z(n7892) );
  XNOR U9357 ( .A(a[586]), .B(n7895), .Z(n466) );
  IV U9358 ( .A(n7893), .Z(n7895) );
  XNOR U9359 ( .A(b[586]), .B(n7893), .Z(n7894) );
  XOR U9360 ( .A(n7896), .B(n7897), .Z(n7893) );
  ANDN U9361 ( .B(n7898), .A(n467), .Z(n7896) );
  XNOR U9362 ( .A(a[585]), .B(n7899), .Z(n467) );
  IV U9363 ( .A(n7897), .Z(n7899) );
  XNOR U9364 ( .A(b[585]), .B(n7897), .Z(n7898) );
  XOR U9365 ( .A(n7900), .B(n7901), .Z(n7897) );
  ANDN U9366 ( .B(n7902), .A(n468), .Z(n7900) );
  XNOR U9367 ( .A(a[584]), .B(n7903), .Z(n468) );
  IV U9368 ( .A(n7901), .Z(n7903) );
  XNOR U9369 ( .A(b[584]), .B(n7901), .Z(n7902) );
  XOR U9370 ( .A(n7904), .B(n7905), .Z(n7901) );
  ANDN U9371 ( .B(n7906), .A(n469), .Z(n7904) );
  XNOR U9372 ( .A(a[583]), .B(n7907), .Z(n469) );
  IV U9373 ( .A(n7905), .Z(n7907) );
  XNOR U9374 ( .A(b[583]), .B(n7905), .Z(n7906) );
  XOR U9375 ( .A(n7908), .B(n7909), .Z(n7905) );
  ANDN U9376 ( .B(n7910), .A(n470), .Z(n7908) );
  XNOR U9377 ( .A(a[582]), .B(n7911), .Z(n470) );
  IV U9378 ( .A(n7909), .Z(n7911) );
  XNOR U9379 ( .A(b[582]), .B(n7909), .Z(n7910) );
  XOR U9380 ( .A(n7912), .B(n7913), .Z(n7909) );
  ANDN U9381 ( .B(n7914), .A(n471), .Z(n7912) );
  XNOR U9382 ( .A(a[581]), .B(n7915), .Z(n471) );
  IV U9383 ( .A(n7913), .Z(n7915) );
  XNOR U9384 ( .A(b[581]), .B(n7913), .Z(n7914) );
  XOR U9385 ( .A(n7916), .B(n7917), .Z(n7913) );
  ANDN U9386 ( .B(n7918), .A(n472), .Z(n7916) );
  XNOR U9387 ( .A(a[580]), .B(n7919), .Z(n472) );
  IV U9388 ( .A(n7917), .Z(n7919) );
  XNOR U9389 ( .A(b[580]), .B(n7917), .Z(n7918) );
  XOR U9390 ( .A(n7920), .B(n7921), .Z(n7917) );
  ANDN U9391 ( .B(n7922), .A(n474), .Z(n7920) );
  XNOR U9392 ( .A(a[579]), .B(n7923), .Z(n474) );
  IV U9393 ( .A(n7921), .Z(n7923) );
  XNOR U9394 ( .A(b[579]), .B(n7921), .Z(n7922) );
  XOR U9395 ( .A(n7924), .B(n7925), .Z(n7921) );
  ANDN U9396 ( .B(n7926), .A(n475), .Z(n7924) );
  XNOR U9397 ( .A(a[578]), .B(n7927), .Z(n475) );
  IV U9398 ( .A(n7925), .Z(n7927) );
  XNOR U9399 ( .A(b[578]), .B(n7925), .Z(n7926) );
  XOR U9400 ( .A(n7928), .B(n7929), .Z(n7925) );
  ANDN U9401 ( .B(n7930), .A(n476), .Z(n7928) );
  XNOR U9402 ( .A(a[577]), .B(n7931), .Z(n476) );
  IV U9403 ( .A(n7929), .Z(n7931) );
  XNOR U9404 ( .A(b[577]), .B(n7929), .Z(n7930) );
  XOR U9405 ( .A(n7932), .B(n7933), .Z(n7929) );
  ANDN U9406 ( .B(n7934), .A(n477), .Z(n7932) );
  XNOR U9407 ( .A(a[576]), .B(n7935), .Z(n477) );
  IV U9408 ( .A(n7933), .Z(n7935) );
  XNOR U9409 ( .A(b[576]), .B(n7933), .Z(n7934) );
  XOR U9410 ( .A(n7936), .B(n7937), .Z(n7933) );
  ANDN U9411 ( .B(n7938), .A(n478), .Z(n7936) );
  XNOR U9412 ( .A(a[575]), .B(n7939), .Z(n478) );
  IV U9413 ( .A(n7937), .Z(n7939) );
  XNOR U9414 ( .A(b[575]), .B(n7937), .Z(n7938) );
  XOR U9415 ( .A(n7940), .B(n7941), .Z(n7937) );
  ANDN U9416 ( .B(n7942), .A(n479), .Z(n7940) );
  XNOR U9417 ( .A(a[574]), .B(n7943), .Z(n479) );
  IV U9418 ( .A(n7941), .Z(n7943) );
  XNOR U9419 ( .A(b[574]), .B(n7941), .Z(n7942) );
  XOR U9420 ( .A(n7944), .B(n7945), .Z(n7941) );
  ANDN U9421 ( .B(n7946), .A(n480), .Z(n7944) );
  XNOR U9422 ( .A(a[573]), .B(n7947), .Z(n480) );
  IV U9423 ( .A(n7945), .Z(n7947) );
  XNOR U9424 ( .A(b[573]), .B(n7945), .Z(n7946) );
  XOR U9425 ( .A(n7948), .B(n7949), .Z(n7945) );
  ANDN U9426 ( .B(n7950), .A(n481), .Z(n7948) );
  XNOR U9427 ( .A(a[572]), .B(n7951), .Z(n481) );
  IV U9428 ( .A(n7949), .Z(n7951) );
  XNOR U9429 ( .A(b[572]), .B(n7949), .Z(n7950) );
  XOR U9430 ( .A(n7952), .B(n7953), .Z(n7949) );
  ANDN U9431 ( .B(n7954), .A(n482), .Z(n7952) );
  XNOR U9432 ( .A(a[571]), .B(n7955), .Z(n482) );
  IV U9433 ( .A(n7953), .Z(n7955) );
  XNOR U9434 ( .A(b[571]), .B(n7953), .Z(n7954) );
  XOR U9435 ( .A(n7956), .B(n7957), .Z(n7953) );
  ANDN U9436 ( .B(n7958), .A(n483), .Z(n7956) );
  XNOR U9437 ( .A(a[570]), .B(n7959), .Z(n483) );
  IV U9438 ( .A(n7957), .Z(n7959) );
  XNOR U9439 ( .A(b[570]), .B(n7957), .Z(n7958) );
  XOR U9440 ( .A(n7960), .B(n7961), .Z(n7957) );
  ANDN U9441 ( .B(n7962), .A(n485), .Z(n7960) );
  XNOR U9442 ( .A(a[569]), .B(n7963), .Z(n485) );
  IV U9443 ( .A(n7961), .Z(n7963) );
  XNOR U9444 ( .A(b[569]), .B(n7961), .Z(n7962) );
  XOR U9445 ( .A(n7964), .B(n7965), .Z(n7961) );
  ANDN U9446 ( .B(n7966), .A(n486), .Z(n7964) );
  XNOR U9447 ( .A(a[568]), .B(n7967), .Z(n486) );
  IV U9448 ( .A(n7965), .Z(n7967) );
  XNOR U9449 ( .A(b[568]), .B(n7965), .Z(n7966) );
  XOR U9450 ( .A(n7968), .B(n7969), .Z(n7965) );
  ANDN U9451 ( .B(n7970), .A(n487), .Z(n7968) );
  XNOR U9452 ( .A(a[567]), .B(n7971), .Z(n487) );
  IV U9453 ( .A(n7969), .Z(n7971) );
  XNOR U9454 ( .A(b[567]), .B(n7969), .Z(n7970) );
  XOR U9455 ( .A(n7972), .B(n7973), .Z(n7969) );
  ANDN U9456 ( .B(n7974), .A(n488), .Z(n7972) );
  XNOR U9457 ( .A(a[566]), .B(n7975), .Z(n488) );
  IV U9458 ( .A(n7973), .Z(n7975) );
  XNOR U9459 ( .A(b[566]), .B(n7973), .Z(n7974) );
  XOR U9460 ( .A(n7976), .B(n7977), .Z(n7973) );
  ANDN U9461 ( .B(n7978), .A(n489), .Z(n7976) );
  XNOR U9462 ( .A(a[565]), .B(n7979), .Z(n489) );
  IV U9463 ( .A(n7977), .Z(n7979) );
  XNOR U9464 ( .A(b[565]), .B(n7977), .Z(n7978) );
  XOR U9465 ( .A(n7980), .B(n7981), .Z(n7977) );
  ANDN U9466 ( .B(n7982), .A(n490), .Z(n7980) );
  XNOR U9467 ( .A(a[564]), .B(n7983), .Z(n490) );
  IV U9468 ( .A(n7981), .Z(n7983) );
  XNOR U9469 ( .A(b[564]), .B(n7981), .Z(n7982) );
  XOR U9470 ( .A(n7984), .B(n7985), .Z(n7981) );
  ANDN U9471 ( .B(n7986), .A(n491), .Z(n7984) );
  XNOR U9472 ( .A(a[563]), .B(n7987), .Z(n491) );
  IV U9473 ( .A(n7985), .Z(n7987) );
  XNOR U9474 ( .A(b[563]), .B(n7985), .Z(n7986) );
  XOR U9475 ( .A(n7988), .B(n7989), .Z(n7985) );
  ANDN U9476 ( .B(n7990), .A(n492), .Z(n7988) );
  XNOR U9477 ( .A(a[562]), .B(n7991), .Z(n492) );
  IV U9478 ( .A(n7989), .Z(n7991) );
  XNOR U9479 ( .A(b[562]), .B(n7989), .Z(n7990) );
  XOR U9480 ( .A(n7992), .B(n7993), .Z(n7989) );
  ANDN U9481 ( .B(n7994), .A(n493), .Z(n7992) );
  XNOR U9482 ( .A(a[561]), .B(n7995), .Z(n493) );
  IV U9483 ( .A(n7993), .Z(n7995) );
  XNOR U9484 ( .A(b[561]), .B(n7993), .Z(n7994) );
  XOR U9485 ( .A(n7996), .B(n7997), .Z(n7993) );
  ANDN U9486 ( .B(n7998), .A(n494), .Z(n7996) );
  XNOR U9487 ( .A(a[560]), .B(n7999), .Z(n494) );
  IV U9488 ( .A(n7997), .Z(n7999) );
  XNOR U9489 ( .A(b[560]), .B(n7997), .Z(n7998) );
  XOR U9490 ( .A(n8000), .B(n8001), .Z(n7997) );
  ANDN U9491 ( .B(n8002), .A(n496), .Z(n8000) );
  XNOR U9492 ( .A(a[559]), .B(n8003), .Z(n496) );
  IV U9493 ( .A(n8001), .Z(n8003) );
  XNOR U9494 ( .A(b[559]), .B(n8001), .Z(n8002) );
  XOR U9495 ( .A(n8004), .B(n8005), .Z(n8001) );
  ANDN U9496 ( .B(n8006), .A(n497), .Z(n8004) );
  XNOR U9497 ( .A(a[558]), .B(n8007), .Z(n497) );
  IV U9498 ( .A(n8005), .Z(n8007) );
  XNOR U9499 ( .A(b[558]), .B(n8005), .Z(n8006) );
  XOR U9500 ( .A(n8008), .B(n8009), .Z(n8005) );
  ANDN U9501 ( .B(n8010), .A(n498), .Z(n8008) );
  XNOR U9502 ( .A(a[557]), .B(n8011), .Z(n498) );
  IV U9503 ( .A(n8009), .Z(n8011) );
  XNOR U9504 ( .A(b[557]), .B(n8009), .Z(n8010) );
  XOR U9505 ( .A(n8012), .B(n8013), .Z(n8009) );
  ANDN U9506 ( .B(n8014), .A(n499), .Z(n8012) );
  XNOR U9507 ( .A(a[556]), .B(n8015), .Z(n499) );
  IV U9508 ( .A(n8013), .Z(n8015) );
  XNOR U9509 ( .A(b[556]), .B(n8013), .Z(n8014) );
  XOR U9510 ( .A(n8016), .B(n8017), .Z(n8013) );
  ANDN U9511 ( .B(n8018), .A(n500), .Z(n8016) );
  XNOR U9512 ( .A(a[555]), .B(n8019), .Z(n500) );
  IV U9513 ( .A(n8017), .Z(n8019) );
  XNOR U9514 ( .A(b[555]), .B(n8017), .Z(n8018) );
  XOR U9515 ( .A(n8020), .B(n8021), .Z(n8017) );
  ANDN U9516 ( .B(n8022), .A(n501), .Z(n8020) );
  XNOR U9517 ( .A(a[554]), .B(n8023), .Z(n501) );
  IV U9518 ( .A(n8021), .Z(n8023) );
  XNOR U9519 ( .A(b[554]), .B(n8021), .Z(n8022) );
  XOR U9520 ( .A(n8024), .B(n8025), .Z(n8021) );
  ANDN U9521 ( .B(n8026), .A(n502), .Z(n8024) );
  XNOR U9522 ( .A(a[553]), .B(n8027), .Z(n502) );
  IV U9523 ( .A(n8025), .Z(n8027) );
  XNOR U9524 ( .A(b[553]), .B(n8025), .Z(n8026) );
  XOR U9525 ( .A(n8028), .B(n8029), .Z(n8025) );
  ANDN U9526 ( .B(n8030), .A(n503), .Z(n8028) );
  XNOR U9527 ( .A(a[552]), .B(n8031), .Z(n503) );
  IV U9528 ( .A(n8029), .Z(n8031) );
  XNOR U9529 ( .A(b[552]), .B(n8029), .Z(n8030) );
  XOR U9530 ( .A(n8032), .B(n8033), .Z(n8029) );
  ANDN U9531 ( .B(n8034), .A(n504), .Z(n8032) );
  XNOR U9532 ( .A(a[551]), .B(n8035), .Z(n504) );
  IV U9533 ( .A(n8033), .Z(n8035) );
  XNOR U9534 ( .A(b[551]), .B(n8033), .Z(n8034) );
  XOR U9535 ( .A(n8036), .B(n8037), .Z(n8033) );
  ANDN U9536 ( .B(n8038), .A(n505), .Z(n8036) );
  XNOR U9537 ( .A(a[550]), .B(n8039), .Z(n505) );
  IV U9538 ( .A(n8037), .Z(n8039) );
  XNOR U9539 ( .A(b[550]), .B(n8037), .Z(n8038) );
  XOR U9540 ( .A(n8040), .B(n8041), .Z(n8037) );
  ANDN U9541 ( .B(n8042), .A(n507), .Z(n8040) );
  XNOR U9542 ( .A(a[549]), .B(n8043), .Z(n507) );
  IV U9543 ( .A(n8041), .Z(n8043) );
  XNOR U9544 ( .A(b[549]), .B(n8041), .Z(n8042) );
  XOR U9545 ( .A(n8044), .B(n8045), .Z(n8041) );
  ANDN U9546 ( .B(n8046), .A(n508), .Z(n8044) );
  XNOR U9547 ( .A(a[548]), .B(n8047), .Z(n508) );
  IV U9548 ( .A(n8045), .Z(n8047) );
  XNOR U9549 ( .A(b[548]), .B(n8045), .Z(n8046) );
  XOR U9550 ( .A(n8048), .B(n8049), .Z(n8045) );
  ANDN U9551 ( .B(n8050), .A(n509), .Z(n8048) );
  XNOR U9552 ( .A(a[547]), .B(n8051), .Z(n509) );
  IV U9553 ( .A(n8049), .Z(n8051) );
  XNOR U9554 ( .A(b[547]), .B(n8049), .Z(n8050) );
  XOR U9555 ( .A(n8052), .B(n8053), .Z(n8049) );
  ANDN U9556 ( .B(n8054), .A(n510), .Z(n8052) );
  XNOR U9557 ( .A(a[546]), .B(n8055), .Z(n510) );
  IV U9558 ( .A(n8053), .Z(n8055) );
  XNOR U9559 ( .A(b[546]), .B(n8053), .Z(n8054) );
  XOR U9560 ( .A(n8056), .B(n8057), .Z(n8053) );
  ANDN U9561 ( .B(n8058), .A(n511), .Z(n8056) );
  XNOR U9562 ( .A(a[545]), .B(n8059), .Z(n511) );
  IV U9563 ( .A(n8057), .Z(n8059) );
  XNOR U9564 ( .A(b[545]), .B(n8057), .Z(n8058) );
  XOR U9565 ( .A(n8060), .B(n8061), .Z(n8057) );
  ANDN U9566 ( .B(n8062), .A(n512), .Z(n8060) );
  XNOR U9567 ( .A(a[544]), .B(n8063), .Z(n512) );
  IV U9568 ( .A(n8061), .Z(n8063) );
  XNOR U9569 ( .A(b[544]), .B(n8061), .Z(n8062) );
  XOR U9570 ( .A(n8064), .B(n8065), .Z(n8061) );
  ANDN U9571 ( .B(n8066), .A(n513), .Z(n8064) );
  XNOR U9572 ( .A(a[543]), .B(n8067), .Z(n513) );
  IV U9573 ( .A(n8065), .Z(n8067) );
  XNOR U9574 ( .A(b[543]), .B(n8065), .Z(n8066) );
  XOR U9575 ( .A(n8068), .B(n8069), .Z(n8065) );
  ANDN U9576 ( .B(n8070), .A(n514), .Z(n8068) );
  XNOR U9577 ( .A(a[542]), .B(n8071), .Z(n514) );
  IV U9578 ( .A(n8069), .Z(n8071) );
  XNOR U9579 ( .A(b[542]), .B(n8069), .Z(n8070) );
  XOR U9580 ( .A(n8072), .B(n8073), .Z(n8069) );
  ANDN U9581 ( .B(n8074), .A(n515), .Z(n8072) );
  XNOR U9582 ( .A(a[541]), .B(n8075), .Z(n515) );
  IV U9583 ( .A(n8073), .Z(n8075) );
  XNOR U9584 ( .A(b[541]), .B(n8073), .Z(n8074) );
  XOR U9585 ( .A(n8076), .B(n8077), .Z(n8073) );
  ANDN U9586 ( .B(n8078), .A(n516), .Z(n8076) );
  XNOR U9587 ( .A(a[540]), .B(n8079), .Z(n516) );
  IV U9588 ( .A(n8077), .Z(n8079) );
  XNOR U9589 ( .A(b[540]), .B(n8077), .Z(n8078) );
  XOR U9590 ( .A(n8080), .B(n8081), .Z(n8077) );
  ANDN U9591 ( .B(n8082), .A(n518), .Z(n8080) );
  XNOR U9592 ( .A(a[539]), .B(n8083), .Z(n518) );
  IV U9593 ( .A(n8081), .Z(n8083) );
  XNOR U9594 ( .A(b[539]), .B(n8081), .Z(n8082) );
  XOR U9595 ( .A(n8084), .B(n8085), .Z(n8081) );
  ANDN U9596 ( .B(n8086), .A(n519), .Z(n8084) );
  XNOR U9597 ( .A(a[538]), .B(n8087), .Z(n519) );
  IV U9598 ( .A(n8085), .Z(n8087) );
  XNOR U9599 ( .A(b[538]), .B(n8085), .Z(n8086) );
  XOR U9600 ( .A(n8088), .B(n8089), .Z(n8085) );
  ANDN U9601 ( .B(n8090), .A(n520), .Z(n8088) );
  XNOR U9602 ( .A(a[537]), .B(n8091), .Z(n520) );
  IV U9603 ( .A(n8089), .Z(n8091) );
  XNOR U9604 ( .A(b[537]), .B(n8089), .Z(n8090) );
  XOR U9605 ( .A(n8092), .B(n8093), .Z(n8089) );
  ANDN U9606 ( .B(n8094), .A(n521), .Z(n8092) );
  XNOR U9607 ( .A(a[536]), .B(n8095), .Z(n521) );
  IV U9608 ( .A(n8093), .Z(n8095) );
  XNOR U9609 ( .A(b[536]), .B(n8093), .Z(n8094) );
  XOR U9610 ( .A(n8096), .B(n8097), .Z(n8093) );
  ANDN U9611 ( .B(n8098), .A(n522), .Z(n8096) );
  XNOR U9612 ( .A(a[535]), .B(n8099), .Z(n522) );
  IV U9613 ( .A(n8097), .Z(n8099) );
  XNOR U9614 ( .A(b[535]), .B(n8097), .Z(n8098) );
  XOR U9615 ( .A(n8100), .B(n8101), .Z(n8097) );
  ANDN U9616 ( .B(n8102), .A(n523), .Z(n8100) );
  XNOR U9617 ( .A(a[534]), .B(n8103), .Z(n523) );
  IV U9618 ( .A(n8101), .Z(n8103) );
  XNOR U9619 ( .A(b[534]), .B(n8101), .Z(n8102) );
  XOR U9620 ( .A(n8104), .B(n8105), .Z(n8101) );
  ANDN U9621 ( .B(n8106), .A(n524), .Z(n8104) );
  XNOR U9622 ( .A(a[533]), .B(n8107), .Z(n524) );
  IV U9623 ( .A(n8105), .Z(n8107) );
  XNOR U9624 ( .A(b[533]), .B(n8105), .Z(n8106) );
  XOR U9625 ( .A(n8108), .B(n8109), .Z(n8105) );
  ANDN U9626 ( .B(n8110), .A(n525), .Z(n8108) );
  XNOR U9627 ( .A(a[532]), .B(n8111), .Z(n525) );
  IV U9628 ( .A(n8109), .Z(n8111) );
  XNOR U9629 ( .A(b[532]), .B(n8109), .Z(n8110) );
  XOR U9630 ( .A(n8112), .B(n8113), .Z(n8109) );
  ANDN U9631 ( .B(n8114), .A(n526), .Z(n8112) );
  XNOR U9632 ( .A(a[531]), .B(n8115), .Z(n526) );
  IV U9633 ( .A(n8113), .Z(n8115) );
  XNOR U9634 ( .A(b[531]), .B(n8113), .Z(n8114) );
  XOR U9635 ( .A(n8116), .B(n8117), .Z(n8113) );
  ANDN U9636 ( .B(n8118), .A(n527), .Z(n8116) );
  XNOR U9637 ( .A(a[530]), .B(n8119), .Z(n527) );
  IV U9638 ( .A(n8117), .Z(n8119) );
  XNOR U9639 ( .A(b[530]), .B(n8117), .Z(n8118) );
  XOR U9640 ( .A(n8120), .B(n8121), .Z(n8117) );
  ANDN U9641 ( .B(n8122), .A(n529), .Z(n8120) );
  XNOR U9642 ( .A(a[529]), .B(n8123), .Z(n529) );
  IV U9643 ( .A(n8121), .Z(n8123) );
  XNOR U9644 ( .A(b[529]), .B(n8121), .Z(n8122) );
  XOR U9645 ( .A(n8124), .B(n8125), .Z(n8121) );
  ANDN U9646 ( .B(n8126), .A(n530), .Z(n8124) );
  XNOR U9647 ( .A(a[528]), .B(n8127), .Z(n530) );
  IV U9648 ( .A(n8125), .Z(n8127) );
  XNOR U9649 ( .A(b[528]), .B(n8125), .Z(n8126) );
  XOR U9650 ( .A(n8128), .B(n8129), .Z(n8125) );
  ANDN U9651 ( .B(n8130), .A(n531), .Z(n8128) );
  XNOR U9652 ( .A(a[527]), .B(n8131), .Z(n531) );
  IV U9653 ( .A(n8129), .Z(n8131) );
  XNOR U9654 ( .A(b[527]), .B(n8129), .Z(n8130) );
  XOR U9655 ( .A(n8132), .B(n8133), .Z(n8129) );
  ANDN U9656 ( .B(n8134), .A(n532), .Z(n8132) );
  XNOR U9657 ( .A(a[526]), .B(n8135), .Z(n532) );
  IV U9658 ( .A(n8133), .Z(n8135) );
  XNOR U9659 ( .A(b[526]), .B(n8133), .Z(n8134) );
  XOR U9660 ( .A(n8136), .B(n8137), .Z(n8133) );
  ANDN U9661 ( .B(n8138), .A(n533), .Z(n8136) );
  XNOR U9662 ( .A(a[525]), .B(n8139), .Z(n533) );
  IV U9663 ( .A(n8137), .Z(n8139) );
  XNOR U9664 ( .A(b[525]), .B(n8137), .Z(n8138) );
  XOR U9665 ( .A(n8140), .B(n8141), .Z(n8137) );
  ANDN U9666 ( .B(n8142), .A(n534), .Z(n8140) );
  XNOR U9667 ( .A(a[524]), .B(n8143), .Z(n534) );
  IV U9668 ( .A(n8141), .Z(n8143) );
  XNOR U9669 ( .A(b[524]), .B(n8141), .Z(n8142) );
  XOR U9670 ( .A(n8144), .B(n8145), .Z(n8141) );
  ANDN U9671 ( .B(n8146), .A(n535), .Z(n8144) );
  XNOR U9672 ( .A(a[523]), .B(n8147), .Z(n535) );
  IV U9673 ( .A(n8145), .Z(n8147) );
  XNOR U9674 ( .A(b[523]), .B(n8145), .Z(n8146) );
  XOR U9675 ( .A(n8148), .B(n8149), .Z(n8145) );
  ANDN U9676 ( .B(n8150), .A(n536), .Z(n8148) );
  XNOR U9677 ( .A(a[522]), .B(n8151), .Z(n536) );
  IV U9678 ( .A(n8149), .Z(n8151) );
  XNOR U9679 ( .A(b[522]), .B(n8149), .Z(n8150) );
  XOR U9680 ( .A(n8152), .B(n8153), .Z(n8149) );
  ANDN U9681 ( .B(n8154), .A(n537), .Z(n8152) );
  XNOR U9682 ( .A(a[521]), .B(n8155), .Z(n537) );
  IV U9683 ( .A(n8153), .Z(n8155) );
  XNOR U9684 ( .A(b[521]), .B(n8153), .Z(n8154) );
  XOR U9685 ( .A(n8156), .B(n8157), .Z(n8153) );
  ANDN U9686 ( .B(n8158), .A(n538), .Z(n8156) );
  XNOR U9687 ( .A(a[520]), .B(n8159), .Z(n538) );
  IV U9688 ( .A(n8157), .Z(n8159) );
  XNOR U9689 ( .A(b[520]), .B(n8157), .Z(n8158) );
  XOR U9690 ( .A(n8160), .B(n8161), .Z(n8157) );
  ANDN U9691 ( .B(n8162), .A(n540), .Z(n8160) );
  XNOR U9692 ( .A(a[519]), .B(n8163), .Z(n540) );
  IV U9693 ( .A(n8161), .Z(n8163) );
  XNOR U9694 ( .A(b[519]), .B(n8161), .Z(n8162) );
  XOR U9695 ( .A(n8164), .B(n8165), .Z(n8161) );
  ANDN U9696 ( .B(n8166), .A(n541), .Z(n8164) );
  XNOR U9697 ( .A(a[518]), .B(n8167), .Z(n541) );
  IV U9698 ( .A(n8165), .Z(n8167) );
  XNOR U9699 ( .A(b[518]), .B(n8165), .Z(n8166) );
  XOR U9700 ( .A(n8168), .B(n8169), .Z(n8165) );
  ANDN U9701 ( .B(n8170), .A(n542), .Z(n8168) );
  XNOR U9702 ( .A(a[517]), .B(n8171), .Z(n542) );
  IV U9703 ( .A(n8169), .Z(n8171) );
  XNOR U9704 ( .A(b[517]), .B(n8169), .Z(n8170) );
  XOR U9705 ( .A(n8172), .B(n8173), .Z(n8169) );
  ANDN U9706 ( .B(n8174), .A(n543), .Z(n8172) );
  XNOR U9707 ( .A(a[516]), .B(n8175), .Z(n543) );
  IV U9708 ( .A(n8173), .Z(n8175) );
  XNOR U9709 ( .A(b[516]), .B(n8173), .Z(n8174) );
  XOR U9710 ( .A(n8176), .B(n8177), .Z(n8173) );
  ANDN U9711 ( .B(n8178), .A(n544), .Z(n8176) );
  XNOR U9712 ( .A(a[515]), .B(n8179), .Z(n544) );
  IV U9713 ( .A(n8177), .Z(n8179) );
  XNOR U9714 ( .A(b[515]), .B(n8177), .Z(n8178) );
  XOR U9715 ( .A(n8180), .B(n8181), .Z(n8177) );
  ANDN U9716 ( .B(n8182), .A(n545), .Z(n8180) );
  XNOR U9717 ( .A(a[514]), .B(n8183), .Z(n545) );
  IV U9718 ( .A(n8181), .Z(n8183) );
  XNOR U9719 ( .A(b[514]), .B(n8181), .Z(n8182) );
  XOR U9720 ( .A(n8184), .B(n8185), .Z(n8181) );
  ANDN U9721 ( .B(n8186), .A(n546), .Z(n8184) );
  XNOR U9722 ( .A(a[513]), .B(n8187), .Z(n546) );
  IV U9723 ( .A(n8185), .Z(n8187) );
  XNOR U9724 ( .A(b[513]), .B(n8185), .Z(n8186) );
  XOR U9725 ( .A(n8188), .B(n8189), .Z(n8185) );
  ANDN U9726 ( .B(n8190), .A(n547), .Z(n8188) );
  XNOR U9727 ( .A(a[512]), .B(n8191), .Z(n547) );
  IV U9728 ( .A(n8189), .Z(n8191) );
  XNOR U9729 ( .A(b[512]), .B(n8189), .Z(n8190) );
  XOR U9730 ( .A(n8192), .B(n8193), .Z(n8189) );
  ANDN U9731 ( .B(n8194), .A(n548), .Z(n8192) );
  XNOR U9732 ( .A(a[511]), .B(n8195), .Z(n548) );
  IV U9733 ( .A(n8193), .Z(n8195) );
  XNOR U9734 ( .A(b[511]), .B(n8193), .Z(n8194) );
  XOR U9735 ( .A(n8196), .B(n8197), .Z(n8193) );
  ANDN U9736 ( .B(n8198), .A(n549), .Z(n8196) );
  XNOR U9737 ( .A(a[510]), .B(n8199), .Z(n549) );
  IV U9738 ( .A(n8197), .Z(n8199) );
  XNOR U9739 ( .A(b[510]), .B(n8197), .Z(n8198) );
  XOR U9740 ( .A(n8200), .B(n8201), .Z(n8197) );
  ANDN U9741 ( .B(n8202), .A(n551), .Z(n8200) );
  XNOR U9742 ( .A(a[509]), .B(n8203), .Z(n551) );
  IV U9743 ( .A(n8201), .Z(n8203) );
  XNOR U9744 ( .A(b[509]), .B(n8201), .Z(n8202) );
  XOR U9745 ( .A(n8204), .B(n8205), .Z(n8201) );
  ANDN U9746 ( .B(n8206), .A(n552), .Z(n8204) );
  XNOR U9747 ( .A(a[508]), .B(n8207), .Z(n552) );
  IV U9748 ( .A(n8205), .Z(n8207) );
  XNOR U9749 ( .A(b[508]), .B(n8205), .Z(n8206) );
  XOR U9750 ( .A(n8208), .B(n8209), .Z(n8205) );
  ANDN U9751 ( .B(n8210), .A(n553), .Z(n8208) );
  XNOR U9752 ( .A(a[507]), .B(n8211), .Z(n553) );
  IV U9753 ( .A(n8209), .Z(n8211) );
  XNOR U9754 ( .A(b[507]), .B(n8209), .Z(n8210) );
  XOR U9755 ( .A(n8212), .B(n8213), .Z(n8209) );
  ANDN U9756 ( .B(n8214), .A(n554), .Z(n8212) );
  XNOR U9757 ( .A(a[506]), .B(n8215), .Z(n554) );
  IV U9758 ( .A(n8213), .Z(n8215) );
  XNOR U9759 ( .A(b[506]), .B(n8213), .Z(n8214) );
  XOR U9760 ( .A(n8216), .B(n8217), .Z(n8213) );
  ANDN U9761 ( .B(n8218), .A(n555), .Z(n8216) );
  XNOR U9762 ( .A(a[505]), .B(n8219), .Z(n555) );
  IV U9763 ( .A(n8217), .Z(n8219) );
  XNOR U9764 ( .A(b[505]), .B(n8217), .Z(n8218) );
  XOR U9765 ( .A(n8220), .B(n8221), .Z(n8217) );
  ANDN U9766 ( .B(n8222), .A(n556), .Z(n8220) );
  XNOR U9767 ( .A(a[504]), .B(n8223), .Z(n556) );
  IV U9768 ( .A(n8221), .Z(n8223) );
  XNOR U9769 ( .A(b[504]), .B(n8221), .Z(n8222) );
  XOR U9770 ( .A(n8224), .B(n8225), .Z(n8221) );
  ANDN U9771 ( .B(n8226), .A(n557), .Z(n8224) );
  XNOR U9772 ( .A(a[503]), .B(n8227), .Z(n557) );
  IV U9773 ( .A(n8225), .Z(n8227) );
  XNOR U9774 ( .A(b[503]), .B(n8225), .Z(n8226) );
  XOR U9775 ( .A(n8228), .B(n8229), .Z(n8225) );
  ANDN U9776 ( .B(n8230), .A(n558), .Z(n8228) );
  XNOR U9777 ( .A(a[502]), .B(n8231), .Z(n558) );
  IV U9778 ( .A(n8229), .Z(n8231) );
  XNOR U9779 ( .A(b[502]), .B(n8229), .Z(n8230) );
  XOR U9780 ( .A(n8232), .B(n8233), .Z(n8229) );
  ANDN U9781 ( .B(n8234), .A(n559), .Z(n8232) );
  XNOR U9782 ( .A(a[501]), .B(n8235), .Z(n559) );
  IV U9783 ( .A(n8233), .Z(n8235) );
  XNOR U9784 ( .A(b[501]), .B(n8233), .Z(n8234) );
  XOR U9785 ( .A(n8236), .B(n8237), .Z(n8233) );
  ANDN U9786 ( .B(n8238), .A(n560), .Z(n8236) );
  XNOR U9787 ( .A(a[500]), .B(n8239), .Z(n560) );
  IV U9788 ( .A(n8237), .Z(n8239) );
  XNOR U9789 ( .A(b[500]), .B(n8237), .Z(n8238) );
  XOR U9790 ( .A(n8240), .B(n8241), .Z(n8237) );
  ANDN U9791 ( .B(n8242), .A(n563), .Z(n8240) );
  XNOR U9792 ( .A(a[499]), .B(n8243), .Z(n563) );
  IV U9793 ( .A(n8241), .Z(n8243) );
  XNOR U9794 ( .A(b[499]), .B(n8241), .Z(n8242) );
  XOR U9795 ( .A(n8244), .B(n8245), .Z(n8241) );
  ANDN U9796 ( .B(n8246), .A(n564), .Z(n8244) );
  XNOR U9797 ( .A(a[498]), .B(n8247), .Z(n564) );
  IV U9798 ( .A(n8245), .Z(n8247) );
  XNOR U9799 ( .A(b[498]), .B(n8245), .Z(n8246) );
  XOR U9800 ( .A(n8248), .B(n8249), .Z(n8245) );
  ANDN U9801 ( .B(n8250), .A(n565), .Z(n8248) );
  XNOR U9802 ( .A(a[497]), .B(n8251), .Z(n565) );
  IV U9803 ( .A(n8249), .Z(n8251) );
  XNOR U9804 ( .A(b[497]), .B(n8249), .Z(n8250) );
  XOR U9805 ( .A(n8252), .B(n8253), .Z(n8249) );
  ANDN U9806 ( .B(n8254), .A(n566), .Z(n8252) );
  XNOR U9807 ( .A(a[496]), .B(n8255), .Z(n566) );
  IV U9808 ( .A(n8253), .Z(n8255) );
  XNOR U9809 ( .A(b[496]), .B(n8253), .Z(n8254) );
  XOR U9810 ( .A(n8256), .B(n8257), .Z(n8253) );
  ANDN U9811 ( .B(n8258), .A(n567), .Z(n8256) );
  XNOR U9812 ( .A(a[495]), .B(n8259), .Z(n567) );
  IV U9813 ( .A(n8257), .Z(n8259) );
  XNOR U9814 ( .A(b[495]), .B(n8257), .Z(n8258) );
  XOR U9815 ( .A(n8260), .B(n8261), .Z(n8257) );
  ANDN U9816 ( .B(n8262), .A(n568), .Z(n8260) );
  XNOR U9817 ( .A(a[494]), .B(n8263), .Z(n568) );
  IV U9818 ( .A(n8261), .Z(n8263) );
  XNOR U9819 ( .A(b[494]), .B(n8261), .Z(n8262) );
  XOR U9820 ( .A(n8264), .B(n8265), .Z(n8261) );
  ANDN U9821 ( .B(n8266), .A(n569), .Z(n8264) );
  XNOR U9822 ( .A(a[493]), .B(n8267), .Z(n569) );
  IV U9823 ( .A(n8265), .Z(n8267) );
  XNOR U9824 ( .A(b[493]), .B(n8265), .Z(n8266) );
  XOR U9825 ( .A(n8268), .B(n8269), .Z(n8265) );
  ANDN U9826 ( .B(n8270), .A(n570), .Z(n8268) );
  XNOR U9827 ( .A(a[492]), .B(n8271), .Z(n570) );
  IV U9828 ( .A(n8269), .Z(n8271) );
  XNOR U9829 ( .A(b[492]), .B(n8269), .Z(n8270) );
  XOR U9830 ( .A(n8272), .B(n8273), .Z(n8269) );
  ANDN U9831 ( .B(n8274), .A(n571), .Z(n8272) );
  XNOR U9832 ( .A(a[491]), .B(n8275), .Z(n571) );
  IV U9833 ( .A(n8273), .Z(n8275) );
  XNOR U9834 ( .A(b[491]), .B(n8273), .Z(n8274) );
  XOR U9835 ( .A(n8276), .B(n8277), .Z(n8273) );
  ANDN U9836 ( .B(n8278), .A(n572), .Z(n8276) );
  XNOR U9837 ( .A(a[490]), .B(n8279), .Z(n572) );
  IV U9838 ( .A(n8277), .Z(n8279) );
  XNOR U9839 ( .A(b[490]), .B(n8277), .Z(n8278) );
  XOR U9840 ( .A(n8280), .B(n8281), .Z(n8277) );
  ANDN U9841 ( .B(n8282), .A(n574), .Z(n8280) );
  XNOR U9842 ( .A(a[489]), .B(n8283), .Z(n574) );
  IV U9843 ( .A(n8281), .Z(n8283) );
  XNOR U9844 ( .A(b[489]), .B(n8281), .Z(n8282) );
  XOR U9845 ( .A(n8284), .B(n8285), .Z(n8281) );
  ANDN U9846 ( .B(n8286), .A(n575), .Z(n8284) );
  XNOR U9847 ( .A(a[488]), .B(n8287), .Z(n575) );
  IV U9848 ( .A(n8285), .Z(n8287) );
  XNOR U9849 ( .A(b[488]), .B(n8285), .Z(n8286) );
  XOR U9850 ( .A(n8288), .B(n8289), .Z(n8285) );
  ANDN U9851 ( .B(n8290), .A(n576), .Z(n8288) );
  XNOR U9852 ( .A(a[487]), .B(n8291), .Z(n576) );
  IV U9853 ( .A(n8289), .Z(n8291) );
  XNOR U9854 ( .A(b[487]), .B(n8289), .Z(n8290) );
  XOR U9855 ( .A(n8292), .B(n8293), .Z(n8289) );
  ANDN U9856 ( .B(n8294), .A(n577), .Z(n8292) );
  XNOR U9857 ( .A(a[486]), .B(n8295), .Z(n577) );
  IV U9858 ( .A(n8293), .Z(n8295) );
  XNOR U9859 ( .A(b[486]), .B(n8293), .Z(n8294) );
  XOR U9860 ( .A(n8296), .B(n8297), .Z(n8293) );
  ANDN U9861 ( .B(n8298), .A(n578), .Z(n8296) );
  XNOR U9862 ( .A(a[485]), .B(n8299), .Z(n578) );
  IV U9863 ( .A(n8297), .Z(n8299) );
  XNOR U9864 ( .A(b[485]), .B(n8297), .Z(n8298) );
  XOR U9865 ( .A(n8300), .B(n8301), .Z(n8297) );
  ANDN U9866 ( .B(n8302), .A(n579), .Z(n8300) );
  XNOR U9867 ( .A(a[484]), .B(n8303), .Z(n579) );
  IV U9868 ( .A(n8301), .Z(n8303) );
  XNOR U9869 ( .A(b[484]), .B(n8301), .Z(n8302) );
  XOR U9870 ( .A(n8304), .B(n8305), .Z(n8301) );
  ANDN U9871 ( .B(n8306), .A(n580), .Z(n8304) );
  XNOR U9872 ( .A(a[483]), .B(n8307), .Z(n580) );
  IV U9873 ( .A(n8305), .Z(n8307) );
  XNOR U9874 ( .A(b[483]), .B(n8305), .Z(n8306) );
  XOR U9875 ( .A(n8308), .B(n8309), .Z(n8305) );
  ANDN U9876 ( .B(n8310), .A(n581), .Z(n8308) );
  XNOR U9877 ( .A(a[482]), .B(n8311), .Z(n581) );
  IV U9878 ( .A(n8309), .Z(n8311) );
  XNOR U9879 ( .A(b[482]), .B(n8309), .Z(n8310) );
  XOR U9880 ( .A(n8312), .B(n8313), .Z(n8309) );
  ANDN U9881 ( .B(n8314), .A(n582), .Z(n8312) );
  XNOR U9882 ( .A(a[481]), .B(n8315), .Z(n582) );
  IV U9883 ( .A(n8313), .Z(n8315) );
  XNOR U9884 ( .A(b[481]), .B(n8313), .Z(n8314) );
  XOR U9885 ( .A(n8316), .B(n8317), .Z(n8313) );
  ANDN U9886 ( .B(n8318), .A(n583), .Z(n8316) );
  XNOR U9887 ( .A(a[480]), .B(n8319), .Z(n583) );
  IV U9888 ( .A(n8317), .Z(n8319) );
  XNOR U9889 ( .A(b[480]), .B(n8317), .Z(n8318) );
  XOR U9890 ( .A(n8320), .B(n8321), .Z(n8317) );
  ANDN U9891 ( .B(n8322), .A(n585), .Z(n8320) );
  XNOR U9892 ( .A(a[479]), .B(n8323), .Z(n585) );
  IV U9893 ( .A(n8321), .Z(n8323) );
  XNOR U9894 ( .A(b[479]), .B(n8321), .Z(n8322) );
  XOR U9895 ( .A(n8324), .B(n8325), .Z(n8321) );
  ANDN U9896 ( .B(n8326), .A(n586), .Z(n8324) );
  XNOR U9897 ( .A(a[478]), .B(n8327), .Z(n586) );
  IV U9898 ( .A(n8325), .Z(n8327) );
  XNOR U9899 ( .A(b[478]), .B(n8325), .Z(n8326) );
  XOR U9900 ( .A(n8328), .B(n8329), .Z(n8325) );
  ANDN U9901 ( .B(n8330), .A(n587), .Z(n8328) );
  XNOR U9902 ( .A(a[477]), .B(n8331), .Z(n587) );
  IV U9903 ( .A(n8329), .Z(n8331) );
  XNOR U9904 ( .A(b[477]), .B(n8329), .Z(n8330) );
  XOR U9905 ( .A(n8332), .B(n8333), .Z(n8329) );
  ANDN U9906 ( .B(n8334), .A(n588), .Z(n8332) );
  XNOR U9907 ( .A(a[476]), .B(n8335), .Z(n588) );
  IV U9908 ( .A(n8333), .Z(n8335) );
  XNOR U9909 ( .A(b[476]), .B(n8333), .Z(n8334) );
  XOR U9910 ( .A(n8336), .B(n8337), .Z(n8333) );
  ANDN U9911 ( .B(n8338), .A(n589), .Z(n8336) );
  XNOR U9912 ( .A(a[475]), .B(n8339), .Z(n589) );
  IV U9913 ( .A(n8337), .Z(n8339) );
  XNOR U9914 ( .A(b[475]), .B(n8337), .Z(n8338) );
  XOR U9915 ( .A(n8340), .B(n8341), .Z(n8337) );
  ANDN U9916 ( .B(n8342), .A(n590), .Z(n8340) );
  XNOR U9917 ( .A(a[474]), .B(n8343), .Z(n590) );
  IV U9918 ( .A(n8341), .Z(n8343) );
  XNOR U9919 ( .A(b[474]), .B(n8341), .Z(n8342) );
  XOR U9920 ( .A(n8344), .B(n8345), .Z(n8341) );
  ANDN U9921 ( .B(n8346), .A(n591), .Z(n8344) );
  XNOR U9922 ( .A(a[473]), .B(n8347), .Z(n591) );
  IV U9923 ( .A(n8345), .Z(n8347) );
  XNOR U9924 ( .A(b[473]), .B(n8345), .Z(n8346) );
  XOR U9925 ( .A(n8348), .B(n8349), .Z(n8345) );
  ANDN U9926 ( .B(n8350), .A(n592), .Z(n8348) );
  XNOR U9927 ( .A(a[472]), .B(n8351), .Z(n592) );
  IV U9928 ( .A(n8349), .Z(n8351) );
  XNOR U9929 ( .A(b[472]), .B(n8349), .Z(n8350) );
  XOR U9930 ( .A(n8352), .B(n8353), .Z(n8349) );
  ANDN U9931 ( .B(n8354), .A(n593), .Z(n8352) );
  XNOR U9932 ( .A(a[471]), .B(n8355), .Z(n593) );
  IV U9933 ( .A(n8353), .Z(n8355) );
  XNOR U9934 ( .A(b[471]), .B(n8353), .Z(n8354) );
  XOR U9935 ( .A(n8356), .B(n8357), .Z(n8353) );
  ANDN U9936 ( .B(n8358), .A(n594), .Z(n8356) );
  XNOR U9937 ( .A(a[470]), .B(n8359), .Z(n594) );
  IV U9938 ( .A(n8357), .Z(n8359) );
  XNOR U9939 ( .A(b[470]), .B(n8357), .Z(n8358) );
  XOR U9940 ( .A(n8360), .B(n8361), .Z(n8357) );
  ANDN U9941 ( .B(n8362), .A(n596), .Z(n8360) );
  XNOR U9942 ( .A(a[469]), .B(n8363), .Z(n596) );
  IV U9943 ( .A(n8361), .Z(n8363) );
  XNOR U9944 ( .A(b[469]), .B(n8361), .Z(n8362) );
  XOR U9945 ( .A(n8364), .B(n8365), .Z(n8361) );
  ANDN U9946 ( .B(n8366), .A(n597), .Z(n8364) );
  XNOR U9947 ( .A(a[468]), .B(n8367), .Z(n597) );
  IV U9948 ( .A(n8365), .Z(n8367) );
  XNOR U9949 ( .A(b[468]), .B(n8365), .Z(n8366) );
  XOR U9950 ( .A(n8368), .B(n8369), .Z(n8365) );
  ANDN U9951 ( .B(n8370), .A(n598), .Z(n8368) );
  XNOR U9952 ( .A(a[467]), .B(n8371), .Z(n598) );
  IV U9953 ( .A(n8369), .Z(n8371) );
  XNOR U9954 ( .A(b[467]), .B(n8369), .Z(n8370) );
  XOR U9955 ( .A(n8372), .B(n8373), .Z(n8369) );
  ANDN U9956 ( .B(n8374), .A(n599), .Z(n8372) );
  XNOR U9957 ( .A(a[466]), .B(n8375), .Z(n599) );
  IV U9958 ( .A(n8373), .Z(n8375) );
  XNOR U9959 ( .A(b[466]), .B(n8373), .Z(n8374) );
  XOR U9960 ( .A(n8376), .B(n8377), .Z(n8373) );
  ANDN U9961 ( .B(n8378), .A(n600), .Z(n8376) );
  XNOR U9962 ( .A(a[465]), .B(n8379), .Z(n600) );
  IV U9963 ( .A(n8377), .Z(n8379) );
  XNOR U9964 ( .A(b[465]), .B(n8377), .Z(n8378) );
  XOR U9965 ( .A(n8380), .B(n8381), .Z(n8377) );
  ANDN U9966 ( .B(n8382), .A(n601), .Z(n8380) );
  XNOR U9967 ( .A(a[464]), .B(n8383), .Z(n601) );
  IV U9968 ( .A(n8381), .Z(n8383) );
  XNOR U9969 ( .A(b[464]), .B(n8381), .Z(n8382) );
  XOR U9970 ( .A(n8384), .B(n8385), .Z(n8381) );
  ANDN U9971 ( .B(n8386), .A(n602), .Z(n8384) );
  XNOR U9972 ( .A(a[463]), .B(n8387), .Z(n602) );
  IV U9973 ( .A(n8385), .Z(n8387) );
  XNOR U9974 ( .A(b[463]), .B(n8385), .Z(n8386) );
  XOR U9975 ( .A(n8388), .B(n8389), .Z(n8385) );
  ANDN U9976 ( .B(n8390), .A(n603), .Z(n8388) );
  XNOR U9977 ( .A(a[462]), .B(n8391), .Z(n603) );
  IV U9978 ( .A(n8389), .Z(n8391) );
  XNOR U9979 ( .A(b[462]), .B(n8389), .Z(n8390) );
  XOR U9980 ( .A(n8392), .B(n8393), .Z(n8389) );
  ANDN U9981 ( .B(n8394), .A(n604), .Z(n8392) );
  XNOR U9982 ( .A(a[461]), .B(n8395), .Z(n604) );
  IV U9983 ( .A(n8393), .Z(n8395) );
  XNOR U9984 ( .A(b[461]), .B(n8393), .Z(n8394) );
  XOR U9985 ( .A(n8396), .B(n8397), .Z(n8393) );
  ANDN U9986 ( .B(n8398), .A(n605), .Z(n8396) );
  XNOR U9987 ( .A(a[460]), .B(n8399), .Z(n605) );
  IV U9988 ( .A(n8397), .Z(n8399) );
  XNOR U9989 ( .A(b[460]), .B(n8397), .Z(n8398) );
  XOR U9990 ( .A(n8400), .B(n8401), .Z(n8397) );
  ANDN U9991 ( .B(n8402), .A(n607), .Z(n8400) );
  XNOR U9992 ( .A(a[459]), .B(n8403), .Z(n607) );
  IV U9993 ( .A(n8401), .Z(n8403) );
  XNOR U9994 ( .A(b[459]), .B(n8401), .Z(n8402) );
  XOR U9995 ( .A(n8404), .B(n8405), .Z(n8401) );
  ANDN U9996 ( .B(n8406), .A(n608), .Z(n8404) );
  XNOR U9997 ( .A(a[458]), .B(n8407), .Z(n608) );
  IV U9998 ( .A(n8405), .Z(n8407) );
  XNOR U9999 ( .A(b[458]), .B(n8405), .Z(n8406) );
  XOR U10000 ( .A(n8408), .B(n8409), .Z(n8405) );
  ANDN U10001 ( .B(n8410), .A(n609), .Z(n8408) );
  XNOR U10002 ( .A(a[457]), .B(n8411), .Z(n609) );
  IV U10003 ( .A(n8409), .Z(n8411) );
  XNOR U10004 ( .A(b[457]), .B(n8409), .Z(n8410) );
  XOR U10005 ( .A(n8412), .B(n8413), .Z(n8409) );
  ANDN U10006 ( .B(n8414), .A(n610), .Z(n8412) );
  XNOR U10007 ( .A(a[456]), .B(n8415), .Z(n610) );
  IV U10008 ( .A(n8413), .Z(n8415) );
  XNOR U10009 ( .A(b[456]), .B(n8413), .Z(n8414) );
  XOR U10010 ( .A(n8416), .B(n8417), .Z(n8413) );
  ANDN U10011 ( .B(n8418), .A(n611), .Z(n8416) );
  XNOR U10012 ( .A(a[455]), .B(n8419), .Z(n611) );
  IV U10013 ( .A(n8417), .Z(n8419) );
  XNOR U10014 ( .A(b[455]), .B(n8417), .Z(n8418) );
  XOR U10015 ( .A(n8420), .B(n8421), .Z(n8417) );
  ANDN U10016 ( .B(n8422), .A(n612), .Z(n8420) );
  XNOR U10017 ( .A(a[454]), .B(n8423), .Z(n612) );
  IV U10018 ( .A(n8421), .Z(n8423) );
  XNOR U10019 ( .A(b[454]), .B(n8421), .Z(n8422) );
  XOR U10020 ( .A(n8424), .B(n8425), .Z(n8421) );
  ANDN U10021 ( .B(n8426), .A(n613), .Z(n8424) );
  XNOR U10022 ( .A(a[453]), .B(n8427), .Z(n613) );
  IV U10023 ( .A(n8425), .Z(n8427) );
  XNOR U10024 ( .A(b[453]), .B(n8425), .Z(n8426) );
  XOR U10025 ( .A(n8428), .B(n8429), .Z(n8425) );
  ANDN U10026 ( .B(n8430), .A(n614), .Z(n8428) );
  XNOR U10027 ( .A(a[452]), .B(n8431), .Z(n614) );
  IV U10028 ( .A(n8429), .Z(n8431) );
  XNOR U10029 ( .A(b[452]), .B(n8429), .Z(n8430) );
  XOR U10030 ( .A(n8432), .B(n8433), .Z(n8429) );
  ANDN U10031 ( .B(n8434), .A(n615), .Z(n8432) );
  XNOR U10032 ( .A(a[451]), .B(n8435), .Z(n615) );
  IV U10033 ( .A(n8433), .Z(n8435) );
  XNOR U10034 ( .A(b[451]), .B(n8433), .Z(n8434) );
  XOR U10035 ( .A(n8436), .B(n8437), .Z(n8433) );
  ANDN U10036 ( .B(n8438), .A(n616), .Z(n8436) );
  XNOR U10037 ( .A(a[450]), .B(n8439), .Z(n616) );
  IV U10038 ( .A(n8437), .Z(n8439) );
  XNOR U10039 ( .A(b[450]), .B(n8437), .Z(n8438) );
  XOR U10040 ( .A(n8440), .B(n8441), .Z(n8437) );
  ANDN U10041 ( .B(n8442), .A(n618), .Z(n8440) );
  XNOR U10042 ( .A(a[449]), .B(n8443), .Z(n618) );
  IV U10043 ( .A(n8441), .Z(n8443) );
  XNOR U10044 ( .A(b[449]), .B(n8441), .Z(n8442) );
  XOR U10045 ( .A(n8444), .B(n8445), .Z(n8441) );
  ANDN U10046 ( .B(n8446), .A(n619), .Z(n8444) );
  XNOR U10047 ( .A(a[448]), .B(n8447), .Z(n619) );
  IV U10048 ( .A(n8445), .Z(n8447) );
  XNOR U10049 ( .A(b[448]), .B(n8445), .Z(n8446) );
  XOR U10050 ( .A(n8448), .B(n8449), .Z(n8445) );
  ANDN U10051 ( .B(n8450), .A(n620), .Z(n8448) );
  XNOR U10052 ( .A(a[447]), .B(n8451), .Z(n620) );
  IV U10053 ( .A(n8449), .Z(n8451) );
  XNOR U10054 ( .A(b[447]), .B(n8449), .Z(n8450) );
  XOR U10055 ( .A(n8452), .B(n8453), .Z(n8449) );
  ANDN U10056 ( .B(n8454), .A(n621), .Z(n8452) );
  XNOR U10057 ( .A(a[446]), .B(n8455), .Z(n621) );
  IV U10058 ( .A(n8453), .Z(n8455) );
  XNOR U10059 ( .A(b[446]), .B(n8453), .Z(n8454) );
  XOR U10060 ( .A(n8456), .B(n8457), .Z(n8453) );
  ANDN U10061 ( .B(n8458), .A(n622), .Z(n8456) );
  XNOR U10062 ( .A(a[445]), .B(n8459), .Z(n622) );
  IV U10063 ( .A(n8457), .Z(n8459) );
  XNOR U10064 ( .A(b[445]), .B(n8457), .Z(n8458) );
  XOR U10065 ( .A(n8460), .B(n8461), .Z(n8457) );
  ANDN U10066 ( .B(n8462), .A(n623), .Z(n8460) );
  XNOR U10067 ( .A(a[444]), .B(n8463), .Z(n623) );
  IV U10068 ( .A(n8461), .Z(n8463) );
  XNOR U10069 ( .A(b[444]), .B(n8461), .Z(n8462) );
  XOR U10070 ( .A(n8464), .B(n8465), .Z(n8461) );
  ANDN U10071 ( .B(n8466), .A(n624), .Z(n8464) );
  XNOR U10072 ( .A(a[443]), .B(n8467), .Z(n624) );
  IV U10073 ( .A(n8465), .Z(n8467) );
  XNOR U10074 ( .A(b[443]), .B(n8465), .Z(n8466) );
  XOR U10075 ( .A(n8468), .B(n8469), .Z(n8465) );
  ANDN U10076 ( .B(n8470), .A(n625), .Z(n8468) );
  XNOR U10077 ( .A(a[442]), .B(n8471), .Z(n625) );
  IV U10078 ( .A(n8469), .Z(n8471) );
  XNOR U10079 ( .A(b[442]), .B(n8469), .Z(n8470) );
  XOR U10080 ( .A(n8472), .B(n8473), .Z(n8469) );
  ANDN U10081 ( .B(n8474), .A(n626), .Z(n8472) );
  XNOR U10082 ( .A(a[441]), .B(n8475), .Z(n626) );
  IV U10083 ( .A(n8473), .Z(n8475) );
  XNOR U10084 ( .A(b[441]), .B(n8473), .Z(n8474) );
  XOR U10085 ( .A(n8476), .B(n8477), .Z(n8473) );
  ANDN U10086 ( .B(n8478), .A(n627), .Z(n8476) );
  XNOR U10087 ( .A(a[440]), .B(n8479), .Z(n627) );
  IV U10088 ( .A(n8477), .Z(n8479) );
  XNOR U10089 ( .A(b[440]), .B(n8477), .Z(n8478) );
  XOR U10090 ( .A(n8480), .B(n8481), .Z(n8477) );
  ANDN U10091 ( .B(n8482), .A(n629), .Z(n8480) );
  XNOR U10092 ( .A(a[439]), .B(n8483), .Z(n629) );
  IV U10093 ( .A(n8481), .Z(n8483) );
  XNOR U10094 ( .A(b[439]), .B(n8481), .Z(n8482) );
  XOR U10095 ( .A(n8484), .B(n8485), .Z(n8481) );
  ANDN U10096 ( .B(n8486), .A(n630), .Z(n8484) );
  XNOR U10097 ( .A(a[438]), .B(n8487), .Z(n630) );
  IV U10098 ( .A(n8485), .Z(n8487) );
  XNOR U10099 ( .A(b[438]), .B(n8485), .Z(n8486) );
  XOR U10100 ( .A(n8488), .B(n8489), .Z(n8485) );
  ANDN U10101 ( .B(n8490), .A(n631), .Z(n8488) );
  XNOR U10102 ( .A(a[437]), .B(n8491), .Z(n631) );
  IV U10103 ( .A(n8489), .Z(n8491) );
  XNOR U10104 ( .A(b[437]), .B(n8489), .Z(n8490) );
  XOR U10105 ( .A(n8492), .B(n8493), .Z(n8489) );
  ANDN U10106 ( .B(n8494), .A(n632), .Z(n8492) );
  XNOR U10107 ( .A(a[436]), .B(n8495), .Z(n632) );
  IV U10108 ( .A(n8493), .Z(n8495) );
  XNOR U10109 ( .A(b[436]), .B(n8493), .Z(n8494) );
  XOR U10110 ( .A(n8496), .B(n8497), .Z(n8493) );
  ANDN U10111 ( .B(n8498), .A(n633), .Z(n8496) );
  XNOR U10112 ( .A(a[435]), .B(n8499), .Z(n633) );
  IV U10113 ( .A(n8497), .Z(n8499) );
  XNOR U10114 ( .A(b[435]), .B(n8497), .Z(n8498) );
  XOR U10115 ( .A(n8500), .B(n8501), .Z(n8497) );
  ANDN U10116 ( .B(n8502), .A(n634), .Z(n8500) );
  XNOR U10117 ( .A(a[434]), .B(n8503), .Z(n634) );
  IV U10118 ( .A(n8501), .Z(n8503) );
  XNOR U10119 ( .A(b[434]), .B(n8501), .Z(n8502) );
  XOR U10120 ( .A(n8504), .B(n8505), .Z(n8501) );
  ANDN U10121 ( .B(n8506), .A(n635), .Z(n8504) );
  XNOR U10122 ( .A(a[433]), .B(n8507), .Z(n635) );
  IV U10123 ( .A(n8505), .Z(n8507) );
  XNOR U10124 ( .A(b[433]), .B(n8505), .Z(n8506) );
  XOR U10125 ( .A(n8508), .B(n8509), .Z(n8505) );
  ANDN U10126 ( .B(n8510), .A(n636), .Z(n8508) );
  XNOR U10127 ( .A(a[432]), .B(n8511), .Z(n636) );
  IV U10128 ( .A(n8509), .Z(n8511) );
  XNOR U10129 ( .A(b[432]), .B(n8509), .Z(n8510) );
  XOR U10130 ( .A(n8512), .B(n8513), .Z(n8509) );
  ANDN U10131 ( .B(n8514), .A(n637), .Z(n8512) );
  XNOR U10132 ( .A(a[431]), .B(n8515), .Z(n637) );
  IV U10133 ( .A(n8513), .Z(n8515) );
  XNOR U10134 ( .A(b[431]), .B(n8513), .Z(n8514) );
  XOR U10135 ( .A(n8516), .B(n8517), .Z(n8513) );
  ANDN U10136 ( .B(n8518), .A(n638), .Z(n8516) );
  XNOR U10137 ( .A(a[430]), .B(n8519), .Z(n638) );
  IV U10138 ( .A(n8517), .Z(n8519) );
  XNOR U10139 ( .A(b[430]), .B(n8517), .Z(n8518) );
  XOR U10140 ( .A(n8520), .B(n8521), .Z(n8517) );
  ANDN U10141 ( .B(n8522), .A(n640), .Z(n8520) );
  XNOR U10142 ( .A(a[429]), .B(n8523), .Z(n640) );
  IV U10143 ( .A(n8521), .Z(n8523) );
  XNOR U10144 ( .A(b[429]), .B(n8521), .Z(n8522) );
  XOR U10145 ( .A(n8524), .B(n8525), .Z(n8521) );
  ANDN U10146 ( .B(n8526), .A(n641), .Z(n8524) );
  XNOR U10147 ( .A(a[428]), .B(n8527), .Z(n641) );
  IV U10148 ( .A(n8525), .Z(n8527) );
  XNOR U10149 ( .A(b[428]), .B(n8525), .Z(n8526) );
  XOR U10150 ( .A(n8528), .B(n8529), .Z(n8525) );
  ANDN U10151 ( .B(n8530), .A(n642), .Z(n8528) );
  XNOR U10152 ( .A(a[427]), .B(n8531), .Z(n642) );
  IV U10153 ( .A(n8529), .Z(n8531) );
  XNOR U10154 ( .A(b[427]), .B(n8529), .Z(n8530) );
  XOR U10155 ( .A(n8532), .B(n8533), .Z(n8529) );
  ANDN U10156 ( .B(n8534), .A(n643), .Z(n8532) );
  XNOR U10157 ( .A(a[426]), .B(n8535), .Z(n643) );
  IV U10158 ( .A(n8533), .Z(n8535) );
  XNOR U10159 ( .A(b[426]), .B(n8533), .Z(n8534) );
  XOR U10160 ( .A(n8536), .B(n8537), .Z(n8533) );
  ANDN U10161 ( .B(n8538), .A(n644), .Z(n8536) );
  XNOR U10162 ( .A(a[425]), .B(n8539), .Z(n644) );
  IV U10163 ( .A(n8537), .Z(n8539) );
  XNOR U10164 ( .A(b[425]), .B(n8537), .Z(n8538) );
  XOR U10165 ( .A(n8540), .B(n8541), .Z(n8537) );
  ANDN U10166 ( .B(n8542), .A(n645), .Z(n8540) );
  XNOR U10167 ( .A(a[424]), .B(n8543), .Z(n645) );
  IV U10168 ( .A(n8541), .Z(n8543) );
  XNOR U10169 ( .A(b[424]), .B(n8541), .Z(n8542) );
  XOR U10170 ( .A(n8544), .B(n8545), .Z(n8541) );
  ANDN U10171 ( .B(n8546), .A(n646), .Z(n8544) );
  XNOR U10172 ( .A(a[423]), .B(n8547), .Z(n646) );
  IV U10173 ( .A(n8545), .Z(n8547) );
  XNOR U10174 ( .A(b[423]), .B(n8545), .Z(n8546) );
  XOR U10175 ( .A(n8548), .B(n8549), .Z(n8545) );
  ANDN U10176 ( .B(n8550), .A(n647), .Z(n8548) );
  XNOR U10177 ( .A(a[422]), .B(n8551), .Z(n647) );
  IV U10178 ( .A(n8549), .Z(n8551) );
  XNOR U10179 ( .A(b[422]), .B(n8549), .Z(n8550) );
  XOR U10180 ( .A(n8552), .B(n8553), .Z(n8549) );
  ANDN U10181 ( .B(n8554), .A(n648), .Z(n8552) );
  XNOR U10182 ( .A(a[421]), .B(n8555), .Z(n648) );
  IV U10183 ( .A(n8553), .Z(n8555) );
  XNOR U10184 ( .A(b[421]), .B(n8553), .Z(n8554) );
  XOR U10185 ( .A(n8556), .B(n8557), .Z(n8553) );
  ANDN U10186 ( .B(n8558), .A(n649), .Z(n8556) );
  XNOR U10187 ( .A(a[420]), .B(n8559), .Z(n649) );
  IV U10188 ( .A(n8557), .Z(n8559) );
  XNOR U10189 ( .A(b[420]), .B(n8557), .Z(n8558) );
  XOR U10190 ( .A(n8560), .B(n8561), .Z(n8557) );
  ANDN U10191 ( .B(n8562), .A(n651), .Z(n8560) );
  XNOR U10192 ( .A(a[419]), .B(n8563), .Z(n651) );
  IV U10193 ( .A(n8561), .Z(n8563) );
  XNOR U10194 ( .A(b[419]), .B(n8561), .Z(n8562) );
  XOR U10195 ( .A(n8564), .B(n8565), .Z(n8561) );
  ANDN U10196 ( .B(n8566), .A(n652), .Z(n8564) );
  XNOR U10197 ( .A(a[418]), .B(n8567), .Z(n652) );
  IV U10198 ( .A(n8565), .Z(n8567) );
  XNOR U10199 ( .A(b[418]), .B(n8565), .Z(n8566) );
  XOR U10200 ( .A(n8568), .B(n8569), .Z(n8565) );
  ANDN U10201 ( .B(n8570), .A(n653), .Z(n8568) );
  XNOR U10202 ( .A(a[417]), .B(n8571), .Z(n653) );
  IV U10203 ( .A(n8569), .Z(n8571) );
  XNOR U10204 ( .A(b[417]), .B(n8569), .Z(n8570) );
  XOR U10205 ( .A(n8572), .B(n8573), .Z(n8569) );
  ANDN U10206 ( .B(n8574), .A(n654), .Z(n8572) );
  XNOR U10207 ( .A(a[416]), .B(n8575), .Z(n654) );
  IV U10208 ( .A(n8573), .Z(n8575) );
  XNOR U10209 ( .A(b[416]), .B(n8573), .Z(n8574) );
  XOR U10210 ( .A(n8576), .B(n8577), .Z(n8573) );
  ANDN U10211 ( .B(n8578), .A(n655), .Z(n8576) );
  XNOR U10212 ( .A(a[415]), .B(n8579), .Z(n655) );
  IV U10213 ( .A(n8577), .Z(n8579) );
  XNOR U10214 ( .A(b[415]), .B(n8577), .Z(n8578) );
  XOR U10215 ( .A(n8580), .B(n8581), .Z(n8577) );
  ANDN U10216 ( .B(n8582), .A(n656), .Z(n8580) );
  XNOR U10217 ( .A(a[414]), .B(n8583), .Z(n656) );
  IV U10218 ( .A(n8581), .Z(n8583) );
  XNOR U10219 ( .A(b[414]), .B(n8581), .Z(n8582) );
  XOR U10220 ( .A(n8584), .B(n8585), .Z(n8581) );
  ANDN U10221 ( .B(n8586), .A(n657), .Z(n8584) );
  XNOR U10222 ( .A(a[413]), .B(n8587), .Z(n657) );
  IV U10223 ( .A(n8585), .Z(n8587) );
  XNOR U10224 ( .A(b[413]), .B(n8585), .Z(n8586) );
  XOR U10225 ( .A(n8588), .B(n8589), .Z(n8585) );
  ANDN U10226 ( .B(n8590), .A(n658), .Z(n8588) );
  XNOR U10227 ( .A(a[412]), .B(n8591), .Z(n658) );
  IV U10228 ( .A(n8589), .Z(n8591) );
  XNOR U10229 ( .A(b[412]), .B(n8589), .Z(n8590) );
  XOR U10230 ( .A(n8592), .B(n8593), .Z(n8589) );
  ANDN U10231 ( .B(n8594), .A(n659), .Z(n8592) );
  XNOR U10232 ( .A(a[411]), .B(n8595), .Z(n659) );
  IV U10233 ( .A(n8593), .Z(n8595) );
  XNOR U10234 ( .A(b[411]), .B(n8593), .Z(n8594) );
  XOR U10235 ( .A(n8596), .B(n8597), .Z(n8593) );
  ANDN U10236 ( .B(n8598), .A(n660), .Z(n8596) );
  XNOR U10237 ( .A(a[410]), .B(n8599), .Z(n660) );
  IV U10238 ( .A(n8597), .Z(n8599) );
  XNOR U10239 ( .A(b[410]), .B(n8597), .Z(n8598) );
  XOR U10240 ( .A(n8600), .B(n8601), .Z(n8597) );
  ANDN U10241 ( .B(n8602), .A(n662), .Z(n8600) );
  XNOR U10242 ( .A(a[409]), .B(n8603), .Z(n662) );
  IV U10243 ( .A(n8601), .Z(n8603) );
  XNOR U10244 ( .A(b[409]), .B(n8601), .Z(n8602) );
  XOR U10245 ( .A(n8604), .B(n8605), .Z(n8601) );
  ANDN U10246 ( .B(n8606), .A(n663), .Z(n8604) );
  XNOR U10247 ( .A(a[408]), .B(n8607), .Z(n663) );
  IV U10248 ( .A(n8605), .Z(n8607) );
  XNOR U10249 ( .A(b[408]), .B(n8605), .Z(n8606) );
  XOR U10250 ( .A(n8608), .B(n8609), .Z(n8605) );
  ANDN U10251 ( .B(n8610), .A(n664), .Z(n8608) );
  XNOR U10252 ( .A(a[407]), .B(n8611), .Z(n664) );
  IV U10253 ( .A(n8609), .Z(n8611) );
  XNOR U10254 ( .A(b[407]), .B(n8609), .Z(n8610) );
  XOR U10255 ( .A(n8612), .B(n8613), .Z(n8609) );
  ANDN U10256 ( .B(n8614), .A(n665), .Z(n8612) );
  XNOR U10257 ( .A(a[406]), .B(n8615), .Z(n665) );
  IV U10258 ( .A(n8613), .Z(n8615) );
  XNOR U10259 ( .A(b[406]), .B(n8613), .Z(n8614) );
  XOR U10260 ( .A(n8616), .B(n8617), .Z(n8613) );
  ANDN U10261 ( .B(n8618), .A(n666), .Z(n8616) );
  XNOR U10262 ( .A(a[405]), .B(n8619), .Z(n666) );
  IV U10263 ( .A(n8617), .Z(n8619) );
  XNOR U10264 ( .A(b[405]), .B(n8617), .Z(n8618) );
  XOR U10265 ( .A(n8620), .B(n8621), .Z(n8617) );
  ANDN U10266 ( .B(n8622), .A(n667), .Z(n8620) );
  XNOR U10267 ( .A(a[404]), .B(n8623), .Z(n667) );
  IV U10268 ( .A(n8621), .Z(n8623) );
  XNOR U10269 ( .A(b[404]), .B(n8621), .Z(n8622) );
  XOR U10270 ( .A(n8624), .B(n8625), .Z(n8621) );
  ANDN U10271 ( .B(n8626), .A(n668), .Z(n8624) );
  XNOR U10272 ( .A(a[403]), .B(n8627), .Z(n668) );
  IV U10273 ( .A(n8625), .Z(n8627) );
  XNOR U10274 ( .A(b[403]), .B(n8625), .Z(n8626) );
  XOR U10275 ( .A(n8628), .B(n8629), .Z(n8625) );
  ANDN U10276 ( .B(n8630), .A(n669), .Z(n8628) );
  XNOR U10277 ( .A(a[402]), .B(n8631), .Z(n669) );
  IV U10278 ( .A(n8629), .Z(n8631) );
  XNOR U10279 ( .A(b[402]), .B(n8629), .Z(n8630) );
  XOR U10280 ( .A(n8632), .B(n8633), .Z(n8629) );
  ANDN U10281 ( .B(n8634), .A(n670), .Z(n8632) );
  XNOR U10282 ( .A(a[401]), .B(n8635), .Z(n670) );
  IV U10283 ( .A(n8633), .Z(n8635) );
  XNOR U10284 ( .A(b[401]), .B(n8633), .Z(n8634) );
  XOR U10285 ( .A(n8636), .B(n8637), .Z(n8633) );
  ANDN U10286 ( .B(n8638), .A(n671), .Z(n8636) );
  XNOR U10287 ( .A(a[400]), .B(n8639), .Z(n671) );
  IV U10288 ( .A(n8637), .Z(n8639) );
  XNOR U10289 ( .A(b[400]), .B(n8637), .Z(n8638) );
  XOR U10290 ( .A(n8640), .B(n8641), .Z(n8637) );
  ANDN U10291 ( .B(n8642), .A(n674), .Z(n8640) );
  XNOR U10292 ( .A(a[399]), .B(n8643), .Z(n674) );
  IV U10293 ( .A(n8641), .Z(n8643) );
  XNOR U10294 ( .A(b[399]), .B(n8641), .Z(n8642) );
  XOR U10295 ( .A(n8644), .B(n8645), .Z(n8641) );
  ANDN U10296 ( .B(n8646), .A(n675), .Z(n8644) );
  XNOR U10297 ( .A(a[398]), .B(n8647), .Z(n675) );
  IV U10298 ( .A(n8645), .Z(n8647) );
  XNOR U10299 ( .A(b[398]), .B(n8645), .Z(n8646) );
  XOR U10300 ( .A(n8648), .B(n8649), .Z(n8645) );
  ANDN U10301 ( .B(n8650), .A(n676), .Z(n8648) );
  XNOR U10302 ( .A(a[397]), .B(n8651), .Z(n676) );
  IV U10303 ( .A(n8649), .Z(n8651) );
  XNOR U10304 ( .A(b[397]), .B(n8649), .Z(n8650) );
  XOR U10305 ( .A(n8652), .B(n8653), .Z(n8649) );
  ANDN U10306 ( .B(n8654), .A(n677), .Z(n8652) );
  XNOR U10307 ( .A(a[396]), .B(n8655), .Z(n677) );
  IV U10308 ( .A(n8653), .Z(n8655) );
  XNOR U10309 ( .A(b[396]), .B(n8653), .Z(n8654) );
  XOR U10310 ( .A(n8656), .B(n8657), .Z(n8653) );
  ANDN U10311 ( .B(n8658), .A(n678), .Z(n8656) );
  XNOR U10312 ( .A(a[395]), .B(n8659), .Z(n678) );
  IV U10313 ( .A(n8657), .Z(n8659) );
  XNOR U10314 ( .A(b[395]), .B(n8657), .Z(n8658) );
  XOR U10315 ( .A(n8660), .B(n8661), .Z(n8657) );
  ANDN U10316 ( .B(n8662), .A(n679), .Z(n8660) );
  XNOR U10317 ( .A(a[394]), .B(n8663), .Z(n679) );
  IV U10318 ( .A(n8661), .Z(n8663) );
  XNOR U10319 ( .A(b[394]), .B(n8661), .Z(n8662) );
  XOR U10320 ( .A(n8664), .B(n8665), .Z(n8661) );
  ANDN U10321 ( .B(n8666), .A(n680), .Z(n8664) );
  XNOR U10322 ( .A(a[393]), .B(n8667), .Z(n680) );
  IV U10323 ( .A(n8665), .Z(n8667) );
  XNOR U10324 ( .A(b[393]), .B(n8665), .Z(n8666) );
  XOR U10325 ( .A(n8668), .B(n8669), .Z(n8665) );
  ANDN U10326 ( .B(n8670), .A(n681), .Z(n8668) );
  XNOR U10327 ( .A(a[392]), .B(n8671), .Z(n681) );
  IV U10328 ( .A(n8669), .Z(n8671) );
  XNOR U10329 ( .A(b[392]), .B(n8669), .Z(n8670) );
  XOR U10330 ( .A(n8672), .B(n8673), .Z(n8669) );
  ANDN U10331 ( .B(n8674), .A(n682), .Z(n8672) );
  XNOR U10332 ( .A(a[391]), .B(n8675), .Z(n682) );
  IV U10333 ( .A(n8673), .Z(n8675) );
  XNOR U10334 ( .A(b[391]), .B(n8673), .Z(n8674) );
  XOR U10335 ( .A(n8676), .B(n8677), .Z(n8673) );
  ANDN U10336 ( .B(n8678), .A(n683), .Z(n8676) );
  XNOR U10337 ( .A(a[390]), .B(n8679), .Z(n683) );
  IV U10338 ( .A(n8677), .Z(n8679) );
  XNOR U10339 ( .A(b[390]), .B(n8677), .Z(n8678) );
  XOR U10340 ( .A(n8680), .B(n8681), .Z(n8677) );
  ANDN U10341 ( .B(n8682), .A(n685), .Z(n8680) );
  XNOR U10342 ( .A(a[389]), .B(n8683), .Z(n685) );
  IV U10343 ( .A(n8681), .Z(n8683) );
  XNOR U10344 ( .A(b[389]), .B(n8681), .Z(n8682) );
  XOR U10345 ( .A(n8684), .B(n8685), .Z(n8681) );
  ANDN U10346 ( .B(n8686), .A(n686), .Z(n8684) );
  XNOR U10347 ( .A(a[388]), .B(n8687), .Z(n686) );
  IV U10348 ( .A(n8685), .Z(n8687) );
  XNOR U10349 ( .A(b[388]), .B(n8685), .Z(n8686) );
  XOR U10350 ( .A(n8688), .B(n8689), .Z(n8685) );
  ANDN U10351 ( .B(n8690), .A(n687), .Z(n8688) );
  XNOR U10352 ( .A(a[387]), .B(n8691), .Z(n687) );
  IV U10353 ( .A(n8689), .Z(n8691) );
  XNOR U10354 ( .A(b[387]), .B(n8689), .Z(n8690) );
  XOR U10355 ( .A(n8692), .B(n8693), .Z(n8689) );
  ANDN U10356 ( .B(n8694), .A(n688), .Z(n8692) );
  XNOR U10357 ( .A(a[386]), .B(n8695), .Z(n688) );
  IV U10358 ( .A(n8693), .Z(n8695) );
  XNOR U10359 ( .A(b[386]), .B(n8693), .Z(n8694) );
  XOR U10360 ( .A(n8696), .B(n8697), .Z(n8693) );
  ANDN U10361 ( .B(n8698), .A(n689), .Z(n8696) );
  XNOR U10362 ( .A(a[385]), .B(n8699), .Z(n689) );
  IV U10363 ( .A(n8697), .Z(n8699) );
  XNOR U10364 ( .A(b[385]), .B(n8697), .Z(n8698) );
  XOR U10365 ( .A(n8700), .B(n8701), .Z(n8697) );
  ANDN U10366 ( .B(n8702), .A(n690), .Z(n8700) );
  XNOR U10367 ( .A(a[384]), .B(n8703), .Z(n690) );
  IV U10368 ( .A(n8701), .Z(n8703) );
  XNOR U10369 ( .A(b[384]), .B(n8701), .Z(n8702) );
  XOR U10370 ( .A(n8704), .B(n8705), .Z(n8701) );
  ANDN U10371 ( .B(n8706), .A(n691), .Z(n8704) );
  XNOR U10372 ( .A(a[383]), .B(n8707), .Z(n691) );
  IV U10373 ( .A(n8705), .Z(n8707) );
  XNOR U10374 ( .A(b[383]), .B(n8705), .Z(n8706) );
  XOR U10375 ( .A(n8708), .B(n8709), .Z(n8705) );
  ANDN U10376 ( .B(n8710), .A(n692), .Z(n8708) );
  XNOR U10377 ( .A(a[382]), .B(n8711), .Z(n692) );
  IV U10378 ( .A(n8709), .Z(n8711) );
  XNOR U10379 ( .A(b[382]), .B(n8709), .Z(n8710) );
  XOR U10380 ( .A(n8712), .B(n8713), .Z(n8709) );
  ANDN U10381 ( .B(n8714), .A(n693), .Z(n8712) );
  XNOR U10382 ( .A(a[381]), .B(n8715), .Z(n693) );
  IV U10383 ( .A(n8713), .Z(n8715) );
  XNOR U10384 ( .A(b[381]), .B(n8713), .Z(n8714) );
  XOR U10385 ( .A(n8716), .B(n8717), .Z(n8713) );
  ANDN U10386 ( .B(n8718), .A(n694), .Z(n8716) );
  XNOR U10387 ( .A(a[380]), .B(n8719), .Z(n694) );
  IV U10388 ( .A(n8717), .Z(n8719) );
  XNOR U10389 ( .A(b[380]), .B(n8717), .Z(n8718) );
  XOR U10390 ( .A(n8720), .B(n8721), .Z(n8717) );
  ANDN U10391 ( .B(n8722), .A(n696), .Z(n8720) );
  XNOR U10392 ( .A(a[379]), .B(n8723), .Z(n696) );
  IV U10393 ( .A(n8721), .Z(n8723) );
  XNOR U10394 ( .A(b[379]), .B(n8721), .Z(n8722) );
  XOR U10395 ( .A(n8724), .B(n8725), .Z(n8721) );
  ANDN U10396 ( .B(n8726), .A(n697), .Z(n8724) );
  XNOR U10397 ( .A(a[378]), .B(n8727), .Z(n697) );
  IV U10398 ( .A(n8725), .Z(n8727) );
  XNOR U10399 ( .A(b[378]), .B(n8725), .Z(n8726) );
  XOR U10400 ( .A(n8728), .B(n8729), .Z(n8725) );
  ANDN U10401 ( .B(n8730), .A(n698), .Z(n8728) );
  XNOR U10402 ( .A(a[377]), .B(n8731), .Z(n698) );
  IV U10403 ( .A(n8729), .Z(n8731) );
  XNOR U10404 ( .A(b[377]), .B(n8729), .Z(n8730) );
  XOR U10405 ( .A(n8732), .B(n8733), .Z(n8729) );
  ANDN U10406 ( .B(n8734), .A(n699), .Z(n8732) );
  XNOR U10407 ( .A(a[376]), .B(n8735), .Z(n699) );
  IV U10408 ( .A(n8733), .Z(n8735) );
  XNOR U10409 ( .A(b[376]), .B(n8733), .Z(n8734) );
  XOR U10410 ( .A(n8736), .B(n8737), .Z(n8733) );
  ANDN U10411 ( .B(n8738), .A(n700), .Z(n8736) );
  XNOR U10412 ( .A(a[375]), .B(n8739), .Z(n700) );
  IV U10413 ( .A(n8737), .Z(n8739) );
  XNOR U10414 ( .A(b[375]), .B(n8737), .Z(n8738) );
  XOR U10415 ( .A(n8740), .B(n8741), .Z(n8737) );
  ANDN U10416 ( .B(n8742), .A(n701), .Z(n8740) );
  XNOR U10417 ( .A(a[374]), .B(n8743), .Z(n701) );
  IV U10418 ( .A(n8741), .Z(n8743) );
  XNOR U10419 ( .A(b[374]), .B(n8741), .Z(n8742) );
  XOR U10420 ( .A(n8744), .B(n8745), .Z(n8741) );
  ANDN U10421 ( .B(n8746), .A(n702), .Z(n8744) );
  XNOR U10422 ( .A(a[373]), .B(n8747), .Z(n702) );
  IV U10423 ( .A(n8745), .Z(n8747) );
  XNOR U10424 ( .A(b[373]), .B(n8745), .Z(n8746) );
  XOR U10425 ( .A(n8748), .B(n8749), .Z(n8745) );
  ANDN U10426 ( .B(n8750), .A(n703), .Z(n8748) );
  XNOR U10427 ( .A(a[372]), .B(n8751), .Z(n703) );
  IV U10428 ( .A(n8749), .Z(n8751) );
  XNOR U10429 ( .A(b[372]), .B(n8749), .Z(n8750) );
  XOR U10430 ( .A(n8752), .B(n8753), .Z(n8749) );
  ANDN U10431 ( .B(n8754), .A(n704), .Z(n8752) );
  XNOR U10432 ( .A(a[371]), .B(n8755), .Z(n704) );
  IV U10433 ( .A(n8753), .Z(n8755) );
  XNOR U10434 ( .A(b[371]), .B(n8753), .Z(n8754) );
  XOR U10435 ( .A(n8756), .B(n8757), .Z(n8753) );
  ANDN U10436 ( .B(n8758), .A(n705), .Z(n8756) );
  XNOR U10437 ( .A(a[370]), .B(n8759), .Z(n705) );
  IV U10438 ( .A(n8757), .Z(n8759) );
  XNOR U10439 ( .A(b[370]), .B(n8757), .Z(n8758) );
  XOR U10440 ( .A(n8760), .B(n8761), .Z(n8757) );
  ANDN U10441 ( .B(n8762), .A(n707), .Z(n8760) );
  XNOR U10442 ( .A(a[369]), .B(n8763), .Z(n707) );
  IV U10443 ( .A(n8761), .Z(n8763) );
  XNOR U10444 ( .A(b[369]), .B(n8761), .Z(n8762) );
  XOR U10445 ( .A(n8764), .B(n8765), .Z(n8761) );
  ANDN U10446 ( .B(n8766), .A(n708), .Z(n8764) );
  XNOR U10447 ( .A(a[368]), .B(n8767), .Z(n708) );
  IV U10448 ( .A(n8765), .Z(n8767) );
  XNOR U10449 ( .A(b[368]), .B(n8765), .Z(n8766) );
  XOR U10450 ( .A(n8768), .B(n8769), .Z(n8765) );
  ANDN U10451 ( .B(n8770), .A(n709), .Z(n8768) );
  XNOR U10452 ( .A(a[367]), .B(n8771), .Z(n709) );
  IV U10453 ( .A(n8769), .Z(n8771) );
  XNOR U10454 ( .A(b[367]), .B(n8769), .Z(n8770) );
  XOR U10455 ( .A(n8772), .B(n8773), .Z(n8769) );
  ANDN U10456 ( .B(n8774), .A(n710), .Z(n8772) );
  XNOR U10457 ( .A(a[366]), .B(n8775), .Z(n710) );
  IV U10458 ( .A(n8773), .Z(n8775) );
  XNOR U10459 ( .A(b[366]), .B(n8773), .Z(n8774) );
  XOR U10460 ( .A(n8776), .B(n8777), .Z(n8773) );
  ANDN U10461 ( .B(n8778), .A(n711), .Z(n8776) );
  XNOR U10462 ( .A(a[365]), .B(n8779), .Z(n711) );
  IV U10463 ( .A(n8777), .Z(n8779) );
  XNOR U10464 ( .A(b[365]), .B(n8777), .Z(n8778) );
  XOR U10465 ( .A(n8780), .B(n8781), .Z(n8777) );
  ANDN U10466 ( .B(n8782), .A(n712), .Z(n8780) );
  XNOR U10467 ( .A(a[364]), .B(n8783), .Z(n712) );
  IV U10468 ( .A(n8781), .Z(n8783) );
  XNOR U10469 ( .A(b[364]), .B(n8781), .Z(n8782) );
  XOR U10470 ( .A(n8784), .B(n8785), .Z(n8781) );
  ANDN U10471 ( .B(n8786), .A(n713), .Z(n8784) );
  XNOR U10472 ( .A(a[363]), .B(n8787), .Z(n713) );
  IV U10473 ( .A(n8785), .Z(n8787) );
  XNOR U10474 ( .A(b[363]), .B(n8785), .Z(n8786) );
  XOR U10475 ( .A(n8788), .B(n8789), .Z(n8785) );
  ANDN U10476 ( .B(n8790), .A(n714), .Z(n8788) );
  XNOR U10477 ( .A(a[362]), .B(n8791), .Z(n714) );
  IV U10478 ( .A(n8789), .Z(n8791) );
  XNOR U10479 ( .A(b[362]), .B(n8789), .Z(n8790) );
  XOR U10480 ( .A(n8792), .B(n8793), .Z(n8789) );
  ANDN U10481 ( .B(n8794), .A(n715), .Z(n8792) );
  XNOR U10482 ( .A(a[361]), .B(n8795), .Z(n715) );
  IV U10483 ( .A(n8793), .Z(n8795) );
  XNOR U10484 ( .A(b[361]), .B(n8793), .Z(n8794) );
  XOR U10485 ( .A(n8796), .B(n8797), .Z(n8793) );
  ANDN U10486 ( .B(n8798), .A(n716), .Z(n8796) );
  XNOR U10487 ( .A(a[360]), .B(n8799), .Z(n716) );
  IV U10488 ( .A(n8797), .Z(n8799) );
  XNOR U10489 ( .A(b[360]), .B(n8797), .Z(n8798) );
  XOR U10490 ( .A(n8800), .B(n8801), .Z(n8797) );
  ANDN U10491 ( .B(n8802), .A(n718), .Z(n8800) );
  XNOR U10492 ( .A(a[359]), .B(n8803), .Z(n718) );
  IV U10493 ( .A(n8801), .Z(n8803) );
  XNOR U10494 ( .A(b[359]), .B(n8801), .Z(n8802) );
  XOR U10495 ( .A(n8804), .B(n8805), .Z(n8801) );
  ANDN U10496 ( .B(n8806), .A(n719), .Z(n8804) );
  XNOR U10497 ( .A(a[358]), .B(n8807), .Z(n719) );
  IV U10498 ( .A(n8805), .Z(n8807) );
  XNOR U10499 ( .A(b[358]), .B(n8805), .Z(n8806) );
  XOR U10500 ( .A(n8808), .B(n8809), .Z(n8805) );
  ANDN U10501 ( .B(n8810), .A(n720), .Z(n8808) );
  XNOR U10502 ( .A(a[357]), .B(n8811), .Z(n720) );
  IV U10503 ( .A(n8809), .Z(n8811) );
  XNOR U10504 ( .A(b[357]), .B(n8809), .Z(n8810) );
  XOR U10505 ( .A(n8812), .B(n8813), .Z(n8809) );
  ANDN U10506 ( .B(n8814), .A(n721), .Z(n8812) );
  XNOR U10507 ( .A(a[356]), .B(n8815), .Z(n721) );
  IV U10508 ( .A(n8813), .Z(n8815) );
  XNOR U10509 ( .A(b[356]), .B(n8813), .Z(n8814) );
  XOR U10510 ( .A(n8816), .B(n8817), .Z(n8813) );
  ANDN U10511 ( .B(n8818), .A(n722), .Z(n8816) );
  XNOR U10512 ( .A(a[355]), .B(n8819), .Z(n722) );
  IV U10513 ( .A(n8817), .Z(n8819) );
  XNOR U10514 ( .A(b[355]), .B(n8817), .Z(n8818) );
  XOR U10515 ( .A(n8820), .B(n8821), .Z(n8817) );
  ANDN U10516 ( .B(n8822), .A(n723), .Z(n8820) );
  XNOR U10517 ( .A(a[354]), .B(n8823), .Z(n723) );
  IV U10518 ( .A(n8821), .Z(n8823) );
  XNOR U10519 ( .A(b[354]), .B(n8821), .Z(n8822) );
  XOR U10520 ( .A(n8824), .B(n8825), .Z(n8821) );
  ANDN U10521 ( .B(n8826), .A(n724), .Z(n8824) );
  XNOR U10522 ( .A(a[353]), .B(n8827), .Z(n724) );
  IV U10523 ( .A(n8825), .Z(n8827) );
  XNOR U10524 ( .A(b[353]), .B(n8825), .Z(n8826) );
  XOR U10525 ( .A(n8828), .B(n8829), .Z(n8825) );
  ANDN U10526 ( .B(n8830), .A(n725), .Z(n8828) );
  XNOR U10527 ( .A(a[352]), .B(n8831), .Z(n725) );
  IV U10528 ( .A(n8829), .Z(n8831) );
  XNOR U10529 ( .A(b[352]), .B(n8829), .Z(n8830) );
  XOR U10530 ( .A(n8832), .B(n8833), .Z(n8829) );
  ANDN U10531 ( .B(n8834), .A(n726), .Z(n8832) );
  XNOR U10532 ( .A(a[351]), .B(n8835), .Z(n726) );
  IV U10533 ( .A(n8833), .Z(n8835) );
  XNOR U10534 ( .A(b[351]), .B(n8833), .Z(n8834) );
  XOR U10535 ( .A(n8836), .B(n8837), .Z(n8833) );
  ANDN U10536 ( .B(n8838), .A(n727), .Z(n8836) );
  XNOR U10537 ( .A(a[350]), .B(n8839), .Z(n727) );
  IV U10538 ( .A(n8837), .Z(n8839) );
  XNOR U10539 ( .A(b[350]), .B(n8837), .Z(n8838) );
  XOR U10540 ( .A(n8840), .B(n8841), .Z(n8837) );
  ANDN U10541 ( .B(n8842), .A(n729), .Z(n8840) );
  XNOR U10542 ( .A(a[349]), .B(n8843), .Z(n729) );
  IV U10543 ( .A(n8841), .Z(n8843) );
  XNOR U10544 ( .A(b[349]), .B(n8841), .Z(n8842) );
  XOR U10545 ( .A(n8844), .B(n8845), .Z(n8841) );
  ANDN U10546 ( .B(n8846), .A(n730), .Z(n8844) );
  XNOR U10547 ( .A(a[348]), .B(n8847), .Z(n730) );
  IV U10548 ( .A(n8845), .Z(n8847) );
  XNOR U10549 ( .A(b[348]), .B(n8845), .Z(n8846) );
  XOR U10550 ( .A(n8848), .B(n8849), .Z(n8845) );
  ANDN U10551 ( .B(n8850), .A(n731), .Z(n8848) );
  XNOR U10552 ( .A(a[347]), .B(n8851), .Z(n731) );
  IV U10553 ( .A(n8849), .Z(n8851) );
  XNOR U10554 ( .A(b[347]), .B(n8849), .Z(n8850) );
  XOR U10555 ( .A(n8852), .B(n8853), .Z(n8849) );
  ANDN U10556 ( .B(n8854), .A(n732), .Z(n8852) );
  XNOR U10557 ( .A(a[346]), .B(n8855), .Z(n732) );
  IV U10558 ( .A(n8853), .Z(n8855) );
  XNOR U10559 ( .A(b[346]), .B(n8853), .Z(n8854) );
  XOR U10560 ( .A(n8856), .B(n8857), .Z(n8853) );
  ANDN U10561 ( .B(n8858), .A(n733), .Z(n8856) );
  XNOR U10562 ( .A(a[345]), .B(n8859), .Z(n733) );
  IV U10563 ( .A(n8857), .Z(n8859) );
  XNOR U10564 ( .A(b[345]), .B(n8857), .Z(n8858) );
  XOR U10565 ( .A(n8860), .B(n8861), .Z(n8857) );
  ANDN U10566 ( .B(n8862), .A(n734), .Z(n8860) );
  XNOR U10567 ( .A(a[344]), .B(n8863), .Z(n734) );
  IV U10568 ( .A(n8861), .Z(n8863) );
  XNOR U10569 ( .A(b[344]), .B(n8861), .Z(n8862) );
  XOR U10570 ( .A(n8864), .B(n8865), .Z(n8861) );
  ANDN U10571 ( .B(n8866), .A(n735), .Z(n8864) );
  XNOR U10572 ( .A(a[343]), .B(n8867), .Z(n735) );
  IV U10573 ( .A(n8865), .Z(n8867) );
  XNOR U10574 ( .A(b[343]), .B(n8865), .Z(n8866) );
  XOR U10575 ( .A(n8868), .B(n8869), .Z(n8865) );
  ANDN U10576 ( .B(n8870), .A(n736), .Z(n8868) );
  XNOR U10577 ( .A(a[342]), .B(n8871), .Z(n736) );
  IV U10578 ( .A(n8869), .Z(n8871) );
  XNOR U10579 ( .A(b[342]), .B(n8869), .Z(n8870) );
  XOR U10580 ( .A(n8872), .B(n8873), .Z(n8869) );
  ANDN U10581 ( .B(n8874), .A(n737), .Z(n8872) );
  XNOR U10582 ( .A(a[341]), .B(n8875), .Z(n737) );
  IV U10583 ( .A(n8873), .Z(n8875) );
  XNOR U10584 ( .A(b[341]), .B(n8873), .Z(n8874) );
  XOR U10585 ( .A(n8876), .B(n8877), .Z(n8873) );
  ANDN U10586 ( .B(n8878), .A(n738), .Z(n8876) );
  XNOR U10587 ( .A(a[340]), .B(n8879), .Z(n738) );
  IV U10588 ( .A(n8877), .Z(n8879) );
  XNOR U10589 ( .A(b[340]), .B(n8877), .Z(n8878) );
  XOR U10590 ( .A(n8880), .B(n8881), .Z(n8877) );
  ANDN U10591 ( .B(n8882), .A(n740), .Z(n8880) );
  XNOR U10592 ( .A(a[339]), .B(n8883), .Z(n740) );
  IV U10593 ( .A(n8881), .Z(n8883) );
  XNOR U10594 ( .A(b[339]), .B(n8881), .Z(n8882) );
  XOR U10595 ( .A(n8884), .B(n8885), .Z(n8881) );
  ANDN U10596 ( .B(n8886), .A(n741), .Z(n8884) );
  XNOR U10597 ( .A(a[338]), .B(n8887), .Z(n741) );
  IV U10598 ( .A(n8885), .Z(n8887) );
  XNOR U10599 ( .A(b[338]), .B(n8885), .Z(n8886) );
  XOR U10600 ( .A(n8888), .B(n8889), .Z(n8885) );
  ANDN U10601 ( .B(n8890), .A(n742), .Z(n8888) );
  XNOR U10602 ( .A(a[337]), .B(n8891), .Z(n742) );
  IV U10603 ( .A(n8889), .Z(n8891) );
  XNOR U10604 ( .A(b[337]), .B(n8889), .Z(n8890) );
  XOR U10605 ( .A(n8892), .B(n8893), .Z(n8889) );
  ANDN U10606 ( .B(n8894), .A(n743), .Z(n8892) );
  XNOR U10607 ( .A(a[336]), .B(n8895), .Z(n743) );
  IV U10608 ( .A(n8893), .Z(n8895) );
  XNOR U10609 ( .A(b[336]), .B(n8893), .Z(n8894) );
  XOR U10610 ( .A(n8896), .B(n8897), .Z(n8893) );
  ANDN U10611 ( .B(n8898), .A(n744), .Z(n8896) );
  XNOR U10612 ( .A(a[335]), .B(n8899), .Z(n744) );
  IV U10613 ( .A(n8897), .Z(n8899) );
  XNOR U10614 ( .A(b[335]), .B(n8897), .Z(n8898) );
  XOR U10615 ( .A(n8900), .B(n8901), .Z(n8897) );
  ANDN U10616 ( .B(n8902), .A(n745), .Z(n8900) );
  XNOR U10617 ( .A(a[334]), .B(n8903), .Z(n745) );
  IV U10618 ( .A(n8901), .Z(n8903) );
  XNOR U10619 ( .A(b[334]), .B(n8901), .Z(n8902) );
  XOR U10620 ( .A(n8904), .B(n8905), .Z(n8901) );
  ANDN U10621 ( .B(n8906), .A(n746), .Z(n8904) );
  XNOR U10622 ( .A(a[333]), .B(n8907), .Z(n746) );
  IV U10623 ( .A(n8905), .Z(n8907) );
  XNOR U10624 ( .A(b[333]), .B(n8905), .Z(n8906) );
  XOR U10625 ( .A(n8908), .B(n8909), .Z(n8905) );
  ANDN U10626 ( .B(n8910), .A(n747), .Z(n8908) );
  XNOR U10627 ( .A(a[332]), .B(n8911), .Z(n747) );
  IV U10628 ( .A(n8909), .Z(n8911) );
  XNOR U10629 ( .A(b[332]), .B(n8909), .Z(n8910) );
  XOR U10630 ( .A(n8912), .B(n8913), .Z(n8909) );
  ANDN U10631 ( .B(n8914), .A(n748), .Z(n8912) );
  XNOR U10632 ( .A(a[331]), .B(n8915), .Z(n748) );
  IV U10633 ( .A(n8913), .Z(n8915) );
  XNOR U10634 ( .A(b[331]), .B(n8913), .Z(n8914) );
  XOR U10635 ( .A(n8916), .B(n8917), .Z(n8913) );
  ANDN U10636 ( .B(n8918), .A(n749), .Z(n8916) );
  XNOR U10637 ( .A(a[330]), .B(n8919), .Z(n749) );
  IV U10638 ( .A(n8917), .Z(n8919) );
  XNOR U10639 ( .A(b[330]), .B(n8917), .Z(n8918) );
  XOR U10640 ( .A(n8920), .B(n8921), .Z(n8917) );
  ANDN U10641 ( .B(n8922), .A(n751), .Z(n8920) );
  XNOR U10642 ( .A(a[329]), .B(n8923), .Z(n751) );
  IV U10643 ( .A(n8921), .Z(n8923) );
  XNOR U10644 ( .A(b[329]), .B(n8921), .Z(n8922) );
  XOR U10645 ( .A(n8924), .B(n8925), .Z(n8921) );
  ANDN U10646 ( .B(n8926), .A(n752), .Z(n8924) );
  XNOR U10647 ( .A(a[328]), .B(n8927), .Z(n752) );
  IV U10648 ( .A(n8925), .Z(n8927) );
  XNOR U10649 ( .A(b[328]), .B(n8925), .Z(n8926) );
  XOR U10650 ( .A(n8928), .B(n8929), .Z(n8925) );
  ANDN U10651 ( .B(n8930), .A(n753), .Z(n8928) );
  XNOR U10652 ( .A(a[327]), .B(n8931), .Z(n753) );
  IV U10653 ( .A(n8929), .Z(n8931) );
  XNOR U10654 ( .A(b[327]), .B(n8929), .Z(n8930) );
  XOR U10655 ( .A(n8932), .B(n8933), .Z(n8929) );
  ANDN U10656 ( .B(n8934), .A(n754), .Z(n8932) );
  XNOR U10657 ( .A(a[326]), .B(n8935), .Z(n754) );
  IV U10658 ( .A(n8933), .Z(n8935) );
  XNOR U10659 ( .A(b[326]), .B(n8933), .Z(n8934) );
  XOR U10660 ( .A(n8936), .B(n8937), .Z(n8933) );
  ANDN U10661 ( .B(n8938), .A(n755), .Z(n8936) );
  XNOR U10662 ( .A(a[325]), .B(n8939), .Z(n755) );
  IV U10663 ( .A(n8937), .Z(n8939) );
  XNOR U10664 ( .A(b[325]), .B(n8937), .Z(n8938) );
  XOR U10665 ( .A(n8940), .B(n8941), .Z(n8937) );
  ANDN U10666 ( .B(n8942), .A(n756), .Z(n8940) );
  XNOR U10667 ( .A(a[324]), .B(n8943), .Z(n756) );
  IV U10668 ( .A(n8941), .Z(n8943) );
  XNOR U10669 ( .A(b[324]), .B(n8941), .Z(n8942) );
  XOR U10670 ( .A(n8944), .B(n8945), .Z(n8941) );
  ANDN U10671 ( .B(n8946), .A(n757), .Z(n8944) );
  XNOR U10672 ( .A(a[323]), .B(n8947), .Z(n757) );
  IV U10673 ( .A(n8945), .Z(n8947) );
  XNOR U10674 ( .A(b[323]), .B(n8945), .Z(n8946) );
  XOR U10675 ( .A(n8948), .B(n8949), .Z(n8945) );
  ANDN U10676 ( .B(n8950), .A(n758), .Z(n8948) );
  XNOR U10677 ( .A(a[322]), .B(n8951), .Z(n758) );
  IV U10678 ( .A(n8949), .Z(n8951) );
  XNOR U10679 ( .A(b[322]), .B(n8949), .Z(n8950) );
  XOR U10680 ( .A(n8952), .B(n8953), .Z(n8949) );
  ANDN U10681 ( .B(n8954), .A(n759), .Z(n8952) );
  XNOR U10682 ( .A(a[321]), .B(n8955), .Z(n759) );
  IV U10683 ( .A(n8953), .Z(n8955) );
  XNOR U10684 ( .A(b[321]), .B(n8953), .Z(n8954) );
  XOR U10685 ( .A(n8956), .B(n8957), .Z(n8953) );
  ANDN U10686 ( .B(n8958), .A(n760), .Z(n8956) );
  XNOR U10687 ( .A(a[320]), .B(n8959), .Z(n760) );
  IV U10688 ( .A(n8957), .Z(n8959) );
  XNOR U10689 ( .A(b[320]), .B(n8957), .Z(n8958) );
  XOR U10690 ( .A(n8960), .B(n8961), .Z(n8957) );
  ANDN U10691 ( .B(n8962), .A(n762), .Z(n8960) );
  XNOR U10692 ( .A(a[319]), .B(n8963), .Z(n762) );
  IV U10693 ( .A(n8961), .Z(n8963) );
  XNOR U10694 ( .A(b[319]), .B(n8961), .Z(n8962) );
  XOR U10695 ( .A(n8964), .B(n8965), .Z(n8961) );
  ANDN U10696 ( .B(n8966), .A(n763), .Z(n8964) );
  XNOR U10697 ( .A(a[318]), .B(n8967), .Z(n763) );
  IV U10698 ( .A(n8965), .Z(n8967) );
  XNOR U10699 ( .A(b[318]), .B(n8965), .Z(n8966) );
  XOR U10700 ( .A(n8968), .B(n8969), .Z(n8965) );
  ANDN U10701 ( .B(n8970), .A(n764), .Z(n8968) );
  XNOR U10702 ( .A(a[317]), .B(n8971), .Z(n764) );
  IV U10703 ( .A(n8969), .Z(n8971) );
  XNOR U10704 ( .A(b[317]), .B(n8969), .Z(n8970) );
  XOR U10705 ( .A(n8972), .B(n8973), .Z(n8969) );
  ANDN U10706 ( .B(n8974), .A(n765), .Z(n8972) );
  XNOR U10707 ( .A(a[316]), .B(n8975), .Z(n765) );
  IV U10708 ( .A(n8973), .Z(n8975) );
  XNOR U10709 ( .A(b[316]), .B(n8973), .Z(n8974) );
  XOR U10710 ( .A(n8976), .B(n8977), .Z(n8973) );
  ANDN U10711 ( .B(n8978), .A(n766), .Z(n8976) );
  XNOR U10712 ( .A(a[315]), .B(n8979), .Z(n766) );
  IV U10713 ( .A(n8977), .Z(n8979) );
  XNOR U10714 ( .A(b[315]), .B(n8977), .Z(n8978) );
  XOR U10715 ( .A(n8980), .B(n8981), .Z(n8977) );
  ANDN U10716 ( .B(n8982), .A(n767), .Z(n8980) );
  XNOR U10717 ( .A(a[314]), .B(n8983), .Z(n767) );
  IV U10718 ( .A(n8981), .Z(n8983) );
  XNOR U10719 ( .A(b[314]), .B(n8981), .Z(n8982) );
  XOR U10720 ( .A(n8984), .B(n8985), .Z(n8981) );
  ANDN U10721 ( .B(n8986), .A(n768), .Z(n8984) );
  XNOR U10722 ( .A(a[313]), .B(n8987), .Z(n768) );
  IV U10723 ( .A(n8985), .Z(n8987) );
  XNOR U10724 ( .A(b[313]), .B(n8985), .Z(n8986) );
  XOR U10725 ( .A(n8988), .B(n8989), .Z(n8985) );
  ANDN U10726 ( .B(n8990), .A(n769), .Z(n8988) );
  XNOR U10727 ( .A(a[312]), .B(n8991), .Z(n769) );
  IV U10728 ( .A(n8989), .Z(n8991) );
  XNOR U10729 ( .A(b[312]), .B(n8989), .Z(n8990) );
  XOR U10730 ( .A(n8992), .B(n8993), .Z(n8989) );
  ANDN U10731 ( .B(n8994), .A(n770), .Z(n8992) );
  XNOR U10732 ( .A(a[311]), .B(n8995), .Z(n770) );
  IV U10733 ( .A(n8993), .Z(n8995) );
  XNOR U10734 ( .A(b[311]), .B(n8993), .Z(n8994) );
  XOR U10735 ( .A(n8996), .B(n8997), .Z(n8993) );
  ANDN U10736 ( .B(n8998), .A(n771), .Z(n8996) );
  XNOR U10737 ( .A(a[310]), .B(n8999), .Z(n771) );
  IV U10738 ( .A(n8997), .Z(n8999) );
  XNOR U10739 ( .A(b[310]), .B(n8997), .Z(n8998) );
  XOR U10740 ( .A(n9000), .B(n9001), .Z(n8997) );
  ANDN U10741 ( .B(n9002), .A(n773), .Z(n9000) );
  XNOR U10742 ( .A(a[309]), .B(n9003), .Z(n773) );
  IV U10743 ( .A(n9001), .Z(n9003) );
  XNOR U10744 ( .A(b[309]), .B(n9001), .Z(n9002) );
  XOR U10745 ( .A(n9004), .B(n9005), .Z(n9001) );
  ANDN U10746 ( .B(n9006), .A(n774), .Z(n9004) );
  XNOR U10747 ( .A(a[308]), .B(n9007), .Z(n774) );
  IV U10748 ( .A(n9005), .Z(n9007) );
  XNOR U10749 ( .A(b[308]), .B(n9005), .Z(n9006) );
  XOR U10750 ( .A(n9008), .B(n9009), .Z(n9005) );
  ANDN U10751 ( .B(n9010), .A(n775), .Z(n9008) );
  XNOR U10752 ( .A(a[307]), .B(n9011), .Z(n775) );
  IV U10753 ( .A(n9009), .Z(n9011) );
  XNOR U10754 ( .A(b[307]), .B(n9009), .Z(n9010) );
  XOR U10755 ( .A(n9012), .B(n9013), .Z(n9009) );
  ANDN U10756 ( .B(n9014), .A(n776), .Z(n9012) );
  XNOR U10757 ( .A(a[306]), .B(n9015), .Z(n776) );
  IV U10758 ( .A(n9013), .Z(n9015) );
  XNOR U10759 ( .A(b[306]), .B(n9013), .Z(n9014) );
  XOR U10760 ( .A(n9016), .B(n9017), .Z(n9013) );
  ANDN U10761 ( .B(n9018), .A(n777), .Z(n9016) );
  XNOR U10762 ( .A(a[305]), .B(n9019), .Z(n777) );
  IV U10763 ( .A(n9017), .Z(n9019) );
  XNOR U10764 ( .A(b[305]), .B(n9017), .Z(n9018) );
  XOR U10765 ( .A(n9020), .B(n9021), .Z(n9017) );
  ANDN U10766 ( .B(n9022), .A(n778), .Z(n9020) );
  XNOR U10767 ( .A(a[304]), .B(n9023), .Z(n778) );
  IV U10768 ( .A(n9021), .Z(n9023) );
  XNOR U10769 ( .A(b[304]), .B(n9021), .Z(n9022) );
  XOR U10770 ( .A(n9024), .B(n9025), .Z(n9021) );
  ANDN U10771 ( .B(n9026), .A(n779), .Z(n9024) );
  XNOR U10772 ( .A(a[303]), .B(n9027), .Z(n779) );
  IV U10773 ( .A(n9025), .Z(n9027) );
  XNOR U10774 ( .A(b[303]), .B(n9025), .Z(n9026) );
  XOR U10775 ( .A(n9028), .B(n9029), .Z(n9025) );
  ANDN U10776 ( .B(n9030), .A(n780), .Z(n9028) );
  XNOR U10777 ( .A(a[302]), .B(n9031), .Z(n780) );
  IV U10778 ( .A(n9029), .Z(n9031) );
  XNOR U10779 ( .A(b[302]), .B(n9029), .Z(n9030) );
  XOR U10780 ( .A(n9032), .B(n9033), .Z(n9029) );
  ANDN U10781 ( .B(n9034), .A(n781), .Z(n9032) );
  XNOR U10782 ( .A(a[301]), .B(n9035), .Z(n781) );
  IV U10783 ( .A(n9033), .Z(n9035) );
  XNOR U10784 ( .A(b[301]), .B(n9033), .Z(n9034) );
  XOR U10785 ( .A(n9036), .B(n9037), .Z(n9033) );
  ANDN U10786 ( .B(n9038), .A(n782), .Z(n9036) );
  XNOR U10787 ( .A(a[300]), .B(n9039), .Z(n782) );
  IV U10788 ( .A(n9037), .Z(n9039) );
  XNOR U10789 ( .A(b[300]), .B(n9037), .Z(n9038) );
  XOR U10790 ( .A(n9040), .B(n9041), .Z(n9037) );
  ANDN U10791 ( .B(n9042), .A(n785), .Z(n9040) );
  XNOR U10792 ( .A(a[299]), .B(n9043), .Z(n785) );
  IV U10793 ( .A(n9041), .Z(n9043) );
  XNOR U10794 ( .A(b[299]), .B(n9041), .Z(n9042) );
  XOR U10795 ( .A(n9044), .B(n9045), .Z(n9041) );
  ANDN U10796 ( .B(n9046), .A(n786), .Z(n9044) );
  XNOR U10797 ( .A(a[298]), .B(n9047), .Z(n786) );
  IV U10798 ( .A(n9045), .Z(n9047) );
  XNOR U10799 ( .A(b[298]), .B(n9045), .Z(n9046) );
  XOR U10800 ( .A(n9048), .B(n9049), .Z(n9045) );
  ANDN U10801 ( .B(n9050), .A(n787), .Z(n9048) );
  XNOR U10802 ( .A(a[297]), .B(n9051), .Z(n787) );
  IV U10803 ( .A(n9049), .Z(n9051) );
  XNOR U10804 ( .A(b[297]), .B(n9049), .Z(n9050) );
  XOR U10805 ( .A(n9052), .B(n9053), .Z(n9049) );
  ANDN U10806 ( .B(n9054), .A(n788), .Z(n9052) );
  XNOR U10807 ( .A(a[296]), .B(n9055), .Z(n788) );
  IV U10808 ( .A(n9053), .Z(n9055) );
  XNOR U10809 ( .A(b[296]), .B(n9053), .Z(n9054) );
  XOR U10810 ( .A(n9056), .B(n9057), .Z(n9053) );
  ANDN U10811 ( .B(n9058), .A(n789), .Z(n9056) );
  XNOR U10812 ( .A(a[295]), .B(n9059), .Z(n789) );
  IV U10813 ( .A(n9057), .Z(n9059) );
  XNOR U10814 ( .A(b[295]), .B(n9057), .Z(n9058) );
  XOR U10815 ( .A(n9060), .B(n9061), .Z(n9057) );
  ANDN U10816 ( .B(n9062), .A(n790), .Z(n9060) );
  XNOR U10817 ( .A(a[294]), .B(n9063), .Z(n790) );
  IV U10818 ( .A(n9061), .Z(n9063) );
  XNOR U10819 ( .A(b[294]), .B(n9061), .Z(n9062) );
  XOR U10820 ( .A(n9064), .B(n9065), .Z(n9061) );
  ANDN U10821 ( .B(n9066), .A(n791), .Z(n9064) );
  XNOR U10822 ( .A(a[293]), .B(n9067), .Z(n791) );
  IV U10823 ( .A(n9065), .Z(n9067) );
  XNOR U10824 ( .A(b[293]), .B(n9065), .Z(n9066) );
  XOR U10825 ( .A(n9068), .B(n9069), .Z(n9065) );
  ANDN U10826 ( .B(n9070), .A(n792), .Z(n9068) );
  XNOR U10827 ( .A(a[292]), .B(n9071), .Z(n792) );
  IV U10828 ( .A(n9069), .Z(n9071) );
  XNOR U10829 ( .A(b[292]), .B(n9069), .Z(n9070) );
  XOR U10830 ( .A(n9072), .B(n9073), .Z(n9069) );
  ANDN U10831 ( .B(n9074), .A(n793), .Z(n9072) );
  XNOR U10832 ( .A(a[291]), .B(n9075), .Z(n793) );
  IV U10833 ( .A(n9073), .Z(n9075) );
  XNOR U10834 ( .A(b[291]), .B(n9073), .Z(n9074) );
  XOR U10835 ( .A(n9076), .B(n9077), .Z(n9073) );
  ANDN U10836 ( .B(n9078), .A(n794), .Z(n9076) );
  XNOR U10837 ( .A(a[290]), .B(n9079), .Z(n794) );
  IV U10838 ( .A(n9077), .Z(n9079) );
  XNOR U10839 ( .A(b[290]), .B(n9077), .Z(n9078) );
  XOR U10840 ( .A(n9080), .B(n9081), .Z(n9077) );
  ANDN U10841 ( .B(n9082), .A(n796), .Z(n9080) );
  XNOR U10842 ( .A(a[289]), .B(n9083), .Z(n796) );
  IV U10843 ( .A(n9081), .Z(n9083) );
  XNOR U10844 ( .A(b[289]), .B(n9081), .Z(n9082) );
  XOR U10845 ( .A(n9084), .B(n9085), .Z(n9081) );
  ANDN U10846 ( .B(n9086), .A(n797), .Z(n9084) );
  XNOR U10847 ( .A(a[288]), .B(n9087), .Z(n797) );
  IV U10848 ( .A(n9085), .Z(n9087) );
  XNOR U10849 ( .A(b[288]), .B(n9085), .Z(n9086) );
  XOR U10850 ( .A(n9088), .B(n9089), .Z(n9085) );
  ANDN U10851 ( .B(n9090), .A(n798), .Z(n9088) );
  XNOR U10852 ( .A(a[287]), .B(n9091), .Z(n798) );
  IV U10853 ( .A(n9089), .Z(n9091) );
  XNOR U10854 ( .A(b[287]), .B(n9089), .Z(n9090) );
  XOR U10855 ( .A(n9092), .B(n9093), .Z(n9089) );
  ANDN U10856 ( .B(n9094), .A(n799), .Z(n9092) );
  XNOR U10857 ( .A(a[286]), .B(n9095), .Z(n799) );
  IV U10858 ( .A(n9093), .Z(n9095) );
  XNOR U10859 ( .A(b[286]), .B(n9093), .Z(n9094) );
  XOR U10860 ( .A(n9096), .B(n9097), .Z(n9093) );
  ANDN U10861 ( .B(n9098), .A(n800), .Z(n9096) );
  XNOR U10862 ( .A(a[285]), .B(n9099), .Z(n800) );
  IV U10863 ( .A(n9097), .Z(n9099) );
  XNOR U10864 ( .A(b[285]), .B(n9097), .Z(n9098) );
  XOR U10865 ( .A(n9100), .B(n9101), .Z(n9097) );
  ANDN U10866 ( .B(n9102), .A(n801), .Z(n9100) );
  XNOR U10867 ( .A(a[284]), .B(n9103), .Z(n801) );
  IV U10868 ( .A(n9101), .Z(n9103) );
  XNOR U10869 ( .A(b[284]), .B(n9101), .Z(n9102) );
  XOR U10870 ( .A(n9104), .B(n9105), .Z(n9101) );
  ANDN U10871 ( .B(n9106), .A(n802), .Z(n9104) );
  XNOR U10872 ( .A(a[283]), .B(n9107), .Z(n802) );
  IV U10873 ( .A(n9105), .Z(n9107) );
  XNOR U10874 ( .A(b[283]), .B(n9105), .Z(n9106) );
  XOR U10875 ( .A(n9108), .B(n9109), .Z(n9105) );
  ANDN U10876 ( .B(n9110), .A(n803), .Z(n9108) );
  XNOR U10877 ( .A(a[282]), .B(n9111), .Z(n803) );
  IV U10878 ( .A(n9109), .Z(n9111) );
  XNOR U10879 ( .A(b[282]), .B(n9109), .Z(n9110) );
  XOR U10880 ( .A(n9112), .B(n9113), .Z(n9109) );
  ANDN U10881 ( .B(n9114), .A(n804), .Z(n9112) );
  XNOR U10882 ( .A(a[281]), .B(n9115), .Z(n804) );
  IV U10883 ( .A(n9113), .Z(n9115) );
  XNOR U10884 ( .A(b[281]), .B(n9113), .Z(n9114) );
  XOR U10885 ( .A(n9116), .B(n9117), .Z(n9113) );
  ANDN U10886 ( .B(n9118), .A(n805), .Z(n9116) );
  XNOR U10887 ( .A(a[280]), .B(n9119), .Z(n805) );
  IV U10888 ( .A(n9117), .Z(n9119) );
  XNOR U10889 ( .A(b[280]), .B(n9117), .Z(n9118) );
  XOR U10890 ( .A(n9120), .B(n9121), .Z(n9117) );
  ANDN U10891 ( .B(n9122), .A(n807), .Z(n9120) );
  XNOR U10892 ( .A(a[279]), .B(n9123), .Z(n807) );
  IV U10893 ( .A(n9121), .Z(n9123) );
  XNOR U10894 ( .A(b[279]), .B(n9121), .Z(n9122) );
  XOR U10895 ( .A(n9124), .B(n9125), .Z(n9121) );
  ANDN U10896 ( .B(n9126), .A(n808), .Z(n9124) );
  XNOR U10897 ( .A(a[278]), .B(n9127), .Z(n808) );
  IV U10898 ( .A(n9125), .Z(n9127) );
  XNOR U10899 ( .A(b[278]), .B(n9125), .Z(n9126) );
  XOR U10900 ( .A(n9128), .B(n9129), .Z(n9125) );
  ANDN U10901 ( .B(n9130), .A(n809), .Z(n9128) );
  XNOR U10902 ( .A(a[277]), .B(n9131), .Z(n809) );
  IV U10903 ( .A(n9129), .Z(n9131) );
  XNOR U10904 ( .A(b[277]), .B(n9129), .Z(n9130) );
  XOR U10905 ( .A(n9132), .B(n9133), .Z(n9129) );
  ANDN U10906 ( .B(n9134), .A(n810), .Z(n9132) );
  XNOR U10907 ( .A(a[276]), .B(n9135), .Z(n810) );
  IV U10908 ( .A(n9133), .Z(n9135) );
  XNOR U10909 ( .A(b[276]), .B(n9133), .Z(n9134) );
  XOR U10910 ( .A(n9136), .B(n9137), .Z(n9133) );
  ANDN U10911 ( .B(n9138), .A(n811), .Z(n9136) );
  XNOR U10912 ( .A(a[275]), .B(n9139), .Z(n811) );
  IV U10913 ( .A(n9137), .Z(n9139) );
  XNOR U10914 ( .A(b[275]), .B(n9137), .Z(n9138) );
  XOR U10915 ( .A(n9140), .B(n9141), .Z(n9137) );
  ANDN U10916 ( .B(n9142), .A(n812), .Z(n9140) );
  XNOR U10917 ( .A(a[274]), .B(n9143), .Z(n812) );
  IV U10918 ( .A(n9141), .Z(n9143) );
  XNOR U10919 ( .A(b[274]), .B(n9141), .Z(n9142) );
  XOR U10920 ( .A(n9144), .B(n9145), .Z(n9141) );
  ANDN U10921 ( .B(n9146), .A(n813), .Z(n9144) );
  XNOR U10922 ( .A(a[273]), .B(n9147), .Z(n813) );
  IV U10923 ( .A(n9145), .Z(n9147) );
  XNOR U10924 ( .A(b[273]), .B(n9145), .Z(n9146) );
  XOR U10925 ( .A(n9148), .B(n9149), .Z(n9145) );
  ANDN U10926 ( .B(n9150), .A(n814), .Z(n9148) );
  XNOR U10927 ( .A(a[272]), .B(n9151), .Z(n814) );
  IV U10928 ( .A(n9149), .Z(n9151) );
  XNOR U10929 ( .A(b[272]), .B(n9149), .Z(n9150) );
  XOR U10930 ( .A(n9152), .B(n9153), .Z(n9149) );
  ANDN U10931 ( .B(n9154), .A(n815), .Z(n9152) );
  XNOR U10932 ( .A(a[271]), .B(n9155), .Z(n815) );
  IV U10933 ( .A(n9153), .Z(n9155) );
  XNOR U10934 ( .A(b[271]), .B(n9153), .Z(n9154) );
  XOR U10935 ( .A(n9156), .B(n9157), .Z(n9153) );
  ANDN U10936 ( .B(n9158), .A(n816), .Z(n9156) );
  XNOR U10937 ( .A(a[270]), .B(n9159), .Z(n816) );
  IV U10938 ( .A(n9157), .Z(n9159) );
  XNOR U10939 ( .A(b[270]), .B(n9157), .Z(n9158) );
  XOR U10940 ( .A(n9160), .B(n9161), .Z(n9157) );
  ANDN U10941 ( .B(n9162), .A(n818), .Z(n9160) );
  XNOR U10942 ( .A(a[269]), .B(n9163), .Z(n818) );
  IV U10943 ( .A(n9161), .Z(n9163) );
  XNOR U10944 ( .A(b[269]), .B(n9161), .Z(n9162) );
  XOR U10945 ( .A(n9164), .B(n9165), .Z(n9161) );
  ANDN U10946 ( .B(n9166), .A(n819), .Z(n9164) );
  XNOR U10947 ( .A(a[268]), .B(n9167), .Z(n819) );
  IV U10948 ( .A(n9165), .Z(n9167) );
  XNOR U10949 ( .A(b[268]), .B(n9165), .Z(n9166) );
  XOR U10950 ( .A(n9168), .B(n9169), .Z(n9165) );
  ANDN U10951 ( .B(n9170), .A(n820), .Z(n9168) );
  XNOR U10952 ( .A(a[267]), .B(n9171), .Z(n820) );
  IV U10953 ( .A(n9169), .Z(n9171) );
  XNOR U10954 ( .A(b[267]), .B(n9169), .Z(n9170) );
  XOR U10955 ( .A(n9172), .B(n9173), .Z(n9169) );
  ANDN U10956 ( .B(n9174), .A(n821), .Z(n9172) );
  XNOR U10957 ( .A(a[266]), .B(n9175), .Z(n821) );
  IV U10958 ( .A(n9173), .Z(n9175) );
  XNOR U10959 ( .A(b[266]), .B(n9173), .Z(n9174) );
  XOR U10960 ( .A(n9176), .B(n9177), .Z(n9173) );
  ANDN U10961 ( .B(n9178), .A(n822), .Z(n9176) );
  XNOR U10962 ( .A(a[265]), .B(n9179), .Z(n822) );
  IV U10963 ( .A(n9177), .Z(n9179) );
  XNOR U10964 ( .A(b[265]), .B(n9177), .Z(n9178) );
  XOR U10965 ( .A(n9180), .B(n9181), .Z(n9177) );
  ANDN U10966 ( .B(n9182), .A(n823), .Z(n9180) );
  XNOR U10967 ( .A(a[264]), .B(n9183), .Z(n823) );
  IV U10968 ( .A(n9181), .Z(n9183) );
  XNOR U10969 ( .A(b[264]), .B(n9181), .Z(n9182) );
  XOR U10970 ( .A(n9184), .B(n9185), .Z(n9181) );
  ANDN U10971 ( .B(n9186), .A(n824), .Z(n9184) );
  XNOR U10972 ( .A(a[263]), .B(n9187), .Z(n824) );
  IV U10973 ( .A(n9185), .Z(n9187) );
  XNOR U10974 ( .A(b[263]), .B(n9185), .Z(n9186) );
  XOR U10975 ( .A(n9188), .B(n9189), .Z(n9185) );
  ANDN U10976 ( .B(n9190), .A(n825), .Z(n9188) );
  XNOR U10977 ( .A(a[262]), .B(n9191), .Z(n825) );
  IV U10978 ( .A(n9189), .Z(n9191) );
  XNOR U10979 ( .A(b[262]), .B(n9189), .Z(n9190) );
  XOR U10980 ( .A(n9192), .B(n9193), .Z(n9189) );
  ANDN U10981 ( .B(n9194), .A(n826), .Z(n9192) );
  XNOR U10982 ( .A(a[261]), .B(n9195), .Z(n826) );
  IV U10983 ( .A(n9193), .Z(n9195) );
  XNOR U10984 ( .A(b[261]), .B(n9193), .Z(n9194) );
  XOR U10985 ( .A(n9196), .B(n9197), .Z(n9193) );
  ANDN U10986 ( .B(n9198), .A(n827), .Z(n9196) );
  XNOR U10987 ( .A(a[260]), .B(n9199), .Z(n827) );
  IV U10988 ( .A(n9197), .Z(n9199) );
  XNOR U10989 ( .A(b[260]), .B(n9197), .Z(n9198) );
  XOR U10990 ( .A(n9200), .B(n9201), .Z(n9197) );
  ANDN U10991 ( .B(n9202), .A(n829), .Z(n9200) );
  XNOR U10992 ( .A(a[259]), .B(n9203), .Z(n829) );
  IV U10993 ( .A(n9201), .Z(n9203) );
  XNOR U10994 ( .A(b[259]), .B(n9201), .Z(n9202) );
  XOR U10995 ( .A(n9204), .B(n9205), .Z(n9201) );
  ANDN U10996 ( .B(n9206), .A(n830), .Z(n9204) );
  XNOR U10997 ( .A(a[258]), .B(n9207), .Z(n830) );
  IV U10998 ( .A(n9205), .Z(n9207) );
  XNOR U10999 ( .A(b[258]), .B(n9205), .Z(n9206) );
  XOR U11000 ( .A(n9208), .B(n9209), .Z(n9205) );
  ANDN U11001 ( .B(n9210), .A(n831), .Z(n9208) );
  XNOR U11002 ( .A(a[257]), .B(n9211), .Z(n831) );
  IV U11003 ( .A(n9209), .Z(n9211) );
  XNOR U11004 ( .A(b[257]), .B(n9209), .Z(n9210) );
  XOR U11005 ( .A(n9212), .B(n9213), .Z(n9209) );
  ANDN U11006 ( .B(n9214), .A(n832), .Z(n9212) );
  XNOR U11007 ( .A(a[256]), .B(n9215), .Z(n832) );
  IV U11008 ( .A(n9213), .Z(n9215) );
  XNOR U11009 ( .A(b[256]), .B(n9213), .Z(n9214) );
  XOR U11010 ( .A(n9216), .B(n9217), .Z(n9213) );
  ANDN U11011 ( .B(n9218), .A(n833), .Z(n9216) );
  XNOR U11012 ( .A(a[255]), .B(n9219), .Z(n833) );
  IV U11013 ( .A(n9217), .Z(n9219) );
  XNOR U11014 ( .A(b[255]), .B(n9217), .Z(n9218) );
  XOR U11015 ( .A(n9220), .B(n9221), .Z(n9217) );
  ANDN U11016 ( .B(n9222), .A(n834), .Z(n9220) );
  XNOR U11017 ( .A(a[254]), .B(n9223), .Z(n834) );
  IV U11018 ( .A(n9221), .Z(n9223) );
  XNOR U11019 ( .A(b[254]), .B(n9221), .Z(n9222) );
  XOR U11020 ( .A(n9224), .B(n9225), .Z(n9221) );
  ANDN U11021 ( .B(n9226), .A(n835), .Z(n9224) );
  XNOR U11022 ( .A(a[253]), .B(n9227), .Z(n835) );
  IV U11023 ( .A(n9225), .Z(n9227) );
  XNOR U11024 ( .A(b[253]), .B(n9225), .Z(n9226) );
  XOR U11025 ( .A(n9228), .B(n9229), .Z(n9225) );
  ANDN U11026 ( .B(n9230), .A(n836), .Z(n9228) );
  XNOR U11027 ( .A(a[252]), .B(n9231), .Z(n836) );
  IV U11028 ( .A(n9229), .Z(n9231) );
  XNOR U11029 ( .A(b[252]), .B(n9229), .Z(n9230) );
  XOR U11030 ( .A(n9232), .B(n9233), .Z(n9229) );
  ANDN U11031 ( .B(n9234), .A(n837), .Z(n9232) );
  XNOR U11032 ( .A(a[251]), .B(n9235), .Z(n837) );
  IV U11033 ( .A(n9233), .Z(n9235) );
  XNOR U11034 ( .A(b[251]), .B(n9233), .Z(n9234) );
  XOR U11035 ( .A(n9236), .B(n9237), .Z(n9233) );
  ANDN U11036 ( .B(n9238), .A(n838), .Z(n9236) );
  XNOR U11037 ( .A(a[250]), .B(n9239), .Z(n838) );
  IV U11038 ( .A(n9237), .Z(n9239) );
  XNOR U11039 ( .A(b[250]), .B(n9237), .Z(n9238) );
  XOR U11040 ( .A(n9240), .B(n9241), .Z(n9237) );
  ANDN U11041 ( .B(n9242), .A(n840), .Z(n9240) );
  XNOR U11042 ( .A(a[249]), .B(n9243), .Z(n840) );
  IV U11043 ( .A(n9241), .Z(n9243) );
  XNOR U11044 ( .A(b[249]), .B(n9241), .Z(n9242) );
  XOR U11045 ( .A(n9244), .B(n9245), .Z(n9241) );
  ANDN U11046 ( .B(n9246), .A(n841), .Z(n9244) );
  XNOR U11047 ( .A(a[248]), .B(n9247), .Z(n841) );
  IV U11048 ( .A(n9245), .Z(n9247) );
  XNOR U11049 ( .A(b[248]), .B(n9245), .Z(n9246) );
  XOR U11050 ( .A(n9248), .B(n9249), .Z(n9245) );
  ANDN U11051 ( .B(n9250), .A(n842), .Z(n9248) );
  XNOR U11052 ( .A(a[247]), .B(n9251), .Z(n842) );
  IV U11053 ( .A(n9249), .Z(n9251) );
  XNOR U11054 ( .A(b[247]), .B(n9249), .Z(n9250) );
  XOR U11055 ( .A(n9252), .B(n9253), .Z(n9249) );
  ANDN U11056 ( .B(n9254), .A(n843), .Z(n9252) );
  XNOR U11057 ( .A(a[246]), .B(n9255), .Z(n843) );
  IV U11058 ( .A(n9253), .Z(n9255) );
  XNOR U11059 ( .A(b[246]), .B(n9253), .Z(n9254) );
  XOR U11060 ( .A(n9256), .B(n9257), .Z(n9253) );
  ANDN U11061 ( .B(n9258), .A(n844), .Z(n9256) );
  XNOR U11062 ( .A(a[245]), .B(n9259), .Z(n844) );
  IV U11063 ( .A(n9257), .Z(n9259) );
  XNOR U11064 ( .A(b[245]), .B(n9257), .Z(n9258) );
  XOR U11065 ( .A(n9260), .B(n9261), .Z(n9257) );
  ANDN U11066 ( .B(n9262), .A(n845), .Z(n9260) );
  XNOR U11067 ( .A(a[244]), .B(n9263), .Z(n845) );
  IV U11068 ( .A(n9261), .Z(n9263) );
  XNOR U11069 ( .A(b[244]), .B(n9261), .Z(n9262) );
  XOR U11070 ( .A(n9264), .B(n9265), .Z(n9261) );
  ANDN U11071 ( .B(n9266), .A(n846), .Z(n9264) );
  XNOR U11072 ( .A(a[243]), .B(n9267), .Z(n846) );
  IV U11073 ( .A(n9265), .Z(n9267) );
  XNOR U11074 ( .A(b[243]), .B(n9265), .Z(n9266) );
  XOR U11075 ( .A(n9268), .B(n9269), .Z(n9265) );
  ANDN U11076 ( .B(n9270), .A(n847), .Z(n9268) );
  XNOR U11077 ( .A(a[242]), .B(n9271), .Z(n847) );
  IV U11078 ( .A(n9269), .Z(n9271) );
  XNOR U11079 ( .A(b[242]), .B(n9269), .Z(n9270) );
  XOR U11080 ( .A(n9272), .B(n9273), .Z(n9269) );
  ANDN U11081 ( .B(n9274), .A(n848), .Z(n9272) );
  XNOR U11082 ( .A(a[241]), .B(n9275), .Z(n848) );
  IV U11083 ( .A(n9273), .Z(n9275) );
  XNOR U11084 ( .A(b[241]), .B(n9273), .Z(n9274) );
  XOR U11085 ( .A(n9276), .B(n9277), .Z(n9273) );
  ANDN U11086 ( .B(n9278), .A(n849), .Z(n9276) );
  XNOR U11087 ( .A(a[240]), .B(n9279), .Z(n849) );
  IV U11088 ( .A(n9277), .Z(n9279) );
  XNOR U11089 ( .A(b[240]), .B(n9277), .Z(n9278) );
  XOR U11090 ( .A(n9280), .B(n9281), .Z(n9277) );
  ANDN U11091 ( .B(n9282), .A(n851), .Z(n9280) );
  XNOR U11092 ( .A(a[239]), .B(n9283), .Z(n851) );
  IV U11093 ( .A(n9281), .Z(n9283) );
  XNOR U11094 ( .A(b[239]), .B(n9281), .Z(n9282) );
  XOR U11095 ( .A(n9284), .B(n9285), .Z(n9281) );
  ANDN U11096 ( .B(n9286), .A(n852), .Z(n9284) );
  XNOR U11097 ( .A(a[238]), .B(n9287), .Z(n852) );
  IV U11098 ( .A(n9285), .Z(n9287) );
  XNOR U11099 ( .A(b[238]), .B(n9285), .Z(n9286) );
  XOR U11100 ( .A(n9288), .B(n9289), .Z(n9285) );
  ANDN U11101 ( .B(n9290), .A(n853), .Z(n9288) );
  XNOR U11102 ( .A(a[237]), .B(n9291), .Z(n853) );
  IV U11103 ( .A(n9289), .Z(n9291) );
  XNOR U11104 ( .A(b[237]), .B(n9289), .Z(n9290) );
  XOR U11105 ( .A(n9292), .B(n9293), .Z(n9289) );
  ANDN U11106 ( .B(n9294), .A(n854), .Z(n9292) );
  XNOR U11107 ( .A(a[236]), .B(n9295), .Z(n854) );
  IV U11108 ( .A(n9293), .Z(n9295) );
  XNOR U11109 ( .A(b[236]), .B(n9293), .Z(n9294) );
  XOR U11110 ( .A(n9296), .B(n9297), .Z(n9293) );
  ANDN U11111 ( .B(n9298), .A(n855), .Z(n9296) );
  XNOR U11112 ( .A(a[235]), .B(n9299), .Z(n855) );
  IV U11113 ( .A(n9297), .Z(n9299) );
  XNOR U11114 ( .A(b[235]), .B(n9297), .Z(n9298) );
  XOR U11115 ( .A(n9300), .B(n9301), .Z(n9297) );
  ANDN U11116 ( .B(n9302), .A(n856), .Z(n9300) );
  XNOR U11117 ( .A(a[234]), .B(n9303), .Z(n856) );
  IV U11118 ( .A(n9301), .Z(n9303) );
  XNOR U11119 ( .A(b[234]), .B(n9301), .Z(n9302) );
  XOR U11120 ( .A(n9304), .B(n9305), .Z(n9301) );
  ANDN U11121 ( .B(n9306), .A(n857), .Z(n9304) );
  XNOR U11122 ( .A(a[233]), .B(n9307), .Z(n857) );
  IV U11123 ( .A(n9305), .Z(n9307) );
  XNOR U11124 ( .A(b[233]), .B(n9305), .Z(n9306) );
  XOR U11125 ( .A(n9308), .B(n9309), .Z(n9305) );
  ANDN U11126 ( .B(n9310), .A(n858), .Z(n9308) );
  XNOR U11127 ( .A(a[232]), .B(n9311), .Z(n858) );
  IV U11128 ( .A(n9309), .Z(n9311) );
  XNOR U11129 ( .A(b[232]), .B(n9309), .Z(n9310) );
  XOR U11130 ( .A(n9312), .B(n9313), .Z(n9309) );
  ANDN U11131 ( .B(n9314), .A(n859), .Z(n9312) );
  XNOR U11132 ( .A(a[231]), .B(n9315), .Z(n859) );
  IV U11133 ( .A(n9313), .Z(n9315) );
  XNOR U11134 ( .A(b[231]), .B(n9313), .Z(n9314) );
  XOR U11135 ( .A(n9316), .B(n9317), .Z(n9313) );
  ANDN U11136 ( .B(n9318), .A(n860), .Z(n9316) );
  XNOR U11137 ( .A(a[230]), .B(n9319), .Z(n860) );
  IV U11138 ( .A(n9317), .Z(n9319) );
  XNOR U11139 ( .A(b[230]), .B(n9317), .Z(n9318) );
  XOR U11140 ( .A(n9320), .B(n9321), .Z(n9317) );
  ANDN U11141 ( .B(n9322), .A(n862), .Z(n9320) );
  XNOR U11142 ( .A(a[229]), .B(n9323), .Z(n862) );
  IV U11143 ( .A(n9321), .Z(n9323) );
  XNOR U11144 ( .A(b[229]), .B(n9321), .Z(n9322) );
  XOR U11145 ( .A(n9324), .B(n9325), .Z(n9321) );
  ANDN U11146 ( .B(n9326), .A(n863), .Z(n9324) );
  XNOR U11147 ( .A(a[228]), .B(n9327), .Z(n863) );
  IV U11148 ( .A(n9325), .Z(n9327) );
  XNOR U11149 ( .A(b[228]), .B(n9325), .Z(n9326) );
  XOR U11150 ( .A(n9328), .B(n9329), .Z(n9325) );
  ANDN U11151 ( .B(n9330), .A(n864), .Z(n9328) );
  XNOR U11152 ( .A(a[227]), .B(n9331), .Z(n864) );
  IV U11153 ( .A(n9329), .Z(n9331) );
  XNOR U11154 ( .A(b[227]), .B(n9329), .Z(n9330) );
  XOR U11155 ( .A(n9332), .B(n9333), .Z(n9329) );
  ANDN U11156 ( .B(n9334), .A(n865), .Z(n9332) );
  XNOR U11157 ( .A(a[226]), .B(n9335), .Z(n865) );
  IV U11158 ( .A(n9333), .Z(n9335) );
  XNOR U11159 ( .A(b[226]), .B(n9333), .Z(n9334) );
  XOR U11160 ( .A(n9336), .B(n9337), .Z(n9333) );
  ANDN U11161 ( .B(n9338), .A(n866), .Z(n9336) );
  XNOR U11162 ( .A(a[225]), .B(n9339), .Z(n866) );
  IV U11163 ( .A(n9337), .Z(n9339) );
  XNOR U11164 ( .A(b[225]), .B(n9337), .Z(n9338) );
  XOR U11165 ( .A(n9340), .B(n9341), .Z(n9337) );
  ANDN U11166 ( .B(n9342), .A(n867), .Z(n9340) );
  XNOR U11167 ( .A(a[224]), .B(n9343), .Z(n867) );
  IV U11168 ( .A(n9341), .Z(n9343) );
  XNOR U11169 ( .A(b[224]), .B(n9341), .Z(n9342) );
  XOR U11170 ( .A(n9344), .B(n9345), .Z(n9341) );
  ANDN U11171 ( .B(n9346), .A(n868), .Z(n9344) );
  XNOR U11172 ( .A(a[223]), .B(n9347), .Z(n868) );
  IV U11173 ( .A(n9345), .Z(n9347) );
  XNOR U11174 ( .A(b[223]), .B(n9345), .Z(n9346) );
  XOR U11175 ( .A(n9348), .B(n9349), .Z(n9345) );
  ANDN U11176 ( .B(n9350), .A(n869), .Z(n9348) );
  XNOR U11177 ( .A(a[222]), .B(n9351), .Z(n869) );
  IV U11178 ( .A(n9349), .Z(n9351) );
  XNOR U11179 ( .A(b[222]), .B(n9349), .Z(n9350) );
  XOR U11180 ( .A(n9352), .B(n9353), .Z(n9349) );
  ANDN U11181 ( .B(n9354), .A(n870), .Z(n9352) );
  XNOR U11182 ( .A(a[221]), .B(n9355), .Z(n870) );
  IV U11183 ( .A(n9353), .Z(n9355) );
  XNOR U11184 ( .A(b[221]), .B(n9353), .Z(n9354) );
  XOR U11185 ( .A(n9356), .B(n9357), .Z(n9353) );
  ANDN U11186 ( .B(n9358), .A(n871), .Z(n9356) );
  XNOR U11187 ( .A(a[220]), .B(n9359), .Z(n871) );
  IV U11188 ( .A(n9357), .Z(n9359) );
  XNOR U11189 ( .A(b[220]), .B(n9357), .Z(n9358) );
  XOR U11190 ( .A(n9360), .B(n9361), .Z(n9357) );
  ANDN U11191 ( .B(n9362), .A(n873), .Z(n9360) );
  XNOR U11192 ( .A(a[219]), .B(n9363), .Z(n873) );
  IV U11193 ( .A(n9361), .Z(n9363) );
  XNOR U11194 ( .A(b[219]), .B(n9361), .Z(n9362) );
  XOR U11195 ( .A(n9364), .B(n9365), .Z(n9361) );
  ANDN U11196 ( .B(n9366), .A(n874), .Z(n9364) );
  XNOR U11197 ( .A(a[218]), .B(n9367), .Z(n874) );
  IV U11198 ( .A(n9365), .Z(n9367) );
  XNOR U11199 ( .A(b[218]), .B(n9365), .Z(n9366) );
  XOR U11200 ( .A(n9368), .B(n9369), .Z(n9365) );
  ANDN U11201 ( .B(n9370), .A(n875), .Z(n9368) );
  XNOR U11202 ( .A(a[217]), .B(n9371), .Z(n875) );
  IV U11203 ( .A(n9369), .Z(n9371) );
  XNOR U11204 ( .A(b[217]), .B(n9369), .Z(n9370) );
  XOR U11205 ( .A(n9372), .B(n9373), .Z(n9369) );
  ANDN U11206 ( .B(n9374), .A(n876), .Z(n9372) );
  XNOR U11207 ( .A(a[216]), .B(n9375), .Z(n876) );
  IV U11208 ( .A(n9373), .Z(n9375) );
  XNOR U11209 ( .A(b[216]), .B(n9373), .Z(n9374) );
  XOR U11210 ( .A(n9376), .B(n9377), .Z(n9373) );
  ANDN U11211 ( .B(n9378), .A(n877), .Z(n9376) );
  XNOR U11212 ( .A(a[215]), .B(n9379), .Z(n877) );
  IV U11213 ( .A(n9377), .Z(n9379) );
  XNOR U11214 ( .A(b[215]), .B(n9377), .Z(n9378) );
  XOR U11215 ( .A(n9380), .B(n9381), .Z(n9377) );
  ANDN U11216 ( .B(n9382), .A(n878), .Z(n9380) );
  XNOR U11217 ( .A(a[214]), .B(n9383), .Z(n878) );
  IV U11218 ( .A(n9381), .Z(n9383) );
  XNOR U11219 ( .A(b[214]), .B(n9381), .Z(n9382) );
  XOR U11220 ( .A(n9384), .B(n9385), .Z(n9381) );
  ANDN U11221 ( .B(n9386), .A(n879), .Z(n9384) );
  XNOR U11222 ( .A(a[213]), .B(n9387), .Z(n879) );
  IV U11223 ( .A(n9385), .Z(n9387) );
  XNOR U11224 ( .A(b[213]), .B(n9385), .Z(n9386) );
  XOR U11225 ( .A(n9388), .B(n9389), .Z(n9385) );
  ANDN U11226 ( .B(n9390), .A(n880), .Z(n9388) );
  XNOR U11227 ( .A(a[212]), .B(n9391), .Z(n880) );
  IV U11228 ( .A(n9389), .Z(n9391) );
  XNOR U11229 ( .A(b[212]), .B(n9389), .Z(n9390) );
  XOR U11230 ( .A(n9392), .B(n9393), .Z(n9389) );
  ANDN U11231 ( .B(n9394), .A(n881), .Z(n9392) );
  XNOR U11232 ( .A(a[211]), .B(n9395), .Z(n881) );
  IV U11233 ( .A(n9393), .Z(n9395) );
  XNOR U11234 ( .A(b[211]), .B(n9393), .Z(n9394) );
  XOR U11235 ( .A(n9396), .B(n9397), .Z(n9393) );
  ANDN U11236 ( .B(n9398), .A(n882), .Z(n9396) );
  XNOR U11237 ( .A(a[210]), .B(n9399), .Z(n882) );
  IV U11238 ( .A(n9397), .Z(n9399) );
  XNOR U11239 ( .A(b[210]), .B(n9397), .Z(n9398) );
  XOR U11240 ( .A(n9400), .B(n9401), .Z(n9397) );
  ANDN U11241 ( .B(n9402), .A(n884), .Z(n9400) );
  XNOR U11242 ( .A(a[209]), .B(n9403), .Z(n884) );
  IV U11243 ( .A(n9401), .Z(n9403) );
  XNOR U11244 ( .A(b[209]), .B(n9401), .Z(n9402) );
  XOR U11245 ( .A(n9404), .B(n9405), .Z(n9401) );
  ANDN U11246 ( .B(n9406), .A(n885), .Z(n9404) );
  XNOR U11247 ( .A(a[208]), .B(n9407), .Z(n885) );
  IV U11248 ( .A(n9405), .Z(n9407) );
  XNOR U11249 ( .A(b[208]), .B(n9405), .Z(n9406) );
  XOR U11250 ( .A(n9408), .B(n9409), .Z(n9405) );
  ANDN U11251 ( .B(n9410), .A(n886), .Z(n9408) );
  XNOR U11252 ( .A(a[207]), .B(n9411), .Z(n886) );
  IV U11253 ( .A(n9409), .Z(n9411) );
  XNOR U11254 ( .A(b[207]), .B(n9409), .Z(n9410) );
  XOR U11255 ( .A(n9412), .B(n9413), .Z(n9409) );
  ANDN U11256 ( .B(n9414), .A(n887), .Z(n9412) );
  XNOR U11257 ( .A(a[206]), .B(n9415), .Z(n887) );
  IV U11258 ( .A(n9413), .Z(n9415) );
  XNOR U11259 ( .A(b[206]), .B(n9413), .Z(n9414) );
  XOR U11260 ( .A(n9416), .B(n9417), .Z(n9413) );
  ANDN U11261 ( .B(n9418), .A(n888), .Z(n9416) );
  XNOR U11262 ( .A(a[205]), .B(n9419), .Z(n888) );
  IV U11263 ( .A(n9417), .Z(n9419) );
  XNOR U11264 ( .A(b[205]), .B(n9417), .Z(n9418) );
  XOR U11265 ( .A(n9420), .B(n9421), .Z(n9417) );
  ANDN U11266 ( .B(n9422), .A(n889), .Z(n9420) );
  XNOR U11267 ( .A(a[204]), .B(n9423), .Z(n889) );
  IV U11268 ( .A(n9421), .Z(n9423) );
  XNOR U11269 ( .A(b[204]), .B(n9421), .Z(n9422) );
  XOR U11270 ( .A(n9424), .B(n9425), .Z(n9421) );
  ANDN U11271 ( .B(n9426), .A(n929), .Z(n9424) );
  XNOR U11272 ( .A(a[203]), .B(n9427), .Z(n929) );
  IV U11273 ( .A(n9425), .Z(n9427) );
  XNOR U11274 ( .A(b[203]), .B(n9425), .Z(n9426) );
  XOR U11275 ( .A(n9428), .B(n9429), .Z(n9425) );
  ANDN U11276 ( .B(n9430), .A(n980), .Z(n9428) );
  XNOR U11277 ( .A(a[202]), .B(n9431), .Z(n980) );
  IV U11278 ( .A(n9429), .Z(n9431) );
  XNOR U11279 ( .A(b[202]), .B(n9429), .Z(n9430) );
  XOR U11280 ( .A(n9432), .B(n9433), .Z(n9429) );
  ANDN U11281 ( .B(n9434), .A(n1031), .Z(n9432) );
  XNOR U11282 ( .A(a[201]), .B(n9435), .Z(n1031) );
  IV U11283 ( .A(n9433), .Z(n9435) );
  XNOR U11284 ( .A(b[201]), .B(n9433), .Z(n9434) );
  XOR U11285 ( .A(n9436), .B(n9437), .Z(n9433) );
  ANDN U11286 ( .B(n9438), .A(n1082), .Z(n9436) );
  XNOR U11287 ( .A(a[200]), .B(n9439), .Z(n1082) );
  IV U11288 ( .A(n9437), .Z(n9439) );
  XNOR U11289 ( .A(b[200]), .B(n9437), .Z(n9438) );
  XOR U11290 ( .A(n9440), .B(n9441), .Z(n9437) );
  ANDN U11291 ( .B(n9442), .A(n1135), .Z(n9440) );
  XNOR U11292 ( .A(a[199]), .B(n9443), .Z(n1135) );
  IV U11293 ( .A(n9441), .Z(n9443) );
  XNOR U11294 ( .A(b[199]), .B(n9441), .Z(n9442) );
  XOR U11295 ( .A(n9444), .B(n9445), .Z(n9441) );
  ANDN U11296 ( .B(n9446), .A(n1186), .Z(n9444) );
  XNOR U11297 ( .A(a[198]), .B(n9447), .Z(n1186) );
  IV U11298 ( .A(n9445), .Z(n9447) );
  XNOR U11299 ( .A(b[198]), .B(n9445), .Z(n9446) );
  XOR U11300 ( .A(n9448), .B(n9449), .Z(n9445) );
  ANDN U11301 ( .B(n9450), .A(n1237), .Z(n9448) );
  XNOR U11302 ( .A(a[197]), .B(n9451), .Z(n1237) );
  IV U11303 ( .A(n9449), .Z(n9451) );
  XNOR U11304 ( .A(b[197]), .B(n9449), .Z(n9450) );
  XOR U11305 ( .A(n9452), .B(n9453), .Z(n9449) );
  ANDN U11306 ( .B(n9454), .A(n1288), .Z(n9452) );
  XNOR U11307 ( .A(a[196]), .B(n9455), .Z(n1288) );
  IV U11308 ( .A(n9453), .Z(n9455) );
  XNOR U11309 ( .A(b[196]), .B(n9453), .Z(n9454) );
  XOR U11310 ( .A(n9456), .B(n9457), .Z(n9453) );
  ANDN U11311 ( .B(n9458), .A(n1339), .Z(n9456) );
  XNOR U11312 ( .A(a[195]), .B(n9459), .Z(n1339) );
  IV U11313 ( .A(n9457), .Z(n9459) );
  XNOR U11314 ( .A(b[195]), .B(n9457), .Z(n9458) );
  XOR U11315 ( .A(n9460), .B(n9461), .Z(n9457) );
  ANDN U11316 ( .B(n9462), .A(n1390), .Z(n9460) );
  XNOR U11317 ( .A(a[194]), .B(n9463), .Z(n1390) );
  IV U11318 ( .A(n9461), .Z(n9463) );
  XNOR U11319 ( .A(b[194]), .B(n9461), .Z(n9462) );
  XOR U11320 ( .A(n9464), .B(n9465), .Z(n9461) );
  ANDN U11321 ( .B(n9466), .A(n1441), .Z(n9464) );
  XNOR U11322 ( .A(a[193]), .B(n9467), .Z(n1441) );
  IV U11323 ( .A(n9465), .Z(n9467) );
  XNOR U11324 ( .A(b[193]), .B(n9465), .Z(n9466) );
  XOR U11325 ( .A(n9468), .B(n9469), .Z(n9465) );
  ANDN U11326 ( .B(n9470), .A(n1492), .Z(n9468) );
  XNOR U11327 ( .A(a[192]), .B(n9471), .Z(n1492) );
  IV U11328 ( .A(n9469), .Z(n9471) );
  XNOR U11329 ( .A(b[192]), .B(n9469), .Z(n9470) );
  XOR U11330 ( .A(n9472), .B(n9473), .Z(n9469) );
  ANDN U11331 ( .B(n9474), .A(n1543), .Z(n9472) );
  XNOR U11332 ( .A(a[191]), .B(n9475), .Z(n1543) );
  IV U11333 ( .A(n9473), .Z(n9475) );
  XNOR U11334 ( .A(b[191]), .B(n9473), .Z(n9474) );
  XOR U11335 ( .A(n9476), .B(n9477), .Z(n9473) );
  ANDN U11336 ( .B(n9478), .A(n1594), .Z(n9476) );
  XNOR U11337 ( .A(a[190]), .B(n9479), .Z(n1594) );
  IV U11338 ( .A(n9477), .Z(n9479) );
  XNOR U11339 ( .A(b[190]), .B(n9477), .Z(n9478) );
  XOR U11340 ( .A(n9480), .B(n9481), .Z(n9477) );
  ANDN U11341 ( .B(n9482), .A(n1646), .Z(n9480) );
  XNOR U11342 ( .A(a[189]), .B(n9483), .Z(n1646) );
  IV U11343 ( .A(n9481), .Z(n9483) );
  XNOR U11344 ( .A(b[189]), .B(n9481), .Z(n9482) );
  XOR U11345 ( .A(n9484), .B(n9485), .Z(n9481) );
  ANDN U11346 ( .B(n9486), .A(n1697), .Z(n9484) );
  XNOR U11347 ( .A(a[188]), .B(n9487), .Z(n1697) );
  IV U11348 ( .A(n9485), .Z(n9487) );
  XNOR U11349 ( .A(b[188]), .B(n9485), .Z(n9486) );
  XOR U11350 ( .A(n9488), .B(n9489), .Z(n9485) );
  ANDN U11351 ( .B(n9490), .A(n1748), .Z(n9488) );
  XNOR U11352 ( .A(a[187]), .B(n9491), .Z(n1748) );
  IV U11353 ( .A(n9489), .Z(n9491) );
  XNOR U11354 ( .A(b[187]), .B(n9489), .Z(n9490) );
  XOR U11355 ( .A(n9492), .B(n9493), .Z(n9489) );
  ANDN U11356 ( .B(n9494), .A(n1799), .Z(n9492) );
  XNOR U11357 ( .A(a[186]), .B(n9495), .Z(n1799) );
  IV U11358 ( .A(n9493), .Z(n9495) );
  XNOR U11359 ( .A(b[186]), .B(n9493), .Z(n9494) );
  XOR U11360 ( .A(n9496), .B(n9497), .Z(n9493) );
  ANDN U11361 ( .B(n9498), .A(n1850), .Z(n9496) );
  XNOR U11362 ( .A(a[185]), .B(n9499), .Z(n1850) );
  IV U11363 ( .A(n9497), .Z(n9499) );
  XNOR U11364 ( .A(b[185]), .B(n9497), .Z(n9498) );
  XOR U11365 ( .A(n9500), .B(n9501), .Z(n9497) );
  ANDN U11366 ( .B(n9502), .A(n1901), .Z(n9500) );
  XNOR U11367 ( .A(a[184]), .B(n9503), .Z(n1901) );
  IV U11368 ( .A(n9501), .Z(n9503) );
  XNOR U11369 ( .A(b[184]), .B(n9501), .Z(n9502) );
  XOR U11370 ( .A(n9504), .B(n9505), .Z(n9501) );
  ANDN U11371 ( .B(n9506), .A(n1952), .Z(n9504) );
  XNOR U11372 ( .A(a[183]), .B(n9507), .Z(n1952) );
  IV U11373 ( .A(n9505), .Z(n9507) );
  XNOR U11374 ( .A(b[183]), .B(n9505), .Z(n9506) );
  XOR U11375 ( .A(n9508), .B(n9509), .Z(n9505) );
  ANDN U11376 ( .B(n9510), .A(n2003), .Z(n9508) );
  XNOR U11377 ( .A(a[182]), .B(n9511), .Z(n2003) );
  IV U11378 ( .A(n9509), .Z(n9511) );
  XNOR U11379 ( .A(b[182]), .B(n9509), .Z(n9510) );
  XOR U11380 ( .A(n9512), .B(n9513), .Z(n9509) );
  ANDN U11381 ( .B(n9514), .A(n2054), .Z(n9512) );
  XNOR U11382 ( .A(a[181]), .B(n9515), .Z(n2054) );
  IV U11383 ( .A(n9513), .Z(n9515) );
  XNOR U11384 ( .A(b[181]), .B(n9513), .Z(n9514) );
  XOR U11385 ( .A(n9516), .B(n9517), .Z(n9513) );
  ANDN U11386 ( .B(n9518), .A(n2105), .Z(n9516) );
  XNOR U11387 ( .A(a[180]), .B(n9519), .Z(n2105) );
  IV U11388 ( .A(n9517), .Z(n9519) );
  XNOR U11389 ( .A(b[180]), .B(n9517), .Z(n9518) );
  XOR U11390 ( .A(n9520), .B(n9521), .Z(n9517) );
  ANDN U11391 ( .B(n9522), .A(n2157), .Z(n9520) );
  XNOR U11392 ( .A(a[179]), .B(n9523), .Z(n2157) );
  IV U11393 ( .A(n9521), .Z(n9523) );
  XNOR U11394 ( .A(b[179]), .B(n9521), .Z(n9522) );
  XOR U11395 ( .A(n9524), .B(n9525), .Z(n9521) );
  ANDN U11396 ( .B(n9526), .A(n2208), .Z(n9524) );
  XNOR U11397 ( .A(a[178]), .B(n9527), .Z(n2208) );
  IV U11398 ( .A(n9525), .Z(n9527) );
  XNOR U11399 ( .A(b[178]), .B(n9525), .Z(n9526) );
  XOR U11400 ( .A(n9528), .B(n9529), .Z(n9525) );
  ANDN U11401 ( .B(n9530), .A(n2259), .Z(n9528) );
  XNOR U11402 ( .A(a[177]), .B(n9531), .Z(n2259) );
  IV U11403 ( .A(n9529), .Z(n9531) );
  XNOR U11404 ( .A(b[177]), .B(n9529), .Z(n9530) );
  XOR U11405 ( .A(n9532), .B(n9533), .Z(n9529) );
  ANDN U11406 ( .B(n9534), .A(n2310), .Z(n9532) );
  XNOR U11407 ( .A(a[176]), .B(n9535), .Z(n2310) );
  IV U11408 ( .A(n9533), .Z(n9535) );
  XNOR U11409 ( .A(b[176]), .B(n9533), .Z(n9534) );
  XOR U11410 ( .A(n9536), .B(n9537), .Z(n9533) );
  ANDN U11411 ( .B(n9538), .A(n2361), .Z(n9536) );
  XNOR U11412 ( .A(a[175]), .B(n9539), .Z(n2361) );
  IV U11413 ( .A(n9537), .Z(n9539) );
  XNOR U11414 ( .A(b[175]), .B(n9537), .Z(n9538) );
  XOR U11415 ( .A(n9540), .B(n9541), .Z(n9537) );
  ANDN U11416 ( .B(n9542), .A(n2412), .Z(n9540) );
  XNOR U11417 ( .A(a[174]), .B(n9543), .Z(n2412) );
  IV U11418 ( .A(n9541), .Z(n9543) );
  XNOR U11419 ( .A(b[174]), .B(n9541), .Z(n9542) );
  XOR U11420 ( .A(n9544), .B(n9545), .Z(n9541) );
  ANDN U11421 ( .B(n9546), .A(n2463), .Z(n9544) );
  XNOR U11422 ( .A(a[173]), .B(n9547), .Z(n2463) );
  IV U11423 ( .A(n9545), .Z(n9547) );
  XNOR U11424 ( .A(b[173]), .B(n9545), .Z(n9546) );
  XOR U11425 ( .A(n9548), .B(n9549), .Z(n9545) );
  ANDN U11426 ( .B(n9550), .A(n2514), .Z(n9548) );
  XNOR U11427 ( .A(a[172]), .B(n9551), .Z(n2514) );
  IV U11428 ( .A(n9549), .Z(n9551) );
  XNOR U11429 ( .A(b[172]), .B(n9549), .Z(n9550) );
  XOR U11430 ( .A(n9552), .B(n9553), .Z(n9549) );
  ANDN U11431 ( .B(n9554), .A(n2565), .Z(n9552) );
  XNOR U11432 ( .A(a[171]), .B(n9555), .Z(n2565) );
  IV U11433 ( .A(n9553), .Z(n9555) );
  XNOR U11434 ( .A(b[171]), .B(n9553), .Z(n9554) );
  XOR U11435 ( .A(n9556), .B(n9557), .Z(n9553) );
  ANDN U11436 ( .B(n9558), .A(n2616), .Z(n9556) );
  XNOR U11437 ( .A(a[170]), .B(n9559), .Z(n2616) );
  IV U11438 ( .A(n9557), .Z(n9559) );
  XNOR U11439 ( .A(b[170]), .B(n9557), .Z(n9558) );
  XOR U11440 ( .A(n9560), .B(n9561), .Z(n9557) );
  ANDN U11441 ( .B(n9562), .A(n2668), .Z(n9560) );
  XNOR U11442 ( .A(a[169]), .B(n9563), .Z(n2668) );
  IV U11443 ( .A(n9561), .Z(n9563) );
  XNOR U11444 ( .A(b[169]), .B(n9561), .Z(n9562) );
  XOR U11445 ( .A(n9564), .B(n9565), .Z(n9561) );
  ANDN U11446 ( .B(n9566), .A(n2719), .Z(n9564) );
  XNOR U11447 ( .A(a[168]), .B(n9567), .Z(n2719) );
  IV U11448 ( .A(n9565), .Z(n9567) );
  XNOR U11449 ( .A(b[168]), .B(n9565), .Z(n9566) );
  XOR U11450 ( .A(n9568), .B(n9569), .Z(n9565) );
  ANDN U11451 ( .B(n9570), .A(n2770), .Z(n9568) );
  XNOR U11452 ( .A(a[167]), .B(n9571), .Z(n2770) );
  IV U11453 ( .A(n9569), .Z(n9571) );
  XNOR U11454 ( .A(b[167]), .B(n9569), .Z(n9570) );
  XOR U11455 ( .A(n9572), .B(n9573), .Z(n9569) );
  ANDN U11456 ( .B(n9574), .A(n2821), .Z(n9572) );
  XNOR U11457 ( .A(a[166]), .B(n9575), .Z(n2821) );
  IV U11458 ( .A(n9573), .Z(n9575) );
  XNOR U11459 ( .A(b[166]), .B(n9573), .Z(n9574) );
  XOR U11460 ( .A(n9576), .B(n9577), .Z(n9573) );
  ANDN U11461 ( .B(n9578), .A(n2872), .Z(n9576) );
  XNOR U11462 ( .A(a[165]), .B(n9579), .Z(n2872) );
  IV U11463 ( .A(n9577), .Z(n9579) );
  XNOR U11464 ( .A(b[165]), .B(n9577), .Z(n9578) );
  XOR U11465 ( .A(n9580), .B(n9581), .Z(n9577) );
  ANDN U11466 ( .B(n9582), .A(n2923), .Z(n9580) );
  XNOR U11467 ( .A(a[164]), .B(n9583), .Z(n2923) );
  IV U11468 ( .A(n9581), .Z(n9583) );
  XNOR U11469 ( .A(b[164]), .B(n9581), .Z(n9582) );
  XOR U11470 ( .A(n9584), .B(n9585), .Z(n9581) );
  ANDN U11471 ( .B(n9586), .A(n2974), .Z(n9584) );
  XNOR U11472 ( .A(a[163]), .B(n9587), .Z(n2974) );
  IV U11473 ( .A(n9585), .Z(n9587) );
  XNOR U11474 ( .A(b[163]), .B(n9585), .Z(n9586) );
  XOR U11475 ( .A(n9588), .B(n9589), .Z(n9585) );
  ANDN U11476 ( .B(n9590), .A(n3025), .Z(n9588) );
  XNOR U11477 ( .A(a[162]), .B(n9591), .Z(n3025) );
  IV U11478 ( .A(n9589), .Z(n9591) );
  XNOR U11479 ( .A(b[162]), .B(n9589), .Z(n9590) );
  XOR U11480 ( .A(n9592), .B(n9593), .Z(n9589) );
  ANDN U11481 ( .B(n9594), .A(n3076), .Z(n9592) );
  XNOR U11482 ( .A(a[161]), .B(n9595), .Z(n3076) );
  IV U11483 ( .A(n9593), .Z(n9595) );
  XNOR U11484 ( .A(b[161]), .B(n9593), .Z(n9594) );
  XOR U11485 ( .A(n9596), .B(n9597), .Z(n9593) );
  ANDN U11486 ( .B(n9598), .A(n3127), .Z(n9596) );
  XNOR U11487 ( .A(a[160]), .B(n9599), .Z(n3127) );
  IV U11488 ( .A(n9597), .Z(n9599) );
  XNOR U11489 ( .A(b[160]), .B(n9597), .Z(n9598) );
  XOR U11490 ( .A(n9600), .B(n9601), .Z(n9597) );
  ANDN U11491 ( .B(n9602), .A(n3179), .Z(n9600) );
  XNOR U11492 ( .A(a[159]), .B(n9603), .Z(n3179) );
  IV U11493 ( .A(n9601), .Z(n9603) );
  XNOR U11494 ( .A(b[159]), .B(n9601), .Z(n9602) );
  XOR U11495 ( .A(n9604), .B(n9605), .Z(n9601) );
  ANDN U11496 ( .B(n9606), .A(n3230), .Z(n9604) );
  XNOR U11497 ( .A(a[158]), .B(n9607), .Z(n3230) );
  IV U11498 ( .A(n9605), .Z(n9607) );
  XNOR U11499 ( .A(b[158]), .B(n9605), .Z(n9606) );
  XOR U11500 ( .A(n9608), .B(n9609), .Z(n9605) );
  ANDN U11501 ( .B(n9610), .A(n3281), .Z(n9608) );
  XNOR U11502 ( .A(a[157]), .B(n9611), .Z(n3281) );
  IV U11503 ( .A(n9609), .Z(n9611) );
  XNOR U11504 ( .A(b[157]), .B(n9609), .Z(n9610) );
  XOR U11505 ( .A(n9612), .B(n9613), .Z(n9609) );
  ANDN U11506 ( .B(n9614), .A(n3332), .Z(n9612) );
  XNOR U11507 ( .A(a[156]), .B(n9615), .Z(n3332) );
  IV U11508 ( .A(n9613), .Z(n9615) );
  XNOR U11509 ( .A(b[156]), .B(n9613), .Z(n9614) );
  XOR U11510 ( .A(n9616), .B(n9617), .Z(n9613) );
  ANDN U11511 ( .B(n9618), .A(n3383), .Z(n9616) );
  XNOR U11512 ( .A(a[155]), .B(n9619), .Z(n3383) );
  IV U11513 ( .A(n9617), .Z(n9619) );
  XNOR U11514 ( .A(b[155]), .B(n9617), .Z(n9618) );
  XOR U11515 ( .A(n9620), .B(n9621), .Z(n9617) );
  ANDN U11516 ( .B(n9622), .A(n3434), .Z(n9620) );
  XNOR U11517 ( .A(a[154]), .B(n9623), .Z(n3434) );
  IV U11518 ( .A(n9621), .Z(n9623) );
  XNOR U11519 ( .A(b[154]), .B(n9621), .Z(n9622) );
  XOR U11520 ( .A(n9624), .B(n9625), .Z(n9621) );
  ANDN U11521 ( .B(n9626), .A(n3485), .Z(n9624) );
  XNOR U11522 ( .A(a[153]), .B(n9627), .Z(n3485) );
  IV U11523 ( .A(n9625), .Z(n9627) );
  XNOR U11524 ( .A(b[153]), .B(n9625), .Z(n9626) );
  XOR U11525 ( .A(n9628), .B(n9629), .Z(n9625) );
  ANDN U11526 ( .B(n9630), .A(n3536), .Z(n9628) );
  XNOR U11527 ( .A(a[152]), .B(n9631), .Z(n3536) );
  IV U11528 ( .A(n9629), .Z(n9631) );
  XNOR U11529 ( .A(b[152]), .B(n9629), .Z(n9630) );
  XOR U11530 ( .A(n9632), .B(n9633), .Z(n9629) );
  ANDN U11531 ( .B(n9634), .A(n3587), .Z(n9632) );
  XNOR U11532 ( .A(a[151]), .B(n9635), .Z(n3587) );
  IV U11533 ( .A(n9633), .Z(n9635) );
  XNOR U11534 ( .A(b[151]), .B(n9633), .Z(n9634) );
  XOR U11535 ( .A(n9636), .B(n9637), .Z(n9633) );
  ANDN U11536 ( .B(n9638), .A(n3638), .Z(n9636) );
  XNOR U11537 ( .A(a[150]), .B(n9639), .Z(n3638) );
  IV U11538 ( .A(n9637), .Z(n9639) );
  XNOR U11539 ( .A(b[150]), .B(n9637), .Z(n9638) );
  XOR U11540 ( .A(n9640), .B(n9641), .Z(n9637) );
  ANDN U11541 ( .B(n9642), .A(n3690), .Z(n9640) );
  XNOR U11542 ( .A(a[149]), .B(n9643), .Z(n3690) );
  IV U11543 ( .A(n9641), .Z(n9643) );
  XNOR U11544 ( .A(b[149]), .B(n9641), .Z(n9642) );
  XOR U11545 ( .A(n9644), .B(n9645), .Z(n9641) );
  ANDN U11546 ( .B(n9646), .A(n3741), .Z(n9644) );
  XNOR U11547 ( .A(a[148]), .B(n9647), .Z(n3741) );
  IV U11548 ( .A(n9645), .Z(n9647) );
  XNOR U11549 ( .A(b[148]), .B(n9645), .Z(n9646) );
  XOR U11550 ( .A(n9648), .B(n9649), .Z(n9645) );
  ANDN U11551 ( .B(n9650), .A(n3792), .Z(n9648) );
  XNOR U11552 ( .A(a[147]), .B(n9651), .Z(n3792) );
  IV U11553 ( .A(n9649), .Z(n9651) );
  XNOR U11554 ( .A(b[147]), .B(n9649), .Z(n9650) );
  XOR U11555 ( .A(n9652), .B(n9653), .Z(n9649) );
  ANDN U11556 ( .B(n9654), .A(n3843), .Z(n9652) );
  XNOR U11557 ( .A(a[146]), .B(n9655), .Z(n3843) );
  IV U11558 ( .A(n9653), .Z(n9655) );
  XNOR U11559 ( .A(b[146]), .B(n9653), .Z(n9654) );
  XOR U11560 ( .A(n9656), .B(n9657), .Z(n9653) );
  ANDN U11561 ( .B(n9658), .A(n3894), .Z(n9656) );
  XNOR U11562 ( .A(a[145]), .B(n9659), .Z(n3894) );
  IV U11563 ( .A(n9657), .Z(n9659) );
  XNOR U11564 ( .A(b[145]), .B(n9657), .Z(n9658) );
  XOR U11565 ( .A(n9660), .B(n9661), .Z(n9657) );
  ANDN U11566 ( .B(n9662), .A(n3945), .Z(n9660) );
  XNOR U11567 ( .A(a[144]), .B(n9663), .Z(n3945) );
  IV U11568 ( .A(n9661), .Z(n9663) );
  XNOR U11569 ( .A(b[144]), .B(n9661), .Z(n9662) );
  XOR U11570 ( .A(n9664), .B(n9665), .Z(n9661) );
  ANDN U11571 ( .B(n9666), .A(n3996), .Z(n9664) );
  XNOR U11572 ( .A(a[143]), .B(n9667), .Z(n3996) );
  IV U11573 ( .A(n9665), .Z(n9667) );
  XNOR U11574 ( .A(b[143]), .B(n9665), .Z(n9666) );
  XOR U11575 ( .A(n9668), .B(n9669), .Z(n9665) );
  ANDN U11576 ( .B(n9670), .A(n4047), .Z(n9668) );
  XNOR U11577 ( .A(a[142]), .B(n9671), .Z(n4047) );
  IV U11578 ( .A(n9669), .Z(n9671) );
  XNOR U11579 ( .A(b[142]), .B(n9669), .Z(n9670) );
  XOR U11580 ( .A(n9672), .B(n9673), .Z(n9669) );
  ANDN U11581 ( .B(n9674), .A(n4098), .Z(n9672) );
  XNOR U11582 ( .A(a[141]), .B(n9675), .Z(n4098) );
  IV U11583 ( .A(n9673), .Z(n9675) );
  XNOR U11584 ( .A(b[141]), .B(n9673), .Z(n9674) );
  XOR U11585 ( .A(n9676), .B(n9677), .Z(n9673) );
  ANDN U11586 ( .B(n9678), .A(n4149), .Z(n9676) );
  XNOR U11587 ( .A(a[140]), .B(n9679), .Z(n4149) );
  IV U11588 ( .A(n9677), .Z(n9679) );
  XNOR U11589 ( .A(b[140]), .B(n9677), .Z(n9678) );
  XOR U11590 ( .A(n9680), .B(n9681), .Z(n9677) );
  ANDN U11591 ( .B(n9682), .A(n4201), .Z(n9680) );
  XNOR U11592 ( .A(a[139]), .B(n9683), .Z(n4201) );
  IV U11593 ( .A(n9681), .Z(n9683) );
  XNOR U11594 ( .A(b[139]), .B(n9681), .Z(n9682) );
  XOR U11595 ( .A(n9684), .B(n9685), .Z(n9681) );
  ANDN U11596 ( .B(n9686), .A(n4252), .Z(n9684) );
  XNOR U11597 ( .A(a[138]), .B(n9687), .Z(n4252) );
  IV U11598 ( .A(n9685), .Z(n9687) );
  XNOR U11599 ( .A(b[138]), .B(n9685), .Z(n9686) );
  XOR U11600 ( .A(n9688), .B(n9689), .Z(n9685) );
  ANDN U11601 ( .B(n9690), .A(n4303), .Z(n9688) );
  XNOR U11602 ( .A(a[137]), .B(n9691), .Z(n4303) );
  IV U11603 ( .A(n9689), .Z(n9691) );
  XNOR U11604 ( .A(b[137]), .B(n9689), .Z(n9690) );
  XOR U11605 ( .A(n9692), .B(n9693), .Z(n9689) );
  ANDN U11606 ( .B(n9694), .A(n4354), .Z(n9692) );
  XNOR U11607 ( .A(a[136]), .B(n9695), .Z(n4354) );
  IV U11608 ( .A(n9693), .Z(n9695) );
  XNOR U11609 ( .A(b[136]), .B(n9693), .Z(n9694) );
  XOR U11610 ( .A(n9696), .B(n9697), .Z(n9693) );
  ANDN U11611 ( .B(n9698), .A(n4405), .Z(n9696) );
  XNOR U11612 ( .A(a[135]), .B(n9699), .Z(n4405) );
  IV U11613 ( .A(n9697), .Z(n9699) );
  XNOR U11614 ( .A(b[135]), .B(n9697), .Z(n9698) );
  XOR U11615 ( .A(n9700), .B(n9701), .Z(n9697) );
  ANDN U11616 ( .B(n9702), .A(n4456), .Z(n9700) );
  XNOR U11617 ( .A(a[134]), .B(n9703), .Z(n4456) );
  IV U11618 ( .A(n9701), .Z(n9703) );
  XNOR U11619 ( .A(b[134]), .B(n9701), .Z(n9702) );
  XOR U11620 ( .A(n9704), .B(n9705), .Z(n9701) );
  ANDN U11621 ( .B(n9706), .A(n4507), .Z(n9704) );
  XNOR U11622 ( .A(a[133]), .B(n9707), .Z(n4507) );
  IV U11623 ( .A(n9705), .Z(n9707) );
  XNOR U11624 ( .A(b[133]), .B(n9705), .Z(n9706) );
  XOR U11625 ( .A(n9708), .B(n9709), .Z(n9705) );
  ANDN U11626 ( .B(n9710), .A(n4558), .Z(n9708) );
  XNOR U11627 ( .A(a[132]), .B(n9711), .Z(n4558) );
  IV U11628 ( .A(n9709), .Z(n9711) );
  XNOR U11629 ( .A(b[132]), .B(n9709), .Z(n9710) );
  XOR U11630 ( .A(n9712), .B(n9713), .Z(n9709) );
  ANDN U11631 ( .B(n9714), .A(n4609), .Z(n9712) );
  XNOR U11632 ( .A(a[131]), .B(n9715), .Z(n4609) );
  IV U11633 ( .A(n9713), .Z(n9715) );
  XNOR U11634 ( .A(b[131]), .B(n9713), .Z(n9714) );
  XOR U11635 ( .A(n9716), .B(n9717), .Z(n9713) );
  ANDN U11636 ( .B(n9718), .A(n4660), .Z(n9716) );
  XNOR U11637 ( .A(a[130]), .B(n9719), .Z(n4660) );
  IV U11638 ( .A(n9717), .Z(n9719) );
  XNOR U11639 ( .A(b[130]), .B(n9717), .Z(n9718) );
  XOR U11640 ( .A(n9720), .B(n9721), .Z(n9717) );
  ANDN U11641 ( .B(n9722), .A(n4712), .Z(n9720) );
  XNOR U11642 ( .A(a[129]), .B(n9723), .Z(n4712) );
  IV U11643 ( .A(n9721), .Z(n9723) );
  XNOR U11644 ( .A(b[129]), .B(n9721), .Z(n9722) );
  XOR U11645 ( .A(n9724), .B(n9725), .Z(n9721) );
  ANDN U11646 ( .B(n9726), .A(n4763), .Z(n9724) );
  XNOR U11647 ( .A(a[128]), .B(n9727), .Z(n4763) );
  IV U11648 ( .A(n9725), .Z(n9727) );
  XNOR U11649 ( .A(b[128]), .B(n9725), .Z(n9726) );
  XOR U11650 ( .A(n9728), .B(n9729), .Z(n9725) );
  ANDN U11651 ( .B(n9730), .A(n4814), .Z(n9728) );
  XNOR U11652 ( .A(a[127]), .B(n9731), .Z(n4814) );
  IV U11653 ( .A(n9729), .Z(n9731) );
  XNOR U11654 ( .A(b[127]), .B(n9729), .Z(n9730) );
  XOR U11655 ( .A(n9732), .B(n9733), .Z(n9729) );
  ANDN U11656 ( .B(n9734), .A(n4865), .Z(n9732) );
  XNOR U11657 ( .A(a[126]), .B(n9735), .Z(n4865) );
  IV U11658 ( .A(n9733), .Z(n9735) );
  XNOR U11659 ( .A(b[126]), .B(n9733), .Z(n9734) );
  XOR U11660 ( .A(n9736), .B(n9737), .Z(n9733) );
  ANDN U11661 ( .B(n9738), .A(n4916), .Z(n9736) );
  XNOR U11662 ( .A(a[125]), .B(n9739), .Z(n4916) );
  IV U11663 ( .A(n9737), .Z(n9739) );
  XNOR U11664 ( .A(b[125]), .B(n9737), .Z(n9738) );
  XOR U11665 ( .A(n9740), .B(n9741), .Z(n9737) );
  ANDN U11666 ( .B(n9742), .A(n4967), .Z(n9740) );
  XNOR U11667 ( .A(a[124]), .B(n9743), .Z(n4967) );
  IV U11668 ( .A(n9741), .Z(n9743) );
  XNOR U11669 ( .A(b[124]), .B(n9741), .Z(n9742) );
  XOR U11670 ( .A(n9744), .B(n9745), .Z(n9741) );
  ANDN U11671 ( .B(n9746), .A(n5018), .Z(n9744) );
  XNOR U11672 ( .A(a[123]), .B(n9747), .Z(n5018) );
  IV U11673 ( .A(n9745), .Z(n9747) );
  XNOR U11674 ( .A(b[123]), .B(n9745), .Z(n9746) );
  XOR U11675 ( .A(n9748), .B(n9749), .Z(n9745) );
  ANDN U11676 ( .B(n9750), .A(n5069), .Z(n9748) );
  XNOR U11677 ( .A(a[122]), .B(n9751), .Z(n5069) );
  IV U11678 ( .A(n9749), .Z(n9751) );
  XNOR U11679 ( .A(b[122]), .B(n9749), .Z(n9750) );
  XOR U11680 ( .A(n9752), .B(n9753), .Z(n9749) );
  ANDN U11681 ( .B(n9754), .A(n5120), .Z(n9752) );
  XNOR U11682 ( .A(a[121]), .B(n9755), .Z(n5120) );
  IV U11683 ( .A(n9753), .Z(n9755) );
  XNOR U11684 ( .A(b[121]), .B(n9753), .Z(n9754) );
  XOR U11685 ( .A(n9756), .B(n9757), .Z(n9753) );
  ANDN U11686 ( .B(n9758), .A(n5171), .Z(n9756) );
  XNOR U11687 ( .A(a[120]), .B(n9759), .Z(n5171) );
  IV U11688 ( .A(n9757), .Z(n9759) );
  XNOR U11689 ( .A(b[120]), .B(n9757), .Z(n9758) );
  XOR U11690 ( .A(n9760), .B(n9761), .Z(n9757) );
  ANDN U11691 ( .B(n9762), .A(n5223), .Z(n9760) );
  XNOR U11692 ( .A(a[119]), .B(n9763), .Z(n5223) );
  IV U11693 ( .A(n9761), .Z(n9763) );
  XNOR U11694 ( .A(b[119]), .B(n9761), .Z(n9762) );
  XOR U11695 ( .A(n9764), .B(n9765), .Z(n9761) );
  ANDN U11696 ( .B(n9766), .A(n5274), .Z(n9764) );
  XNOR U11697 ( .A(a[118]), .B(n9767), .Z(n5274) );
  IV U11698 ( .A(n9765), .Z(n9767) );
  XNOR U11699 ( .A(b[118]), .B(n9765), .Z(n9766) );
  XOR U11700 ( .A(n9768), .B(n9769), .Z(n9765) );
  ANDN U11701 ( .B(n9770), .A(n5325), .Z(n9768) );
  XNOR U11702 ( .A(a[117]), .B(n9771), .Z(n5325) );
  IV U11703 ( .A(n9769), .Z(n9771) );
  XNOR U11704 ( .A(b[117]), .B(n9769), .Z(n9770) );
  XOR U11705 ( .A(n9772), .B(n9773), .Z(n9769) );
  ANDN U11706 ( .B(n9774), .A(n5376), .Z(n9772) );
  XNOR U11707 ( .A(a[116]), .B(n9775), .Z(n5376) );
  IV U11708 ( .A(n9773), .Z(n9775) );
  XNOR U11709 ( .A(b[116]), .B(n9773), .Z(n9774) );
  XOR U11710 ( .A(n9776), .B(n9777), .Z(n9773) );
  ANDN U11711 ( .B(n9778), .A(n5427), .Z(n9776) );
  XNOR U11712 ( .A(a[115]), .B(n9779), .Z(n5427) );
  IV U11713 ( .A(n9777), .Z(n9779) );
  XNOR U11714 ( .A(b[115]), .B(n9777), .Z(n9778) );
  XOR U11715 ( .A(n9780), .B(n9781), .Z(n9777) );
  ANDN U11716 ( .B(n9782), .A(n5478), .Z(n9780) );
  XNOR U11717 ( .A(a[114]), .B(n9783), .Z(n5478) );
  IV U11718 ( .A(n9781), .Z(n9783) );
  XNOR U11719 ( .A(b[114]), .B(n9781), .Z(n9782) );
  XOR U11720 ( .A(n9784), .B(n9785), .Z(n9781) );
  ANDN U11721 ( .B(n9786), .A(n5529), .Z(n9784) );
  XNOR U11722 ( .A(a[113]), .B(n9787), .Z(n5529) );
  IV U11723 ( .A(n9785), .Z(n9787) );
  XNOR U11724 ( .A(b[113]), .B(n9785), .Z(n9786) );
  XOR U11725 ( .A(n9788), .B(n9789), .Z(n9785) );
  ANDN U11726 ( .B(n9790), .A(n5580), .Z(n9788) );
  XNOR U11727 ( .A(a[112]), .B(n9791), .Z(n5580) );
  IV U11728 ( .A(n9789), .Z(n9791) );
  XNOR U11729 ( .A(b[112]), .B(n9789), .Z(n9790) );
  XOR U11730 ( .A(n9792), .B(n9793), .Z(n9789) );
  ANDN U11731 ( .B(n9794), .A(n5631), .Z(n9792) );
  XNOR U11732 ( .A(a[111]), .B(n9795), .Z(n5631) );
  IV U11733 ( .A(n9793), .Z(n9795) );
  XNOR U11734 ( .A(b[111]), .B(n9793), .Z(n9794) );
  XOR U11735 ( .A(n9796), .B(n9797), .Z(n9793) );
  ANDN U11736 ( .B(n9798), .A(n5682), .Z(n9796) );
  XNOR U11737 ( .A(a[110]), .B(n9799), .Z(n5682) );
  IV U11738 ( .A(n9797), .Z(n9799) );
  XNOR U11739 ( .A(b[110]), .B(n9797), .Z(n9798) );
  XOR U11740 ( .A(n9800), .B(n9801), .Z(n9797) );
  ANDN U11741 ( .B(n9802), .A(n5734), .Z(n9800) );
  XNOR U11742 ( .A(a[109]), .B(n9803), .Z(n5734) );
  IV U11743 ( .A(n9801), .Z(n9803) );
  XNOR U11744 ( .A(b[109]), .B(n9801), .Z(n9802) );
  XOR U11745 ( .A(n9804), .B(n9805), .Z(n9801) );
  ANDN U11746 ( .B(n9806), .A(n5785), .Z(n9804) );
  XNOR U11747 ( .A(a[108]), .B(n9807), .Z(n5785) );
  IV U11748 ( .A(n9805), .Z(n9807) );
  XNOR U11749 ( .A(b[108]), .B(n9805), .Z(n9806) );
  XOR U11750 ( .A(n9808), .B(n9809), .Z(n9805) );
  ANDN U11751 ( .B(n9810), .A(n5836), .Z(n9808) );
  XNOR U11752 ( .A(a[107]), .B(n9811), .Z(n5836) );
  IV U11753 ( .A(n9809), .Z(n9811) );
  XNOR U11754 ( .A(b[107]), .B(n9809), .Z(n9810) );
  XOR U11755 ( .A(n9812), .B(n9813), .Z(n9809) );
  ANDN U11756 ( .B(n9814), .A(n5887), .Z(n9812) );
  XNOR U11757 ( .A(a[106]), .B(n9815), .Z(n5887) );
  IV U11758 ( .A(n9813), .Z(n9815) );
  XNOR U11759 ( .A(b[106]), .B(n9813), .Z(n9814) );
  XOR U11760 ( .A(n9816), .B(n9817), .Z(n9813) );
  ANDN U11761 ( .B(n9818), .A(n5938), .Z(n9816) );
  XNOR U11762 ( .A(a[105]), .B(n9819), .Z(n5938) );
  IV U11763 ( .A(n9817), .Z(n9819) );
  XNOR U11764 ( .A(b[105]), .B(n9817), .Z(n9818) );
  XOR U11765 ( .A(n9820), .B(n9821), .Z(n9817) );
  ANDN U11766 ( .B(n9822), .A(n5989), .Z(n9820) );
  XNOR U11767 ( .A(a[104]), .B(n9823), .Z(n5989) );
  IV U11768 ( .A(n9821), .Z(n9823) );
  XNOR U11769 ( .A(b[104]), .B(n9821), .Z(n9822) );
  XOR U11770 ( .A(n9824), .B(n9825), .Z(n9821) );
  ANDN U11771 ( .B(n9826), .A(n6040), .Z(n9824) );
  XNOR U11772 ( .A(a[103]), .B(n9827), .Z(n6040) );
  IV U11773 ( .A(n9825), .Z(n9827) );
  XNOR U11774 ( .A(b[103]), .B(n9825), .Z(n9826) );
  XOR U11775 ( .A(n9828), .B(n9829), .Z(n9825) );
  ANDN U11776 ( .B(n9830), .A(n6091), .Z(n9828) );
  XNOR U11777 ( .A(a[102]), .B(n9831), .Z(n6091) );
  IV U11778 ( .A(n9829), .Z(n9831) );
  XNOR U11779 ( .A(b[102]), .B(n9829), .Z(n9830) );
  XOR U11780 ( .A(n9832), .B(n9833), .Z(n9829) );
  ANDN U11781 ( .B(n9834), .A(n6142), .Z(n9832) );
  XNOR U11782 ( .A(a[101]), .B(n9835), .Z(n6142) );
  IV U11783 ( .A(n9833), .Z(n9835) );
  XNOR U11784 ( .A(b[101]), .B(n9833), .Z(n9834) );
  XOR U11785 ( .A(n9836), .B(n9837), .Z(n9833) );
  ANDN U11786 ( .B(n9838), .A(n6193), .Z(n9836) );
  XNOR U11787 ( .A(a[100]), .B(n9839), .Z(n6193) );
  IV U11788 ( .A(n9837), .Z(n9839) );
  XNOR U11789 ( .A(b[100]), .B(n9837), .Z(n9838) );
  XOR U11790 ( .A(n9840), .B(n9841), .Z(n9837) );
  ANDN U11791 ( .B(n9842), .A(n7), .Z(n9840) );
  XNOR U11792 ( .A(a[99]), .B(n9843), .Z(n7) );
  IV U11793 ( .A(n9841), .Z(n9843) );
  XNOR U11794 ( .A(b[99]), .B(n9841), .Z(n9842) );
  XOR U11795 ( .A(n9844), .B(n9845), .Z(n9841) );
  ANDN U11796 ( .B(n9846), .A(n18), .Z(n9844) );
  XNOR U11797 ( .A(a[98]), .B(n9847), .Z(n18) );
  IV U11798 ( .A(n9845), .Z(n9847) );
  XNOR U11799 ( .A(b[98]), .B(n9845), .Z(n9846) );
  XOR U11800 ( .A(n9848), .B(n9849), .Z(n9845) );
  ANDN U11801 ( .B(n9850), .A(n29), .Z(n9848) );
  XNOR U11802 ( .A(a[97]), .B(n9851), .Z(n29) );
  IV U11803 ( .A(n9849), .Z(n9851) );
  XNOR U11804 ( .A(b[97]), .B(n9849), .Z(n9850) );
  XOR U11805 ( .A(n9852), .B(n9853), .Z(n9849) );
  ANDN U11806 ( .B(n9854), .A(n40), .Z(n9852) );
  XNOR U11807 ( .A(a[96]), .B(n9855), .Z(n40) );
  IV U11808 ( .A(n9853), .Z(n9855) );
  XNOR U11809 ( .A(b[96]), .B(n9853), .Z(n9854) );
  XOR U11810 ( .A(n9856), .B(n9857), .Z(n9853) );
  ANDN U11811 ( .B(n9858), .A(n51), .Z(n9856) );
  XNOR U11812 ( .A(a[95]), .B(n9859), .Z(n51) );
  IV U11813 ( .A(n9857), .Z(n9859) );
  XNOR U11814 ( .A(b[95]), .B(n9857), .Z(n9858) );
  XOR U11815 ( .A(n9860), .B(n9861), .Z(n9857) );
  ANDN U11816 ( .B(n9862), .A(n62), .Z(n9860) );
  XNOR U11817 ( .A(a[94]), .B(n9863), .Z(n62) );
  IV U11818 ( .A(n9861), .Z(n9863) );
  XNOR U11819 ( .A(b[94]), .B(n9861), .Z(n9862) );
  XOR U11820 ( .A(n9864), .B(n9865), .Z(n9861) );
  ANDN U11821 ( .B(n9866), .A(n73), .Z(n9864) );
  XNOR U11822 ( .A(a[93]), .B(n9867), .Z(n73) );
  IV U11823 ( .A(n9865), .Z(n9867) );
  XNOR U11824 ( .A(b[93]), .B(n9865), .Z(n9866) );
  XOR U11825 ( .A(n9868), .B(n9869), .Z(n9865) );
  ANDN U11826 ( .B(n9870), .A(n84), .Z(n9868) );
  XNOR U11827 ( .A(a[92]), .B(n9871), .Z(n84) );
  IV U11828 ( .A(n9869), .Z(n9871) );
  XNOR U11829 ( .A(b[92]), .B(n9869), .Z(n9870) );
  XOR U11830 ( .A(n9872), .B(n9873), .Z(n9869) );
  ANDN U11831 ( .B(n9874), .A(n95), .Z(n9872) );
  XNOR U11832 ( .A(a[91]), .B(n9875), .Z(n95) );
  IV U11833 ( .A(n9873), .Z(n9875) );
  XNOR U11834 ( .A(b[91]), .B(n9873), .Z(n9874) );
  XOR U11835 ( .A(n9876), .B(n9877), .Z(n9873) );
  ANDN U11836 ( .B(n9878), .A(n106), .Z(n9876) );
  XNOR U11837 ( .A(a[90]), .B(n9879), .Z(n106) );
  IV U11838 ( .A(n9877), .Z(n9879) );
  XNOR U11839 ( .A(b[90]), .B(n9877), .Z(n9878) );
  XOR U11840 ( .A(n9880), .B(n9881), .Z(n9877) );
  ANDN U11841 ( .B(n9882), .A(n118), .Z(n9880) );
  XNOR U11842 ( .A(a[89]), .B(n9883), .Z(n118) );
  IV U11843 ( .A(n9881), .Z(n9883) );
  XNOR U11844 ( .A(b[89]), .B(n9881), .Z(n9882) );
  XOR U11845 ( .A(n9884), .B(n9885), .Z(n9881) );
  ANDN U11846 ( .B(n9886), .A(n129), .Z(n9884) );
  XNOR U11847 ( .A(a[88]), .B(n9887), .Z(n129) );
  IV U11848 ( .A(n9885), .Z(n9887) );
  XNOR U11849 ( .A(b[88]), .B(n9885), .Z(n9886) );
  XOR U11850 ( .A(n9888), .B(n9889), .Z(n9885) );
  ANDN U11851 ( .B(n9890), .A(n140), .Z(n9888) );
  XNOR U11852 ( .A(a[87]), .B(n9891), .Z(n140) );
  IV U11853 ( .A(n9889), .Z(n9891) );
  XNOR U11854 ( .A(b[87]), .B(n9889), .Z(n9890) );
  XOR U11855 ( .A(n9892), .B(n9893), .Z(n9889) );
  ANDN U11856 ( .B(n9894), .A(n151), .Z(n9892) );
  XNOR U11857 ( .A(a[86]), .B(n9895), .Z(n151) );
  IV U11858 ( .A(n9893), .Z(n9895) );
  XNOR U11859 ( .A(b[86]), .B(n9893), .Z(n9894) );
  XOR U11860 ( .A(n9896), .B(n9897), .Z(n9893) );
  ANDN U11861 ( .B(n9898), .A(n162), .Z(n9896) );
  XNOR U11862 ( .A(a[85]), .B(n9899), .Z(n162) );
  IV U11863 ( .A(n9897), .Z(n9899) );
  XNOR U11864 ( .A(b[85]), .B(n9897), .Z(n9898) );
  XOR U11865 ( .A(n9900), .B(n9901), .Z(n9897) );
  ANDN U11866 ( .B(n9902), .A(n173), .Z(n9900) );
  XNOR U11867 ( .A(a[84]), .B(n9903), .Z(n173) );
  IV U11868 ( .A(n9901), .Z(n9903) );
  XNOR U11869 ( .A(b[84]), .B(n9901), .Z(n9902) );
  XOR U11870 ( .A(n9904), .B(n9905), .Z(n9901) );
  ANDN U11871 ( .B(n9906), .A(n184), .Z(n9904) );
  XNOR U11872 ( .A(a[83]), .B(n9907), .Z(n184) );
  IV U11873 ( .A(n9905), .Z(n9907) );
  XNOR U11874 ( .A(b[83]), .B(n9905), .Z(n9906) );
  XOR U11875 ( .A(n9908), .B(n9909), .Z(n9905) );
  ANDN U11876 ( .B(n9910), .A(n195), .Z(n9908) );
  XNOR U11877 ( .A(a[82]), .B(n9911), .Z(n195) );
  IV U11878 ( .A(n9909), .Z(n9911) );
  XNOR U11879 ( .A(b[82]), .B(n9909), .Z(n9910) );
  XOR U11880 ( .A(n9912), .B(n9913), .Z(n9909) );
  ANDN U11881 ( .B(n9914), .A(n206), .Z(n9912) );
  XNOR U11882 ( .A(a[81]), .B(n9915), .Z(n206) );
  IV U11883 ( .A(n9913), .Z(n9915) );
  XNOR U11884 ( .A(b[81]), .B(n9913), .Z(n9914) );
  XOR U11885 ( .A(n9916), .B(n9917), .Z(n9913) );
  ANDN U11886 ( .B(n9918), .A(n217), .Z(n9916) );
  XNOR U11887 ( .A(a[80]), .B(n9919), .Z(n217) );
  IV U11888 ( .A(n9917), .Z(n9919) );
  XNOR U11889 ( .A(b[80]), .B(n9917), .Z(n9918) );
  XOR U11890 ( .A(n9920), .B(n9921), .Z(n9917) );
  ANDN U11891 ( .B(n9922), .A(n229), .Z(n9920) );
  XNOR U11892 ( .A(a[79]), .B(n9923), .Z(n229) );
  IV U11893 ( .A(n9921), .Z(n9923) );
  XNOR U11894 ( .A(b[79]), .B(n9921), .Z(n9922) );
  XOR U11895 ( .A(n9924), .B(n9925), .Z(n9921) );
  ANDN U11896 ( .B(n9926), .A(n240), .Z(n9924) );
  XNOR U11897 ( .A(a[78]), .B(n9927), .Z(n240) );
  IV U11898 ( .A(n9925), .Z(n9927) );
  XNOR U11899 ( .A(b[78]), .B(n9925), .Z(n9926) );
  XOR U11900 ( .A(n9928), .B(n9929), .Z(n9925) );
  ANDN U11901 ( .B(n9930), .A(n251), .Z(n9928) );
  XNOR U11902 ( .A(a[77]), .B(n9931), .Z(n251) );
  IV U11903 ( .A(n9929), .Z(n9931) );
  XNOR U11904 ( .A(b[77]), .B(n9929), .Z(n9930) );
  XOR U11905 ( .A(n9932), .B(n9933), .Z(n9929) );
  ANDN U11906 ( .B(n9934), .A(n262), .Z(n9932) );
  XNOR U11907 ( .A(a[76]), .B(n9935), .Z(n262) );
  IV U11908 ( .A(n9933), .Z(n9935) );
  XNOR U11909 ( .A(b[76]), .B(n9933), .Z(n9934) );
  XOR U11910 ( .A(n9936), .B(n9937), .Z(n9933) );
  ANDN U11911 ( .B(n9938), .A(n273), .Z(n9936) );
  XNOR U11912 ( .A(a[75]), .B(n9939), .Z(n273) );
  IV U11913 ( .A(n9937), .Z(n9939) );
  XNOR U11914 ( .A(b[75]), .B(n9937), .Z(n9938) );
  XOR U11915 ( .A(n9940), .B(n9941), .Z(n9937) );
  ANDN U11916 ( .B(n9942), .A(n284), .Z(n9940) );
  XNOR U11917 ( .A(a[74]), .B(n9943), .Z(n284) );
  IV U11918 ( .A(n9941), .Z(n9943) );
  XNOR U11919 ( .A(b[74]), .B(n9941), .Z(n9942) );
  XOR U11920 ( .A(n9944), .B(n9945), .Z(n9941) );
  ANDN U11921 ( .B(n9946), .A(n295), .Z(n9944) );
  XNOR U11922 ( .A(a[73]), .B(n9947), .Z(n295) );
  IV U11923 ( .A(n9945), .Z(n9947) );
  XNOR U11924 ( .A(b[73]), .B(n9945), .Z(n9946) );
  XOR U11925 ( .A(n9948), .B(n9949), .Z(n9945) );
  ANDN U11926 ( .B(n9950), .A(n306), .Z(n9948) );
  XNOR U11927 ( .A(a[72]), .B(n9951), .Z(n306) );
  IV U11928 ( .A(n9949), .Z(n9951) );
  XNOR U11929 ( .A(b[72]), .B(n9949), .Z(n9950) );
  XOR U11930 ( .A(n9952), .B(n9953), .Z(n9949) );
  ANDN U11931 ( .B(n9954), .A(n317), .Z(n9952) );
  XNOR U11932 ( .A(a[71]), .B(n9955), .Z(n317) );
  IV U11933 ( .A(n9953), .Z(n9955) );
  XNOR U11934 ( .A(b[71]), .B(n9953), .Z(n9954) );
  XOR U11935 ( .A(n9956), .B(n9957), .Z(n9953) );
  ANDN U11936 ( .B(n9958), .A(n328), .Z(n9956) );
  XNOR U11937 ( .A(a[70]), .B(n9959), .Z(n328) );
  IV U11938 ( .A(n9957), .Z(n9959) );
  XNOR U11939 ( .A(b[70]), .B(n9957), .Z(n9958) );
  XOR U11940 ( .A(n9960), .B(n9961), .Z(n9957) );
  ANDN U11941 ( .B(n9962), .A(n340), .Z(n9960) );
  XNOR U11942 ( .A(a[69]), .B(n9963), .Z(n340) );
  IV U11943 ( .A(n9961), .Z(n9963) );
  XNOR U11944 ( .A(b[69]), .B(n9961), .Z(n9962) );
  XOR U11945 ( .A(n9964), .B(n9965), .Z(n9961) );
  ANDN U11946 ( .B(n9966), .A(n351), .Z(n9964) );
  XNOR U11947 ( .A(a[68]), .B(n9967), .Z(n351) );
  IV U11948 ( .A(n9965), .Z(n9967) );
  XNOR U11949 ( .A(b[68]), .B(n9965), .Z(n9966) );
  XOR U11950 ( .A(n9968), .B(n9969), .Z(n9965) );
  ANDN U11951 ( .B(n9970), .A(n362), .Z(n9968) );
  XNOR U11952 ( .A(a[67]), .B(n9971), .Z(n362) );
  IV U11953 ( .A(n9969), .Z(n9971) );
  XNOR U11954 ( .A(b[67]), .B(n9969), .Z(n9970) );
  XOR U11955 ( .A(n9972), .B(n9973), .Z(n9969) );
  ANDN U11956 ( .B(n9974), .A(n373), .Z(n9972) );
  XNOR U11957 ( .A(a[66]), .B(n9975), .Z(n373) );
  IV U11958 ( .A(n9973), .Z(n9975) );
  XNOR U11959 ( .A(b[66]), .B(n9973), .Z(n9974) );
  XOR U11960 ( .A(n9976), .B(n9977), .Z(n9973) );
  ANDN U11961 ( .B(n9978), .A(n384), .Z(n9976) );
  XNOR U11962 ( .A(a[65]), .B(n9979), .Z(n384) );
  IV U11963 ( .A(n9977), .Z(n9979) );
  XNOR U11964 ( .A(b[65]), .B(n9977), .Z(n9978) );
  XOR U11965 ( .A(n9980), .B(n9981), .Z(n9977) );
  ANDN U11966 ( .B(n9982), .A(n395), .Z(n9980) );
  XNOR U11967 ( .A(a[64]), .B(n9983), .Z(n395) );
  IV U11968 ( .A(n9981), .Z(n9983) );
  XNOR U11969 ( .A(b[64]), .B(n9981), .Z(n9982) );
  XOR U11970 ( .A(n9984), .B(n9985), .Z(n9981) );
  ANDN U11971 ( .B(n9986), .A(n406), .Z(n9984) );
  XNOR U11972 ( .A(a[63]), .B(n9987), .Z(n406) );
  IV U11973 ( .A(n9985), .Z(n9987) );
  XNOR U11974 ( .A(b[63]), .B(n9985), .Z(n9986) );
  XOR U11975 ( .A(n9988), .B(n9989), .Z(n9985) );
  ANDN U11976 ( .B(n9990), .A(n417), .Z(n9988) );
  XNOR U11977 ( .A(a[62]), .B(n9991), .Z(n417) );
  IV U11978 ( .A(n9989), .Z(n9991) );
  XNOR U11979 ( .A(b[62]), .B(n9989), .Z(n9990) );
  XOR U11980 ( .A(n9992), .B(n9993), .Z(n9989) );
  ANDN U11981 ( .B(n9994), .A(n428), .Z(n9992) );
  XNOR U11982 ( .A(a[61]), .B(n9995), .Z(n428) );
  IV U11983 ( .A(n9993), .Z(n9995) );
  XNOR U11984 ( .A(b[61]), .B(n9993), .Z(n9994) );
  XOR U11985 ( .A(n9996), .B(n9997), .Z(n9993) );
  ANDN U11986 ( .B(n9998), .A(n439), .Z(n9996) );
  XNOR U11987 ( .A(a[60]), .B(n9999), .Z(n439) );
  IV U11988 ( .A(n9997), .Z(n9999) );
  XNOR U11989 ( .A(b[60]), .B(n9997), .Z(n9998) );
  XOR U11990 ( .A(n10000), .B(n10001), .Z(n9997) );
  ANDN U11991 ( .B(n10002), .A(n451), .Z(n10000) );
  XNOR U11992 ( .A(a[59]), .B(n10003), .Z(n451) );
  IV U11993 ( .A(n10001), .Z(n10003) );
  XNOR U11994 ( .A(b[59]), .B(n10001), .Z(n10002) );
  XOR U11995 ( .A(n10004), .B(n10005), .Z(n10001) );
  ANDN U11996 ( .B(n10006), .A(n462), .Z(n10004) );
  XNOR U11997 ( .A(a[58]), .B(n10007), .Z(n462) );
  IV U11998 ( .A(n10005), .Z(n10007) );
  XNOR U11999 ( .A(b[58]), .B(n10005), .Z(n10006) );
  XOR U12000 ( .A(n10008), .B(n10009), .Z(n10005) );
  ANDN U12001 ( .B(n10010), .A(n473), .Z(n10008) );
  XNOR U12002 ( .A(a[57]), .B(n10011), .Z(n473) );
  IV U12003 ( .A(n10009), .Z(n10011) );
  XNOR U12004 ( .A(b[57]), .B(n10009), .Z(n10010) );
  XOR U12005 ( .A(n10012), .B(n10013), .Z(n10009) );
  ANDN U12006 ( .B(n10014), .A(n484), .Z(n10012) );
  XNOR U12007 ( .A(a[56]), .B(n10015), .Z(n484) );
  IV U12008 ( .A(n10013), .Z(n10015) );
  XNOR U12009 ( .A(b[56]), .B(n10013), .Z(n10014) );
  XOR U12010 ( .A(n10016), .B(n10017), .Z(n10013) );
  ANDN U12011 ( .B(n10018), .A(n495), .Z(n10016) );
  XNOR U12012 ( .A(a[55]), .B(n10019), .Z(n495) );
  IV U12013 ( .A(n10017), .Z(n10019) );
  XNOR U12014 ( .A(b[55]), .B(n10017), .Z(n10018) );
  XOR U12015 ( .A(n10020), .B(n10021), .Z(n10017) );
  ANDN U12016 ( .B(n10022), .A(n506), .Z(n10020) );
  XNOR U12017 ( .A(a[54]), .B(n10023), .Z(n506) );
  IV U12018 ( .A(n10021), .Z(n10023) );
  XNOR U12019 ( .A(b[54]), .B(n10021), .Z(n10022) );
  XOR U12020 ( .A(n10024), .B(n10025), .Z(n10021) );
  ANDN U12021 ( .B(n10026), .A(n517), .Z(n10024) );
  XNOR U12022 ( .A(a[53]), .B(n10027), .Z(n517) );
  IV U12023 ( .A(n10025), .Z(n10027) );
  XNOR U12024 ( .A(b[53]), .B(n10025), .Z(n10026) );
  XOR U12025 ( .A(n10028), .B(n10029), .Z(n10025) );
  ANDN U12026 ( .B(n10030), .A(n528), .Z(n10028) );
  XNOR U12027 ( .A(a[52]), .B(n10031), .Z(n528) );
  IV U12028 ( .A(n10029), .Z(n10031) );
  XNOR U12029 ( .A(b[52]), .B(n10029), .Z(n10030) );
  XOR U12030 ( .A(n10032), .B(n10033), .Z(n10029) );
  ANDN U12031 ( .B(n10034), .A(n539), .Z(n10032) );
  XNOR U12032 ( .A(a[51]), .B(n10035), .Z(n539) );
  IV U12033 ( .A(n10033), .Z(n10035) );
  XNOR U12034 ( .A(b[51]), .B(n10033), .Z(n10034) );
  XOR U12035 ( .A(n10036), .B(n10037), .Z(n10033) );
  ANDN U12036 ( .B(n10038), .A(n550), .Z(n10036) );
  XNOR U12037 ( .A(a[50]), .B(n10039), .Z(n550) );
  IV U12038 ( .A(n10037), .Z(n10039) );
  XNOR U12039 ( .A(b[50]), .B(n10037), .Z(n10038) );
  XOR U12040 ( .A(n10040), .B(n10041), .Z(n10037) );
  ANDN U12041 ( .B(n10042), .A(n562), .Z(n10040) );
  XNOR U12042 ( .A(a[49]), .B(n10043), .Z(n562) );
  IV U12043 ( .A(n10041), .Z(n10043) );
  XNOR U12044 ( .A(b[49]), .B(n10041), .Z(n10042) );
  XOR U12045 ( .A(n10044), .B(n10045), .Z(n10041) );
  ANDN U12046 ( .B(n10046), .A(n573), .Z(n10044) );
  XNOR U12047 ( .A(a[48]), .B(n10047), .Z(n573) );
  IV U12048 ( .A(n10045), .Z(n10047) );
  XNOR U12049 ( .A(b[48]), .B(n10045), .Z(n10046) );
  XOR U12050 ( .A(n10048), .B(n10049), .Z(n10045) );
  ANDN U12051 ( .B(n10050), .A(n584), .Z(n10048) );
  XNOR U12052 ( .A(a[47]), .B(n10051), .Z(n584) );
  IV U12053 ( .A(n10049), .Z(n10051) );
  XNOR U12054 ( .A(b[47]), .B(n10049), .Z(n10050) );
  XOR U12055 ( .A(n10052), .B(n10053), .Z(n10049) );
  ANDN U12056 ( .B(n10054), .A(n595), .Z(n10052) );
  XNOR U12057 ( .A(a[46]), .B(n10055), .Z(n595) );
  IV U12058 ( .A(n10053), .Z(n10055) );
  XNOR U12059 ( .A(b[46]), .B(n10053), .Z(n10054) );
  XOR U12060 ( .A(n10056), .B(n10057), .Z(n10053) );
  ANDN U12061 ( .B(n10058), .A(n606), .Z(n10056) );
  XNOR U12062 ( .A(a[45]), .B(n10059), .Z(n606) );
  IV U12063 ( .A(n10057), .Z(n10059) );
  XNOR U12064 ( .A(b[45]), .B(n10057), .Z(n10058) );
  XOR U12065 ( .A(n10060), .B(n10061), .Z(n10057) );
  ANDN U12066 ( .B(n10062), .A(n617), .Z(n10060) );
  XNOR U12067 ( .A(a[44]), .B(n10063), .Z(n617) );
  IV U12068 ( .A(n10061), .Z(n10063) );
  XNOR U12069 ( .A(b[44]), .B(n10061), .Z(n10062) );
  XOR U12070 ( .A(n10064), .B(n10065), .Z(n10061) );
  ANDN U12071 ( .B(n10066), .A(n628), .Z(n10064) );
  XNOR U12072 ( .A(a[43]), .B(n10067), .Z(n628) );
  IV U12073 ( .A(n10065), .Z(n10067) );
  XNOR U12074 ( .A(b[43]), .B(n10065), .Z(n10066) );
  XOR U12075 ( .A(n10068), .B(n10069), .Z(n10065) );
  ANDN U12076 ( .B(n10070), .A(n639), .Z(n10068) );
  XNOR U12077 ( .A(a[42]), .B(n10071), .Z(n639) );
  IV U12078 ( .A(n10069), .Z(n10071) );
  XNOR U12079 ( .A(b[42]), .B(n10069), .Z(n10070) );
  XOR U12080 ( .A(n10072), .B(n10073), .Z(n10069) );
  ANDN U12081 ( .B(n10074), .A(n650), .Z(n10072) );
  XNOR U12082 ( .A(a[41]), .B(n10075), .Z(n650) );
  IV U12083 ( .A(n10073), .Z(n10075) );
  XNOR U12084 ( .A(b[41]), .B(n10073), .Z(n10074) );
  XOR U12085 ( .A(n10076), .B(n10077), .Z(n10073) );
  ANDN U12086 ( .B(n10078), .A(n661), .Z(n10076) );
  XNOR U12087 ( .A(a[40]), .B(n10079), .Z(n661) );
  IV U12088 ( .A(n10077), .Z(n10079) );
  XNOR U12089 ( .A(b[40]), .B(n10077), .Z(n10078) );
  XOR U12090 ( .A(n10080), .B(n10081), .Z(n10077) );
  ANDN U12091 ( .B(n10082), .A(n673), .Z(n10080) );
  XNOR U12092 ( .A(a[39]), .B(n10083), .Z(n673) );
  IV U12093 ( .A(n10081), .Z(n10083) );
  XNOR U12094 ( .A(b[39]), .B(n10081), .Z(n10082) );
  XOR U12095 ( .A(n10084), .B(n10085), .Z(n10081) );
  ANDN U12096 ( .B(n10086), .A(n684), .Z(n10084) );
  XNOR U12097 ( .A(a[38]), .B(n10087), .Z(n684) );
  IV U12098 ( .A(n10085), .Z(n10087) );
  XNOR U12099 ( .A(b[38]), .B(n10085), .Z(n10086) );
  XOR U12100 ( .A(n10088), .B(n10089), .Z(n10085) );
  ANDN U12101 ( .B(n10090), .A(n695), .Z(n10088) );
  XNOR U12102 ( .A(a[37]), .B(n10091), .Z(n695) );
  IV U12103 ( .A(n10089), .Z(n10091) );
  XNOR U12104 ( .A(b[37]), .B(n10089), .Z(n10090) );
  XOR U12105 ( .A(n10092), .B(n10093), .Z(n10089) );
  ANDN U12106 ( .B(n10094), .A(n706), .Z(n10092) );
  XNOR U12107 ( .A(a[36]), .B(n10095), .Z(n706) );
  IV U12108 ( .A(n10093), .Z(n10095) );
  XNOR U12109 ( .A(b[36]), .B(n10093), .Z(n10094) );
  XOR U12110 ( .A(n10096), .B(n10097), .Z(n10093) );
  ANDN U12111 ( .B(n10098), .A(n717), .Z(n10096) );
  XNOR U12112 ( .A(a[35]), .B(n10099), .Z(n717) );
  IV U12113 ( .A(n10097), .Z(n10099) );
  XNOR U12114 ( .A(b[35]), .B(n10097), .Z(n10098) );
  XOR U12115 ( .A(n10100), .B(n10101), .Z(n10097) );
  ANDN U12116 ( .B(n10102), .A(n728), .Z(n10100) );
  XNOR U12117 ( .A(a[34]), .B(n10103), .Z(n728) );
  IV U12118 ( .A(n10101), .Z(n10103) );
  XNOR U12119 ( .A(b[34]), .B(n10101), .Z(n10102) );
  XOR U12120 ( .A(n10104), .B(n10105), .Z(n10101) );
  ANDN U12121 ( .B(n10106), .A(n739), .Z(n10104) );
  XNOR U12122 ( .A(a[33]), .B(n10107), .Z(n739) );
  IV U12123 ( .A(n10105), .Z(n10107) );
  XNOR U12124 ( .A(b[33]), .B(n10105), .Z(n10106) );
  XOR U12125 ( .A(n10108), .B(n10109), .Z(n10105) );
  ANDN U12126 ( .B(n10110), .A(n750), .Z(n10108) );
  XNOR U12127 ( .A(a[32]), .B(n10111), .Z(n750) );
  IV U12128 ( .A(n10109), .Z(n10111) );
  XNOR U12129 ( .A(b[32]), .B(n10109), .Z(n10110) );
  XOR U12130 ( .A(n10112), .B(n10113), .Z(n10109) );
  ANDN U12131 ( .B(n10114), .A(n761), .Z(n10112) );
  XNOR U12132 ( .A(a[31]), .B(n10115), .Z(n761) );
  IV U12133 ( .A(n10113), .Z(n10115) );
  XNOR U12134 ( .A(b[31]), .B(n10113), .Z(n10114) );
  XOR U12135 ( .A(n10116), .B(n10117), .Z(n10113) );
  ANDN U12136 ( .B(n10118), .A(n772), .Z(n10116) );
  XNOR U12137 ( .A(a[30]), .B(n10119), .Z(n772) );
  IV U12138 ( .A(n10117), .Z(n10119) );
  XNOR U12139 ( .A(b[30]), .B(n10117), .Z(n10118) );
  XOR U12140 ( .A(n10120), .B(n10121), .Z(n10117) );
  ANDN U12141 ( .B(n10122), .A(n784), .Z(n10120) );
  XNOR U12142 ( .A(a[29]), .B(n10123), .Z(n784) );
  IV U12143 ( .A(n10121), .Z(n10123) );
  XNOR U12144 ( .A(b[29]), .B(n10121), .Z(n10122) );
  XOR U12145 ( .A(n10124), .B(n10125), .Z(n10121) );
  ANDN U12146 ( .B(n10126), .A(n795), .Z(n10124) );
  XNOR U12147 ( .A(a[28]), .B(n10127), .Z(n795) );
  IV U12148 ( .A(n10125), .Z(n10127) );
  XNOR U12149 ( .A(b[28]), .B(n10125), .Z(n10126) );
  XOR U12150 ( .A(n10128), .B(n10129), .Z(n10125) );
  ANDN U12151 ( .B(n10130), .A(n806), .Z(n10128) );
  XNOR U12152 ( .A(a[27]), .B(n10131), .Z(n806) );
  IV U12153 ( .A(n10129), .Z(n10131) );
  XNOR U12154 ( .A(b[27]), .B(n10129), .Z(n10130) );
  XOR U12155 ( .A(n10132), .B(n10133), .Z(n10129) );
  ANDN U12156 ( .B(n10134), .A(n817), .Z(n10132) );
  XNOR U12157 ( .A(a[26]), .B(n10135), .Z(n817) );
  IV U12158 ( .A(n10133), .Z(n10135) );
  XNOR U12159 ( .A(b[26]), .B(n10133), .Z(n10134) );
  XOR U12160 ( .A(n10136), .B(n10137), .Z(n10133) );
  ANDN U12161 ( .B(n10138), .A(n828), .Z(n10136) );
  XNOR U12162 ( .A(a[25]), .B(n10139), .Z(n828) );
  IV U12163 ( .A(n10137), .Z(n10139) );
  XNOR U12164 ( .A(b[25]), .B(n10137), .Z(n10138) );
  XOR U12165 ( .A(n10140), .B(n10141), .Z(n10137) );
  ANDN U12166 ( .B(n10142), .A(n839), .Z(n10140) );
  XNOR U12167 ( .A(a[24]), .B(n10143), .Z(n839) );
  IV U12168 ( .A(n10141), .Z(n10143) );
  XNOR U12169 ( .A(b[24]), .B(n10141), .Z(n10142) );
  XOR U12170 ( .A(n10144), .B(n10145), .Z(n10141) );
  ANDN U12171 ( .B(n10146), .A(n850), .Z(n10144) );
  XNOR U12172 ( .A(a[23]), .B(n10147), .Z(n850) );
  IV U12173 ( .A(n10145), .Z(n10147) );
  XNOR U12174 ( .A(b[23]), .B(n10145), .Z(n10146) );
  XOR U12175 ( .A(n10148), .B(n10149), .Z(n10145) );
  ANDN U12176 ( .B(n10150), .A(n861), .Z(n10148) );
  XNOR U12177 ( .A(a[22]), .B(n10151), .Z(n861) );
  IV U12178 ( .A(n10149), .Z(n10151) );
  XNOR U12179 ( .A(b[22]), .B(n10149), .Z(n10150) );
  XOR U12180 ( .A(n10152), .B(n10153), .Z(n10149) );
  ANDN U12181 ( .B(n10154), .A(n872), .Z(n10152) );
  XNOR U12182 ( .A(a[21]), .B(n10155), .Z(n872) );
  IV U12183 ( .A(n10153), .Z(n10155) );
  XNOR U12184 ( .A(b[21]), .B(n10153), .Z(n10154) );
  XOR U12185 ( .A(n10156), .B(n10157), .Z(n10153) );
  ANDN U12186 ( .B(n10158), .A(n883), .Z(n10156) );
  XNOR U12187 ( .A(a[20]), .B(n10159), .Z(n883) );
  IV U12188 ( .A(n10157), .Z(n10159) );
  XNOR U12189 ( .A(b[20]), .B(n10157), .Z(n10158) );
  XOR U12190 ( .A(n10160), .B(n10161), .Z(n10157) );
  ANDN U12191 ( .B(n10162), .A(n1134), .Z(n10160) );
  XNOR U12192 ( .A(a[19]), .B(n10163), .Z(n1134) );
  IV U12193 ( .A(n10161), .Z(n10163) );
  XNOR U12194 ( .A(b[19]), .B(n10161), .Z(n10162) );
  XOR U12195 ( .A(n10164), .B(n10165), .Z(n10161) );
  ANDN U12196 ( .B(n10166), .A(n1645), .Z(n10164) );
  XNOR U12197 ( .A(a[18]), .B(n10167), .Z(n1645) );
  IV U12198 ( .A(n10165), .Z(n10167) );
  XNOR U12199 ( .A(b[18]), .B(n10165), .Z(n10166) );
  XOR U12200 ( .A(n10168), .B(n10169), .Z(n10165) );
  ANDN U12201 ( .B(n10170), .A(n2156), .Z(n10168) );
  XNOR U12202 ( .A(a[17]), .B(n10171), .Z(n2156) );
  IV U12203 ( .A(n10169), .Z(n10171) );
  XNOR U12204 ( .A(b[17]), .B(n10169), .Z(n10170) );
  XOR U12205 ( .A(n10172), .B(n10173), .Z(n10169) );
  ANDN U12206 ( .B(n10174), .A(n2667), .Z(n10172) );
  XNOR U12207 ( .A(a[16]), .B(n10175), .Z(n2667) );
  IV U12208 ( .A(n10173), .Z(n10175) );
  XNOR U12209 ( .A(b[16]), .B(n10173), .Z(n10174) );
  XOR U12210 ( .A(n10176), .B(n10177), .Z(n10173) );
  ANDN U12211 ( .B(n10178), .A(n3178), .Z(n10176) );
  XNOR U12212 ( .A(a[15]), .B(n10179), .Z(n3178) );
  IV U12213 ( .A(n10177), .Z(n10179) );
  XNOR U12214 ( .A(b[15]), .B(n10177), .Z(n10178) );
  XOR U12215 ( .A(n10180), .B(n10181), .Z(n10177) );
  ANDN U12216 ( .B(n10182), .A(n3689), .Z(n10180) );
  XNOR U12217 ( .A(a[14]), .B(n10183), .Z(n3689) );
  IV U12218 ( .A(n10181), .Z(n10183) );
  XNOR U12219 ( .A(b[14]), .B(n10181), .Z(n10182) );
  XOR U12220 ( .A(n10184), .B(n10185), .Z(n10181) );
  ANDN U12221 ( .B(n10186), .A(n4200), .Z(n10184) );
  XNOR U12222 ( .A(a[13]), .B(n10187), .Z(n4200) );
  IV U12223 ( .A(n10185), .Z(n10187) );
  XNOR U12224 ( .A(b[13]), .B(n10185), .Z(n10186) );
  XOR U12225 ( .A(n10188), .B(n10189), .Z(n10185) );
  ANDN U12226 ( .B(n10190), .A(n4711), .Z(n10188) );
  XNOR U12227 ( .A(a[12]), .B(n10191), .Z(n4711) );
  IV U12228 ( .A(n10189), .Z(n10191) );
  XNOR U12229 ( .A(b[12]), .B(n10189), .Z(n10190) );
  XOR U12230 ( .A(n10192), .B(n10193), .Z(n10189) );
  ANDN U12231 ( .B(n10194), .A(n5222), .Z(n10192) );
  XNOR U12232 ( .A(a[11]), .B(n10195), .Z(n5222) );
  IV U12233 ( .A(n10193), .Z(n10195) );
  XNOR U12234 ( .A(b[11]), .B(n10193), .Z(n10194) );
  XOR U12235 ( .A(n10196), .B(n10197), .Z(n10193) );
  ANDN U12236 ( .B(n10198), .A(n5733), .Z(n10196) );
  XNOR U12237 ( .A(a[10]), .B(n10199), .Z(n5733) );
  IV U12238 ( .A(n10197), .Z(n10199) );
  XNOR U12239 ( .A(b[10]), .B(n10197), .Z(n10198) );
  XOR U12240 ( .A(n10200), .B(n10201), .Z(n10197) );
  ANDN U12241 ( .B(n10202), .A(n6), .Z(n10200) );
  XNOR U12242 ( .A(a[9]), .B(n10203), .Z(n6) );
  IV U12243 ( .A(n10201), .Z(n10203) );
  XNOR U12244 ( .A(b[9]), .B(n10201), .Z(n10202) );
  XOR U12245 ( .A(n10204), .B(n10205), .Z(n10201) );
  ANDN U12246 ( .B(n10206), .A(n117), .Z(n10204) );
  XNOR U12247 ( .A(a[8]), .B(n10207), .Z(n117) );
  IV U12248 ( .A(n10205), .Z(n10207) );
  XNOR U12249 ( .A(b[8]), .B(n10205), .Z(n10206) );
  XOR U12250 ( .A(n10208), .B(n10209), .Z(n10205) );
  ANDN U12251 ( .B(n10210), .A(n228), .Z(n10208) );
  XNOR U12252 ( .A(a[7]), .B(n10211), .Z(n228) );
  IV U12253 ( .A(n10209), .Z(n10211) );
  XNOR U12254 ( .A(b[7]), .B(n10209), .Z(n10210) );
  XOR U12255 ( .A(n10212), .B(n10213), .Z(n10209) );
  ANDN U12256 ( .B(n10214), .A(n339), .Z(n10212) );
  XNOR U12257 ( .A(a[6]), .B(n10215), .Z(n339) );
  IV U12258 ( .A(n10213), .Z(n10215) );
  XNOR U12259 ( .A(b[6]), .B(n10213), .Z(n10214) );
  XOR U12260 ( .A(n10216), .B(n10217), .Z(n10213) );
  ANDN U12261 ( .B(n10218), .A(n450), .Z(n10216) );
  XNOR U12262 ( .A(a[5]), .B(n10219), .Z(n450) );
  IV U12263 ( .A(n10217), .Z(n10219) );
  XNOR U12264 ( .A(b[5]), .B(n10217), .Z(n10218) );
  XOR U12265 ( .A(n10220), .B(n10221), .Z(n10217) );
  ANDN U12266 ( .B(n10222), .A(n561), .Z(n10220) );
  XNOR U12267 ( .A(a[4]), .B(n10223), .Z(n561) );
  IV U12268 ( .A(n10221), .Z(n10223) );
  XNOR U12269 ( .A(b[4]), .B(n10221), .Z(n10222) );
  XOR U12270 ( .A(n10224), .B(n10225), .Z(n10221) );
  ANDN U12271 ( .B(n10226), .A(n672), .Z(n10224) );
  XNOR U12272 ( .A(a[3]), .B(n10227), .Z(n672) );
  IV U12273 ( .A(n10225), .Z(n10227) );
  XNOR U12274 ( .A(b[3]), .B(n10225), .Z(n10226) );
  XOR U12275 ( .A(n10228), .B(n10229), .Z(n10225) );
  ANDN U12276 ( .B(n10230), .A(n783), .Z(n10228) );
  XNOR U12277 ( .A(a[2]), .B(n10231), .Z(n783) );
  IV U12278 ( .A(n10229), .Z(n10231) );
  XNOR U12279 ( .A(b[2]), .B(n10229), .Z(n10230) );
  XOR U12280 ( .A(n10232), .B(n10233), .Z(n10229) );
  ANDN U12281 ( .B(n10234), .A(n1133), .Z(n10232) );
  XNOR U12282 ( .A(a[1]), .B(n10235), .Z(n1133) );
  IV U12283 ( .A(n10233), .Z(n10235) );
  XNOR U12284 ( .A(b[1]), .B(n10233), .Z(n10234) );
  XOR U12285 ( .A(carry_on), .B(n10236), .Z(n10233) );
  NANDN U12286 ( .A(n10237), .B(n10238), .Z(n10236) );
  XOR U12287 ( .A(carry_on), .B(b[0]), .Z(n10238) );
  XNOR U12288 ( .A(b[0]), .B(n10237), .Z(c[0]) );
  XNOR U12289 ( .A(a[0]), .B(carry_on), .Z(n10237) );
endmodule

