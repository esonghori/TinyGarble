
module aes_seq_CC2 ( clk, rst, msg, key, out );
  input [127:0] msg;
  input [639:0] key;
  output [127:0] out;
  input clk, rst;
  wire   \w0[4][127] , \w0[4][126] , \w0[4][125] , \w0[4][124] , \w0[4][123] ,
         \w0[4][122] , \w0[4][121] , \w0[4][120] , \w0[4][119] , \w0[4][118] ,
         \w0[4][117] , \w0[4][116] , \w0[4][115] , \w0[4][114] , \w0[4][113] ,
         \w0[4][112] , \w0[4][111] , \w0[4][110] , \w0[4][109] , \w0[4][108] ,
         \w0[4][107] , \w0[4][106] , \w0[4][105] , \w0[4][104] , \w0[4][103] ,
         \w0[4][102] , \w0[4][101] , \w0[4][100] , \w0[4][99] , \w0[4][98] ,
         \w0[4][97] , \w0[4][96] , \w0[4][95] , \w0[4][94] , \w0[4][93] ,
         \w0[4][92] , \w0[4][91] , \w0[4][90] , \w0[4][89] , \w0[4][88] ,
         \w0[4][87] , \w0[4][86] , \w0[4][85] , \w0[4][84] , \w0[4][83] ,
         \w0[4][82] , \w0[4][81] , \w0[4][80] , \w0[4][79] , \w0[4][78] ,
         \w0[4][77] , \w0[4][76] , \w0[4][75] , \w0[4][74] , \w0[4][73] ,
         \w0[4][72] , \w0[4][71] , \w0[4][70] , \w0[4][69] , \w0[4][68] ,
         \w0[4][67] , \w0[4][66] , \w0[4][65] , \w0[4][64] , \w0[4][63] ,
         \w0[4][62] , \w0[4][61] , \w0[4][60] , \w0[4][59] , \w0[4][58] ,
         \w0[4][57] , \w0[4][56] , \w0[4][55] , \w0[4][54] , \w0[4][53] ,
         \w0[4][52] , \w0[4][51] , \w0[4][50] , \w0[4][49] , \w0[4][48] ,
         \w0[4][47] , \w0[4][46] , \w0[4][45] , \w0[4][44] , \w0[4][43] ,
         \w0[4][42] , \w0[4][41] , \w0[4][40] , \w0[4][39] , \w0[4][38] ,
         \w0[4][37] , \w0[4][36] , \w0[4][35] , \w0[4][34] , \w0[4][33] ,
         \w0[4][32] , \w0[4][31] , \w0[4][30] , \w0[4][29] , \w0[4][28] ,
         \w0[4][27] , \w0[4][26] , \w0[4][25] , \w0[4][24] , \w0[4][23] ,
         \w0[4][22] , \w0[4][21] , \w0[4][20] , \w0[4][19] , \w0[4][18] ,
         \w0[4][17] , \w0[4][16] , \w0[4][15] , \w0[4][14] , \w0[4][13] ,
         \w0[4][12] , \w0[4][11] , \w0[4][10] , \w0[4][9] , \w0[4][8] ,
         \w0[4][7] , \w0[4][6] , \w0[4][5] , \w0[4][4] , \w0[4][3] ,
         \w0[4][2] , \w0[4][1] , \w0[4][0] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474;
  wire   [127:0] state;

  DFF \state_reg[0]  ( .D(\w0[4][0] ), .CLK(clk), .RST(rst), .I(msg[0]), .Q(
        state[0]) );
  DFF \state_reg[1]  ( .D(\w0[4][1] ), .CLK(clk), .RST(rst), .I(msg[1]), .Q(
        state[1]) );
  DFF \state_reg[2]  ( .D(\w0[4][2] ), .CLK(clk), .RST(rst), .I(msg[2]), .Q(
        state[2]) );
  DFF \state_reg[3]  ( .D(\w0[4][3] ), .CLK(clk), .RST(rst), .I(msg[3]), .Q(
        state[3]) );
  DFF \state_reg[4]  ( .D(\w0[4][4] ), .CLK(clk), .RST(rst), .I(msg[4]), .Q(
        state[4]) );
  DFF \state_reg[5]  ( .D(\w0[4][5] ), .CLK(clk), .RST(rst), .I(msg[5]), .Q(
        state[5]) );
  DFF \state_reg[6]  ( .D(\w0[4][6] ), .CLK(clk), .RST(rst), .I(msg[6]), .Q(
        state[6]) );
  DFF \state_reg[7]  ( .D(\w0[4][7] ), .CLK(clk), .RST(rst), .I(msg[7]), .Q(
        state[7]) );
  DFF \state_reg[8]  ( .D(\w0[4][8] ), .CLK(clk), .RST(rst), .I(msg[8]), .Q(
        state[8]) );
  DFF \state_reg[9]  ( .D(\w0[4][9] ), .CLK(clk), .RST(rst), .I(msg[9]), .Q(
        state[9]) );
  DFF \state_reg[10]  ( .D(\w0[4][10] ), .CLK(clk), .RST(rst), .I(msg[10]), 
        .Q(state[10]) );
  DFF \state_reg[11]  ( .D(\w0[4][11] ), .CLK(clk), .RST(rst), .I(msg[11]), 
        .Q(state[11]) );
  DFF \state_reg[12]  ( .D(\w0[4][12] ), .CLK(clk), .RST(rst), .I(msg[12]), 
        .Q(state[12]) );
  DFF \state_reg[13]  ( .D(\w0[4][13] ), .CLK(clk), .RST(rst), .I(msg[13]), 
        .Q(state[13]) );
  DFF \state_reg[14]  ( .D(\w0[4][14] ), .CLK(clk), .RST(rst), .I(msg[14]), 
        .Q(state[14]) );
  DFF \state_reg[15]  ( .D(\w0[4][15] ), .CLK(clk), .RST(rst), .I(msg[15]), 
        .Q(state[15]) );
  DFF \state_reg[16]  ( .D(\w0[4][16] ), .CLK(clk), .RST(rst), .I(msg[16]), 
        .Q(state[16]) );
  DFF \state_reg[17]  ( .D(\w0[4][17] ), .CLK(clk), .RST(rst), .I(msg[17]), 
        .Q(state[17]) );
  DFF \state_reg[18]  ( .D(\w0[4][18] ), .CLK(clk), .RST(rst), .I(msg[18]), 
        .Q(state[18]) );
  DFF \state_reg[19]  ( .D(\w0[4][19] ), .CLK(clk), .RST(rst), .I(msg[19]), 
        .Q(state[19]) );
  DFF \state_reg[20]  ( .D(\w0[4][20] ), .CLK(clk), .RST(rst), .I(msg[20]), 
        .Q(state[20]) );
  DFF \state_reg[21]  ( .D(\w0[4][21] ), .CLK(clk), .RST(rst), .I(msg[21]), 
        .Q(state[21]) );
  DFF \state_reg[22]  ( .D(\w0[4][22] ), .CLK(clk), .RST(rst), .I(msg[22]), 
        .Q(state[22]) );
  DFF \state_reg[23]  ( .D(\w0[4][23] ), .CLK(clk), .RST(rst), .I(msg[23]), 
        .Q(state[23]) );
  DFF \state_reg[24]  ( .D(\w0[4][24] ), .CLK(clk), .RST(rst), .I(msg[24]), 
        .Q(state[24]) );
  DFF \state_reg[25]  ( .D(\w0[4][25] ), .CLK(clk), .RST(rst), .I(msg[25]), 
        .Q(state[25]) );
  DFF \state_reg[26]  ( .D(\w0[4][26] ), .CLK(clk), .RST(rst), .I(msg[26]), 
        .Q(state[26]) );
  DFF \state_reg[27]  ( .D(\w0[4][27] ), .CLK(clk), .RST(rst), .I(msg[27]), 
        .Q(state[27]) );
  DFF \state_reg[28]  ( .D(\w0[4][28] ), .CLK(clk), .RST(rst), .I(msg[28]), 
        .Q(state[28]) );
  DFF \state_reg[29]  ( .D(\w0[4][29] ), .CLK(clk), .RST(rst), .I(msg[29]), 
        .Q(state[29]) );
  DFF \state_reg[30]  ( .D(\w0[4][30] ), .CLK(clk), .RST(rst), .I(msg[30]), 
        .Q(state[30]) );
  DFF \state_reg[31]  ( .D(\w0[4][31] ), .CLK(clk), .RST(rst), .I(msg[31]), 
        .Q(state[31]) );
  DFF \state_reg[32]  ( .D(\w0[4][32] ), .CLK(clk), .RST(rst), .I(msg[32]), 
        .Q(state[32]) );
  DFF \state_reg[33]  ( .D(\w0[4][33] ), .CLK(clk), .RST(rst), .I(msg[33]), 
        .Q(state[33]) );
  DFF \state_reg[34]  ( .D(\w0[4][34] ), .CLK(clk), .RST(rst), .I(msg[34]), 
        .Q(state[34]) );
  DFF \state_reg[35]  ( .D(\w0[4][35] ), .CLK(clk), .RST(rst), .I(msg[35]), 
        .Q(state[35]) );
  DFF \state_reg[36]  ( .D(\w0[4][36] ), .CLK(clk), .RST(rst), .I(msg[36]), 
        .Q(state[36]) );
  DFF \state_reg[37]  ( .D(\w0[4][37] ), .CLK(clk), .RST(rst), .I(msg[37]), 
        .Q(state[37]) );
  DFF \state_reg[38]  ( .D(\w0[4][38] ), .CLK(clk), .RST(rst), .I(msg[38]), 
        .Q(state[38]) );
  DFF \state_reg[39]  ( .D(\w0[4][39] ), .CLK(clk), .RST(rst), .I(msg[39]), 
        .Q(state[39]) );
  DFF \state_reg[40]  ( .D(\w0[4][40] ), .CLK(clk), .RST(rst), .I(msg[40]), 
        .Q(state[40]) );
  DFF \state_reg[41]  ( .D(\w0[4][41] ), .CLK(clk), .RST(rst), .I(msg[41]), 
        .Q(state[41]) );
  DFF \state_reg[42]  ( .D(\w0[4][42] ), .CLK(clk), .RST(rst), .I(msg[42]), 
        .Q(state[42]) );
  DFF \state_reg[43]  ( .D(\w0[4][43] ), .CLK(clk), .RST(rst), .I(msg[43]), 
        .Q(state[43]) );
  DFF \state_reg[44]  ( .D(\w0[4][44] ), .CLK(clk), .RST(rst), .I(msg[44]), 
        .Q(state[44]) );
  DFF \state_reg[45]  ( .D(\w0[4][45] ), .CLK(clk), .RST(rst), .I(msg[45]), 
        .Q(state[45]) );
  DFF \state_reg[46]  ( .D(\w0[4][46] ), .CLK(clk), .RST(rst), .I(msg[46]), 
        .Q(state[46]) );
  DFF \state_reg[47]  ( .D(\w0[4][47] ), .CLK(clk), .RST(rst), .I(msg[47]), 
        .Q(state[47]) );
  DFF \state_reg[48]  ( .D(\w0[4][48] ), .CLK(clk), .RST(rst), .I(msg[48]), 
        .Q(state[48]) );
  DFF \state_reg[49]  ( .D(\w0[4][49] ), .CLK(clk), .RST(rst), .I(msg[49]), 
        .Q(state[49]) );
  DFF \state_reg[50]  ( .D(\w0[4][50] ), .CLK(clk), .RST(rst), .I(msg[50]), 
        .Q(state[50]) );
  DFF \state_reg[51]  ( .D(\w0[4][51] ), .CLK(clk), .RST(rst), .I(msg[51]), 
        .Q(state[51]) );
  DFF \state_reg[52]  ( .D(\w0[4][52] ), .CLK(clk), .RST(rst), .I(msg[52]), 
        .Q(state[52]) );
  DFF \state_reg[53]  ( .D(\w0[4][53] ), .CLK(clk), .RST(rst), .I(msg[53]), 
        .Q(state[53]) );
  DFF \state_reg[54]  ( .D(\w0[4][54] ), .CLK(clk), .RST(rst), .I(msg[54]), 
        .Q(state[54]) );
  DFF \state_reg[55]  ( .D(\w0[4][55] ), .CLK(clk), .RST(rst), .I(msg[55]), 
        .Q(state[55]) );
  DFF \state_reg[56]  ( .D(\w0[4][56] ), .CLK(clk), .RST(rst), .I(msg[56]), 
        .Q(state[56]) );
  DFF \state_reg[57]  ( .D(\w0[4][57] ), .CLK(clk), .RST(rst), .I(msg[57]), 
        .Q(state[57]) );
  DFF \state_reg[58]  ( .D(\w0[4][58] ), .CLK(clk), .RST(rst), .I(msg[58]), 
        .Q(state[58]) );
  DFF \state_reg[59]  ( .D(\w0[4][59] ), .CLK(clk), .RST(rst), .I(msg[59]), 
        .Q(state[59]) );
  DFF \state_reg[60]  ( .D(\w0[4][60] ), .CLK(clk), .RST(rst), .I(msg[60]), 
        .Q(state[60]) );
  DFF \state_reg[61]  ( .D(\w0[4][61] ), .CLK(clk), .RST(rst), .I(msg[61]), 
        .Q(state[61]) );
  DFF \state_reg[62]  ( .D(\w0[4][62] ), .CLK(clk), .RST(rst), .I(msg[62]), 
        .Q(state[62]) );
  DFF \state_reg[63]  ( .D(\w0[4][63] ), .CLK(clk), .RST(rst), .I(msg[63]), 
        .Q(state[63]) );
  DFF \state_reg[64]  ( .D(\w0[4][64] ), .CLK(clk), .RST(rst), .I(msg[64]), 
        .Q(state[64]) );
  DFF \state_reg[65]  ( .D(\w0[4][65] ), .CLK(clk), .RST(rst), .I(msg[65]), 
        .Q(state[65]) );
  DFF \state_reg[66]  ( .D(\w0[4][66] ), .CLK(clk), .RST(rst), .I(msg[66]), 
        .Q(state[66]) );
  DFF \state_reg[67]  ( .D(\w0[4][67] ), .CLK(clk), .RST(rst), .I(msg[67]), 
        .Q(state[67]) );
  DFF \state_reg[68]  ( .D(\w0[4][68] ), .CLK(clk), .RST(rst), .I(msg[68]), 
        .Q(state[68]) );
  DFF \state_reg[69]  ( .D(\w0[4][69] ), .CLK(clk), .RST(rst), .I(msg[69]), 
        .Q(state[69]) );
  DFF \state_reg[70]  ( .D(\w0[4][70] ), .CLK(clk), .RST(rst), .I(msg[70]), 
        .Q(state[70]) );
  DFF \state_reg[71]  ( .D(\w0[4][71] ), .CLK(clk), .RST(rst), .I(msg[71]), 
        .Q(state[71]) );
  DFF \state_reg[72]  ( .D(\w0[4][72] ), .CLK(clk), .RST(rst), .I(msg[72]), 
        .Q(state[72]) );
  DFF \state_reg[73]  ( .D(\w0[4][73] ), .CLK(clk), .RST(rst), .I(msg[73]), 
        .Q(state[73]) );
  DFF \state_reg[74]  ( .D(\w0[4][74] ), .CLK(clk), .RST(rst), .I(msg[74]), 
        .Q(state[74]) );
  DFF \state_reg[75]  ( .D(\w0[4][75] ), .CLK(clk), .RST(rst), .I(msg[75]), 
        .Q(state[75]) );
  DFF \state_reg[76]  ( .D(\w0[4][76] ), .CLK(clk), .RST(rst), .I(msg[76]), 
        .Q(state[76]) );
  DFF \state_reg[77]  ( .D(\w0[4][77] ), .CLK(clk), .RST(rst), .I(msg[77]), 
        .Q(state[77]) );
  DFF \state_reg[78]  ( .D(\w0[4][78] ), .CLK(clk), .RST(rst), .I(msg[78]), 
        .Q(state[78]) );
  DFF \state_reg[79]  ( .D(\w0[4][79] ), .CLK(clk), .RST(rst), .I(msg[79]), 
        .Q(state[79]) );
  DFF \state_reg[80]  ( .D(\w0[4][80] ), .CLK(clk), .RST(rst), .I(msg[80]), 
        .Q(state[80]) );
  DFF \state_reg[81]  ( .D(\w0[4][81] ), .CLK(clk), .RST(rst), .I(msg[81]), 
        .Q(state[81]) );
  DFF \state_reg[82]  ( .D(\w0[4][82] ), .CLK(clk), .RST(rst), .I(msg[82]), 
        .Q(state[82]) );
  DFF \state_reg[83]  ( .D(\w0[4][83] ), .CLK(clk), .RST(rst), .I(msg[83]), 
        .Q(state[83]) );
  DFF \state_reg[84]  ( .D(\w0[4][84] ), .CLK(clk), .RST(rst), .I(msg[84]), 
        .Q(state[84]) );
  DFF \state_reg[85]  ( .D(\w0[4][85] ), .CLK(clk), .RST(rst), .I(msg[85]), 
        .Q(state[85]) );
  DFF \state_reg[86]  ( .D(\w0[4][86] ), .CLK(clk), .RST(rst), .I(msg[86]), 
        .Q(state[86]) );
  DFF \state_reg[87]  ( .D(\w0[4][87] ), .CLK(clk), .RST(rst), .I(msg[87]), 
        .Q(state[87]) );
  DFF \state_reg[88]  ( .D(\w0[4][88] ), .CLK(clk), .RST(rst), .I(msg[88]), 
        .Q(state[88]) );
  DFF \state_reg[89]  ( .D(\w0[4][89] ), .CLK(clk), .RST(rst), .I(msg[89]), 
        .Q(state[89]) );
  DFF \state_reg[90]  ( .D(\w0[4][90] ), .CLK(clk), .RST(rst), .I(msg[90]), 
        .Q(state[90]) );
  DFF \state_reg[91]  ( .D(\w0[4][91] ), .CLK(clk), .RST(rst), .I(msg[91]), 
        .Q(state[91]) );
  DFF \state_reg[92]  ( .D(\w0[4][92] ), .CLK(clk), .RST(rst), .I(msg[92]), 
        .Q(state[92]) );
  DFF \state_reg[93]  ( .D(\w0[4][93] ), .CLK(clk), .RST(rst), .I(msg[93]), 
        .Q(state[93]) );
  DFF \state_reg[94]  ( .D(\w0[4][94] ), .CLK(clk), .RST(rst), .I(msg[94]), 
        .Q(state[94]) );
  DFF \state_reg[95]  ( .D(\w0[4][95] ), .CLK(clk), .RST(rst), .I(msg[95]), 
        .Q(state[95]) );
  DFF \state_reg[96]  ( .D(\w0[4][96] ), .CLK(clk), .RST(rst), .I(msg[96]), 
        .Q(state[96]) );
  DFF \state_reg[97]  ( .D(\w0[4][97] ), .CLK(clk), .RST(rst), .I(msg[97]), 
        .Q(state[97]) );
  DFF \state_reg[98]  ( .D(\w0[4][98] ), .CLK(clk), .RST(rst), .I(msg[98]), 
        .Q(state[98]) );
  DFF \state_reg[99]  ( .D(\w0[4][99] ), .CLK(clk), .RST(rst), .I(msg[99]), 
        .Q(state[99]) );
  DFF \state_reg[100]  ( .D(\w0[4][100] ), .CLK(clk), .RST(rst), .I(msg[100]), 
        .Q(state[100]) );
  DFF \state_reg[101]  ( .D(\w0[4][101] ), .CLK(clk), .RST(rst), .I(msg[101]), 
        .Q(state[101]) );
  DFF \state_reg[102]  ( .D(\w0[4][102] ), .CLK(clk), .RST(rst), .I(msg[102]), 
        .Q(state[102]) );
  DFF \state_reg[103]  ( .D(\w0[4][103] ), .CLK(clk), .RST(rst), .I(msg[103]), 
        .Q(state[103]) );
  DFF \state_reg[104]  ( .D(\w0[4][104] ), .CLK(clk), .RST(rst), .I(msg[104]), 
        .Q(state[104]) );
  DFF \state_reg[105]  ( .D(\w0[4][105] ), .CLK(clk), .RST(rst), .I(msg[105]), 
        .Q(state[105]) );
  DFF \state_reg[106]  ( .D(\w0[4][106] ), .CLK(clk), .RST(rst), .I(msg[106]), 
        .Q(state[106]) );
  DFF \state_reg[107]  ( .D(\w0[4][107] ), .CLK(clk), .RST(rst), .I(msg[107]), 
        .Q(state[107]) );
  DFF \state_reg[108]  ( .D(\w0[4][108] ), .CLK(clk), .RST(rst), .I(msg[108]), 
        .Q(state[108]) );
  DFF \state_reg[109]  ( .D(\w0[4][109] ), .CLK(clk), .RST(rst), .I(msg[109]), 
        .Q(state[109]) );
  DFF \state_reg[110]  ( .D(\w0[4][110] ), .CLK(clk), .RST(rst), .I(msg[110]), 
        .Q(state[110]) );
  DFF \state_reg[111]  ( .D(\w0[4][111] ), .CLK(clk), .RST(rst), .I(msg[111]), 
        .Q(state[111]) );
  DFF \state_reg[112]  ( .D(\w0[4][112] ), .CLK(clk), .RST(rst), .I(msg[112]), 
        .Q(state[112]) );
  DFF \state_reg[113]  ( .D(\w0[4][113] ), .CLK(clk), .RST(rst), .I(msg[113]), 
        .Q(state[113]) );
  DFF \state_reg[114]  ( .D(\w0[4][114] ), .CLK(clk), .RST(rst), .I(msg[114]), 
        .Q(state[114]) );
  DFF \state_reg[115]  ( .D(\w0[4][115] ), .CLK(clk), .RST(rst), .I(msg[115]), 
        .Q(state[115]) );
  DFF \state_reg[116]  ( .D(\w0[4][116] ), .CLK(clk), .RST(rst), .I(msg[116]), 
        .Q(state[116]) );
  DFF \state_reg[117]  ( .D(\w0[4][117] ), .CLK(clk), .RST(rst), .I(msg[117]), 
        .Q(state[117]) );
  DFF \state_reg[118]  ( .D(\w0[4][118] ), .CLK(clk), .RST(rst), .I(msg[118]), 
        .Q(state[118]) );
  DFF \state_reg[119]  ( .D(\w0[4][119] ), .CLK(clk), .RST(rst), .I(msg[119]), 
        .Q(state[119]) );
  DFF \state_reg[120]  ( .D(\w0[4][120] ), .CLK(clk), .RST(rst), .I(msg[120]), 
        .Q(state[120]) );
  DFF \state_reg[121]  ( .D(\w0[4][121] ), .CLK(clk), .RST(rst), .I(msg[121]), 
        .Q(state[121]) );
  DFF \state_reg[122]  ( .D(\w0[4][122] ), .CLK(clk), .RST(rst), .I(msg[122]), 
        .Q(state[122]) );
  DFF \state_reg[123]  ( .D(\w0[4][123] ), .CLK(clk), .RST(rst), .I(msg[123]), 
        .Q(state[123]) );
  DFF \state_reg[124]  ( .D(\w0[4][124] ), .CLK(clk), .RST(rst), .I(msg[124]), 
        .Q(state[124]) );
  DFF \state_reg[125]  ( .D(\w0[4][125] ), .CLK(clk), .RST(rst), .I(msg[125]), 
        .Q(state[125]) );
  DFF \state_reg[126]  ( .D(\w0[4][126] ), .CLK(clk), .RST(rst), .I(msg[126]), 
        .Q(state[126]) );
  DFF \state_reg[127]  ( .D(\w0[4][127] ), .CLK(clk), .RST(rst), .I(msg[127]), 
        .Q(state[127]) );
  XNOR U3 ( .A(n12626), .B(n12616), .Z(n12623) );
  XNOR U4 ( .A(n12937), .B(n12927), .Z(n12934) );
  XNOR U5 ( .A(n13559), .B(n13550), .Z(n13557) );
  XOR U6 ( .A(n12012), .B(n12019), .Z(n12018) );
  NOR U7 ( .A(n12832), .B(n12831), .Z(n12828) );
  XOR U8 ( .A(n8813), .B(n8809), .Z(n8659) );
  NANDN U9 ( .A(n7812), .B(n7813), .Z(n7568) );
  NANDN U10 ( .A(n6307), .B(n5833), .Z(n6141) );
  XOR U11 ( .A(n11306), .B(n11297), .Z(n8506) );
  XNOR U12 ( .A(n6726), .B(n6750), .Z(n6571) );
  ANDN U13 ( .B(n2339), .A(n2751), .Z(n2382) );
  ANDN U14 ( .B(n5441), .A(n7364), .Z(n7340) );
  XNOR U15 ( .A(n13352), .B(n13343), .Z(n13350) );
  XOR U16 ( .A(n12706), .B(n12720), .Z(n12717) );
  XNOR U17 ( .A(n14321), .B(n14312), .Z(n14319) );
  XNOR U18 ( .A(n14231), .B(n14222), .Z(n14229) );
  XOR U19 ( .A(n12823), .B(n12837), .Z(n12834) );
  XNOR U20 ( .A(n11901), .B(n11891), .Z(n11898) );
  XNOR U21 ( .A(n12090), .B(n12081), .Z(n12088) );
  XOR U22 ( .A(n14134), .B(n14148), .Z(n14145) );
  XNOR U23 ( .A(n14411), .B(n14402), .Z(n14409) );
  XNOR U24 ( .A(n13442), .B(n13433), .Z(n13440) );
  XOR U25 ( .A(n12961), .B(n12968), .Z(n12967) );
  XOR U26 ( .A(n12650), .B(n12657), .Z(n12656) );
  XOR U27 ( .A(n12561), .B(n12556), .Z(n12559) );
  NOR U28 ( .A(n13560), .B(n13559), .Z(n13556) );
  XOR U29 ( .A(n13667), .B(n13654), .Z(n13138) );
  NOR U30 ( .A(n12715), .B(n12714), .Z(n12711) );
  NOR U31 ( .A(n14143), .B(n14142), .Z(n14139) );
  XNOR U32 ( .A(n11785), .B(n11810), .Z(n11784) );
  XOR U33 ( .A(n12581), .B(n12784), .Z(n12462) );
  XNOR U34 ( .A(n12497), .B(n12496), .Z(n12397) );
  XNOR U35 ( .A(n10360), .B(n11235), .Z(n9442) );
  XNOR U36 ( .A(n10179), .B(n10182), .Z(n10210) );
  ANDN U37 ( .B(n9962), .A(n9969), .Z(n9715) );
  XOR U38 ( .A(n6999), .B(n7052), .Z(n7051) );
  XNOR U39 ( .A(n8659), .B(n8751), .Z(n8750) );
  XOR U40 ( .A(key[280]), .B(n7048), .Z(n7047) );
  XNOR U41 ( .A(n8178), .B(n8181), .Z(n8206) );
  NANDN U42 ( .A(n7671), .B(n7667), .Z(n7526) );
  NANDN U43 ( .A(n7204), .B(n6746), .Z(n6776) );
  XOR U44 ( .A(n8517), .B(n8513), .Z(n8337) );
  XOR U45 ( .A(n7508), .B(n7503), .Z(n7474) );
  XNOR U46 ( .A(n7494), .B(n7558), .Z(n7557) );
  XOR U47 ( .A(n5674), .B(n5633), .Z(n5795) );
  XNOR U48 ( .A(n5686), .B(n5660), .Z(n6117) );
  XOR U49 ( .A(n6743), .B(n6759), .Z(n6607) );
  XOR U50 ( .A(n6653), .B(n6700), .Z(n6602) );
  XNOR U51 ( .A(n2139), .B(n2096), .Z(n2193) );
  XOR U52 ( .A(key[409]), .B(n2681), .Z(n5088) );
  XOR U53 ( .A(n3622), .B(n2691), .Z(n5075) );
  XOR U54 ( .A(n2743), .B(n2803), .Z(n2761) );
  XOR U55 ( .A(n3546), .B(n3537), .Z(n3419) );
  ANDN U56 ( .B(n5462), .A(n6440), .Z(n5505) );
  NANDN U57 ( .A(n5524), .B(n5452), .Z(n5479) );
  XOR U58 ( .A(n524), .B(n515), .Z(n444) );
  XNOR U59 ( .A(n5312), .B(n5425), .Z(n5327) );
  XNOR U60 ( .A(n5350), .B(n5363), .Z(n5362) );
  XOR U61 ( .A(n425), .B(n1651), .Z(n1082) );
  XNOR U62 ( .A(n785), .B(n2036), .Z(n807) );
  XNOR U63 ( .A(n12210), .B(n12197), .Z(n12205) );
  XNOR U64 ( .A(n13531), .B(n13526), .Z(n13529) );
  XOR U65 ( .A(n13344), .B(n13358), .Z(n13355) );
  XNOR U66 ( .A(n12714), .B(n12705), .Z(n12712) );
  XOR U67 ( .A(n14313), .B(n14327), .Z(n14324) );
  XOR U68 ( .A(n14223), .B(n14237), .Z(n14234) );
  XNOR U69 ( .A(n12831), .B(n12822), .Z(n12829) );
  XOR U70 ( .A(n13657), .B(n13671), .Z(n13668) );
  XOR U71 ( .A(n11925), .B(n11932), .Z(n11931) );
  XOR U72 ( .A(n11842), .B(n11761), .Z(n11840) );
  XOR U73 ( .A(n12082), .B(n12096), .Z(n12093) );
  XNOR U74 ( .A(n12072), .B(n12067), .Z(n12070) );
  XNOR U75 ( .A(n14099), .B(n14094), .Z(n14097) );
  XOR U76 ( .A(n13434), .B(n13448), .Z(n13445) );
  XNOR U77 ( .A(n13661), .B(n13651), .Z(n13653) );
  XNOR U78 ( .A(n14138), .B(n14128), .Z(n14130) );
  XOR U79 ( .A(n11987), .B(n11978), .Z(n11684) );
  NOR U80 ( .A(n14322), .B(n14321), .Z(n14318) );
  NOR U81 ( .A(n14232), .B(n14231), .Z(n14228) );
  NOR U82 ( .A(n13443), .B(n13442), .Z(n13439) );
  NOR U83 ( .A(n13353), .B(n13352), .Z(n13349) );
  NOR U84 ( .A(n13666), .B(n13665), .Z(n13662) );
  XOR U85 ( .A(n13561), .B(n13548), .Z(n13276) );
  NOR U86 ( .A(n12091), .B(n12090), .Z(n12087) );
  OR U87 ( .A(n11965), .B(n11690), .Z(n11964) );
  XOR U88 ( .A(n14144), .B(n14131), .Z(n13898) );
  XOR U89 ( .A(n14413), .B(n14400), .Z(n13978) );
  AND U90 ( .A(n12797), .B(n12798), .Z(n12794) );
  XOR U91 ( .A(n12592), .B(n12895), .Z(n12473) );
  XOR U92 ( .A(n12536), .B(n12548), .Z(n12405) );
  XNOR U93 ( .A(n13038), .B(n13028), .Z(n13035) );
  XNOR U94 ( .A(n11751), .B(n11793), .Z(n11673) );
  XNOR U95 ( .A(n11164), .B(n11154), .Z(n11161) );
  XNOR U96 ( .A(n10340), .B(n10324), .Z(n9417) );
  XNOR U97 ( .A(n13788), .B(n13778), .Z(n13785) );
  XNOR U98 ( .A(n9840), .B(n9830), .Z(n9837) );
  XNOR U99 ( .A(n9044), .B(n9034), .Z(n9041) );
  XNOR U100 ( .A(n12399), .B(n12400), .Z(n12495) );
  XNOR U101 ( .A(n9192), .B(n9182), .Z(n9189) );
  XOR U102 ( .A(n10370), .B(n9442), .Z(n11803) );
  XNOR U103 ( .A(n9603), .B(n9773), .Z(n9782) );
  XNOR U104 ( .A(n8873), .B(n8789), .Z(n8784) );
  XOR U105 ( .A(n12281), .B(n13060), .Z(n13018) );
  XOR U106 ( .A(n11144), .B(n11186), .Z(n11159) );
  XOR U107 ( .A(n8890), .B(n8881), .Z(n8678) );
  XOR U108 ( .A(n13748), .B(n13810), .Z(n13759) );
  NANDN U109 ( .A(n10114), .B(n9766), .Z(n9665) );
  XOR U110 ( .A(n9820), .B(n9862), .Z(n9835) );
  ANDN U111 ( .B(n10863), .A(n10870), .Z(n10668) );
  XOR U112 ( .A(n10680), .B(n10691), .Z(n10520) );
  XOR U113 ( .A(n10860), .B(n10880), .Z(n10577) );
  XNOR U114 ( .A(n6328), .B(n6318), .Z(n6325) );
  XNOR U115 ( .A(n9563), .B(n6296), .Z(n6244) );
  XOR U116 ( .A(n9959), .B(n9979), .Z(n9662) );
  XOR U117 ( .A(n8653), .B(n8658), .Z(n8657) );
  NAND U118 ( .A(n8567), .B(n8573), .Z(n8579) );
  XNOR U119 ( .A(n10482), .B(n10485), .Z(n10565) );
  XNOR U120 ( .A(n5731), .B(n6171), .Z(n6153) );
  XNOR U121 ( .A(n7550), .B(n8112), .Z(n8098) );
  XNOR U122 ( .A(n6822), .B(n6812), .Z(n6819) );
  XOR U123 ( .A(key[281]), .B(n6390), .Z(n7057) );
  XNOR U124 ( .A(n7844), .B(n7643), .Z(n7638) );
  XOR U125 ( .A(n6783), .B(n6577), .Z(n6801) );
  XOR U126 ( .A(n6188), .B(n6179), .Z(n5725) );
  XOR U127 ( .A(n8129), .B(n8120), .Z(n7585) );
  XOR U128 ( .A(n7040), .B(n6400), .Z(n7037) );
  XOR U129 ( .A(n7861), .B(n7852), .Z(n7515) );
  NANDN U130 ( .A(n5980), .B(n5799), .Z(n5805) );
  NANDN U131 ( .A(n6157), .B(n5732), .Z(n5785) );
  NANDN U132 ( .A(n7599), .B(n7600), .Z(n7594) );
  ANDN U133 ( .B(n9472), .A(n9476), .Z(n8407) );
  XOR U134 ( .A(n7577), .B(n7572), .Z(n7494) );
  XNOR U135 ( .A(n2940), .B(n2930), .Z(n2937) );
  XOR U136 ( .A(n5740), .B(n5756), .Z(n5696) );
  XOR U137 ( .A(n5796), .B(n5813), .Z(n5681) );
  XNOR U138 ( .A(n2476), .B(n2466), .Z(n2473) );
  XOR U139 ( .A(n6662), .B(n6679), .Z(n6592) );
  XOR U140 ( .A(n6605), .B(n6572), .Z(n6742) );
  XNOR U141 ( .A(n8274), .B(n8263), .Z(n8271) );
  XOR U142 ( .A(n5684), .B(n5661), .Z(n5829) );
  XOR U143 ( .A(n2538), .B(n3805), .Z(n4938) );
  XNOR U144 ( .A(n8335), .B(n8440), .Z(n3978) );
  XNOR U145 ( .A(n5122), .B(n5112), .Z(n5119) );
  XNOR U146 ( .A(n1880), .B(n867), .Z(n5275) );
  XNOR U147 ( .A(n1920), .B(n1851), .Z(n1974) );
  XNOR U148 ( .A(n1710), .B(n1667), .Z(n1764) );
  XNOR U149 ( .A(n1303), .B(n1260), .Z(n1357) );
  XNOR U150 ( .A(n1110), .B(n1064), .Z(n1164) );
  XNOR U151 ( .A(n907), .B(n848), .Z(n961) );
  XNOR U152 ( .A(n292), .B(n249), .Z(n346) );
  XNOR U153 ( .A(n89), .B(n43), .Z(n143) );
  XNOR U154 ( .A(n2377), .B(n2424), .Z(n2523) );
  XNOR U155 ( .A(n2366), .B(n2902), .Z(n2987) );
  XNOR U156 ( .A(n2563), .B(n3819), .Z(n4925) );
  XNOR U157 ( .A(n4411), .B(n4401), .Z(n4408) );
  XOR U158 ( .A(n2397), .B(n2641), .Z(n2417) );
  ANDN U159 ( .B(n2351), .A(n2598), .Z(n2405) );
  XOR U160 ( .A(n2832), .B(n2826), .Z(n2837) );
  ANDN U161 ( .B(n3454), .A(n3852), .Z(n3459) );
  NANDN U162 ( .A(n4831), .B(n4579), .Z(n4620) );
  XOR U163 ( .A(key[408]), .B(n5067), .Z(n5082) );
  XOR U164 ( .A(n3421), .B(n3416), .Z(n3351) );
  XOR U165 ( .A(n5376), .B(n5371), .Z(n5334) );
  XNOR U166 ( .A(n5416), .B(n5520), .Z(n5366) );
  XOR U167 ( .A(n862), .B(n857), .Z(n423) );
  XOR U168 ( .A(n1846), .B(n1841), .Z(n1830) );
  XOR U169 ( .A(n1662), .B(n1657), .Z(n1645) );
  XOR U170 ( .A(n1466), .B(n1461), .Z(n1450) );
  XOR U171 ( .A(n1255), .B(n1250), .Z(n1239) );
  XOR U172 ( .A(n1059), .B(n1054), .Z(n1043) );
  XOR U173 ( .A(n843), .B(n838), .Z(n827) );
  XOR U174 ( .A(n446), .B(n441), .Z(n428) );
  XOR U175 ( .A(n244), .B(n239), .Z(n228) );
  XOR U176 ( .A(n38), .B(n33), .Z(n22) );
  XOR U177 ( .A(n4156), .B(n4151), .Z(n3264) );
  XOR U178 ( .A(n3094), .B(n3089), .Z(n3078) );
  XOR U179 ( .A(n2091), .B(n2086), .Z(n2075) );
  XNOR U180 ( .A(n2277), .B(n2898), .Z(n2446) );
  XNOR U181 ( .A(n2230), .B(n2379), .Z(n814) );
  XNOR U182 ( .A(n3480), .B(n3372), .Z(n3659) );
  XOR U183 ( .A(n3387), .B(n3386), .Z(n3385) );
  XOR U184 ( .A(n5328), .B(n5311), .Z(n5325) );
  XNOR U185 ( .A(n5344), .B(n5380), .Z(n5377) );
  XNOR U186 ( .A(n1031), .B(n405), .Z(n1022) );
  XOR U187 ( .A(n819), .B(n1408), .Z(n2237) );
  XNOR U188 ( .A(n11965), .B(n11689), .Z(n12005) );
  XNOR U189 ( .A(n11880), .B(n11703), .Z(n11919) );
  XNOR U190 ( .A(n11986), .B(n11976), .Z(n11983) );
  XNOR U191 ( .A(n12569), .B(n12445), .Z(n12644) );
  XNOR U192 ( .A(n12905), .B(n12384), .Z(n12955) );
  XNOR U193 ( .A(n14018), .B(n14006), .Z(n14016) );
  XNOR U194 ( .A(n12533), .B(n12522), .Z(n12531) );
  XNOR U195 ( .A(n12257), .B(n12255), .Z(n12243) );
  XNOR U196 ( .A(n13306), .B(n13295), .Z(n13304) );
  XNOR U197 ( .A(n13264), .B(n13248), .Z(n13262) );
  XOR U198 ( .A(n13551), .B(n13565), .Z(n13562) );
  XNOR U199 ( .A(n13665), .B(n13656), .Z(n13663) );
  XNOR U200 ( .A(n14142), .B(n14133), .Z(n14140) );
  XOR U201 ( .A(n14403), .B(n14417), .Z(n14414) );
  XNOR U202 ( .A(n12797), .B(n12793), .Z(n12796) );
  XNOR U203 ( .A(n14044), .B(n14028), .Z(n14042) );
  NOR U204 ( .A(n11823), .B(n11981), .Z(n11972) );
  XOR U205 ( .A(n12204), .B(n12195), .Z(n11728) );
  XOR U206 ( .A(n13444), .B(n13431), .Z(n13231) );
  XOR U207 ( .A(n12938), .B(n12929), .Z(n12470) );
  NOR U208 ( .A(n14412), .B(n14411), .Z(n14408) );
  XOR U209 ( .A(n13354), .B(n13341), .Z(n13286) );
  XOR U210 ( .A(n12716), .B(n12703), .Z(n12517) );
  XOR U211 ( .A(n14323), .B(n14310), .Z(n13988) );
  XOR U212 ( .A(n14233), .B(n14220), .Z(n14070) );
  XOR U213 ( .A(n12627), .B(n12618), .Z(n12440) );
  XOR U214 ( .A(n12833), .B(n12820), .Z(n12587) );
  XOR U215 ( .A(n11902), .B(n11893), .Z(n11698) );
  XOR U216 ( .A(n12092), .B(n12079), .Z(n11863) );
  XNOR U217 ( .A(n14064), .B(n14085), .Z(n14063) );
  XNOR U218 ( .A(n13270), .B(n13517), .Z(n13269) );
  AND U219 ( .A(n13661), .B(n13641), .Z(n13652) );
  AND U220 ( .A(n14138), .B(n14118), .Z(n14129) );
  XNOR U221 ( .A(n12462), .B(n12463), .Z(n12777) );
  XNOR U222 ( .A(n10074), .B(n8974), .Z(n8989) );
  XNOR U223 ( .A(n9339), .B(n9329), .Z(n9336) );
  XOR U224 ( .A(n13089), .B(n9900), .Z(n13221) );
  XOR U225 ( .A(n12049), .B(n12059), .Z(n11743) );
  XNOR U226 ( .A(n13205), .B(n11105), .Z(n9930) );
  XNOR U227 ( .A(n10902), .B(n10892), .Z(n10899) );
  XNOR U228 ( .A(n10001), .B(n9991), .Z(n9998) );
  XNOR U229 ( .A(n10316), .B(n10319), .Z(n10343) );
  XOR U230 ( .A(n10094), .B(n10851), .Z(n8959) );
  XNOR U231 ( .A(n9617), .B(n9747), .Z(n9756) );
  XNOR U232 ( .A(n13265), .B(n13193), .Z(n9128) );
  XOR U233 ( .A(n9401), .B(n11236), .Z(n11233) );
  XNOR U234 ( .A(n11471), .B(n11528), .Z(n11522) );
  XNOR U235 ( .A(n11097), .B(n11118), .Z(n11113) );
  XNOR U236 ( .A(n10561), .B(n10689), .Z(n10699) );
  XOR U237 ( .A(n9981), .B(n10023), .Z(n9996) );
  XNOR U238 ( .A(n9289), .B(n9290), .Z(n9288) );
  XNOR U239 ( .A(n11483), .B(n11550), .Z(n11545) );
  XOR U240 ( .A(n11588), .B(n11579), .Z(n11436) );
  XOR U241 ( .A(n12316), .B(n12307), .Z(n11450) );
  XOR U242 ( .A(n10173), .B(n10182), .Z(n10195) );
  XOR U243 ( .A(n10130), .B(n10121), .Z(n9596) );
  XOR U244 ( .A(n10267), .B(n10258), .Z(n9610) );
  NANDN U245 ( .A(n8816), .B(n8817), .Z(n8806) );
  NANDN U246 ( .A(n9023), .B(n9019), .Z(n8720) );
  ANDN U247 ( .B(n12287), .A(n12286), .Z(n12268) );
  ANDN U248 ( .B(n11125), .A(n11132), .Z(n10714) );
  NANDN U249 ( .A(n8859), .B(n8860), .Z(n8712) );
  XOR U250 ( .A(key[128]), .B(n10813), .Z(n14072) );
  XOR U251 ( .A(n10882), .B(n10924), .Z(n10897) );
  ANDN U252 ( .B(n11497), .A(n13767), .Z(n13738) );
  ANDN U253 ( .B(n9801), .A(n9808), .Z(n9725) );
  XOR U254 ( .A(n10753), .B(n10744), .Z(n10540) );
  XOR U255 ( .A(n11025), .B(n11016), .Z(n10555) );
  XOR U256 ( .A(n11122), .B(n11142), .Z(n10608) );
  XOR U257 ( .A(n9798), .B(n9818), .Z(n9642) );
  NANDN U258 ( .A(n8841), .B(n8842), .Z(n8744) );
  NANDN U259 ( .A(n12291), .B(n11538), .Z(n11454) );
  XNOR U260 ( .A(n8652), .B(n8660), .Z(n8751) );
  XOR U261 ( .A(n12282), .B(n12278), .Z(n11415) );
  XOR U262 ( .A(n8741), .B(n8736), .Z(n8666) );
  XOR U263 ( .A(n8680), .B(n8675), .Z(n8633) );
  XOR U264 ( .A(n8690), .B(n8685), .Z(n8641) );
  XNOR U265 ( .A(n10571), .B(n10666), .Z(n10665) );
  XOR U266 ( .A(n11494), .B(n13746), .Z(n11388) );
  XNOR U267 ( .A(n7996), .B(n7986), .Z(n7993) );
  XNOR U268 ( .A(n9674), .B(n9554), .Z(n8187) );
  XNOR U269 ( .A(n8569), .B(n8560), .Z(n8568) );
  XNOR U270 ( .A(n7692), .B(n7682), .Z(n7689) );
  XNOR U271 ( .A(n6001), .B(n5991), .Z(n5998) );
  XNOR U272 ( .A(n7092), .B(n7082), .Z(n7089) );
  XNOR U273 ( .A(n7225), .B(n7215), .Z(n7222) );
  XOR U274 ( .A(key[329]), .B(n5972), .Z(n7329) );
  XNOR U275 ( .A(n10382), .B(n10405), .Z(n10401) );
  XOR U276 ( .A(key[314]), .B(n6287), .Z(n8229) );
  XOR U277 ( .A(n6389), .B(n8081), .Z(n8080) );
  XNOR U278 ( .A(n10592), .B(n10489), .Z(n7941) );
  XNOR U279 ( .A(n9547), .B(n9550), .Z(n9630) );
  XOR U280 ( .A(n8398), .B(n8471), .Z(n8565) );
  XOR U281 ( .A(n7575), .B(n7961), .Z(n7975) );
  XNOR U282 ( .A(n5658), .B(n5773), .Z(n5763) );
  XOR U283 ( .A(n7506), .B(n7611), .Z(n7662) );
  XNOR U284 ( .A(n9471), .B(n8492), .Z(n8488) );
  XOR U285 ( .A(n6761), .B(n6748), .Z(n6772) );
  XOR U286 ( .A(n10433), .B(n10424), .Z(n8449) );
  ANDN U287 ( .B(n10386), .A(n10385), .Z(n8453) );
  XOR U288 ( .A(n8198), .B(n8213), .Z(n8210) );
  XNOR U289 ( .A(n6570), .B(n6718), .Z(n6707) );
  NANDN U290 ( .A(n6791), .B(n6645), .Z(n6733) );
  XOR U291 ( .A(n6681), .B(n6667), .Z(n6692) );
  AND U292 ( .A(n11281), .B(n11282), .Z(n11278) );
  XNOR U293 ( .A(n11358), .B(n11425), .Z(n11285) );
  NANDN U294 ( .A(n7830), .B(n7831), .Z(n7538) );
  XOR U295 ( .A(n5867), .B(n5858), .Z(n5693) );
  NANDN U296 ( .A(n5842), .B(n5743), .Z(n5767) );
  NANDN U297 ( .A(n7071), .B(n6665), .Z(n6696) );
  XOR U298 ( .A(n9498), .B(n9489), .Z(n8388) );
  XOR U299 ( .A(n5830), .B(n6124), .Z(n5686) );
  XOR U300 ( .A(n5662), .B(n6146), .Z(n5617) );
  XOR U301 ( .A(n7591), .B(n7587), .Z(n7562) );
  NANDN U302 ( .A(n6931), .B(n6656), .Z(n6711) );
  XOR U303 ( .A(n6956), .B(n6947), .Z(n6599) );
  XOR U304 ( .A(n5043), .B(n3651), .Z(n5085) );
  XOR U305 ( .A(n7517), .B(n7512), .Z(n7480) );
  XNOR U306 ( .A(n2619), .B(n2609), .Z(n2616) );
  XNOR U307 ( .A(n2781), .B(n2771), .Z(n2778) );
  XNOR U308 ( .A(n3713), .B(n3703), .Z(n3710) );
  XNOR U309 ( .A(n8404), .B(n8403), .Z(n3031) );
  XNOR U310 ( .A(n3875), .B(n3865), .Z(n3872) );
  XNOR U311 ( .A(n6466), .B(n6456), .Z(n6463) );
  XNOR U312 ( .A(n7392), .B(n7382), .Z(n7389) );
  XNOR U313 ( .A(n4142), .B(n4099), .Z(n4816) );
  XNOR U314 ( .A(n5550), .B(n5540), .Z(n5547) );
  XOR U315 ( .A(n5188), .B(n3952), .Z(n3026) );
  ANDN U316 ( .B(n5170), .A(n4634), .Z(n5156) );
  XOR U317 ( .A(n3820), .B(n3788), .Z(n4937) );
  XOR U318 ( .A(n6573), .B(n6780), .Z(n6531) );
  XNOR U319 ( .A(n7474), .B(n7475), .Z(n7473) );
  XOR U320 ( .A(n3018), .B(n3019), .Z(n3017) );
  XOR U321 ( .A(n2581), .B(n2579), .Z(n2575) );
  XNOR U322 ( .A(n5681), .B(n5632), .Z(n5751) );
  XOR U323 ( .A(key[506]), .B(n2844), .Z(n2843) );
  XNOR U324 ( .A(n6607), .B(n6571), .Z(n6753) );
  XNOR U325 ( .A(n3470), .B(n4017), .Z(n4004) );
  XNOR U326 ( .A(n4095), .B(n4122), .Z(n4107) );
  XNOR U327 ( .A(n3595), .B(n3598), .Z(n3623) );
  XNOR U328 ( .A(n4487), .B(n4674), .Z(n4664) );
  XNOR U329 ( .A(n4578), .B(n4845), .Z(n4827) );
  XNOR U330 ( .A(n4564), .B(n4972), .Z(n4964) );
  XNOR U331 ( .A(n5250), .B(n5240), .Z(n5247) );
  XNOR U332 ( .A(n1950), .B(n1940), .Z(n1947) );
  XNOR U333 ( .A(n1740), .B(n1730), .Z(n1737) );
  XNOR U334 ( .A(n1544), .B(n1534), .Z(n1541) );
  XNOR U335 ( .A(n1333), .B(n1323), .Z(n1330) );
  XNOR U336 ( .A(n1140), .B(n1130), .Z(n1137) );
  XNOR U337 ( .A(n937), .B(n927), .Z(n934) );
  XNOR U338 ( .A(n780), .B(n800), .Z(n777) );
  XNOR U339 ( .A(n656), .B(n692), .Z(n686) );
  XNOR U340 ( .A(n322), .B(n312), .Z(n319) );
  XNOR U341 ( .A(n119), .B(n109), .Z(n116) );
  XNOR U342 ( .A(n4234), .B(n4224), .Z(n4231) );
  XNOR U343 ( .A(n3172), .B(n3162), .Z(n3169) );
  XNOR U344 ( .A(n2169), .B(n2159), .Z(n2166) );
  XOR U345 ( .A(key[384]), .B(n2728), .Z(n2724) );
  XOR U346 ( .A(n3673), .B(n3735), .Z(n3685) );
  ANDN U347 ( .B(n3485), .A(n3690), .Z(n3477) );
  XOR U348 ( .A(n4043), .B(n4034), .Z(n3998) );
  XOR U349 ( .A(n3835), .B(n3897), .Z(n3847) );
  NANDN U350 ( .A(n8245), .B(n5397), .Z(n5428) );
  NANDN U351 ( .A(n4697), .B(n4600), .Z(n4668) );
  XOR U352 ( .A(n4723), .B(n4714), .Z(n4537) );
  XOR U353 ( .A(n4862), .B(n4853), .Z(n4572) );
  XOR U354 ( .A(n5000), .B(n4991), .Z(n4557) );
  NANDN U355 ( .A(n4968), .B(n4611), .Z(n4687) );
  XOR U356 ( .A(n5123), .B(n5114), .Z(n4593) );
  NANDN U357 ( .A(n5229), .B(n1442), .Z(n1878) );
  NANDN U358 ( .A(n3273), .B(n3053), .Z(n2064) );
  XOR U359 ( .A(n3293), .B(n3284), .Z(n2053) );
  NANDN U360 ( .A(n1929), .B(n1887), .Z(n1918) );
  NANDN U361 ( .A(n1719), .B(n1677), .Z(n1708) );
  NANDN U362 ( .A(n1523), .B(n1481), .Z(n1512) );
  NANDN U363 ( .A(n1312), .B(n1270), .Z(n1301) );
  NANDN U364 ( .A(n1119), .B(n1074), .Z(n1108) );
  NANDN U365 ( .A(n916), .B(n874), .Z(n905) );
  XOR U366 ( .A(n727), .B(n718), .Z(n650) );
  NANDN U367 ( .A(n301), .B(n259), .Z(n290) );
  NANDN U368 ( .A(n98), .B(n53), .Z(n87) );
  NANDN U369 ( .A(n4213), .B(n4171), .Z(n4202) );
  NANDN U370 ( .A(n3151), .B(n3109), .Z(n3140) );
  NANDN U371 ( .A(n2148), .B(n2106), .Z(n2137) );
  XOR U372 ( .A(n2367), .B(n2361), .Z(n2276) );
  XOR U373 ( .A(n2378), .B(n2372), .Z(n2245) );
  XOR U374 ( .A(n2355), .B(n2349), .Z(n2238) );
  XOR U375 ( .A(n2255), .B(n2250), .Z(n2231) );
  XOR U376 ( .A(n3351), .B(n3370), .Z(n3413) );
  XNOR U377 ( .A(n3345), .B(n3364), .Z(n1633) );
  XOR U378 ( .A(n5404), .B(n5399), .Z(n5328) );
  XOR U379 ( .A(n5334), .B(n5370), .Z(n5367) );
  XOR U380 ( .A(n640), .B(n1438), .Z(n422) );
  XOR U381 ( .A(n1835), .B(n1883), .Z(n1829) );
  XOR U382 ( .A(n1650), .B(n1673), .Z(n1644) );
  XOR U383 ( .A(n1455), .B(n1477), .Z(n1449) );
  XOR U384 ( .A(n1244), .B(n1266), .Z(n1238) );
  XOR U385 ( .A(n1048), .B(n1070), .Z(n1042) );
  XOR U386 ( .A(n832), .B(n870), .Z(n826) );
  XNOR U387 ( .A(n469), .B(n457), .Z(n427) );
  XOR U388 ( .A(n233), .B(n255), .Z(n227) );
  XOR U389 ( .A(n27), .B(n49), .Z(n21) );
  XNOR U390 ( .A(n12), .B(n19), .Z(n13) );
  XOR U391 ( .A(n4335), .B(n4342), .Z(n10) );
  XOR U392 ( .A(n3269), .B(n4167), .Z(n3263) );
  XOR U393 ( .A(n3083), .B(n3105), .Z(n3077) );
  XOR U394 ( .A(n2080), .B(n2102), .Z(n2074) );
  XOR U395 ( .A(n3402), .B(n3387), .Z(n178) );
  XOR U396 ( .A(n814), .B(n1392), .Z(n2391) );
  XOR U397 ( .A(n187), .B(n188), .Z(n186) );
  XOR U398 ( .A(n1036), .B(n1035), .Z(n1032) );
  XNOR U399 ( .A(n1224), .B(n1221), .Z(n1815) );
  XOR U400 ( .A(n1), .B(n2), .Z(out[9]) );
  XNOR U401 ( .A(n3), .B(n4), .Z(n2) );
  XOR U402 ( .A(key[521]), .B(n5), .Z(n1) );
  XOR U403 ( .A(n6), .B(n7), .Z(out[99]) );
  XNOR U404 ( .A(n8), .B(n9), .Z(n7) );
  XOR U405 ( .A(n10), .B(n11), .Z(n6) );
  XNOR U406 ( .A(key[611]), .B(n12), .Z(n11) );
  XNOR U407 ( .A(key[610]), .B(n13), .Z(out[98]) );
  XOR U408 ( .A(n14), .B(n15), .Z(out[97]) );
  XNOR U409 ( .A(n8), .B(n16), .Z(n15) );
  XNOR U410 ( .A(key[609]), .B(n12), .Z(n14) );
  XOR U411 ( .A(n17), .B(n18), .Z(out[96]) );
  XNOR U412 ( .A(key[608]), .B(n19), .Z(n18) );
  XOR U413 ( .A(n20), .B(n21), .Z(out[95]) );
  XOR U414 ( .A(n22), .B(n23), .Z(n20) );
  XOR U415 ( .A(key[607]), .B(n24), .Z(n23) );
  XNOR U416 ( .A(n25), .B(n26), .Z(out[94]) );
  XNOR U417 ( .A(key[606]), .B(n27), .Z(n26) );
  XOR U418 ( .A(n28), .B(n29), .Z(out[93]) );
  XNOR U419 ( .A(n30), .B(n31), .Z(n29) );
  XOR U420 ( .A(n22), .B(n32), .Z(n31) );
  XNOR U421 ( .A(n34), .B(n35), .Z(n33) );
  NANDN U422 ( .A(n36), .B(n37), .Z(n35) );
  XOR U423 ( .A(n39), .B(n40), .Z(n28) );
  XOR U424 ( .A(key[605]), .B(n41), .Z(n40) );
  ANDN U425 ( .B(n42), .A(n43), .Z(n39) );
  XNOR U426 ( .A(n44), .B(n45), .Z(out[92]) );
  XNOR U427 ( .A(key[604]), .B(n46), .Z(n45) );
  XOR U428 ( .A(n47), .B(n48), .Z(out[91]) );
  XNOR U429 ( .A(n49), .B(n25), .Z(n48) );
  XNOR U430 ( .A(n50), .B(n51), .Z(n25) );
  XNOR U431 ( .A(n52), .B(n41), .Z(n51) );
  ANDN U432 ( .B(n53), .A(n54), .Z(n41) );
  NOR U433 ( .A(n55), .B(n56), .Z(n52) );
  XNOR U434 ( .A(n57), .B(n58), .Z(n47) );
  XOR U435 ( .A(key[603]), .B(n24), .Z(n58) );
  XOR U436 ( .A(key[602]), .B(n44), .Z(out[90]) );
  XNOR U437 ( .A(n59), .B(n60), .Z(n44) );
  XNOR U438 ( .A(n61), .B(n62), .Z(out[8]) );
  XNOR U439 ( .A(key[520]), .B(n63), .Z(n62) );
  XOR U440 ( .A(n64), .B(n21), .Z(out[89]) );
  XNOR U441 ( .A(n50), .B(n65), .Z(n49) );
  XNOR U442 ( .A(n66), .B(n67), .Z(n65) );
  NANDN U443 ( .A(n68), .B(n37), .Z(n67) );
  XNOR U444 ( .A(n32), .B(n69), .Z(n50) );
  XNOR U445 ( .A(n70), .B(n71), .Z(n69) );
  NANDN U446 ( .A(n72), .B(n73), .Z(n71) );
  XOR U447 ( .A(n60), .B(n57), .Z(n27) );
  XNOR U448 ( .A(n32), .B(n74), .Z(n57) );
  XNOR U449 ( .A(n66), .B(n75), .Z(n74) );
  NANDN U450 ( .A(n76), .B(n77), .Z(n75) );
  OR U451 ( .A(n78), .B(n79), .Z(n66) );
  XOR U452 ( .A(n80), .B(n70), .Z(n32) );
  NANDN U453 ( .A(n81), .B(n82), .Z(n70) );
  ANDN U454 ( .B(n83), .A(n84), .Z(n80) );
  XNOR U455 ( .A(key[601]), .B(n59), .Z(n64) );
  IV U456 ( .A(n24), .Z(n59) );
  XOR U457 ( .A(n85), .B(n86), .Z(n24) );
  XNOR U458 ( .A(n87), .B(n88), .Z(n86) );
  NAND U459 ( .A(n42), .B(n89), .Z(n88) );
  XNOR U460 ( .A(n30), .B(n90), .Z(out[88]) );
  XOR U461 ( .A(key[600]), .B(n60), .Z(n90) );
  XNOR U462 ( .A(n85), .B(n91), .Z(n60) );
  XOR U463 ( .A(n92), .B(n34), .Z(n91) );
  OR U464 ( .A(n93), .B(n78), .Z(n34) );
  XNOR U465 ( .A(n37), .B(n77), .Z(n78) );
  ANDN U466 ( .B(n94), .A(n95), .Z(n92) );
  IV U467 ( .A(n46), .Z(n30) );
  XOR U468 ( .A(n38), .B(n96), .Z(n46) );
  XOR U469 ( .A(n97), .B(n87), .Z(n96) );
  XNOR U470 ( .A(n56), .B(n42), .Z(n53) );
  NOR U471 ( .A(n99), .B(n56), .Z(n97) );
  XNOR U472 ( .A(n85), .B(n100), .Z(n38) );
  XNOR U473 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U474 ( .A(n72), .B(n103), .Z(n102) );
  XOR U475 ( .A(n104), .B(n101), .Z(n85) );
  OR U476 ( .A(n81), .B(n105), .Z(n101) );
  XOR U477 ( .A(n106), .B(n72), .Z(n81) );
  XNOR U478 ( .A(n77), .B(n42), .Z(n72) );
  XOR U479 ( .A(n107), .B(n108), .Z(n42) );
  NANDN U480 ( .A(n109), .B(n110), .Z(n108) );
  IV U481 ( .A(n95), .Z(n77) );
  XNOR U482 ( .A(n111), .B(n112), .Z(n95) );
  NANDN U483 ( .A(n109), .B(n113), .Z(n112) );
  ANDN U484 ( .B(n106), .A(n114), .Z(n104) );
  IV U485 ( .A(n84), .Z(n106) );
  XOR U486 ( .A(n56), .B(n37), .Z(n84) );
  XNOR U487 ( .A(n115), .B(n111), .Z(n37) );
  NANDN U488 ( .A(n116), .B(n117), .Z(n111) );
  XOR U489 ( .A(n113), .B(n118), .Z(n117) );
  ANDN U490 ( .B(n118), .A(n119), .Z(n115) );
  XOR U491 ( .A(n120), .B(n107), .Z(n56) );
  NANDN U492 ( .A(n116), .B(n121), .Z(n107) );
  XOR U493 ( .A(n122), .B(n110), .Z(n121) );
  XNOR U494 ( .A(n123), .B(n124), .Z(n109) );
  XOR U495 ( .A(n125), .B(n126), .Z(n124) );
  XNOR U496 ( .A(n127), .B(n128), .Z(n123) );
  XNOR U497 ( .A(n129), .B(n130), .Z(n128) );
  ANDN U498 ( .B(n122), .A(n126), .Z(n129) );
  ANDN U499 ( .B(n122), .A(n119), .Z(n120) );
  XNOR U500 ( .A(n125), .B(n131), .Z(n119) );
  XOR U501 ( .A(n132), .B(n130), .Z(n131) );
  NAND U502 ( .A(n133), .B(n134), .Z(n130) );
  XNOR U503 ( .A(n127), .B(n110), .Z(n134) );
  IV U504 ( .A(n122), .Z(n127) );
  XNOR U505 ( .A(n113), .B(n126), .Z(n133) );
  IV U506 ( .A(n118), .Z(n126) );
  XOR U507 ( .A(n135), .B(n136), .Z(n118) );
  XNOR U508 ( .A(n137), .B(n138), .Z(n136) );
  XNOR U509 ( .A(n139), .B(n140), .Z(n135) );
  NOR U510 ( .A(n55), .B(n99), .Z(n139) );
  AND U511 ( .A(n110), .B(n113), .Z(n132) );
  XNOR U512 ( .A(n110), .B(n113), .Z(n125) );
  XNOR U513 ( .A(n141), .B(n142), .Z(n113) );
  XNOR U514 ( .A(n143), .B(n138), .Z(n142) );
  XOR U515 ( .A(n144), .B(n145), .Z(n141) );
  XNOR U516 ( .A(n146), .B(n140), .Z(n145) );
  OR U517 ( .A(n54), .B(n98), .Z(n140) );
  XOR U518 ( .A(n99), .B(n89), .Z(n98) );
  XNOR U519 ( .A(n55), .B(n43), .Z(n54) );
  ANDN U520 ( .B(n89), .A(n43), .Z(n146) );
  XNOR U521 ( .A(n147), .B(n148), .Z(n110) );
  XNOR U522 ( .A(n138), .B(n149), .Z(n148) );
  XOR U523 ( .A(n68), .B(n144), .Z(n149) );
  XNOR U524 ( .A(n99), .B(n150), .Z(n138) );
  XNOR U525 ( .A(n151), .B(n152), .Z(n147) );
  XNOR U526 ( .A(n153), .B(n154), .Z(n152) );
  ANDN U527 ( .B(n94), .A(n76), .Z(n153) );
  XNOR U528 ( .A(n155), .B(n156), .Z(n122) );
  XNOR U529 ( .A(n143), .B(n157), .Z(n156) );
  XNOR U530 ( .A(n76), .B(n137), .Z(n157) );
  XOR U531 ( .A(n144), .B(n158), .Z(n137) );
  XNOR U532 ( .A(n159), .B(n160), .Z(n158) );
  NAND U533 ( .A(n103), .B(n73), .Z(n160) );
  XNOR U534 ( .A(n161), .B(n159), .Z(n144) );
  NANDN U535 ( .A(n105), .B(n82), .Z(n159) );
  XOR U536 ( .A(n83), .B(n73), .Z(n82) );
  XNOR U537 ( .A(n162), .B(n43), .Z(n73) );
  XOR U538 ( .A(n114), .B(n103), .Z(n105) );
  XOR U539 ( .A(n94), .B(n89), .Z(n103) );
  ANDN U540 ( .B(n83), .A(n114), .Z(n161) );
  XOR U541 ( .A(n151), .B(n99), .Z(n114) );
  XOR U542 ( .A(n163), .B(n164), .Z(n99) );
  XOR U543 ( .A(n165), .B(n166), .Z(n164) );
  XOR U544 ( .A(n167), .B(n150), .Z(n83) );
  XNOR U545 ( .A(n168), .B(n169), .Z(n43) );
  XNOR U546 ( .A(n170), .B(n166), .Z(n169) );
  XNOR U547 ( .A(n166), .B(n168), .Z(n89) );
  XNOR U548 ( .A(n94), .B(n171), .Z(n155) );
  XNOR U549 ( .A(n172), .B(n154), .Z(n171) );
  OR U550 ( .A(n79), .B(n93), .Z(n154) );
  XNOR U551 ( .A(n151), .B(n94), .Z(n93) );
  XOR U552 ( .A(n68), .B(n162), .Z(n79) );
  IV U553 ( .A(n76), .Z(n162) );
  XOR U554 ( .A(n150), .B(n173), .Z(n76) );
  XNOR U555 ( .A(n170), .B(n163), .Z(n173) );
  XOR U556 ( .A(key[602]), .B(\w0[4][90] ), .Z(n163) );
  XOR U557 ( .A(n174), .B(n175), .Z(\w0[4][90] ) );
  XOR U558 ( .A(n176), .B(n177), .Z(n175) );
  XOR U559 ( .A(n178), .B(n179), .Z(n174) );
  IV U560 ( .A(n55), .Z(n150) );
  XNOR U561 ( .A(n168), .B(n180), .Z(n55) );
  XNOR U562 ( .A(n166), .B(n181), .Z(n180) );
  ANDN U563 ( .B(n167), .A(n36), .Z(n172) );
  IV U564 ( .A(n68), .Z(n167) );
  XNOR U565 ( .A(n168), .B(n182), .Z(n68) );
  XNOR U566 ( .A(n166), .B(n183), .Z(n182) );
  XOR U567 ( .A(n36), .B(n184), .Z(n166) );
  XOR U568 ( .A(key[606]), .B(\w0[4][94] ), .Z(n184) );
  XNOR U569 ( .A(n185), .B(n186), .Z(\w0[4][94] ) );
  IV U570 ( .A(n151), .Z(n36) );
  XOR U571 ( .A(key[605]), .B(\w0[4][93] ), .Z(n168) );
  XOR U572 ( .A(n189), .B(n190), .Z(\w0[4][93] ) );
  XOR U573 ( .A(n191), .B(n192), .Z(n190) );
  XOR U574 ( .A(n193), .B(n194), .Z(n189) );
  XOR U575 ( .A(n195), .B(n196), .Z(n94) );
  XNOR U576 ( .A(n183), .B(n181), .Z(n196) );
  XOR U577 ( .A(key[607]), .B(\w0[4][95] ), .Z(n181) );
  XNOR U578 ( .A(n197), .B(n198), .Z(\w0[4][95] ) );
  XOR U579 ( .A(n199), .B(n200), .Z(n198) );
  XOR U580 ( .A(key[604]), .B(\w0[4][92] ), .Z(n183) );
  XOR U581 ( .A(n201), .B(n202), .Z(\w0[4][92] ) );
  XOR U582 ( .A(n203), .B(n204), .Z(n202) );
  XOR U583 ( .A(n205), .B(n206), .Z(n201) );
  XNOR U584 ( .A(n151), .B(n165), .Z(n195) );
  XOR U585 ( .A(n170), .B(n207), .Z(n165) );
  XOR U586 ( .A(key[603]), .B(\w0[4][91] ), .Z(n207) );
  XOR U587 ( .A(n208), .B(n209), .Z(\w0[4][91] ) );
  XOR U588 ( .A(n210), .B(n211), .Z(n209) );
  XOR U589 ( .A(n212), .B(n213), .Z(n208) );
  XOR U590 ( .A(key[601]), .B(\w0[4][89] ), .Z(n170) );
  XOR U591 ( .A(n214), .B(n215), .Z(\w0[4][89] ) );
  XOR U592 ( .A(n216), .B(n217), .Z(n215) );
  XOR U593 ( .A(n218), .B(n219), .Z(n214) );
  XOR U594 ( .A(key[600]), .B(\w0[4][88] ), .Z(n151) );
  XOR U595 ( .A(n220), .B(n221), .Z(\w0[4][88] ) );
  XOR U596 ( .A(n222), .B(n223), .Z(n221) );
  XNOR U597 ( .A(n224), .B(n225), .Z(n220) );
  XOR U598 ( .A(n226), .B(n227), .Z(out[87]) );
  XOR U599 ( .A(n228), .B(n229), .Z(n226) );
  XNOR U600 ( .A(key[599]), .B(n230), .Z(n229) );
  XNOR U601 ( .A(n231), .B(n232), .Z(out[86]) );
  XNOR U602 ( .A(key[598]), .B(n233), .Z(n232) );
  XOR U603 ( .A(n234), .B(n235), .Z(out[85]) );
  XNOR U604 ( .A(n236), .B(n237), .Z(n235) );
  XOR U605 ( .A(n228), .B(n238), .Z(n237) );
  XNOR U606 ( .A(n240), .B(n241), .Z(n239) );
  NANDN U607 ( .A(n242), .B(n243), .Z(n241) );
  XOR U608 ( .A(n245), .B(n246), .Z(n234) );
  XOR U609 ( .A(key[597]), .B(n247), .Z(n246) );
  ANDN U610 ( .B(n248), .A(n249), .Z(n245) );
  XNOR U611 ( .A(n250), .B(n251), .Z(out[84]) );
  XNOR U612 ( .A(key[596]), .B(n252), .Z(n251) );
  XOR U613 ( .A(n253), .B(n254), .Z(out[83]) );
  XNOR U614 ( .A(n255), .B(n231), .Z(n254) );
  XNOR U615 ( .A(n256), .B(n257), .Z(n231) );
  XNOR U616 ( .A(n258), .B(n247), .Z(n257) );
  ANDN U617 ( .B(n259), .A(n260), .Z(n247) );
  NOR U618 ( .A(n261), .B(n262), .Z(n258) );
  XNOR U619 ( .A(n263), .B(n264), .Z(n253) );
  XOR U620 ( .A(key[595]), .B(n265), .Z(n264) );
  XOR U621 ( .A(key[594]), .B(n250), .Z(out[82]) );
  XNOR U622 ( .A(n230), .B(n266), .Z(n250) );
  IV U623 ( .A(n265), .Z(n230) );
  XOR U624 ( .A(n267), .B(n227), .Z(out[81]) );
  XNOR U625 ( .A(n256), .B(n268), .Z(n255) );
  XNOR U626 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U627 ( .A(n271), .B(n243), .Z(n270) );
  XNOR U628 ( .A(n238), .B(n272), .Z(n256) );
  XNOR U629 ( .A(n273), .B(n274), .Z(n272) );
  NANDN U630 ( .A(n275), .B(n276), .Z(n274) );
  XOR U631 ( .A(n266), .B(n263), .Z(n233) );
  XNOR U632 ( .A(n238), .B(n277), .Z(n263) );
  XNOR U633 ( .A(n269), .B(n278), .Z(n277) );
  NANDN U634 ( .A(n279), .B(n280), .Z(n278) );
  OR U635 ( .A(n281), .B(n282), .Z(n269) );
  XOR U636 ( .A(n283), .B(n273), .Z(n238) );
  NANDN U637 ( .A(n284), .B(n285), .Z(n273) );
  ANDN U638 ( .B(n286), .A(n287), .Z(n283) );
  XOR U639 ( .A(key[593]), .B(n265), .Z(n267) );
  XOR U640 ( .A(n288), .B(n289), .Z(n265) );
  XNOR U641 ( .A(n290), .B(n291), .Z(n289) );
  NAND U642 ( .A(n248), .B(n292), .Z(n291) );
  XNOR U643 ( .A(n236), .B(n293), .Z(out[80]) );
  XOR U644 ( .A(key[592]), .B(n266), .Z(n293) );
  XNOR U645 ( .A(n288), .B(n294), .Z(n266) );
  XOR U646 ( .A(n295), .B(n240), .Z(n294) );
  OR U647 ( .A(n296), .B(n281), .Z(n240) );
  XNOR U648 ( .A(n243), .B(n280), .Z(n281) );
  ANDN U649 ( .B(n297), .A(n298), .Z(n295) );
  IV U650 ( .A(n252), .Z(n236) );
  XOR U651 ( .A(n244), .B(n299), .Z(n252) );
  XOR U652 ( .A(n300), .B(n290), .Z(n299) );
  XNOR U653 ( .A(n262), .B(n248), .Z(n259) );
  NOR U654 ( .A(n302), .B(n262), .Z(n300) );
  XNOR U655 ( .A(n288), .B(n303), .Z(n244) );
  XNOR U656 ( .A(n304), .B(n305), .Z(n303) );
  NANDN U657 ( .A(n275), .B(n306), .Z(n305) );
  XOR U658 ( .A(n307), .B(n304), .Z(n288) );
  OR U659 ( .A(n284), .B(n308), .Z(n304) );
  XOR U660 ( .A(n309), .B(n275), .Z(n284) );
  XNOR U661 ( .A(n280), .B(n248), .Z(n275) );
  XOR U662 ( .A(n310), .B(n311), .Z(n248) );
  NANDN U663 ( .A(n312), .B(n313), .Z(n311) );
  IV U664 ( .A(n298), .Z(n280) );
  XNOR U665 ( .A(n314), .B(n315), .Z(n298) );
  NANDN U666 ( .A(n312), .B(n316), .Z(n315) );
  ANDN U667 ( .B(n309), .A(n317), .Z(n307) );
  IV U668 ( .A(n287), .Z(n309) );
  XOR U669 ( .A(n262), .B(n243), .Z(n287) );
  XNOR U670 ( .A(n318), .B(n314), .Z(n243) );
  NANDN U671 ( .A(n319), .B(n320), .Z(n314) );
  XOR U672 ( .A(n316), .B(n321), .Z(n320) );
  ANDN U673 ( .B(n321), .A(n322), .Z(n318) );
  XOR U674 ( .A(n323), .B(n310), .Z(n262) );
  NANDN U675 ( .A(n319), .B(n324), .Z(n310) );
  XOR U676 ( .A(n325), .B(n313), .Z(n324) );
  XNOR U677 ( .A(n326), .B(n327), .Z(n312) );
  XOR U678 ( .A(n328), .B(n329), .Z(n327) );
  XNOR U679 ( .A(n330), .B(n331), .Z(n326) );
  XNOR U680 ( .A(n332), .B(n333), .Z(n331) );
  ANDN U681 ( .B(n325), .A(n329), .Z(n332) );
  ANDN U682 ( .B(n325), .A(n322), .Z(n323) );
  XNOR U683 ( .A(n328), .B(n334), .Z(n322) );
  XOR U684 ( .A(n335), .B(n333), .Z(n334) );
  NAND U685 ( .A(n336), .B(n337), .Z(n333) );
  XNOR U686 ( .A(n330), .B(n313), .Z(n337) );
  IV U687 ( .A(n325), .Z(n330) );
  XNOR U688 ( .A(n316), .B(n329), .Z(n336) );
  IV U689 ( .A(n321), .Z(n329) );
  XOR U690 ( .A(n338), .B(n339), .Z(n321) );
  XNOR U691 ( .A(n340), .B(n341), .Z(n339) );
  XNOR U692 ( .A(n342), .B(n343), .Z(n338) );
  NOR U693 ( .A(n261), .B(n302), .Z(n342) );
  AND U694 ( .A(n313), .B(n316), .Z(n335) );
  XNOR U695 ( .A(n313), .B(n316), .Z(n328) );
  XNOR U696 ( .A(n344), .B(n345), .Z(n316) );
  XNOR U697 ( .A(n346), .B(n341), .Z(n345) );
  XOR U698 ( .A(n347), .B(n348), .Z(n344) );
  XNOR U699 ( .A(n349), .B(n343), .Z(n348) );
  OR U700 ( .A(n260), .B(n301), .Z(n343) );
  XOR U701 ( .A(n302), .B(n292), .Z(n301) );
  XNOR U702 ( .A(n261), .B(n249), .Z(n260) );
  ANDN U703 ( .B(n292), .A(n249), .Z(n349) );
  XNOR U704 ( .A(n350), .B(n351), .Z(n313) );
  XNOR U705 ( .A(n341), .B(n352), .Z(n351) );
  XOR U706 ( .A(n271), .B(n347), .Z(n352) );
  XNOR U707 ( .A(n302), .B(n353), .Z(n341) );
  XNOR U708 ( .A(n354), .B(n355), .Z(n350) );
  XNOR U709 ( .A(n356), .B(n357), .Z(n355) );
  ANDN U710 ( .B(n297), .A(n279), .Z(n356) );
  XNOR U711 ( .A(n358), .B(n359), .Z(n325) );
  XNOR U712 ( .A(n346), .B(n360), .Z(n359) );
  XNOR U713 ( .A(n279), .B(n340), .Z(n360) );
  XOR U714 ( .A(n347), .B(n361), .Z(n340) );
  XNOR U715 ( .A(n362), .B(n363), .Z(n361) );
  NAND U716 ( .A(n306), .B(n276), .Z(n363) );
  XNOR U717 ( .A(n364), .B(n362), .Z(n347) );
  NANDN U718 ( .A(n308), .B(n285), .Z(n362) );
  XOR U719 ( .A(n286), .B(n276), .Z(n285) );
  XNOR U720 ( .A(n365), .B(n249), .Z(n276) );
  XOR U721 ( .A(n317), .B(n306), .Z(n308) );
  XOR U722 ( .A(n297), .B(n292), .Z(n306) );
  ANDN U723 ( .B(n286), .A(n317), .Z(n364) );
  XOR U724 ( .A(n354), .B(n302), .Z(n317) );
  XOR U725 ( .A(n366), .B(n367), .Z(n302) );
  XOR U726 ( .A(n368), .B(n369), .Z(n367) );
  XOR U727 ( .A(n370), .B(n353), .Z(n286) );
  XNOR U728 ( .A(n371), .B(n372), .Z(n249) );
  XNOR U729 ( .A(n373), .B(n369), .Z(n372) );
  XNOR U730 ( .A(n369), .B(n371), .Z(n292) );
  XNOR U731 ( .A(n297), .B(n374), .Z(n358) );
  XNOR U732 ( .A(n375), .B(n357), .Z(n374) );
  OR U733 ( .A(n282), .B(n296), .Z(n357) );
  XNOR U734 ( .A(n354), .B(n297), .Z(n296) );
  XOR U735 ( .A(n271), .B(n365), .Z(n282) );
  IV U736 ( .A(n279), .Z(n365) );
  XOR U737 ( .A(n353), .B(n376), .Z(n279) );
  XNOR U738 ( .A(n373), .B(n366), .Z(n376) );
  XOR U739 ( .A(key[562]), .B(\w0[4][50] ), .Z(n366) );
  XNOR U740 ( .A(n377), .B(n378), .Z(\w0[4][50] ) );
  XNOR U741 ( .A(n379), .B(n380), .Z(n378) );
  IV U742 ( .A(n261), .Z(n353) );
  XNOR U743 ( .A(n371), .B(n381), .Z(n261) );
  XNOR U744 ( .A(n369), .B(n382), .Z(n381) );
  ANDN U745 ( .B(n370), .A(n242), .Z(n375) );
  IV U746 ( .A(n271), .Z(n370) );
  XNOR U747 ( .A(n371), .B(n383), .Z(n271) );
  XNOR U748 ( .A(n369), .B(n384), .Z(n383) );
  XOR U749 ( .A(n242), .B(n385), .Z(n369) );
  XOR U750 ( .A(key[566]), .B(\w0[4][54] ), .Z(n385) );
  XNOR U751 ( .A(n386), .B(n387), .Z(\w0[4][54] ) );
  XNOR U752 ( .A(n388), .B(n389), .Z(n387) );
  IV U753 ( .A(n354), .Z(n242) );
  XOR U754 ( .A(key[565]), .B(\w0[4][53] ), .Z(n371) );
  XNOR U755 ( .A(n390), .B(n391), .Z(\w0[4][53] ) );
  XOR U756 ( .A(n392), .B(n393), .Z(n391) );
  XOR U757 ( .A(n394), .B(n395), .Z(n297) );
  XNOR U758 ( .A(n384), .B(n382), .Z(n395) );
  XOR U759 ( .A(key[567]), .B(\w0[4][55] ), .Z(n382) );
  XNOR U760 ( .A(n396), .B(n397), .Z(\w0[4][55] ) );
  XOR U761 ( .A(n398), .B(n399), .Z(n397) );
  XOR U762 ( .A(key[564]), .B(\w0[4][52] ), .Z(n384) );
  XOR U763 ( .A(n400), .B(n401), .Z(\w0[4][52] ) );
  XNOR U764 ( .A(n402), .B(n403), .Z(n401) );
  XOR U765 ( .A(n404), .B(n405), .Z(n400) );
  XNOR U766 ( .A(n354), .B(n368), .Z(n394) );
  XOR U767 ( .A(n373), .B(n406), .Z(n368) );
  XOR U768 ( .A(key[563]), .B(\w0[4][51] ), .Z(n406) );
  XOR U769 ( .A(n407), .B(n408), .Z(\w0[4][51] ) );
  XNOR U770 ( .A(n409), .B(n410), .Z(n408) );
  XOR U771 ( .A(n411), .B(n412), .Z(n407) );
  XOR U772 ( .A(key[561]), .B(\w0[4][49] ), .Z(n373) );
  XNOR U773 ( .A(n413), .B(n414), .Z(\w0[4][49] ) );
  XOR U774 ( .A(n415), .B(n416), .Z(n414) );
  XOR U775 ( .A(key[560]), .B(\w0[4][48] ), .Z(n354) );
  XOR U776 ( .A(n417), .B(n418), .Z(\w0[4][48] ) );
  XNOR U777 ( .A(n419), .B(n420), .Z(n418) );
  XOR U778 ( .A(n421), .B(n422), .Z(out[7]) );
  XOR U779 ( .A(n423), .B(n424), .Z(n421) );
  XOR U780 ( .A(key[519]), .B(n425), .Z(n424) );
  XOR U781 ( .A(n426), .B(n427), .Z(out[79]) );
  XOR U782 ( .A(n428), .B(n429), .Z(n426) );
  XNOR U783 ( .A(key[591]), .B(n430), .Z(n429) );
  XOR U784 ( .A(n431), .B(n432), .Z(out[78]) );
  XNOR U785 ( .A(n433), .B(n434), .Z(n432) );
  XNOR U786 ( .A(key[590]), .B(n435), .Z(n431) );
  XOR U787 ( .A(n436), .B(n437), .Z(out[77]) );
  XNOR U788 ( .A(n438), .B(n439), .Z(n437) );
  XOR U789 ( .A(n428), .B(n440), .Z(n439) );
  XNOR U790 ( .A(n442), .B(n443), .Z(n441) );
  OR U791 ( .A(n444), .B(n445), .Z(n443) );
  XOR U792 ( .A(n447), .B(n448), .Z(n436) );
  XOR U793 ( .A(key[589]), .B(n449), .Z(n448) );
  ANDN U794 ( .B(n450), .A(n451), .Z(n447) );
  XNOR U795 ( .A(n452), .B(n453), .Z(out[76]) );
  XNOR U796 ( .A(key[588]), .B(n454), .Z(n453) );
  XOR U797 ( .A(n455), .B(n456), .Z(out[75]) );
  XNOR U798 ( .A(n457), .B(n434), .Z(n456) );
  XNOR U799 ( .A(n458), .B(n459), .Z(n434) );
  XNOR U800 ( .A(n460), .B(n449), .Z(n459) );
  NOR U801 ( .A(n461), .B(n462), .Z(n449) );
  NOR U802 ( .A(n463), .B(n464), .Z(n460) );
  XOR U803 ( .A(n465), .B(n466), .Z(n455) );
  XOR U804 ( .A(key[587]), .B(n467), .Z(n466) );
  XOR U805 ( .A(key[586]), .B(n452), .Z(out[74]) );
  XNOR U806 ( .A(n430), .B(n435), .Z(n452) );
  XOR U807 ( .A(n468), .B(n427), .Z(out[73]) );
  XNOR U808 ( .A(n458), .B(n470), .Z(n457) );
  XOR U809 ( .A(n471), .B(n472), .Z(n470) );
  ANDN U810 ( .B(n473), .A(n444), .Z(n471) );
  XNOR U811 ( .A(n440), .B(n474), .Z(n458) );
  XNOR U812 ( .A(n475), .B(n476), .Z(n474) );
  NAND U813 ( .A(n477), .B(n478), .Z(n476) );
  XOR U814 ( .A(n435), .B(n465), .Z(n469) );
  IV U815 ( .A(n433), .Z(n465) );
  XNOR U816 ( .A(n440), .B(n479), .Z(n433) );
  XNOR U817 ( .A(n472), .B(n480), .Z(n479) );
  NANDN U818 ( .A(n481), .B(n482), .Z(n480) );
  OR U819 ( .A(n483), .B(n484), .Z(n472) );
  XOR U820 ( .A(n485), .B(n475), .Z(n440) );
  NANDN U821 ( .A(n486), .B(n487), .Z(n475) );
  AND U822 ( .A(n488), .B(n489), .Z(n485) );
  XNOR U823 ( .A(key[585]), .B(n430), .Z(n468) );
  IV U824 ( .A(n467), .Z(n430) );
  XOR U825 ( .A(n490), .B(n491), .Z(n467) );
  XNOR U826 ( .A(n492), .B(n493), .Z(n491) );
  NANDN U827 ( .A(n451), .B(n494), .Z(n493) );
  XNOR U828 ( .A(n438), .B(n495), .Z(out[72]) );
  XOR U829 ( .A(key[584]), .B(n435), .Z(n495) );
  XNOR U830 ( .A(n490), .B(n496), .Z(n435) );
  XOR U831 ( .A(n497), .B(n442), .Z(n496) );
  OR U832 ( .A(n498), .B(n483), .Z(n442) );
  XNOR U833 ( .A(n444), .B(n481), .Z(n483) );
  NOR U834 ( .A(n499), .B(n481), .Z(n497) );
  IV U835 ( .A(n454), .Z(n438) );
  XOR U836 ( .A(n446), .B(n500), .Z(n454) );
  XNOR U837 ( .A(n492), .B(n501), .Z(n500) );
  OR U838 ( .A(n464), .B(n502), .Z(n501) );
  OR U839 ( .A(n503), .B(n461), .Z(n492) );
  XOR U840 ( .A(n464), .B(n504), .Z(n461) );
  XNOR U841 ( .A(n490), .B(n505), .Z(n446) );
  XNOR U842 ( .A(n506), .B(n507), .Z(n505) );
  NAND U843 ( .A(n478), .B(n508), .Z(n507) );
  XOR U844 ( .A(n509), .B(n506), .Z(n490) );
  OR U845 ( .A(n486), .B(n510), .Z(n506) );
  XNOR U846 ( .A(n488), .B(n478), .Z(n486) );
  XOR U847 ( .A(n481), .B(n451), .Z(n478) );
  IV U848 ( .A(n504), .Z(n451) );
  XOR U849 ( .A(n511), .B(n512), .Z(n504) );
  NANDN U850 ( .A(n513), .B(n514), .Z(n512) );
  XNOR U851 ( .A(n515), .B(n516), .Z(n481) );
  OR U852 ( .A(n513), .B(n517), .Z(n516) );
  ANDN U853 ( .B(n488), .A(n518), .Z(n509) );
  XOR U854 ( .A(n444), .B(n464), .Z(n488) );
  XNOR U855 ( .A(n511), .B(n519), .Z(n464) );
  NANDN U856 ( .A(n520), .B(n521), .Z(n519) );
  NANDN U857 ( .A(n522), .B(n523), .Z(n511) );
  OR U858 ( .A(n525), .B(n522), .Z(n515) );
  XOR U859 ( .A(n526), .B(n513), .Z(n522) );
  XNOR U860 ( .A(n527), .B(n528), .Z(n513) );
  XOR U861 ( .A(n529), .B(n521), .Z(n528) );
  XNOR U862 ( .A(n530), .B(n531), .Z(n527) );
  XNOR U863 ( .A(n532), .B(n533), .Z(n531) );
  ANDN U864 ( .B(n521), .A(n534), .Z(n532) );
  IV U865 ( .A(n535), .Z(n521) );
  ANDN U866 ( .B(n526), .A(n534), .Z(n524) );
  IV U867 ( .A(n520), .Z(n526) );
  XNOR U868 ( .A(n529), .B(n536), .Z(n520) );
  XNOR U869 ( .A(n533), .B(n537), .Z(n536) );
  NANDN U870 ( .A(n517), .B(n514), .Z(n537) );
  NANDN U871 ( .A(n525), .B(n523), .Z(n533) );
  XNOR U872 ( .A(n514), .B(n535), .Z(n523) );
  XOR U873 ( .A(n538), .B(n539), .Z(n535) );
  XOR U874 ( .A(n540), .B(n541), .Z(n539) );
  XNOR U875 ( .A(n482), .B(n542), .Z(n541) );
  XNOR U876 ( .A(n543), .B(n544), .Z(n538) );
  XNOR U877 ( .A(n545), .B(n546), .Z(n544) );
  ANDN U878 ( .B(n473), .A(n445), .Z(n545) );
  XNOR U879 ( .A(n534), .B(n517), .Z(n525) );
  IV U880 ( .A(n530), .Z(n534) );
  XOR U881 ( .A(n547), .B(n548), .Z(n530) );
  XNOR U882 ( .A(n549), .B(n542), .Z(n548) );
  XOR U883 ( .A(n550), .B(n551), .Z(n542) );
  XNOR U884 ( .A(n552), .B(n553), .Z(n551) );
  NAND U885 ( .A(n508), .B(n477), .Z(n553) );
  XNOR U886 ( .A(n554), .B(n555), .Z(n547) );
  ANDN U887 ( .B(n556), .A(n502), .Z(n554) );
  XOR U888 ( .A(n517), .B(n514), .Z(n529) );
  XNOR U889 ( .A(n557), .B(n558), .Z(n514) );
  XNOR U890 ( .A(n550), .B(n559), .Z(n558) );
  XNOR U891 ( .A(n549), .B(n473), .Z(n559) );
  XNOR U892 ( .A(n560), .B(n561), .Z(n557) );
  XNOR U893 ( .A(n562), .B(n546), .Z(n561) );
  OR U894 ( .A(n484), .B(n498), .Z(n546) );
  XNOR U895 ( .A(n560), .B(n543), .Z(n498) );
  XNOR U896 ( .A(n473), .B(n482), .Z(n484) );
  ANDN U897 ( .B(n482), .A(n499), .Z(n562) );
  XOR U898 ( .A(n563), .B(n564), .Z(n517) );
  XOR U899 ( .A(n550), .B(n540), .Z(n564) );
  XNOR U900 ( .A(n494), .B(n450), .Z(n540) );
  XOR U901 ( .A(n565), .B(n552), .Z(n550) );
  NANDN U902 ( .A(n510), .B(n487), .Z(n552) );
  XOR U903 ( .A(n489), .B(n477), .Z(n487) );
  XOR U904 ( .A(n450), .B(n482), .Z(n477) );
  XNOR U905 ( .A(n556), .B(n566), .Z(n482) );
  XNOR U906 ( .A(n567), .B(n568), .Z(n566) );
  XOR U907 ( .A(n518), .B(n508), .Z(n510) );
  XNOR U908 ( .A(n499), .B(n494), .Z(n508) );
  IV U909 ( .A(n543), .Z(n499) );
  XOR U910 ( .A(n569), .B(n570), .Z(n543) );
  XNOR U911 ( .A(n571), .B(n572), .Z(n570) );
  XNOR U912 ( .A(n560), .B(n573), .Z(n569) );
  ANDN U913 ( .B(n489), .A(n518), .Z(n565) );
  XNOR U914 ( .A(n560), .B(n574), .Z(n518) );
  XOR U915 ( .A(n556), .B(n473), .Z(n489) );
  XNOR U916 ( .A(n575), .B(n576), .Z(n473) );
  XOR U917 ( .A(n577), .B(n572), .Z(n576) );
  XNOR U918 ( .A(key[524]), .B(\w0[4][12] ), .Z(n572) );
  XNOR U919 ( .A(n578), .B(n579), .Z(\w0[4][12] ) );
  XOR U920 ( .A(n580), .B(n581), .Z(n579) );
  XOR U921 ( .A(n549), .B(n582), .Z(n563) );
  XNOR U922 ( .A(n583), .B(n555), .Z(n582) );
  OR U923 ( .A(n462), .B(n503), .Z(n555) );
  XNOR U924 ( .A(n574), .B(n494), .Z(n503) );
  XNOR U925 ( .A(n556), .B(n450), .Z(n462) );
  IV U926 ( .A(n463), .Z(n556) );
  AND U927 ( .A(n450), .B(n494), .Z(n583) );
  XOR U928 ( .A(n577), .B(n575), .Z(n494) );
  XNOR U929 ( .A(n575), .B(n584), .Z(n450) );
  XOR U930 ( .A(n567), .B(n585), .Z(n584) );
  XNOR U931 ( .A(n502), .B(n463), .Z(n549) );
  XOR U932 ( .A(n575), .B(n586), .Z(n463) );
  XOR U933 ( .A(n577), .B(n571), .Z(n586) );
  XNOR U934 ( .A(key[527]), .B(\w0[4][15] ), .Z(n571) );
  XNOR U935 ( .A(n587), .B(n588), .Z(\w0[4][15] ) );
  XOR U936 ( .A(n589), .B(n590), .Z(n588) );
  XNOR U937 ( .A(key[525]), .B(\w0[4][13] ), .Z(n575) );
  XOR U938 ( .A(n591), .B(n592), .Z(\w0[4][13] ) );
  XOR U939 ( .A(n593), .B(n594), .Z(n592) );
  XNOR U940 ( .A(n595), .B(n596), .Z(n591) );
  IV U941 ( .A(n574), .Z(n502) );
  XNOR U942 ( .A(n568), .B(n597), .Z(n574) );
  XNOR U943 ( .A(n573), .B(n585), .Z(n597) );
  IV U944 ( .A(n577), .Z(n585) );
  XOR U945 ( .A(n445), .B(n598), .Z(n577) );
  XOR U946 ( .A(key[526]), .B(\w0[4][14] ), .Z(n598) );
  XNOR U947 ( .A(n599), .B(n600), .Z(\w0[4][14] ) );
  XNOR U948 ( .A(n601), .B(n602), .Z(n600) );
  IV U949 ( .A(n560), .Z(n445) );
  XOR U950 ( .A(key[520]), .B(\w0[4][8] ), .Z(n560) );
  XOR U951 ( .A(n603), .B(n604), .Z(\w0[4][8] ) );
  XNOR U952 ( .A(n605), .B(n606), .Z(n604) );
  XNOR U953 ( .A(n607), .B(n608), .Z(n603) );
  XOR U954 ( .A(n567), .B(n609), .Z(n573) );
  XOR U955 ( .A(key[523]), .B(\w0[4][11] ), .Z(n609) );
  XOR U956 ( .A(n610), .B(n611), .Z(\w0[4][11] ) );
  XNOR U957 ( .A(n612), .B(n613), .Z(n611) );
  XNOR U958 ( .A(n614), .B(n615), .Z(n610) );
  XOR U959 ( .A(key[521]), .B(\w0[4][9] ), .Z(n567) );
  XOR U960 ( .A(n616), .B(n617), .Z(\w0[4][9] ) );
  XOR U961 ( .A(n618), .B(n619), .Z(n617) );
  XNOR U962 ( .A(n620), .B(n621), .Z(n616) );
  XOR U963 ( .A(key[522]), .B(\w0[4][10] ), .Z(n568) );
  XOR U964 ( .A(n622), .B(n623), .Z(\w0[4][10] ) );
  XNOR U965 ( .A(n624), .B(n625), .Z(n623) );
  XNOR U966 ( .A(n626), .B(n627), .Z(n622) );
  XOR U967 ( .A(n628), .B(n629), .Z(out[71]) );
  XNOR U968 ( .A(n630), .B(n631), .Z(n628) );
  XNOR U969 ( .A(key[583]), .B(n632), .Z(n631) );
  XOR U970 ( .A(n633), .B(n634), .Z(out[70]) );
  XNOR U971 ( .A(n635), .B(n636), .Z(n634) );
  XNOR U972 ( .A(key[582]), .B(n637), .Z(n633) );
  XNOR U973 ( .A(n638), .B(n639), .Z(out[6]) );
  XNOR U974 ( .A(key[518]), .B(n640), .Z(n639) );
  XOR U975 ( .A(n641), .B(n642), .Z(out[69]) );
  XNOR U976 ( .A(n643), .B(n644), .Z(n642) );
  XNOR U977 ( .A(n632), .B(n645), .Z(n644) );
  XNOR U978 ( .A(n646), .B(n647), .Z(n632) );
  XNOR U979 ( .A(n648), .B(n649), .Z(n647) );
  OR U980 ( .A(n650), .B(n651), .Z(n649) );
  XNOR U981 ( .A(n652), .B(n653), .Z(n641) );
  XOR U982 ( .A(key[581]), .B(n654), .Z(n653) );
  ANDN U983 ( .B(n655), .A(n656), .Z(n654) );
  XNOR U984 ( .A(n657), .B(n658), .Z(out[68]) );
  XNOR U985 ( .A(key[580]), .B(n659), .Z(n658) );
  XOR U986 ( .A(n660), .B(n661), .Z(out[67]) );
  XNOR U987 ( .A(n662), .B(n636), .Z(n661) );
  XNOR U988 ( .A(n663), .B(n664), .Z(n636) );
  XNOR U989 ( .A(n652), .B(n665), .Z(n664) );
  OR U990 ( .A(n666), .B(n667), .Z(n665) );
  NANDN U991 ( .A(n668), .B(n669), .Z(n652) );
  XNOR U992 ( .A(n670), .B(n671), .Z(n660) );
  XNOR U993 ( .A(key[579]), .B(n635), .Z(n671) );
  XOR U994 ( .A(key[578]), .B(n657), .Z(out[66]) );
  XNOR U995 ( .A(n637), .B(n662), .Z(n657) );
  XOR U996 ( .A(n672), .B(n629), .Z(out[65]) );
  XNOR U997 ( .A(n670), .B(n662), .Z(n629) );
  XNOR U998 ( .A(n673), .B(n674), .Z(n662) );
  XNOR U999 ( .A(n675), .B(n676), .Z(n674) );
  NAND U1000 ( .A(n677), .B(n655), .Z(n676) );
  XNOR U1001 ( .A(n663), .B(n678), .Z(n670) );
  XNOR U1002 ( .A(n679), .B(n680), .Z(n678) );
  NANDN U1003 ( .A(n650), .B(n681), .Z(n680) );
  XNOR U1004 ( .A(n645), .B(n682), .Z(n663) );
  XNOR U1005 ( .A(n683), .B(n684), .Z(n682) );
  NANDN U1006 ( .A(n685), .B(n686), .Z(n684) );
  XNOR U1007 ( .A(key[577]), .B(n630), .Z(n672) );
  XOR U1008 ( .A(n687), .B(n635), .Z(n630) );
  XNOR U1009 ( .A(n645), .B(n688), .Z(n635) );
  XOR U1010 ( .A(n689), .B(n679), .Z(n688) );
  OR U1011 ( .A(n690), .B(n691), .Z(n679) );
  AND U1012 ( .A(n692), .B(n693), .Z(n689) );
  XOR U1013 ( .A(n694), .B(n683), .Z(n645) );
  NANDN U1014 ( .A(n695), .B(n696), .Z(n683) );
  AND U1015 ( .A(n697), .B(n698), .Z(n694) );
  XNOR U1016 ( .A(n643), .B(n699), .Z(out[64]) );
  XNOR U1017 ( .A(key[576]), .B(n687), .Z(n699) );
  IV U1018 ( .A(n637), .Z(n687) );
  XNOR U1019 ( .A(n673), .B(n700), .Z(n637) );
  XOR U1020 ( .A(n701), .B(n648), .Z(n700) );
  OR U1021 ( .A(n702), .B(n690), .Z(n648) );
  XOR U1022 ( .A(n650), .B(n693), .Z(n690) );
  ANDN U1023 ( .B(n693), .A(n703), .Z(n701) );
  IV U1024 ( .A(n659), .Z(n643) );
  XOR U1025 ( .A(n646), .B(n704), .Z(n659) );
  XOR U1026 ( .A(n705), .B(n675), .Z(n704) );
  NANDN U1027 ( .A(n706), .B(n669), .Z(n675) );
  XNOR U1028 ( .A(n666), .B(n655), .Z(n669) );
  NOR U1029 ( .A(n707), .B(n666), .Z(n705) );
  XNOR U1030 ( .A(n673), .B(n708), .Z(n646) );
  XNOR U1031 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U1032 ( .A(n685), .B(n711), .Z(n710) );
  XOR U1033 ( .A(n712), .B(n709), .Z(n673) );
  OR U1034 ( .A(n695), .B(n713), .Z(n709) );
  XOR U1035 ( .A(n697), .B(n685), .Z(n695) );
  XNOR U1036 ( .A(n693), .B(n655), .Z(n685) );
  XOR U1037 ( .A(n714), .B(n715), .Z(n655) );
  NANDN U1038 ( .A(n716), .B(n717), .Z(n715) );
  XOR U1039 ( .A(n718), .B(n719), .Z(n693) );
  OR U1040 ( .A(n716), .B(n720), .Z(n719) );
  ANDN U1041 ( .B(n697), .A(n721), .Z(n712) );
  XOR U1042 ( .A(n650), .B(n666), .Z(n697) );
  XOR U1043 ( .A(n722), .B(n714), .Z(n666) );
  NANDN U1044 ( .A(n723), .B(n724), .Z(n714) );
  ANDN U1045 ( .B(n725), .A(n726), .Z(n722) );
  NANDN U1046 ( .A(n723), .B(n728), .Z(n718) );
  XOR U1047 ( .A(n729), .B(n716), .Z(n723) );
  XNOR U1048 ( .A(n730), .B(n731), .Z(n716) );
  XOR U1049 ( .A(n732), .B(n725), .Z(n731) );
  XNOR U1050 ( .A(n733), .B(n734), .Z(n730) );
  XNOR U1051 ( .A(n735), .B(n736), .Z(n734) );
  ANDN U1052 ( .B(n725), .A(n737), .Z(n735) );
  IV U1053 ( .A(n738), .Z(n725) );
  ANDN U1054 ( .B(n729), .A(n737), .Z(n727) );
  IV U1055 ( .A(n733), .Z(n737) );
  IV U1056 ( .A(n726), .Z(n729) );
  XNOR U1057 ( .A(n732), .B(n739), .Z(n726) );
  XOR U1058 ( .A(n740), .B(n736), .Z(n739) );
  NAND U1059 ( .A(n728), .B(n724), .Z(n736) );
  XNOR U1060 ( .A(n717), .B(n738), .Z(n724) );
  XOR U1061 ( .A(n741), .B(n742), .Z(n738) );
  XOR U1062 ( .A(n743), .B(n744), .Z(n742) );
  XNOR U1063 ( .A(n692), .B(n745), .Z(n744) );
  XNOR U1064 ( .A(n746), .B(n747), .Z(n741) );
  XNOR U1065 ( .A(n748), .B(n749), .Z(n747) );
  ANDN U1066 ( .B(n681), .A(n651), .Z(n748) );
  XNOR U1067 ( .A(n733), .B(n720), .Z(n728) );
  XOR U1068 ( .A(n750), .B(n751), .Z(n733) );
  XNOR U1069 ( .A(n752), .B(n745), .Z(n751) );
  XOR U1070 ( .A(n753), .B(n754), .Z(n745) );
  XNOR U1071 ( .A(n755), .B(n756), .Z(n754) );
  NAND U1072 ( .A(n711), .B(n686), .Z(n756) );
  XNOR U1073 ( .A(n757), .B(n758), .Z(n750) );
  ANDN U1074 ( .B(n759), .A(n707), .Z(n757) );
  ANDN U1075 ( .B(n717), .A(n720), .Z(n740) );
  XOR U1076 ( .A(n720), .B(n717), .Z(n732) );
  XNOR U1077 ( .A(n760), .B(n761), .Z(n717) );
  XNOR U1078 ( .A(n753), .B(n762), .Z(n761) );
  XNOR U1079 ( .A(n752), .B(n681), .Z(n762) );
  XNOR U1080 ( .A(n763), .B(n764), .Z(n760) );
  XNOR U1081 ( .A(n765), .B(n749), .Z(n764) );
  OR U1082 ( .A(n691), .B(n702), .Z(n749) );
  XNOR U1083 ( .A(n763), .B(n746), .Z(n702) );
  XNOR U1084 ( .A(n681), .B(n692), .Z(n691) );
  ANDN U1085 ( .B(n692), .A(n703), .Z(n765) );
  XOR U1086 ( .A(n766), .B(n767), .Z(n720) );
  XOR U1087 ( .A(n753), .B(n743), .Z(n767) );
  XOR U1088 ( .A(n677), .B(n656), .Z(n743) );
  XOR U1089 ( .A(n768), .B(n755), .Z(n753) );
  NANDN U1090 ( .A(n713), .B(n696), .Z(n755) );
  XOR U1091 ( .A(n698), .B(n686), .Z(n696) );
  XNOR U1092 ( .A(n759), .B(n769), .Z(n692) );
  XOR U1093 ( .A(n770), .B(n771), .Z(n769) );
  XOR U1094 ( .A(n721), .B(n711), .Z(n713) );
  XNOR U1095 ( .A(n703), .B(n677), .Z(n711) );
  IV U1096 ( .A(n746), .Z(n703) );
  XOR U1097 ( .A(n772), .B(n773), .Z(n746) );
  XNOR U1098 ( .A(n774), .B(n775), .Z(n773) );
  XNOR U1099 ( .A(n763), .B(n776), .Z(n772) );
  ANDN U1100 ( .B(n698), .A(n721), .Z(n768) );
  XNOR U1101 ( .A(n763), .B(n777), .Z(n721) );
  XOR U1102 ( .A(n759), .B(n681), .Z(n698) );
  XNOR U1103 ( .A(n778), .B(n779), .Z(n681) );
  XNOR U1104 ( .A(n780), .B(n775), .Z(n779) );
  XOR U1105 ( .A(key[612]), .B(\w0[4][100] ), .Z(n775) );
  XOR U1106 ( .A(n781), .B(n782), .Z(\w0[4][100] ) );
  XNOR U1107 ( .A(n783), .B(n784), .Z(n782) );
  XOR U1108 ( .A(n785), .B(n786), .Z(n781) );
  IV U1109 ( .A(n667), .Z(n759) );
  XOR U1110 ( .A(n752), .B(n787), .Z(n766) );
  XNOR U1111 ( .A(n788), .B(n758), .Z(n787) );
  OR U1112 ( .A(n668), .B(n706), .Z(n758) );
  XNOR U1113 ( .A(n777), .B(n677), .Z(n706) );
  XNOR U1114 ( .A(n667), .B(n656), .Z(n668) );
  ANDN U1115 ( .B(n677), .A(n656), .Z(n788) );
  XOR U1116 ( .A(n778), .B(n789), .Z(n656) );
  XNOR U1117 ( .A(n790), .B(n780), .Z(n789) );
  XOR U1118 ( .A(n780), .B(n778), .Z(n677) );
  XNOR U1119 ( .A(n707), .B(n667), .Z(n752) );
  XOR U1120 ( .A(n778), .B(n791), .Z(n667) );
  XNOR U1121 ( .A(n780), .B(n774), .Z(n791) );
  XOR U1122 ( .A(key[615]), .B(\w0[4][103] ), .Z(n774) );
  XNOR U1123 ( .A(n792), .B(n793), .Z(\w0[4][103] ) );
  XOR U1124 ( .A(n794), .B(n795), .Z(n793) );
  XNOR U1125 ( .A(key[613]), .B(\w0[4][101] ), .Z(n778) );
  XNOR U1126 ( .A(n796), .B(n797), .Z(\w0[4][101] ) );
  XOR U1127 ( .A(n798), .B(n799), .Z(n797) );
  IV U1128 ( .A(n777), .Z(n707) );
  XOR U1129 ( .A(n770), .B(n776), .Z(n800) );
  XNOR U1130 ( .A(n771), .B(n801), .Z(n776) );
  XOR U1131 ( .A(key[611]), .B(\w0[4][99] ), .Z(n801) );
  XOR U1132 ( .A(n802), .B(n803), .Z(\w0[4][99] ) );
  XOR U1133 ( .A(n804), .B(n805), .Z(n803) );
  XOR U1134 ( .A(n806), .B(n807), .Z(n802) );
  IV U1135 ( .A(n790), .Z(n771) );
  XOR U1136 ( .A(key[609]), .B(\w0[4][97] ), .Z(n790) );
  XNOR U1137 ( .A(n808), .B(n809), .Z(\w0[4][97] ) );
  XNOR U1138 ( .A(n810), .B(n811), .Z(n809) );
  XOR U1139 ( .A(key[610]), .B(\w0[4][98] ), .Z(n770) );
  XNOR U1140 ( .A(n812), .B(n813), .Z(\w0[4][98] ) );
  XNOR U1141 ( .A(n814), .B(n815), .Z(n813) );
  XOR U1142 ( .A(n651), .B(n816), .Z(n780) );
  XOR U1143 ( .A(key[614]), .B(\w0[4][102] ), .Z(n816) );
  XNOR U1144 ( .A(n817), .B(n818), .Z(\w0[4][102] ) );
  XNOR U1145 ( .A(n819), .B(n820), .Z(n818) );
  IV U1146 ( .A(n763), .Z(n651) );
  XOR U1147 ( .A(key[608]), .B(\w0[4][96] ), .Z(n763) );
  XNOR U1148 ( .A(n821), .B(n822), .Z(\w0[4][96] ) );
  XOR U1149 ( .A(n823), .B(n824), .Z(n822) );
  XOR U1150 ( .A(n825), .B(n826), .Z(out[63]) );
  XOR U1151 ( .A(n827), .B(n828), .Z(n825) );
  XOR U1152 ( .A(key[575]), .B(n829), .Z(n828) );
  XNOR U1153 ( .A(n830), .B(n831), .Z(out[62]) );
  XNOR U1154 ( .A(key[574]), .B(n832), .Z(n831) );
  XOR U1155 ( .A(n833), .B(n834), .Z(out[61]) );
  XNOR U1156 ( .A(n835), .B(n836), .Z(n834) );
  XOR U1157 ( .A(n827), .B(n837), .Z(n836) );
  XNOR U1158 ( .A(n839), .B(n840), .Z(n838) );
  NANDN U1159 ( .A(n841), .B(n842), .Z(n840) );
  XOR U1160 ( .A(n844), .B(n845), .Z(n833) );
  XOR U1161 ( .A(key[573]), .B(n846), .Z(n845) );
  ANDN U1162 ( .B(n847), .A(n848), .Z(n844) );
  XNOR U1163 ( .A(n849), .B(n850), .Z(out[60]) );
  XNOR U1164 ( .A(key[572]), .B(n851), .Z(n850) );
  XOR U1165 ( .A(n852), .B(n853), .Z(out[5]) );
  XNOR U1166 ( .A(n854), .B(n855), .Z(n853) );
  XOR U1167 ( .A(n423), .B(n856), .Z(n855) );
  XNOR U1168 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U1169 ( .A(n860), .B(n861), .Z(n859) );
  XOR U1170 ( .A(n863), .B(n864), .Z(n852) );
  XOR U1171 ( .A(key[517]), .B(n865), .Z(n864) );
  ANDN U1172 ( .B(n866), .A(n867), .Z(n863) );
  XOR U1173 ( .A(n868), .B(n869), .Z(out[59]) );
  XNOR U1174 ( .A(n870), .B(n830), .Z(n869) );
  XNOR U1175 ( .A(n871), .B(n872), .Z(n830) );
  XNOR U1176 ( .A(n873), .B(n846), .Z(n872) );
  ANDN U1177 ( .B(n874), .A(n875), .Z(n846) );
  NOR U1178 ( .A(n876), .B(n877), .Z(n873) );
  XNOR U1179 ( .A(n878), .B(n879), .Z(n868) );
  XOR U1180 ( .A(key[571]), .B(n829), .Z(n879) );
  XOR U1181 ( .A(key[570]), .B(n849), .Z(out[58]) );
  XNOR U1182 ( .A(n880), .B(n881), .Z(n849) );
  XOR U1183 ( .A(n882), .B(n826), .Z(out[57]) );
  XNOR U1184 ( .A(n871), .B(n883), .Z(n870) );
  XNOR U1185 ( .A(n884), .B(n885), .Z(n883) );
  NANDN U1186 ( .A(n886), .B(n842), .Z(n885) );
  XNOR U1187 ( .A(n837), .B(n887), .Z(n871) );
  XNOR U1188 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U1189 ( .A(n890), .B(n891), .Z(n889) );
  XOR U1190 ( .A(n881), .B(n878), .Z(n832) );
  XNOR U1191 ( .A(n837), .B(n892), .Z(n878) );
  XNOR U1192 ( .A(n884), .B(n893), .Z(n892) );
  NANDN U1193 ( .A(n894), .B(n895), .Z(n893) );
  OR U1194 ( .A(n896), .B(n897), .Z(n884) );
  XOR U1195 ( .A(n898), .B(n888), .Z(n837) );
  NANDN U1196 ( .A(n899), .B(n900), .Z(n888) );
  ANDN U1197 ( .B(n901), .A(n902), .Z(n898) );
  XNOR U1198 ( .A(key[569]), .B(n880), .Z(n882) );
  IV U1199 ( .A(n829), .Z(n880) );
  XOR U1200 ( .A(n903), .B(n904), .Z(n829) );
  XNOR U1201 ( .A(n905), .B(n906), .Z(n904) );
  NAND U1202 ( .A(n847), .B(n907), .Z(n906) );
  XNOR U1203 ( .A(n835), .B(n908), .Z(out[56]) );
  XOR U1204 ( .A(key[568]), .B(n881), .Z(n908) );
  XNOR U1205 ( .A(n903), .B(n909), .Z(n881) );
  XOR U1206 ( .A(n910), .B(n839), .Z(n909) );
  OR U1207 ( .A(n911), .B(n896), .Z(n839) );
  XNOR U1208 ( .A(n842), .B(n895), .Z(n896) );
  ANDN U1209 ( .B(n912), .A(n913), .Z(n910) );
  IV U1210 ( .A(n851), .Z(n835) );
  XOR U1211 ( .A(n843), .B(n914), .Z(n851) );
  XOR U1212 ( .A(n915), .B(n905), .Z(n914) );
  XNOR U1213 ( .A(n877), .B(n847), .Z(n874) );
  NOR U1214 ( .A(n917), .B(n877), .Z(n915) );
  XNOR U1215 ( .A(n903), .B(n918), .Z(n843) );
  XNOR U1216 ( .A(n919), .B(n920), .Z(n918) );
  NANDN U1217 ( .A(n890), .B(n921), .Z(n920) );
  XOR U1218 ( .A(n922), .B(n919), .Z(n903) );
  OR U1219 ( .A(n899), .B(n923), .Z(n919) );
  XOR U1220 ( .A(n924), .B(n890), .Z(n899) );
  XNOR U1221 ( .A(n895), .B(n847), .Z(n890) );
  XOR U1222 ( .A(n925), .B(n926), .Z(n847) );
  NANDN U1223 ( .A(n927), .B(n928), .Z(n926) );
  IV U1224 ( .A(n913), .Z(n895) );
  XNOR U1225 ( .A(n929), .B(n930), .Z(n913) );
  NANDN U1226 ( .A(n927), .B(n931), .Z(n930) );
  ANDN U1227 ( .B(n924), .A(n932), .Z(n922) );
  IV U1228 ( .A(n902), .Z(n924) );
  XOR U1229 ( .A(n877), .B(n842), .Z(n902) );
  XNOR U1230 ( .A(n933), .B(n929), .Z(n842) );
  NANDN U1231 ( .A(n934), .B(n935), .Z(n929) );
  XOR U1232 ( .A(n931), .B(n936), .Z(n935) );
  ANDN U1233 ( .B(n936), .A(n937), .Z(n933) );
  XOR U1234 ( .A(n938), .B(n925), .Z(n877) );
  NANDN U1235 ( .A(n934), .B(n939), .Z(n925) );
  XOR U1236 ( .A(n940), .B(n928), .Z(n939) );
  XNOR U1237 ( .A(n941), .B(n942), .Z(n927) );
  XOR U1238 ( .A(n943), .B(n944), .Z(n942) );
  XNOR U1239 ( .A(n945), .B(n946), .Z(n941) );
  XNOR U1240 ( .A(n947), .B(n948), .Z(n946) );
  ANDN U1241 ( .B(n940), .A(n944), .Z(n947) );
  ANDN U1242 ( .B(n940), .A(n937), .Z(n938) );
  XNOR U1243 ( .A(n943), .B(n949), .Z(n937) );
  XOR U1244 ( .A(n950), .B(n948), .Z(n949) );
  NAND U1245 ( .A(n951), .B(n952), .Z(n948) );
  XNOR U1246 ( .A(n945), .B(n928), .Z(n952) );
  IV U1247 ( .A(n940), .Z(n945) );
  XNOR U1248 ( .A(n931), .B(n944), .Z(n951) );
  IV U1249 ( .A(n936), .Z(n944) );
  XOR U1250 ( .A(n953), .B(n954), .Z(n936) );
  XNOR U1251 ( .A(n955), .B(n956), .Z(n954) );
  XNOR U1252 ( .A(n957), .B(n958), .Z(n953) );
  NOR U1253 ( .A(n876), .B(n917), .Z(n957) );
  AND U1254 ( .A(n928), .B(n931), .Z(n950) );
  XNOR U1255 ( .A(n928), .B(n931), .Z(n943) );
  XNOR U1256 ( .A(n959), .B(n960), .Z(n931) );
  XNOR U1257 ( .A(n961), .B(n956), .Z(n960) );
  XOR U1258 ( .A(n962), .B(n963), .Z(n959) );
  XNOR U1259 ( .A(n964), .B(n958), .Z(n963) );
  OR U1260 ( .A(n875), .B(n916), .Z(n958) );
  XOR U1261 ( .A(n917), .B(n907), .Z(n916) );
  XNOR U1262 ( .A(n876), .B(n848), .Z(n875) );
  ANDN U1263 ( .B(n907), .A(n848), .Z(n964) );
  XNOR U1264 ( .A(n965), .B(n966), .Z(n928) );
  XNOR U1265 ( .A(n956), .B(n967), .Z(n966) );
  XOR U1266 ( .A(n886), .B(n962), .Z(n967) );
  XNOR U1267 ( .A(n917), .B(n968), .Z(n956) );
  XNOR U1268 ( .A(n969), .B(n970), .Z(n965) );
  XNOR U1269 ( .A(n971), .B(n972), .Z(n970) );
  ANDN U1270 ( .B(n912), .A(n894), .Z(n971) );
  XNOR U1271 ( .A(n973), .B(n974), .Z(n940) );
  XNOR U1272 ( .A(n961), .B(n975), .Z(n974) );
  XNOR U1273 ( .A(n894), .B(n955), .Z(n975) );
  XOR U1274 ( .A(n962), .B(n976), .Z(n955) );
  XNOR U1275 ( .A(n977), .B(n978), .Z(n976) );
  NAND U1276 ( .A(n921), .B(n891), .Z(n978) );
  XNOR U1277 ( .A(n979), .B(n977), .Z(n962) );
  NANDN U1278 ( .A(n923), .B(n900), .Z(n977) );
  XOR U1279 ( .A(n901), .B(n891), .Z(n900) );
  XNOR U1280 ( .A(n980), .B(n848), .Z(n891) );
  XOR U1281 ( .A(n932), .B(n921), .Z(n923) );
  XOR U1282 ( .A(n912), .B(n907), .Z(n921) );
  ANDN U1283 ( .B(n901), .A(n932), .Z(n979) );
  XOR U1284 ( .A(n969), .B(n917), .Z(n932) );
  XOR U1285 ( .A(n981), .B(n982), .Z(n917) );
  XOR U1286 ( .A(n983), .B(n984), .Z(n982) );
  XOR U1287 ( .A(n985), .B(n968), .Z(n901) );
  XNOR U1288 ( .A(n986), .B(n987), .Z(n848) );
  XNOR U1289 ( .A(n988), .B(n984), .Z(n987) );
  XNOR U1290 ( .A(n984), .B(n986), .Z(n907) );
  XNOR U1291 ( .A(n912), .B(n989), .Z(n973) );
  XNOR U1292 ( .A(n990), .B(n972), .Z(n989) );
  OR U1293 ( .A(n897), .B(n911), .Z(n972) );
  XNOR U1294 ( .A(n969), .B(n912), .Z(n911) );
  XOR U1295 ( .A(n886), .B(n980), .Z(n897) );
  IV U1296 ( .A(n894), .Z(n980) );
  XOR U1297 ( .A(n968), .B(n991), .Z(n894) );
  XNOR U1298 ( .A(n988), .B(n981), .Z(n991) );
  XOR U1299 ( .A(key[570]), .B(\w0[4][58] ), .Z(n981) );
  XOR U1300 ( .A(n992), .B(n993), .Z(\w0[4][58] ) );
  XOR U1301 ( .A(n415), .B(n994), .Z(n993) );
  IV U1302 ( .A(n995), .Z(n415) );
  XOR U1303 ( .A(n996), .B(n997), .Z(n992) );
  IV U1304 ( .A(n876), .Z(n968) );
  XNOR U1305 ( .A(n986), .B(n998), .Z(n876) );
  XNOR U1306 ( .A(n984), .B(n999), .Z(n998) );
  ANDN U1307 ( .B(n985), .A(n841), .Z(n990) );
  IV U1308 ( .A(n886), .Z(n985) );
  XNOR U1309 ( .A(n986), .B(n1000), .Z(n886) );
  XNOR U1310 ( .A(n984), .B(n1001), .Z(n1000) );
  XOR U1311 ( .A(n841), .B(n1002), .Z(n984) );
  XOR U1312 ( .A(key[574]), .B(\w0[4][62] ), .Z(n1002) );
  XNOR U1313 ( .A(n389), .B(n1003), .Z(\w0[4][62] ) );
  XNOR U1314 ( .A(n1004), .B(n1005), .Z(n1003) );
  XOR U1315 ( .A(n1006), .B(n398), .Z(n389) );
  IV U1316 ( .A(n969), .Z(n841) );
  XOR U1317 ( .A(key[573]), .B(\w0[4][61] ), .Z(n986) );
  XOR U1318 ( .A(n1007), .B(n1008), .Z(\w0[4][61] ) );
  XOR U1319 ( .A(n1009), .B(n1010), .Z(n1008) );
  XOR U1320 ( .A(n1011), .B(n1012), .Z(n1007) );
  XOR U1321 ( .A(n1013), .B(n1014), .Z(n912) );
  XNOR U1322 ( .A(n1001), .B(n999), .Z(n1014) );
  XOR U1323 ( .A(key[575]), .B(\w0[4][63] ), .Z(n999) );
  XNOR U1324 ( .A(n1015), .B(n1016), .Z(\w0[4][63] ) );
  XNOR U1325 ( .A(n1017), .B(n1018), .Z(n1016) );
  XOR U1326 ( .A(key[572]), .B(\w0[4][60] ), .Z(n1001) );
  XOR U1327 ( .A(n1019), .B(n1020), .Z(\w0[4][60] ) );
  XNOR U1328 ( .A(n1021), .B(n1022), .Z(n1020) );
  XOR U1329 ( .A(n1023), .B(n404), .Z(n1019) );
  XNOR U1330 ( .A(n398), .B(n1024), .Z(n404) );
  XNOR U1331 ( .A(n969), .B(n983), .Z(n1013) );
  XOR U1332 ( .A(n988), .B(n1025), .Z(n983) );
  XOR U1333 ( .A(key[571]), .B(\w0[4][59] ), .Z(n1025) );
  XOR U1334 ( .A(n1026), .B(n1027), .Z(\w0[4][59] ) );
  XOR U1335 ( .A(n1028), .B(n1029), .Z(n1027) );
  XOR U1336 ( .A(n1030), .B(n411), .Z(n1026) );
  XOR U1337 ( .A(n398), .B(n1031), .Z(n411) );
  XOR U1338 ( .A(key[569]), .B(\w0[4][57] ), .Z(n988) );
  XOR U1339 ( .A(n1032), .B(n1033), .Z(\w0[4][57] ) );
  XOR U1340 ( .A(n1034), .B(n420), .Z(n1033) );
  XOR U1341 ( .A(key[568]), .B(\w0[4][56] ), .Z(n969) );
  XOR U1342 ( .A(n1037), .B(n1038), .Z(\w0[4][56] ) );
  XOR U1343 ( .A(n417), .B(n1039), .Z(n1038) );
  XNOR U1344 ( .A(n398), .B(n1040), .Z(n1037) );
  XOR U1345 ( .A(n1041), .B(n1042), .Z(out[55]) );
  XOR U1346 ( .A(n1043), .B(n1044), .Z(n1041) );
  XOR U1347 ( .A(key[567]), .B(n1045), .Z(n1044) );
  XNOR U1348 ( .A(n1046), .B(n1047), .Z(out[54]) );
  XNOR U1349 ( .A(key[566]), .B(n1048), .Z(n1047) );
  XOR U1350 ( .A(n1049), .B(n1050), .Z(out[53]) );
  XNOR U1351 ( .A(n1051), .B(n1052), .Z(n1050) );
  XOR U1352 ( .A(n1043), .B(n1053), .Z(n1052) );
  XNOR U1353 ( .A(n1055), .B(n1056), .Z(n1054) );
  NANDN U1354 ( .A(n1057), .B(n1058), .Z(n1056) );
  XOR U1355 ( .A(n1060), .B(n1061), .Z(n1049) );
  XOR U1356 ( .A(key[565]), .B(n1062), .Z(n1061) );
  ANDN U1357 ( .B(n1063), .A(n1064), .Z(n1060) );
  XNOR U1358 ( .A(n1065), .B(n1066), .Z(out[52]) );
  XNOR U1359 ( .A(key[564]), .B(n1067), .Z(n1066) );
  XOR U1360 ( .A(n1068), .B(n1069), .Z(out[51]) );
  XNOR U1361 ( .A(n1070), .B(n1046), .Z(n1069) );
  XNOR U1362 ( .A(n1071), .B(n1072), .Z(n1046) );
  XNOR U1363 ( .A(n1073), .B(n1062), .Z(n1072) );
  ANDN U1364 ( .B(n1074), .A(n1075), .Z(n1062) );
  NOR U1365 ( .A(n1076), .B(n1077), .Z(n1073) );
  XNOR U1366 ( .A(n1078), .B(n1079), .Z(n1068) );
  XOR U1367 ( .A(key[563]), .B(n1045), .Z(n1079) );
  XOR U1368 ( .A(key[562]), .B(n1065), .Z(out[50]) );
  XNOR U1369 ( .A(n1080), .B(n1081), .Z(n1065) );
  XNOR U1370 ( .A(n1082), .B(n1083), .Z(out[4]) );
  XNOR U1371 ( .A(key[516]), .B(n1084), .Z(n1083) );
  XOR U1372 ( .A(n1085), .B(n1042), .Z(out[49]) );
  XNOR U1373 ( .A(n1071), .B(n1086), .Z(n1070) );
  XNOR U1374 ( .A(n1087), .B(n1088), .Z(n1086) );
  NANDN U1375 ( .A(n1089), .B(n1058), .Z(n1088) );
  XNOR U1376 ( .A(n1053), .B(n1090), .Z(n1071) );
  XNOR U1377 ( .A(n1091), .B(n1092), .Z(n1090) );
  NANDN U1378 ( .A(n1093), .B(n1094), .Z(n1092) );
  XOR U1379 ( .A(n1081), .B(n1078), .Z(n1048) );
  XNOR U1380 ( .A(n1053), .B(n1095), .Z(n1078) );
  XNOR U1381 ( .A(n1087), .B(n1096), .Z(n1095) );
  NANDN U1382 ( .A(n1097), .B(n1098), .Z(n1096) );
  OR U1383 ( .A(n1099), .B(n1100), .Z(n1087) );
  XOR U1384 ( .A(n1101), .B(n1091), .Z(n1053) );
  NANDN U1385 ( .A(n1102), .B(n1103), .Z(n1091) );
  ANDN U1386 ( .B(n1104), .A(n1105), .Z(n1101) );
  XNOR U1387 ( .A(key[561]), .B(n1080), .Z(n1085) );
  IV U1388 ( .A(n1045), .Z(n1080) );
  XOR U1389 ( .A(n1106), .B(n1107), .Z(n1045) );
  XNOR U1390 ( .A(n1108), .B(n1109), .Z(n1107) );
  NAND U1391 ( .A(n1063), .B(n1110), .Z(n1109) );
  XNOR U1392 ( .A(n1051), .B(n1111), .Z(out[48]) );
  XOR U1393 ( .A(key[560]), .B(n1081), .Z(n1111) );
  XNOR U1394 ( .A(n1106), .B(n1112), .Z(n1081) );
  XOR U1395 ( .A(n1113), .B(n1055), .Z(n1112) );
  OR U1396 ( .A(n1114), .B(n1099), .Z(n1055) );
  XNOR U1397 ( .A(n1058), .B(n1098), .Z(n1099) );
  ANDN U1398 ( .B(n1115), .A(n1116), .Z(n1113) );
  IV U1399 ( .A(n1067), .Z(n1051) );
  XOR U1400 ( .A(n1059), .B(n1117), .Z(n1067) );
  XOR U1401 ( .A(n1118), .B(n1108), .Z(n1117) );
  XNOR U1402 ( .A(n1077), .B(n1063), .Z(n1074) );
  NOR U1403 ( .A(n1120), .B(n1077), .Z(n1118) );
  XNOR U1404 ( .A(n1106), .B(n1121), .Z(n1059) );
  XNOR U1405 ( .A(n1122), .B(n1123), .Z(n1121) );
  NANDN U1406 ( .A(n1093), .B(n1124), .Z(n1123) );
  XOR U1407 ( .A(n1125), .B(n1122), .Z(n1106) );
  OR U1408 ( .A(n1102), .B(n1126), .Z(n1122) );
  XOR U1409 ( .A(n1127), .B(n1093), .Z(n1102) );
  XNOR U1410 ( .A(n1098), .B(n1063), .Z(n1093) );
  XOR U1411 ( .A(n1128), .B(n1129), .Z(n1063) );
  NANDN U1412 ( .A(n1130), .B(n1131), .Z(n1129) );
  IV U1413 ( .A(n1116), .Z(n1098) );
  XNOR U1414 ( .A(n1132), .B(n1133), .Z(n1116) );
  NANDN U1415 ( .A(n1130), .B(n1134), .Z(n1133) );
  ANDN U1416 ( .B(n1127), .A(n1135), .Z(n1125) );
  IV U1417 ( .A(n1105), .Z(n1127) );
  XOR U1418 ( .A(n1077), .B(n1058), .Z(n1105) );
  XNOR U1419 ( .A(n1136), .B(n1132), .Z(n1058) );
  NANDN U1420 ( .A(n1137), .B(n1138), .Z(n1132) );
  XOR U1421 ( .A(n1134), .B(n1139), .Z(n1138) );
  ANDN U1422 ( .B(n1139), .A(n1140), .Z(n1136) );
  XOR U1423 ( .A(n1141), .B(n1128), .Z(n1077) );
  NANDN U1424 ( .A(n1137), .B(n1142), .Z(n1128) );
  XOR U1425 ( .A(n1143), .B(n1131), .Z(n1142) );
  XNOR U1426 ( .A(n1144), .B(n1145), .Z(n1130) );
  XOR U1427 ( .A(n1146), .B(n1147), .Z(n1145) );
  XNOR U1428 ( .A(n1148), .B(n1149), .Z(n1144) );
  XNOR U1429 ( .A(n1150), .B(n1151), .Z(n1149) );
  ANDN U1430 ( .B(n1143), .A(n1147), .Z(n1150) );
  ANDN U1431 ( .B(n1143), .A(n1140), .Z(n1141) );
  XNOR U1432 ( .A(n1146), .B(n1152), .Z(n1140) );
  XOR U1433 ( .A(n1153), .B(n1151), .Z(n1152) );
  NAND U1434 ( .A(n1154), .B(n1155), .Z(n1151) );
  XNOR U1435 ( .A(n1148), .B(n1131), .Z(n1155) );
  IV U1436 ( .A(n1143), .Z(n1148) );
  XNOR U1437 ( .A(n1134), .B(n1147), .Z(n1154) );
  IV U1438 ( .A(n1139), .Z(n1147) );
  XOR U1439 ( .A(n1156), .B(n1157), .Z(n1139) );
  XNOR U1440 ( .A(n1158), .B(n1159), .Z(n1157) );
  XNOR U1441 ( .A(n1160), .B(n1161), .Z(n1156) );
  NOR U1442 ( .A(n1076), .B(n1120), .Z(n1160) );
  AND U1443 ( .A(n1131), .B(n1134), .Z(n1153) );
  XNOR U1444 ( .A(n1131), .B(n1134), .Z(n1146) );
  XNOR U1445 ( .A(n1162), .B(n1163), .Z(n1134) );
  XNOR U1446 ( .A(n1164), .B(n1159), .Z(n1163) );
  XOR U1447 ( .A(n1165), .B(n1166), .Z(n1162) );
  XNOR U1448 ( .A(n1167), .B(n1161), .Z(n1166) );
  OR U1449 ( .A(n1075), .B(n1119), .Z(n1161) );
  XOR U1450 ( .A(n1120), .B(n1110), .Z(n1119) );
  XNOR U1451 ( .A(n1076), .B(n1064), .Z(n1075) );
  ANDN U1452 ( .B(n1110), .A(n1064), .Z(n1167) );
  XNOR U1453 ( .A(n1168), .B(n1169), .Z(n1131) );
  XNOR U1454 ( .A(n1159), .B(n1170), .Z(n1169) );
  XOR U1455 ( .A(n1089), .B(n1165), .Z(n1170) );
  XNOR U1456 ( .A(n1120), .B(n1171), .Z(n1159) );
  XNOR U1457 ( .A(n1172), .B(n1173), .Z(n1168) );
  XNOR U1458 ( .A(n1174), .B(n1175), .Z(n1173) );
  ANDN U1459 ( .B(n1115), .A(n1097), .Z(n1174) );
  XNOR U1460 ( .A(n1176), .B(n1177), .Z(n1143) );
  XNOR U1461 ( .A(n1164), .B(n1178), .Z(n1177) );
  XNOR U1462 ( .A(n1097), .B(n1158), .Z(n1178) );
  XOR U1463 ( .A(n1165), .B(n1179), .Z(n1158) );
  XNOR U1464 ( .A(n1180), .B(n1181), .Z(n1179) );
  NAND U1465 ( .A(n1124), .B(n1094), .Z(n1181) );
  XNOR U1466 ( .A(n1182), .B(n1180), .Z(n1165) );
  NANDN U1467 ( .A(n1126), .B(n1103), .Z(n1180) );
  XOR U1468 ( .A(n1104), .B(n1094), .Z(n1103) );
  XNOR U1469 ( .A(n1183), .B(n1064), .Z(n1094) );
  XOR U1470 ( .A(n1135), .B(n1124), .Z(n1126) );
  XOR U1471 ( .A(n1115), .B(n1110), .Z(n1124) );
  ANDN U1472 ( .B(n1104), .A(n1135), .Z(n1182) );
  XOR U1473 ( .A(n1172), .B(n1120), .Z(n1135) );
  XOR U1474 ( .A(n1184), .B(n1185), .Z(n1120) );
  XOR U1475 ( .A(n1186), .B(n1187), .Z(n1185) );
  XOR U1476 ( .A(n1188), .B(n1171), .Z(n1104) );
  XNOR U1477 ( .A(n1189), .B(n1190), .Z(n1064) );
  XNOR U1478 ( .A(n1191), .B(n1187), .Z(n1190) );
  XNOR U1479 ( .A(n1187), .B(n1189), .Z(n1110) );
  XNOR U1480 ( .A(n1115), .B(n1192), .Z(n1176) );
  XNOR U1481 ( .A(n1193), .B(n1175), .Z(n1192) );
  OR U1482 ( .A(n1100), .B(n1114), .Z(n1175) );
  XNOR U1483 ( .A(n1172), .B(n1115), .Z(n1114) );
  XOR U1484 ( .A(n1089), .B(n1183), .Z(n1100) );
  IV U1485 ( .A(n1097), .Z(n1183) );
  XOR U1486 ( .A(n1171), .B(n1194), .Z(n1097) );
  XNOR U1487 ( .A(n1191), .B(n1184), .Z(n1194) );
  XOR U1488 ( .A(key[530]), .B(\w0[4][18] ), .Z(n1184) );
  XNOR U1489 ( .A(n625), .B(n1195), .Z(\w0[4][18] ) );
  XOR U1490 ( .A(n621), .B(n1196), .Z(n1195) );
  IV U1491 ( .A(n1076), .Z(n1171) );
  XNOR U1492 ( .A(n1189), .B(n1197), .Z(n1076) );
  XNOR U1493 ( .A(n1187), .B(n1198), .Z(n1197) );
  ANDN U1494 ( .B(n1188), .A(n1057), .Z(n1193) );
  IV U1495 ( .A(n1089), .Z(n1188) );
  XNOR U1496 ( .A(n1189), .B(n1199), .Z(n1089) );
  XNOR U1497 ( .A(n1187), .B(n1200), .Z(n1199) );
  XOR U1498 ( .A(n1057), .B(n1201), .Z(n1187) );
  XOR U1499 ( .A(key[534]), .B(\w0[4][22] ), .Z(n1201) );
  XNOR U1500 ( .A(n599), .B(n1202), .Z(\w0[4][22] ) );
  XNOR U1501 ( .A(n595), .B(n1203), .Z(n1202) );
  XNOR U1502 ( .A(n1204), .B(n1205), .Z(n599) );
  IV U1503 ( .A(n1172), .Z(n1057) );
  XOR U1504 ( .A(key[533]), .B(\w0[4][21] ), .Z(n1189) );
  XNOR U1505 ( .A(n594), .B(n1206), .Z(\w0[4][21] ) );
  XOR U1506 ( .A(n1207), .B(n1208), .Z(n1206) );
  XOR U1507 ( .A(n1209), .B(n1210), .Z(n594) );
  XOR U1508 ( .A(n1211), .B(n1212), .Z(n1115) );
  XNOR U1509 ( .A(n1200), .B(n1198), .Z(n1212) );
  XOR U1510 ( .A(key[535]), .B(\w0[4][23] ), .Z(n1198) );
  XNOR U1511 ( .A(n587), .B(n1213), .Z(\w0[4][23] ) );
  XOR U1512 ( .A(n1214), .B(n1205), .Z(n1213) );
  XOR U1513 ( .A(n1215), .B(n1216), .Z(n1205) );
  XNOR U1514 ( .A(n1217), .B(n1218), .Z(n587) );
  XOR U1515 ( .A(key[532]), .B(\w0[4][20] ), .Z(n1200) );
  XNOR U1516 ( .A(n578), .B(n1219), .Z(\w0[4][20] ) );
  XNOR U1517 ( .A(n1220), .B(n1221), .Z(n1219) );
  XOR U1518 ( .A(n1222), .B(n1223), .Z(n578) );
  XNOR U1519 ( .A(n1224), .B(n1216), .Z(n1223) );
  XNOR U1520 ( .A(n1225), .B(n1226), .Z(n1222) );
  XNOR U1521 ( .A(n1172), .B(n1186), .Z(n1211) );
  XOR U1522 ( .A(n1191), .B(n1227), .Z(n1186) );
  XOR U1523 ( .A(key[531]), .B(\w0[4][19] ), .Z(n1227) );
  XOR U1524 ( .A(n1228), .B(n1229), .Z(\w0[4][19] ) );
  XNOR U1525 ( .A(n1230), .B(n613), .Z(n1229) );
  XOR U1526 ( .A(n1220), .B(n1216), .Z(n613) );
  XOR U1527 ( .A(n627), .B(n1231), .Z(n1228) );
  XOR U1528 ( .A(key[529]), .B(\w0[4][17] ), .Z(n1191) );
  XOR U1529 ( .A(n1232), .B(n1233), .Z(\w0[4][17] ) );
  XOR U1530 ( .A(n620), .B(n606), .Z(n1233) );
  XOR U1531 ( .A(key[528]), .B(\w0[4][16] ), .Z(n1172) );
  XNOR U1532 ( .A(n590), .B(n1234), .Z(\w0[4][16] ) );
  XOR U1533 ( .A(n1235), .B(n1236), .Z(n1234) );
  XOR U1534 ( .A(n1237), .B(n1238), .Z(out[47]) );
  XOR U1535 ( .A(n1239), .B(n1240), .Z(n1237) );
  XNOR U1536 ( .A(key[559]), .B(n1241), .Z(n1240) );
  XNOR U1537 ( .A(n1242), .B(n1243), .Z(out[46]) );
  XNOR U1538 ( .A(key[558]), .B(n1244), .Z(n1243) );
  XOR U1539 ( .A(n1245), .B(n1246), .Z(out[45]) );
  XNOR U1540 ( .A(n1247), .B(n1248), .Z(n1246) );
  XOR U1541 ( .A(n1239), .B(n1249), .Z(n1248) );
  XNOR U1542 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1543 ( .A(n1253), .B(n1254), .Z(n1252) );
  XOR U1544 ( .A(n1256), .B(n1257), .Z(n1245) );
  XOR U1545 ( .A(key[557]), .B(n1258), .Z(n1257) );
  ANDN U1546 ( .B(n1259), .A(n1260), .Z(n1256) );
  XNOR U1547 ( .A(n1261), .B(n1262), .Z(out[44]) );
  XNOR U1548 ( .A(key[556]), .B(n1263), .Z(n1262) );
  XOR U1549 ( .A(n1264), .B(n1265), .Z(out[43]) );
  XNOR U1550 ( .A(n1266), .B(n1242), .Z(n1265) );
  XNOR U1551 ( .A(n1267), .B(n1268), .Z(n1242) );
  XNOR U1552 ( .A(n1269), .B(n1258), .Z(n1268) );
  ANDN U1553 ( .B(n1270), .A(n1271), .Z(n1258) );
  NOR U1554 ( .A(n1272), .B(n1273), .Z(n1269) );
  XNOR U1555 ( .A(n1274), .B(n1275), .Z(n1264) );
  XOR U1556 ( .A(key[555]), .B(n1276), .Z(n1275) );
  XOR U1557 ( .A(key[554]), .B(n1261), .Z(out[42]) );
  XNOR U1558 ( .A(n1241), .B(n1277), .Z(n1261) );
  IV U1559 ( .A(n1276), .Z(n1241) );
  XOR U1560 ( .A(n1278), .B(n1238), .Z(out[41]) );
  XNOR U1561 ( .A(n1267), .B(n1279), .Z(n1266) );
  XNOR U1562 ( .A(n1280), .B(n1281), .Z(n1279) );
  NANDN U1563 ( .A(n1282), .B(n1254), .Z(n1281) );
  XNOR U1564 ( .A(n1249), .B(n1283), .Z(n1267) );
  XNOR U1565 ( .A(n1284), .B(n1285), .Z(n1283) );
  NANDN U1566 ( .A(n1286), .B(n1287), .Z(n1285) );
  XOR U1567 ( .A(n1277), .B(n1274), .Z(n1244) );
  XNOR U1568 ( .A(n1249), .B(n1288), .Z(n1274) );
  XNOR U1569 ( .A(n1280), .B(n1289), .Z(n1288) );
  NANDN U1570 ( .A(n1290), .B(n1291), .Z(n1289) );
  OR U1571 ( .A(n1292), .B(n1293), .Z(n1280) );
  XOR U1572 ( .A(n1294), .B(n1284), .Z(n1249) );
  NANDN U1573 ( .A(n1295), .B(n1296), .Z(n1284) );
  ANDN U1574 ( .B(n1297), .A(n1298), .Z(n1294) );
  XOR U1575 ( .A(key[553]), .B(n1276), .Z(n1278) );
  XOR U1576 ( .A(n1299), .B(n1300), .Z(n1276) );
  XNOR U1577 ( .A(n1301), .B(n1302), .Z(n1300) );
  NAND U1578 ( .A(n1259), .B(n1303), .Z(n1302) );
  XNOR U1579 ( .A(n1247), .B(n1304), .Z(out[40]) );
  XOR U1580 ( .A(key[552]), .B(n1277), .Z(n1304) );
  XNOR U1581 ( .A(n1299), .B(n1305), .Z(n1277) );
  XOR U1582 ( .A(n1306), .B(n1251), .Z(n1305) );
  OR U1583 ( .A(n1307), .B(n1292), .Z(n1251) );
  XNOR U1584 ( .A(n1254), .B(n1291), .Z(n1292) );
  ANDN U1585 ( .B(n1308), .A(n1309), .Z(n1306) );
  IV U1586 ( .A(n1263), .Z(n1247) );
  XOR U1587 ( .A(n1255), .B(n1310), .Z(n1263) );
  XOR U1588 ( .A(n1311), .B(n1301), .Z(n1310) );
  XNOR U1589 ( .A(n1273), .B(n1259), .Z(n1270) );
  NOR U1590 ( .A(n1313), .B(n1273), .Z(n1311) );
  XNOR U1591 ( .A(n1299), .B(n1314), .Z(n1255) );
  XNOR U1592 ( .A(n1315), .B(n1316), .Z(n1314) );
  NANDN U1593 ( .A(n1286), .B(n1317), .Z(n1316) );
  XOR U1594 ( .A(n1318), .B(n1315), .Z(n1299) );
  OR U1595 ( .A(n1295), .B(n1319), .Z(n1315) );
  XOR U1596 ( .A(n1320), .B(n1286), .Z(n1295) );
  XNOR U1597 ( .A(n1291), .B(n1259), .Z(n1286) );
  XOR U1598 ( .A(n1321), .B(n1322), .Z(n1259) );
  NANDN U1599 ( .A(n1323), .B(n1324), .Z(n1322) );
  IV U1600 ( .A(n1309), .Z(n1291) );
  XNOR U1601 ( .A(n1325), .B(n1326), .Z(n1309) );
  NANDN U1602 ( .A(n1323), .B(n1327), .Z(n1326) );
  ANDN U1603 ( .B(n1320), .A(n1328), .Z(n1318) );
  IV U1604 ( .A(n1298), .Z(n1320) );
  XOR U1605 ( .A(n1273), .B(n1254), .Z(n1298) );
  XNOR U1606 ( .A(n1329), .B(n1325), .Z(n1254) );
  NANDN U1607 ( .A(n1330), .B(n1331), .Z(n1325) );
  XOR U1608 ( .A(n1327), .B(n1332), .Z(n1331) );
  ANDN U1609 ( .B(n1332), .A(n1333), .Z(n1329) );
  XOR U1610 ( .A(n1334), .B(n1321), .Z(n1273) );
  NANDN U1611 ( .A(n1330), .B(n1335), .Z(n1321) );
  XOR U1612 ( .A(n1336), .B(n1324), .Z(n1335) );
  XNOR U1613 ( .A(n1337), .B(n1338), .Z(n1323) );
  XOR U1614 ( .A(n1339), .B(n1340), .Z(n1338) );
  XNOR U1615 ( .A(n1341), .B(n1342), .Z(n1337) );
  XNOR U1616 ( .A(n1343), .B(n1344), .Z(n1342) );
  ANDN U1617 ( .B(n1336), .A(n1340), .Z(n1343) );
  ANDN U1618 ( .B(n1336), .A(n1333), .Z(n1334) );
  XNOR U1619 ( .A(n1339), .B(n1345), .Z(n1333) );
  XOR U1620 ( .A(n1346), .B(n1344), .Z(n1345) );
  NAND U1621 ( .A(n1347), .B(n1348), .Z(n1344) );
  XNOR U1622 ( .A(n1341), .B(n1324), .Z(n1348) );
  IV U1623 ( .A(n1336), .Z(n1341) );
  XNOR U1624 ( .A(n1327), .B(n1340), .Z(n1347) );
  IV U1625 ( .A(n1332), .Z(n1340) );
  XOR U1626 ( .A(n1349), .B(n1350), .Z(n1332) );
  XNOR U1627 ( .A(n1351), .B(n1352), .Z(n1350) );
  XNOR U1628 ( .A(n1353), .B(n1354), .Z(n1349) );
  NOR U1629 ( .A(n1272), .B(n1313), .Z(n1353) );
  AND U1630 ( .A(n1324), .B(n1327), .Z(n1346) );
  XNOR U1631 ( .A(n1324), .B(n1327), .Z(n1339) );
  XNOR U1632 ( .A(n1355), .B(n1356), .Z(n1327) );
  XNOR U1633 ( .A(n1357), .B(n1352), .Z(n1356) );
  XOR U1634 ( .A(n1358), .B(n1359), .Z(n1355) );
  XNOR U1635 ( .A(n1360), .B(n1354), .Z(n1359) );
  OR U1636 ( .A(n1271), .B(n1312), .Z(n1354) );
  XOR U1637 ( .A(n1313), .B(n1303), .Z(n1312) );
  XNOR U1638 ( .A(n1272), .B(n1260), .Z(n1271) );
  ANDN U1639 ( .B(n1303), .A(n1260), .Z(n1360) );
  XNOR U1640 ( .A(n1361), .B(n1362), .Z(n1324) );
  XNOR U1641 ( .A(n1352), .B(n1363), .Z(n1362) );
  XOR U1642 ( .A(n1282), .B(n1358), .Z(n1363) );
  XNOR U1643 ( .A(n1313), .B(n1364), .Z(n1352) );
  XNOR U1644 ( .A(n1365), .B(n1366), .Z(n1361) );
  XNOR U1645 ( .A(n1367), .B(n1368), .Z(n1366) );
  ANDN U1646 ( .B(n1308), .A(n1290), .Z(n1367) );
  XNOR U1647 ( .A(n1369), .B(n1370), .Z(n1336) );
  XNOR U1648 ( .A(n1357), .B(n1371), .Z(n1370) );
  XNOR U1649 ( .A(n1290), .B(n1351), .Z(n1371) );
  XOR U1650 ( .A(n1358), .B(n1372), .Z(n1351) );
  XNOR U1651 ( .A(n1373), .B(n1374), .Z(n1372) );
  NAND U1652 ( .A(n1317), .B(n1287), .Z(n1374) );
  XNOR U1653 ( .A(n1375), .B(n1373), .Z(n1358) );
  NANDN U1654 ( .A(n1319), .B(n1296), .Z(n1373) );
  XOR U1655 ( .A(n1297), .B(n1287), .Z(n1296) );
  XNOR U1656 ( .A(n1376), .B(n1260), .Z(n1287) );
  XOR U1657 ( .A(n1328), .B(n1317), .Z(n1319) );
  XOR U1658 ( .A(n1308), .B(n1303), .Z(n1317) );
  ANDN U1659 ( .B(n1297), .A(n1328), .Z(n1375) );
  XOR U1660 ( .A(n1365), .B(n1313), .Z(n1328) );
  XOR U1661 ( .A(n1377), .B(n1378), .Z(n1313) );
  XOR U1662 ( .A(n1379), .B(n1380), .Z(n1378) );
  XOR U1663 ( .A(n1381), .B(n1364), .Z(n1297) );
  XNOR U1664 ( .A(n1382), .B(n1383), .Z(n1260) );
  XNOR U1665 ( .A(n1384), .B(n1380), .Z(n1383) );
  XNOR U1666 ( .A(n1380), .B(n1382), .Z(n1303) );
  XNOR U1667 ( .A(n1308), .B(n1385), .Z(n1369) );
  XNOR U1668 ( .A(n1386), .B(n1368), .Z(n1385) );
  OR U1669 ( .A(n1293), .B(n1307), .Z(n1368) );
  XNOR U1670 ( .A(n1365), .B(n1308), .Z(n1307) );
  XOR U1671 ( .A(n1282), .B(n1376), .Z(n1293) );
  IV U1672 ( .A(n1290), .Z(n1376) );
  XOR U1673 ( .A(n1364), .B(n1387), .Z(n1290) );
  XNOR U1674 ( .A(n1384), .B(n1377), .Z(n1387) );
  XOR U1675 ( .A(key[618]), .B(\w0[4][106] ), .Z(n1377) );
  XOR U1676 ( .A(n1388), .B(n1389), .Z(\w0[4][106] ) );
  XNOR U1677 ( .A(n1390), .B(n811), .Z(n1389) );
  XNOR U1678 ( .A(n1391), .B(n1392), .Z(n1388) );
  IV U1679 ( .A(n1272), .Z(n1364) );
  XNOR U1680 ( .A(n1382), .B(n1393), .Z(n1272) );
  XOR U1681 ( .A(n1380), .B(n1394), .Z(n1393) );
  ANDN U1682 ( .B(n1381), .A(n1253), .Z(n1386) );
  IV U1683 ( .A(n1282), .Z(n1381) );
  XNOR U1684 ( .A(n1382), .B(n1395), .Z(n1282) );
  XNOR U1685 ( .A(n1380), .B(n1396), .Z(n1395) );
  XOR U1686 ( .A(n1253), .B(n1397), .Z(n1380) );
  XOR U1687 ( .A(key[622]), .B(\w0[4][110] ), .Z(n1397) );
  XNOR U1688 ( .A(n817), .B(n1398), .Z(\w0[4][110] ) );
  XNOR U1689 ( .A(n1399), .B(n1400), .Z(n1398) );
  XNOR U1690 ( .A(n1401), .B(n1402), .Z(n817) );
  IV U1691 ( .A(n1365), .Z(n1253) );
  XOR U1692 ( .A(key[621]), .B(\w0[4][109] ), .Z(n1382) );
  XOR U1693 ( .A(n1403), .B(n1404), .Z(\w0[4][109] ) );
  XOR U1694 ( .A(n1405), .B(n1406), .Z(n1404) );
  XNOR U1695 ( .A(n1407), .B(n1408), .Z(n1403) );
  XOR U1696 ( .A(n1409), .B(n1410), .Z(n1308) );
  XOR U1697 ( .A(n1396), .B(n1394), .Z(n1410) );
  XNOR U1698 ( .A(key[623]), .B(\w0[4][111] ), .Z(n1394) );
  XNOR U1699 ( .A(n1411), .B(n1412), .Z(\w0[4][111] ) );
  XOR U1700 ( .A(n1413), .B(n1414), .Z(n1412) );
  XOR U1701 ( .A(key[620]), .B(\w0[4][108] ), .Z(n1396) );
  XOR U1702 ( .A(n1415), .B(n1416), .Z(\w0[4][108] ) );
  XOR U1703 ( .A(n1417), .B(n784), .Z(n1416) );
  XOR U1704 ( .A(n794), .B(n1418), .Z(n784) );
  XOR U1705 ( .A(n1419), .B(n1420), .Z(n1415) );
  XNOR U1706 ( .A(n1365), .B(n1379), .Z(n1409) );
  XOR U1707 ( .A(n1384), .B(n1421), .Z(n1379) );
  XOR U1708 ( .A(key[619]), .B(\w0[4][107] ), .Z(n1421) );
  XOR U1709 ( .A(n1422), .B(n1423), .Z(\w0[4][107] ) );
  XOR U1710 ( .A(n812), .B(n1424), .Z(n1423) );
  XOR U1711 ( .A(n806), .B(n1425), .Z(n1422) );
  XOR U1712 ( .A(n1426), .B(n794), .Z(n806) );
  IV U1713 ( .A(n1401), .Z(n794) );
  XOR U1714 ( .A(key[617]), .B(\w0[4][105] ), .Z(n1384) );
  XOR U1715 ( .A(n1427), .B(n1428), .Z(\w0[4][105] ) );
  XOR U1716 ( .A(n1429), .B(n824), .Z(n1428) );
  XOR U1717 ( .A(n1430), .B(n1431), .Z(n1427) );
  XOR U1718 ( .A(key[616]), .B(\w0[4][104] ), .Z(n1365) );
  XOR U1719 ( .A(n1432), .B(n1433), .Z(\w0[4][104] ) );
  XOR U1720 ( .A(n1434), .B(n821), .Z(n1433) );
  XNOR U1721 ( .A(n1401), .B(n1435), .Z(n1432) );
  XOR U1722 ( .A(n1436), .B(n1437), .Z(out[3]) );
  XNOR U1723 ( .A(n1438), .B(n638), .Z(n1437) );
  XNOR U1724 ( .A(n1439), .B(n1440), .Z(n638) );
  XNOR U1725 ( .A(n1441), .B(n865), .Z(n1440) );
  ANDN U1726 ( .B(n1442), .A(n1443), .Z(n865) );
  NOR U1727 ( .A(n1444), .B(n1445), .Z(n1441) );
  XNOR U1728 ( .A(n1446), .B(n1447), .Z(n1436) );
  XOR U1729 ( .A(key[515]), .B(n425), .Z(n1447) );
  XOR U1730 ( .A(n1448), .B(n1449), .Z(out[39]) );
  XOR U1731 ( .A(n1450), .B(n1451), .Z(n1448) );
  XOR U1732 ( .A(key[551]), .B(n1452), .Z(n1451) );
  XNOR U1733 ( .A(n1453), .B(n1454), .Z(out[38]) );
  XNOR U1734 ( .A(key[550]), .B(n1455), .Z(n1454) );
  XOR U1735 ( .A(n1456), .B(n1457), .Z(out[37]) );
  XNOR U1736 ( .A(n1458), .B(n1459), .Z(n1457) );
  XOR U1737 ( .A(n1450), .B(n1460), .Z(n1459) );
  XNOR U1738 ( .A(n1462), .B(n1463), .Z(n1461) );
  NANDN U1739 ( .A(n1464), .B(n1465), .Z(n1463) );
  XOR U1740 ( .A(n1467), .B(n1468), .Z(n1456) );
  XOR U1741 ( .A(key[549]), .B(n1469), .Z(n1468) );
  ANDN U1742 ( .B(n1470), .A(n1471), .Z(n1467) );
  XNOR U1743 ( .A(n1472), .B(n1473), .Z(out[36]) );
  XNOR U1744 ( .A(key[548]), .B(n1474), .Z(n1473) );
  XOR U1745 ( .A(n1475), .B(n1476), .Z(out[35]) );
  XNOR U1746 ( .A(n1477), .B(n1453), .Z(n1476) );
  XNOR U1747 ( .A(n1478), .B(n1479), .Z(n1453) );
  XNOR U1748 ( .A(n1480), .B(n1469), .Z(n1479) );
  ANDN U1749 ( .B(n1481), .A(n1482), .Z(n1469) );
  NOR U1750 ( .A(n1483), .B(n1484), .Z(n1480) );
  XNOR U1751 ( .A(n1485), .B(n1486), .Z(n1475) );
  XOR U1752 ( .A(key[547]), .B(n1452), .Z(n1486) );
  XOR U1753 ( .A(key[546]), .B(n1472), .Z(out[34]) );
  XNOR U1754 ( .A(n1487), .B(n1488), .Z(n1472) );
  XOR U1755 ( .A(n1489), .B(n1449), .Z(out[33]) );
  XNOR U1756 ( .A(n1478), .B(n1490), .Z(n1477) );
  XNOR U1757 ( .A(n1491), .B(n1492), .Z(n1490) );
  NANDN U1758 ( .A(n1493), .B(n1465), .Z(n1492) );
  XNOR U1759 ( .A(n1460), .B(n1494), .Z(n1478) );
  XNOR U1760 ( .A(n1495), .B(n1496), .Z(n1494) );
  NANDN U1761 ( .A(n1497), .B(n1498), .Z(n1496) );
  XOR U1762 ( .A(n1488), .B(n1485), .Z(n1455) );
  XNOR U1763 ( .A(n1460), .B(n1499), .Z(n1485) );
  XNOR U1764 ( .A(n1491), .B(n1500), .Z(n1499) );
  NANDN U1765 ( .A(n1501), .B(n1502), .Z(n1500) );
  OR U1766 ( .A(n1503), .B(n1504), .Z(n1491) );
  XOR U1767 ( .A(n1505), .B(n1495), .Z(n1460) );
  NANDN U1768 ( .A(n1506), .B(n1507), .Z(n1495) );
  ANDN U1769 ( .B(n1508), .A(n1509), .Z(n1505) );
  XNOR U1770 ( .A(key[545]), .B(n1487), .Z(n1489) );
  IV U1771 ( .A(n1452), .Z(n1487) );
  XOR U1772 ( .A(n1510), .B(n1511), .Z(n1452) );
  XNOR U1773 ( .A(n1512), .B(n1513), .Z(n1511) );
  NANDN U1774 ( .A(n1514), .B(n1470), .Z(n1513) );
  XNOR U1775 ( .A(n1458), .B(n1515), .Z(out[32]) );
  XOR U1776 ( .A(key[544]), .B(n1488), .Z(n1515) );
  XNOR U1777 ( .A(n1510), .B(n1516), .Z(n1488) );
  XOR U1778 ( .A(n1517), .B(n1462), .Z(n1516) );
  OR U1779 ( .A(n1518), .B(n1503), .Z(n1462) );
  XNOR U1780 ( .A(n1465), .B(n1502), .Z(n1503) );
  ANDN U1781 ( .B(n1519), .A(n1520), .Z(n1517) );
  IV U1782 ( .A(n1474), .Z(n1458) );
  XOR U1783 ( .A(n1466), .B(n1521), .Z(n1474) );
  XOR U1784 ( .A(n1522), .B(n1512), .Z(n1521) );
  XNOR U1785 ( .A(n1484), .B(n1470), .Z(n1481) );
  NOR U1786 ( .A(n1524), .B(n1484), .Z(n1522) );
  XNOR U1787 ( .A(n1510), .B(n1525), .Z(n1466) );
  XNOR U1788 ( .A(n1526), .B(n1527), .Z(n1525) );
  NANDN U1789 ( .A(n1497), .B(n1528), .Z(n1527) );
  XOR U1790 ( .A(n1529), .B(n1526), .Z(n1510) );
  OR U1791 ( .A(n1506), .B(n1530), .Z(n1526) );
  XOR U1792 ( .A(n1531), .B(n1497), .Z(n1506) );
  XNOR U1793 ( .A(n1502), .B(n1470), .Z(n1497) );
  XOR U1794 ( .A(n1532), .B(n1533), .Z(n1470) );
  NANDN U1795 ( .A(n1534), .B(n1535), .Z(n1533) );
  IV U1796 ( .A(n1520), .Z(n1502) );
  XNOR U1797 ( .A(n1536), .B(n1537), .Z(n1520) );
  NANDN U1798 ( .A(n1534), .B(n1538), .Z(n1537) );
  ANDN U1799 ( .B(n1531), .A(n1539), .Z(n1529) );
  IV U1800 ( .A(n1509), .Z(n1531) );
  XOR U1801 ( .A(n1484), .B(n1465), .Z(n1509) );
  XNOR U1802 ( .A(n1540), .B(n1536), .Z(n1465) );
  NANDN U1803 ( .A(n1541), .B(n1542), .Z(n1536) );
  XOR U1804 ( .A(n1538), .B(n1543), .Z(n1542) );
  ANDN U1805 ( .B(n1543), .A(n1544), .Z(n1540) );
  XOR U1806 ( .A(n1545), .B(n1532), .Z(n1484) );
  NANDN U1807 ( .A(n1541), .B(n1546), .Z(n1532) );
  XOR U1808 ( .A(n1547), .B(n1535), .Z(n1546) );
  XNOR U1809 ( .A(n1548), .B(n1549), .Z(n1534) );
  XOR U1810 ( .A(n1550), .B(n1551), .Z(n1549) );
  XNOR U1811 ( .A(n1552), .B(n1553), .Z(n1548) );
  XNOR U1812 ( .A(n1554), .B(n1555), .Z(n1553) );
  ANDN U1813 ( .B(n1547), .A(n1551), .Z(n1554) );
  ANDN U1814 ( .B(n1547), .A(n1544), .Z(n1545) );
  XNOR U1815 ( .A(n1550), .B(n1556), .Z(n1544) );
  XOR U1816 ( .A(n1557), .B(n1555), .Z(n1556) );
  NAND U1817 ( .A(n1558), .B(n1559), .Z(n1555) );
  XNOR U1818 ( .A(n1552), .B(n1535), .Z(n1559) );
  IV U1819 ( .A(n1547), .Z(n1552) );
  XNOR U1820 ( .A(n1538), .B(n1551), .Z(n1558) );
  IV U1821 ( .A(n1543), .Z(n1551) );
  XOR U1822 ( .A(n1560), .B(n1561), .Z(n1543) );
  XNOR U1823 ( .A(n1562), .B(n1563), .Z(n1561) );
  XNOR U1824 ( .A(n1564), .B(n1565), .Z(n1560) );
  NOR U1825 ( .A(n1483), .B(n1524), .Z(n1564) );
  AND U1826 ( .A(n1535), .B(n1538), .Z(n1557) );
  XNOR U1827 ( .A(n1535), .B(n1538), .Z(n1550) );
  XNOR U1828 ( .A(n1566), .B(n1567), .Z(n1538) );
  XNOR U1829 ( .A(n1568), .B(n1563), .Z(n1567) );
  XOR U1830 ( .A(n1569), .B(n1570), .Z(n1566) );
  XNOR U1831 ( .A(n1571), .B(n1565), .Z(n1570) );
  OR U1832 ( .A(n1482), .B(n1523), .Z(n1565) );
  XNOR U1833 ( .A(n1524), .B(n1514), .Z(n1523) );
  XNOR U1834 ( .A(n1483), .B(n1471), .Z(n1482) );
  ANDN U1835 ( .B(n1572), .A(n1514), .Z(n1571) );
  XNOR U1836 ( .A(n1573), .B(n1574), .Z(n1535) );
  XNOR U1837 ( .A(n1563), .B(n1575), .Z(n1574) );
  XOR U1838 ( .A(n1493), .B(n1569), .Z(n1575) );
  XNOR U1839 ( .A(n1524), .B(n1576), .Z(n1563) );
  XNOR U1840 ( .A(n1577), .B(n1578), .Z(n1573) );
  XNOR U1841 ( .A(n1579), .B(n1580), .Z(n1578) );
  ANDN U1842 ( .B(n1519), .A(n1501), .Z(n1579) );
  XNOR U1843 ( .A(n1581), .B(n1582), .Z(n1547) );
  XNOR U1844 ( .A(n1568), .B(n1583), .Z(n1582) );
  XNOR U1845 ( .A(n1501), .B(n1562), .Z(n1583) );
  XOR U1846 ( .A(n1569), .B(n1584), .Z(n1562) );
  XNOR U1847 ( .A(n1585), .B(n1586), .Z(n1584) );
  NAND U1848 ( .A(n1528), .B(n1498), .Z(n1586) );
  XNOR U1849 ( .A(n1587), .B(n1585), .Z(n1569) );
  NANDN U1850 ( .A(n1530), .B(n1507), .Z(n1585) );
  XOR U1851 ( .A(n1508), .B(n1498), .Z(n1507) );
  XNOR U1852 ( .A(n1588), .B(n1471), .Z(n1498) );
  XOR U1853 ( .A(n1539), .B(n1528), .Z(n1530) );
  XOR U1854 ( .A(n1519), .B(n1589), .Z(n1528) );
  ANDN U1855 ( .B(n1508), .A(n1539), .Z(n1587) );
  XOR U1856 ( .A(n1577), .B(n1524), .Z(n1539) );
  XOR U1857 ( .A(n1590), .B(n1591), .Z(n1524) );
  XOR U1858 ( .A(n1592), .B(n1593), .Z(n1591) );
  XOR U1859 ( .A(n1594), .B(n1576), .Z(n1508) );
  XOR U1860 ( .A(n1589), .B(n1572), .Z(n1568) );
  IV U1861 ( .A(n1471), .Z(n1572) );
  XOR U1862 ( .A(n1595), .B(n1596), .Z(n1471) );
  XNOR U1863 ( .A(n1597), .B(n1593), .Z(n1596) );
  IV U1864 ( .A(n1514), .Z(n1589) );
  XOR U1865 ( .A(n1593), .B(n1598), .Z(n1514) );
  XNOR U1866 ( .A(n1519), .B(n1599), .Z(n1581) );
  XNOR U1867 ( .A(n1600), .B(n1580), .Z(n1599) );
  OR U1868 ( .A(n1504), .B(n1518), .Z(n1580) );
  XNOR U1869 ( .A(n1577), .B(n1519), .Z(n1518) );
  XOR U1870 ( .A(n1493), .B(n1588), .Z(n1504) );
  IV U1871 ( .A(n1501), .Z(n1588) );
  XOR U1872 ( .A(n1576), .B(n1601), .Z(n1501) );
  XNOR U1873 ( .A(n1597), .B(n1590), .Z(n1601) );
  XOR U1874 ( .A(key[578]), .B(\w0[4][66] ), .Z(n1590) );
  XOR U1875 ( .A(n1602), .B(n1603), .Z(\w0[4][66] ) );
  XNOR U1876 ( .A(n219), .B(n1604), .Z(n1603) );
  IV U1877 ( .A(n1483), .Z(n1576) );
  XOR U1878 ( .A(n1595), .B(n1605), .Z(n1483) );
  XOR U1879 ( .A(n1593), .B(n1606), .Z(n1605) );
  ANDN U1880 ( .B(n1594), .A(n1464), .Z(n1600) );
  IV U1881 ( .A(n1493), .Z(n1594) );
  XOR U1882 ( .A(n1595), .B(n1607), .Z(n1493) );
  XOR U1883 ( .A(n1593), .B(n1608), .Z(n1607) );
  XOR U1884 ( .A(n1464), .B(n1609), .Z(n1593) );
  XOR U1885 ( .A(key[582]), .B(\w0[4][70] ), .Z(n1609) );
  XNOR U1886 ( .A(n1610), .B(n1611), .Z(\w0[4][70] ) );
  XOR U1887 ( .A(n187), .B(n192), .Z(n1611) );
  XNOR U1888 ( .A(n1612), .B(n1613), .Z(n187) );
  IV U1889 ( .A(n1577), .Z(n1464) );
  IV U1890 ( .A(n1598), .Z(n1595) );
  XOR U1891 ( .A(key[581]), .B(\w0[4][69] ), .Z(n1598) );
  XOR U1892 ( .A(n1614), .B(n1615), .Z(\w0[4][69] ) );
  XOR U1893 ( .A(n191), .B(n1616), .Z(n1615) );
  XNOR U1894 ( .A(n1617), .B(n1618), .Z(n191) );
  XOR U1895 ( .A(n1619), .B(n1620), .Z(n1519) );
  XNOR U1896 ( .A(n1608), .B(n1606), .Z(n1620) );
  XNOR U1897 ( .A(key[583]), .B(\w0[4][71] ), .Z(n1606) );
  XOR U1898 ( .A(n1621), .B(n1622), .Z(\w0[4][71] ) );
  XOR U1899 ( .A(n200), .B(n1613), .Z(n1622) );
  XNOR U1900 ( .A(n1623), .B(n1624), .Z(n1613) );
  XOR U1901 ( .A(n1625), .B(n1626), .Z(n200) );
  XNOR U1902 ( .A(key[580]), .B(\w0[4][68] ), .Z(n1608) );
  XOR U1903 ( .A(n1627), .B(n1628), .Z(\w0[4][68] ) );
  XNOR U1904 ( .A(n1629), .B(n1630), .Z(n1628) );
  XNOR U1905 ( .A(n205), .B(n204), .Z(n1627) );
  XNOR U1906 ( .A(n1631), .B(n1632), .Z(n204) );
  XOR U1907 ( .A(n1633), .B(n1616), .Z(n205) );
  XNOR U1908 ( .A(n1577), .B(n1592), .Z(n1619) );
  XOR U1909 ( .A(n1597), .B(n1634), .Z(n1592) );
  XOR U1910 ( .A(key[579]), .B(\w0[4][67] ), .Z(n1634) );
  XOR U1911 ( .A(n1635), .B(n1636), .Z(\w0[4][67] ) );
  XNOR U1912 ( .A(n177), .B(n1637), .Z(n1636) );
  XNOR U1913 ( .A(n212), .B(n211), .Z(n1635) );
  XOR U1914 ( .A(n1633), .B(n1629), .Z(n212) );
  XOR U1915 ( .A(key[577]), .B(\w0[4][65] ), .Z(n1597) );
  XNOR U1916 ( .A(n1638), .B(n1639), .Z(\w0[4][65] ) );
  XOR U1917 ( .A(n217), .B(n223), .Z(n1639) );
  XOR U1918 ( .A(key[576]), .B(\w0[4][64] ), .Z(n1577) );
  XNOR U1919 ( .A(n1640), .B(n1641), .Z(\w0[4][64] ) );
  XNOR U1920 ( .A(n197), .B(n1642), .Z(n1641) );
  XOR U1921 ( .A(n1643), .B(n1644), .Z(out[31]) );
  XOR U1922 ( .A(n1645), .B(n1646), .Z(n1643) );
  XOR U1923 ( .A(key[543]), .B(n1647), .Z(n1646) );
  XNOR U1924 ( .A(n1648), .B(n1649), .Z(out[30]) );
  XNOR U1925 ( .A(key[542]), .B(n1650), .Z(n1649) );
  XOR U1926 ( .A(key[514]), .B(n1082), .Z(out[2]) );
  XOR U1927 ( .A(n1652), .B(n1653), .Z(out[29]) );
  XNOR U1928 ( .A(n1654), .B(n1655), .Z(n1653) );
  XOR U1929 ( .A(n1645), .B(n1656), .Z(n1655) );
  XNOR U1930 ( .A(n1658), .B(n1659), .Z(n1657) );
  NANDN U1931 ( .A(n1660), .B(n1661), .Z(n1659) );
  XOR U1932 ( .A(n1663), .B(n1664), .Z(n1652) );
  XOR U1933 ( .A(key[541]), .B(n1665), .Z(n1664) );
  ANDN U1934 ( .B(n1666), .A(n1667), .Z(n1663) );
  XNOR U1935 ( .A(n1668), .B(n1669), .Z(out[28]) );
  XNOR U1936 ( .A(key[540]), .B(n1670), .Z(n1669) );
  XOR U1937 ( .A(n1671), .B(n1672), .Z(out[27]) );
  XNOR U1938 ( .A(n1673), .B(n1648), .Z(n1672) );
  XNOR U1939 ( .A(n1674), .B(n1675), .Z(n1648) );
  XNOR U1940 ( .A(n1676), .B(n1665), .Z(n1675) );
  ANDN U1941 ( .B(n1677), .A(n1678), .Z(n1665) );
  NOR U1942 ( .A(n1679), .B(n1680), .Z(n1676) );
  XNOR U1943 ( .A(n1681), .B(n1682), .Z(n1671) );
  XOR U1944 ( .A(key[539]), .B(n1647), .Z(n1682) );
  XOR U1945 ( .A(key[538]), .B(n1668), .Z(out[26]) );
  XNOR U1946 ( .A(n1683), .B(n1684), .Z(n1668) );
  XOR U1947 ( .A(n1685), .B(n1644), .Z(out[25]) );
  XNOR U1948 ( .A(n1674), .B(n1686), .Z(n1673) );
  XNOR U1949 ( .A(n1687), .B(n1688), .Z(n1686) );
  NANDN U1950 ( .A(n1689), .B(n1661), .Z(n1688) );
  XNOR U1951 ( .A(n1656), .B(n1690), .Z(n1674) );
  XNOR U1952 ( .A(n1691), .B(n1692), .Z(n1690) );
  NANDN U1953 ( .A(n1693), .B(n1694), .Z(n1692) );
  XOR U1954 ( .A(n1684), .B(n1681), .Z(n1650) );
  XNOR U1955 ( .A(n1656), .B(n1695), .Z(n1681) );
  XNOR U1956 ( .A(n1687), .B(n1696), .Z(n1695) );
  NANDN U1957 ( .A(n1697), .B(n1698), .Z(n1696) );
  OR U1958 ( .A(n1699), .B(n1700), .Z(n1687) );
  XOR U1959 ( .A(n1701), .B(n1691), .Z(n1656) );
  NANDN U1960 ( .A(n1702), .B(n1703), .Z(n1691) );
  ANDN U1961 ( .B(n1704), .A(n1705), .Z(n1701) );
  XNOR U1962 ( .A(key[537]), .B(n1683), .Z(n1685) );
  IV U1963 ( .A(n1647), .Z(n1683) );
  XOR U1964 ( .A(n1706), .B(n1707), .Z(n1647) );
  XNOR U1965 ( .A(n1708), .B(n1709), .Z(n1707) );
  NAND U1966 ( .A(n1666), .B(n1710), .Z(n1709) );
  XNOR U1967 ( .A(n1654), .B(n1711), .Z(out[24]) );
  XOR U1968 ( .A(key[536]), .B(n1684), .Z(n1711) );
  XNOR U1969 ( .A(n1706), .B(n1712), .Z(n1684) );
  XOR U1970 ( .A(n1713), .B(n1658), .Z(n1712) );
  OR U1971 ( .A(n1714), .B(n1699), .Z(n1658) );
  XNOR U1972 ( .A(n1661), .B(n1698), .Z(n1699) );
  ANDN U1973 ( .B(n1715), .A(n1716), .Z(n1713) );
  IV U1974 ( .A(n1670), .Z(n1654) );
  XOR U1975 ( .A(n1662), .B(n1717), .Z(n1670) );
  XOR U1976 ( .A(n1718), .B(n1708), .Z(n1717) );
  XNOR U1977 ( .A(n1680), .B(n1666), .Z(n1677) );
  NOR U1978 ( .A(n1720), .B(n1680), .Z(n1718) );
  XNOR U1979 ( .A(n1706), .B(n1721), .Z(n1662) );
  XNOR U1980 ( .A(n1722), .B(n1723), .Z(n1721) );
  NANDN U1981 ( .A(n1693), .B(n1724), .Z(n1723) );
  XOR U1982 ( .A(n1725), .B(n1722), .Z(n1706) );
  OR U1983 ( .A(n1702), .B(n1726), .Z(n1722) );
  XOR U1984 ( .A(n1727), .B(n1693), .Z(n1702) );
  XNOR U1985 ( .A(n1698), .B(n1666), .Z(n1693) );
  XOR U1986 ( .A(n1728), .B(n1729), .Z(n1666) );
  NANDN U1987 ( .A(n1730), .B(n1731), .Z(n1729) );
  IV U1988 ( .A(n1716), .Z(n1698) );
  XNOR U1989 ( .A(n1732), .B(n1733), .Z(n1716) );
  NANDN U1990 ( .A(n1730), .B(n1734), .Z(n1733) );
  ANDN U1991 ( .B(n1727), .A(n1735), .Z(n1725) );
  IV U1992 ( .A(n1705), .Z(n1727) );
  XOR U1993 ( .A(n1680), .B(n1661), .Z(n1705) );
  XNOR U1994 ( .A(n1736), .B(n1732), .Z(n1661) );
  NANDN U1995 ( .A(n1737), .B(n1738), .Z(n1732) );
  XOR U1996 ( .A(n1734), .B(n1739), .Z(n1738) );
  ANDN U1997 ( .B(n1739), .A(n1740), .Z(n1736) );
  XOR U1998 ( .A(n1741), .B(n1728), .Z(n1680) );
  NANDN U1999 ( .A(n1737), .B(n1742), .Z(n1728) );
  XOR U2000 ( .A(n1743), .B(n1731), .Z(n1742) );
  XNOR U2001 ( .A(n1744), .B(n1745), .Z(n1730) );
  XOR U2002 ( .A(n1746), .B(n1747), .Z(n1745) );
  XNOR U2003 ( .A(n1748), .B(n1749), .Z(n1744) );
  XNOR U2004 ( .A(n1750), .B(n1751), .Z(n1749) );
  ANDN U2005 ( .B(n1743), .A(n1747), .Z(n1750) );
  ANDN U2006 ( .B(n1743), .A(n1740), .Z(n1741) );
  XNOR U2007 ( .A(n1746), .B(n1752), .Z(n1740) );
  XOR U2008 ( .A(n1753), .B(n1751), .Z(n1752) );
  NAND U2009 ( .A(n1754), .B(n1755), .Z(n1751) );
  XNOR U2010 ( .A(n1748), .B(n1731), .Z(n1755) );
  IV U2011 ( .A(n1743), .Z(n1748) );
  XNOR U2012 ( .A(n1734), .B(n1747), .Z(n1754) );
  IV U2013 ( .A(n1739), .Z(n1747) );
  XOR U2014 ( .A(n1756), .B(n1757), .Z(n1739) );
  XNOR U2015 ( .A(n1758), .B(n1759), .Z(n1757) );
  XNOR U2016 ( .A(n1760), .B(n1761), .Z(n1756) );
  NOR U2017 ( .A(n1679), .B(n1720), .Z(n1760) );
  AND U2018 ( .A(n1731), .B(n1734), .Z(n1753) );
  XNOR U2019 ( .A(n1731), .B(n1734), .Z(n1746) );
  XNOR U2020 ( .A(n1762), .B(n1763), .Z(n1734) );
  XNOR U2021 ( .A(n1764), .B(n1759), .Z(n1763) );
  XOR U2022 ( .A(n1765), .B(n1766), .Z(n1762) );
  XNOR U2023 ( .A(n1767), .B(n1761), .Z(n1766) );
  OR U2024 ( .A(n1678), .B(n1719), .Z(n1761) );
  XOR U2025 ( .A(n1720), .B(n1710), .Z(n1719) );
  XNOR U2026 ( .A(n1679), .B(n1667), .Z(n1678) );
  ANDN U2027 ( .B(n1710), .A(n1667), .Z(n1767) );
  XNOR U2028 ( .A(n1768), .B(n1769), .Z(n1731) );
  XNOR U2029 ( .A(n1759), .B(n1770), .Z(n1769) );
  XOR U2030 ( .A(n1689), .B(n1765), .Z(n1770) );
  XNOR U2031 ( .A(n1720), .B(n1771), .Z(n1759) );
  XNOR U2032 ( .A(n1772), .B(n1773), .Z(n1768) );
  XNOR U2033 ( .A(n1774), .B(n1775), .Z(n1773) );
  ANDN U2034 ( .B(n1715), .A(n1697), .Z(n1774) );
  XNOR U2035 ( .A(n1776), .B(n1777), .Z(n1743) );
  XNOR U2036 ( .A(n1764), .B(n1778), .Z(n1777) );
  XNOR U2037 ( .A(n1697), .B(n1758), .Z(n1778) );
  XOR U2038 ( .A(n1765), .B(n1779), .Z(n1758) );
  XNOR U2039 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U2040 ( .A(n1724), .B(n1694), .Z(n1781) );
  XNOR U2041 ( .A(n1782), .B(n1780), .Z(n1765) );
  NANDN U2042 ( .A(n1726), .B(n1703), .Z(n1780) );
  XOR U2043 ( .A(n1704), .B(n1694), .Z(n1703) );
  XNOR U2044 ( .A(n1783), .B(n1667), .Z(n1694) );
  XOR U2045 ( .A(n1735), .B(n1724), .Z(n1726) );
  XOR U2046 ( .A(n1715), .B(n1710), .Z(n1724) );
  ANDN U2047 ( .B(n1704), .A(n1735), .Z(n1782) );
  XOR U2048 ( .A(n1772), .B(n1720), .Z(n1735) );
  XOR U2049 ( .A(n1784), .B(n1785), .Z(n1720) );
  XOR U2050 ( .A(n1786), .B(n1787), .Z(n1785) );
  XOR U2051 ( .A(n1788), .B(n1771), .Z(n1704) );
  XNOR U2052 ( .A(n1789), .B(n1790), .Z(n1667) );
  XNOR U2053 ( .A(n1791), .B(n1787), .Z(n1790) );
  XNOR U2054 ( .A(n1787), .B(n1789), .Z(n1710) );
  XNOR U2055 ( .A(n1715), .B(n1792), .Z(n1776) );
  XNOR U2056 ( .A(n1793), .B(n1775), .Z(n1792) );
  OR U2057 ( .A(n1700), .B(n1714), .Z(n1775) );
  XNOR U2058 ( .A(n1772), .B(n1715), .Z(n1714) );
  XOR U2059 ( .A(n1689), .B(n1783), .Z(n1700) );
  IV U2060 ( .A(n1697), .Z(n1783) );
  XOR U2061 ( .A(n1771), .B(n1794), .Z(n1697) );
  XNOR U2062 ( .A(n1791), .B(n1784), .Z(n1794) );
  XOR U2063 ( .A(key[538]), .B(\w0[4][26] ), .Z(n1784) );
  XOR U2064 ( .A(n1795), .B(n1796), .Z(\w0[4][26] ) );
  XOR U2065 ( .A(n615), .B(n1232), .Z(n1796) );
  XNOR U2066 ( .A(n619), .B(n1797), .Z(n1795) );
  IV U2067 ( .A(n1679), .Z(n1771) );
  XNOR U2068 ( .A(n1789), .B(n1798), .Z(n1679) );
  XNOR U2069 ( .A(n1787), .B(n1799), .Z(n1798) );
  ANDN U2070 ( .B(n1788), .A(n1660), .Z(n1793) );
  IV U2071 ( .A(n1689), .Z(n1788) );
  XNOR U2072 ( .A(n1789), .B(n1800), .Z(n1689) );
  XNOR U2073 ( .A(n1787), .B(n1801), .Z(n1800) );
  XOR U2074 ( .A(n1660), .B(n1802), .Z(n1787) );
  XOR U2075 ( .A(key[542]), .B(\w0[4][30] ), .Z(n1802) );
  XNOR U2076 ( .A(n1203), .B(n1803), .Z(\w0[4][30] ) );
  XNOR U2077 ( .A(n1804), .B(n596), .Z(n1803) );
  XOR U2078 ( .A(n1805), .B(n589), .Z(n1203) );
  IV U2079 ( .A(n1772), .Z(n1660) );
  XOR U2080 ( .A(key[541]), .B(\w0[4][29] ), .Z(n1789) );
  XOR U2081 ( .A(n1806), .B(n1807), .Z(\w0[4][29] ) );
  XOR U2082 ( .A(n1808), .B(n1210), .Z(n1807) );
  XOR U2083 ( .A(n602), .B(n1809), .Z(n1806) );
  XOR U2084 ( .A(n1810), .B(n1811), .Z(n1715) );
  XNOR U2085 ( .A(n1801), .B(n1799), .Z(n1811) );
  XOR U2086 ( .A(key[543]), .B(\w0[4][31] ), .Z(n1799) );
  XNOR U2087 ( .A(n1218), .B(n1812), .Z(\w0[4][31] ) );
  XOR U2088 ( .A(n608), .B(n1813), .Z(n1812) );
  XOR U2089 ( .A(key[540]), .B(\w0[4][28] ), .Z(n1801) );
  XOR U2090 ( .A(n1814), .B(n1815), .Z(\w0[4][28] ) );
  XNOR U2091 ( .A(n1805), .B(n593), .Z(n1221) );
  XNOR U2092 ( .A(n1816), .B(n1817), .Z(n1814) );
  XNOR U2093 ( .A(n1772), .B(n1786), .Z(n1810) );
  XOR U2094 ( .A(n1791), .B(n1818), .Z(n1786) );
  XOR U2095 ( .A(key[539]), .B(\w0[4][27] ), .Z(n1818) );
  XOR U2096 ( .A(n1819), .B(n1820), .Z(\w0[4][27] ) );
  XOR U2097 ( .A(n624), .B(n1230), .Z(n1820) );
  XOR U2098 ( .A(n1214), .B(n581), .Z(n1230) );
  XOR U2099 ( .A(n1821), .B(n1196), .Z(n1819) );
  XOR U2100 ( .A(key[537]), .B(\w0[4][25] ), .Z(n1791) );
  XOR U2101 ( .A(n1822), .B(n1823), .Z(\w0[4][25] ) );
  XOR U2102 ( .A(n626), .B(n1236), .Z(n1823) );
  XOR U2103 ( .A(n607), .B(n1824), .Z(n1822) );
  XOR U2104 ( .A(key[536]), .B(\w0[4][24] ), .Z(n1772) );
  XOR U2105 ( .A(n1825), .B(n1826), .Z(\w0[4][24] ) );
  XNOR U2106 ( .A(n1805), .B(n590), .Z(n1826) );
  XNOR U2107 ( .A(n605), .B(n1216), .Z(n590) );
  XOR U2108 ( .A(n1827), .B(n618), .Z(n1825) );
  XOR U2109 ( .A(n1828), .B(n1829), .Z(out[23]) );
  XOR U2110 ( .A(n1830), .B(n1831), .Z(n1828) );
  XOR U2111 ( .A(key[535]), .B(n1832), .Z(n1831) );
  XNOR U2112 ( .A(n1833), .B(n1834), .Z(out[22]) );
  XNOR U2113 ( .A(key[534]), .B(n1835), .Z(n1834) );
  XOR U2114 ( .A(n1836), .B(n1837), .Z(out[21]) );
  XNOR U2115 ( .A(n1838), .B(n1839), .Z(n1837) );
  XOR U2116 ( .A(n1830), .B(n1840), .Z(n1839) );
  XNOR U2117 ( .A(n1842), .B(n1843), .Z(n1841) );
  NANDN U2118 ( .A(n1844), .B(n1845), .Z(n1843) );
  XOR U2119 ( .A(n1847), .B(n1848), .Z(n1836) );
  XOR U2120 ( .A(key[533]), .B(n1849), .Z(n1848) );
  ANDN U2121 ( .B(n1850), .A(n1851), .Z(n1847) );
  XNOR U2122 ( .A(n1852), .B(n1853), .Z(out[20]) );
  XNOR U2123 ( .A(key[532]), .B(n1854), .Z(n1853) );
  XOR U2124 ( .A(n1855), .B(n422), .Z(out[1]) );
  XNOR U2125 ( .A(n1439), .B(n1856), .Z(n1438) );
  XNOR U2126 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U2127 ( .A(n1859), .B(n861), .Z(n1858) );
  XNOR U2128 ( .A(n856), .B(n1860), .Z(n1439) );
  XNOR U2129 ( .A(n1861), .B(n1862), .Z(n1860) );
  NANDN U2130 ( .A(n1863), .B(n1864), .Z(n1862) );
  XOR U2131 ( .A(n1651), .B(n1446), .Z(n640) );
  XNOR U2132 ( .A(n856), .B(n1865), .Z(n1446) );
  XNOR U2133 ( .A(n1857), .B(n1866), .Z(n1865) );
  NANDN U2134 ( .A(n1867), .B(n1868), .Z(n1866) );
  OR U2135 ( .A(n1869), .B(n1870), .Z(n1857) );
  XOR U2136 ( .A(n1871), .B(n1861), .Z(n856) );
  NANDN U2137 ( .A(n1872), .B(n1873), .Z(n1861) );
  ANDN U2138 ( .B(n1874), .A(n1875), .Z(n1871) );
  XOR U2139 ( .A(key[513]), .B(n425), .Z(n1855) );
  XOR U2140 ( .A(n1876), .B(n1877), .Z(n425) );
  XNOR U2141 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U2142 ( .A(n866), .B(n1880), .Z(n1879) );
  XOR U2143 ( .A(n1881), .B(n1882), .Z(out[19]) );
  XNOR U2144 ( .A(n1883), .B(n1833), .Z(n1882) );
  XNOR U2145 ( .A(n1884), .B(n1885), .Z(n1833) );
  XNOR U2146 ( .A(n1886), .B(n1849), .Z(n1885) );
  ANDN U2147 ( .B(n1887), .A(n1888), .Z(n1849) );
  NOR U2148 ( .A(n1889), .B(n1890), .Z(n1886) );
  XNOR U2149 ( .A(n1891), .B(n1892), .Z(n1881) );
  XOR U2150 ( .A(key[531]), .B(n1832), .Z(n1892) );
  XOR U2151 ( .A(key[530]), .B(n1852), .Z(out[18]) );
  XNOR U2152 ( .A(n1893), .B(n1894), .Z(n1852) );
  XOR U2153 ( .A(n1895), .B(n1829), .Z(out[17]) );
  XNOR U2154 ( .A(n1884), .B(n1896), .Z(n1883) );
  XNOR U2155 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U2156 ( .A(n1899), .B(n1845), .Z(n1898) );
  XNOR U2157 ( .A(n1840), .B(n1900), .Z(n1884) );
  XNOR U2158 ( .A(n1901), .B(n1902), .Z(n1900) );
  NANDN U2159 ( .A(n1903), .B(n1904), .Z(n1902) );
  XOR U2160 ( .A(n1894), .B(n1891), .Z(n1835) );
  XNOR U2161 ( .A(n1840), .B(n1905), .Z(n1891) );
  XNOR U2162 ( .A(n1897), .B(n1906), .Z(n1905) );
  NANDN U2163 ( .A(n1907), .B(n1908), .Z(n1906) );
  OR U2164 ( .A(n1909), .B(n1910), .Z(n1897) );
  XOR U2165 ( .A(n1911), .B(n1901), .Z(n1840) );
  NANDN U2166 ( .A(n1912), .B(n1913), .Z(n1901) );
  ANDN U2167 ( .B(n1914), .A(n1915), .Z(n1911) );
  XNOR U2168 ( .A(key[529]), .B(n1893), .Z(n1895) );
  IV U2169 ( .A(n1832), .Z(n1893) );
  XOR U2170 ( .A(n1916), .B(n1917), .Z(n1832) );
  XNOR U2171 ( .A(n1918), .B(n1919), .Z(n1917) );
  NAND U2172 ( .A(n1850), .B(n1920), .Z(n1919) );
  XNOR U2173 ( .A(n1838), .B(n1921), .Z(out[16]) );
  XOR U2174 ( .A(key[528]), .B(n1894), .Z(n1921) );
  XNOR U2175 ( .A(n1916), .B(n1922), .Z(n1894) );
  XOR U2176 ( .A(n1923), .B(n1842), .Z(n1922) );
  OR U2177 ( .A(n1924), .B(n1909), .Z(n1842) );
  XNOR U2178 ( .A(n1845), .B(n1908), .Z(n1909) );
  ANDN U2179 ( .B(n1925), .A(n1926), .Z(n1923) );
  IV U2180 ( .A(n1854), .Z(n1838) );
  XOR U2181 ( .A(n1846), .B(n1927), .Z(n1854) );
  XOR U2182 ( .A(n1928), .B(n1918), .Z(n1927) );
  XNOR U2183 ( .A(n1890), .B(n1850), .Z(n1887) );
  NOR U2184 ( .A(n1930), .B(n1890), .Z(n1928) );
  XNOR U2185 ( .A(n1916), .B(n1931), .Z(n1846) );
  XNOR U2186 ( .A(n1932), .B(n1933), .Z(n1931) );
  NANDN U2187 ( .A(n1903), .B(n1934), .Z(n1933) );
  XOR U2188 ( .A(n1935), .B(n1932), .Z(n1916) );
  OR U2189 ( .A(n1912), .B(n1936), .Z(n1932) );
  XOR U2190 ( .A(n1937), .B(n1903), .Z(n1912) );
  XNOR U2191 ( .A(n1908), .B(n1850), .Z(n1903) );
  XOR U2192 ( .A(n1938), .B(n1939), .Z(n1850) );
  NANDN U2193 ( .A(n1940), .B(n1941), .Z(n1939) );
  IV U2194 ( .A(n1926), .Z(n1908) );
  XNOR U2195 ( .A(n1942), .B(n1943), .Z(n1926) );
  NANDN U2196 ( .A(n1940), .B(n1944), .Z(n1943) );
  ANDN U2197 ( .B(n1937), .A(n1945), .Z(n1935) );
  IV U2198 ( .A(n1915), .Z(n1937) );
  XOR U2199 ( .A(n1890), .B(n1845), .Z(n1915) );
  XNOR U2200 ( .A(n1946), .B(n1942), .Z(n1845) );
  NANDN U2201 ( .A(n1947), .B(n1948), .Z(n1942) );
  XOR U2202 ( .A(n1944), .B(n1949), .Z(n1948) );
  ANDN U2203 ( .B(n1949), .A(n1950), .Z(n1946) );
  XOR U2204 ( .A(n1951), .B(n1938), .Z(n1890) );
  NANDN U2205 ( .A(n1947), .B(n1952), .Z(n1938) );
  XOR U2206 ( .A(n1953), .B(n1941), .Z(n1952) );
  XNOR U2207 ( .A(n1954), .B(n1955), .Z(n1940) );
  XOR U2208 ( .A(n1956), .B(n1957), .Z(n1955) );
  XNOR U2209 ( .A(n1958), .B(n1959), .Z(n1954) );
  XNOR U2210 ( .A(n1960), .B(n1961), .Z(n1959) );
  ANDN U2211 ( .B(n1953), .A(n1957), .Z(n1960) );
  ANDN U2212 ( .B(n1953), .A(n1950), .Z(n1951) );
  XNOR U2213 ( .A(n1956), .B(n1962), .Z(n1950) );
  XOR U2214 ( .A(n1963), .B(n1961), .Z(n1962) );
  NAND U2215 ( .A(n1964), .B(n1965), .Z(n1961) );
  XNOR U2216 ( .A(n1958), .B(n1941), .Z(n1965) );
  IV U2217 ( .A(n1953), .Z(n1958) );
  XNOR U2218 ( .A(n1944), .B(n1957), .Z(n1964) );
  IV U2219 ( .A(n1949), .Z(n1957) );
  XOR U2220 ( .A(n1966), .B(n1967), .Z(n1949) );
  XNOR U2221 ( .A(n1968), .B(n1969), .Z(n1967) );
  XNOR U2222 ( .A(n1970), .B(n1971), .Z(n1966) );
  NOR U2223 ( .A(n1889), .B(n1930), .Z(n1970) );
  AND U2224 ( .A(n1941), .B(n1944), .Z(n1963) );
  XNOR U2225 ( .A(n1941), .B(n1944), .Z(n1956) );
  XNOR U2226 ( .A(n1972), .B(n1973), .Z(n1944) );
  XNOR U2227 ( .A(n1974), .B(n1969), .Z(n1973) );
  XOR U2228 ( .A(n1975), .B(n1976), .Z(n1972) );
  XNOR U2229 ( .A(n1977), .B(n1971), .Z(n1976) );
  OR U2230 ( .A(n1888), .B(n1929), .Z(n1971) );
  XOR U2231 ( .A(n1930), .B(n1920), .Z(n1929) );
  XNOR U2232 ( .A(n1889), .B(n1851), .Z(n1888) );
  ANDN U2233 ( .B(n1920), .A(n1851), .Z(n1977) );
  XNOR U2234 ( .A(n1978), .B(n1979), .Z(n1941) );
  XNOR U2235 ( .A(n1969), .B(n1980), .Z(n1979) );
  XOR U2236 ( .A(n1899), .B(n1975), .Z(n1980) );
  XNOR U2237 ( .A(n1930), .B(n1981), .Z(n1969) );
  XNOR U2238 ( .A(n1982), .B(n1983), .Z(n1978) );
  XNOR U2239 ( .A(n1984), .B(n1985), .Z(n1983) );
  ANDN U2240 ( .B(n1925), .A(n1907), .Z(n1984) );
  XNOR U2241 ( .A(n1986), .B(n1987), .Z(n1953) );
  XNOR U2242 ( .A(n1974), .B(n1988), .Z(n1987) );
  XNOR U2243 ( .A(n1907), .B(n1968), .Z(n1988) );
  XOR U2244 ( .A(n1975), .B(n1989), .Z(n1968) );
  XNOR U2245 ( .A(n1990), .B(n1991), .Z(n1989) );
  NAND U2246 ( .A(n1934), .B(n1904), .Z(n1991) );
  XNOR U2247 ( .A(n1992), .B(n1990), .Z(n1975) );
  NANDN U2248 ( .A(n1936), .B(n1913), .Z(n1990) );
  XOR U2249 ( .A(n1914), .B(n1904), .Z(n1913) );
  XNOR U2250 ( .A(n1993), .B(n1851), .Z(n1904) );
  XOR U2251 ( .A(n1945), .B(n1934), .Z(n1936) );
  XOR U2252 ( .A(n1925), .B(n1920), .Z(n1934) );
  ANDN U2253 ( .B(n1914), .A(n1945), .Z(n1992) );
  XOR U2254 ( .A(n1982), .B(n1930), .Z(n1945) );
  XOR U2255 ( .A(n1994), .B(n1995), .Z(n1930) );
  XOR U2256 ( .A(n1996), .B(n1997), .Z(n1995) );
  XOR U2257 ( .A(n1998), .B(n1981), .Z(n1914) );
  XNOR U2258 ( .A(n1999), .B(n2000), .Z(n1851) );
  XNOR U2259 ( .A(n2001), .B(n1997), .Z(n2000) );
  XNOR U2260 ( .A(n1997), .B(n1999), .Z(n1920) );
  XNOR U2261 ( .A(n1925), .B(n2002), .Z(n1986) );
  XNOR U2262 ( .A(n2003), .B(n1985), .Z(n2002) );
  OR U2263 ( .A(n1910), .B(n1924), .Z(n1985) );
  XNOR U2264 ( .A(n1982), .B(n1925), .Z(n1924) );
  XOR U2265 ( .A(n1899), .B(n1993), .Z(n1910) );
  IV U2266 ( .A(n1907), .Z(n1993) );
  XOR U2267 ( .A(n1981), .B(n2004), .Z(n1907) );
  XNOR U2268 ( .A(n2001), .B(n1994), .Z(n2004) );
  XOR U2269 ( .A(key[626]), .B(\w0[4][114] ), .Z(n1994) );
  XNOR U2270 ( .A(n811), .B(n2005), .Z(\w0[4][114] ) );
  XOR U2271 ( .A(n2006), .B(n2007), .Z(n2005) );
  XOR U2272 ( .A(n2008), .B(n814), .Z(n811) );
  IV U2273 ( .A(n1889), .Z(n1981) );
  XNOR U2274 ( .A(n1999), .B(n2009), .Z(n1889) );
  XNOR U2275 ( .A(n1997), .B(n2010), .Z(n2009) );
  ANDN U2276 ( .B(n1998), .A(n1844), .Z(n2003) );
  IV U2277 ( .A(n1899), .Z(n1998) );
  XNOR U2278 ( .A(n1999), .B(n2011), .Z(n1899) );
  XNOR U2279 ( .A(n1997), .B(n2012), .Z(n2011) );
  XOR U2280 ( .A(n1844), .B(n2013), .Z(n1997) );
  XOR U2281 ( .A(key[630]), .B(\w0[4][118] ), .Z(n2013) );
  XNOR U2282 ( .A(n1400), .B(n2014), .Z(\w0[4][118] ) );
  XNOR U2283 ( .A(n1407), .B(n2015), .Z(n2014) );
  XNOR U2284 ( .A(n2016), .B(n796), .Z(n1400) );
  XOR U2285 ( .A(n1408), .B(n820), .Z(n796) );
  IV U2286 ( .A(n1982), .Z(n1844) );
  XOR U2287 ( .A(key[629]), .B(\w0[4][117] ), .Z(n1999) );
  XNOR U2288 ( .A(n1406), .B(n2017), .Z(\w0[4][117] ) );
  XOR U2289 ( .A(n2018), .B(n2019), .Z(n2017) );
  XNOR U2290 ( .A(n1418), .B(n799), .Z(n1406) );
  XOR U2291 ( .A(n2020), .B(n2021), .Z(n1925) );
  XNOR U2292 ( .A(n2012), .B(n2010), .Z(n2021) );
  XOR U2293 ( .A(key[631]), .B(\w0[4][119] ), .Z(n2010) );
  XNOR U2294 ( .A(n1411), .B(n2022), .Z(\w0[4][119] ) );
  XOR U2295 ( .A(n2023), .B(n2016), .Z(n2022) );
  XNOR U2296 ( .A(n823), .B(n2024), .Z(n2016) );
  XOR U2297 ( .A(n1402), .B(n2025), .Z(n1411) );
  XOR U2298 ( .A(key[628]), .B(\w0[4][116] ), .Z(n2012) );
  XOR U2299 ( .A(n2026), .B(n2027), .Z(\w0[4][116] ) );
  XOR U2300 ( .A(n1420), .B(n1417), .Z(n2027) );
  XNOR U2301 ( .A(n1426), .B(n785), .Z(n1417) );
  XOR U2302 ( .A(n823), .B(n2019), .Z(n1420) );
  XNOR U2303 ( .A(n2028), .B(n2029), .Z(n2026) );
  XNOR U2304 ( .A(n1982), .B(n1996), .Z(n2020) );
  XOR U2305 ( .A(n2001), .B(n2030), .Z(n1996) );
  XOR U2306 ( .A(key[627]), .B(\w0[4][115] ), .Z(n2030) );
  XOR U2307 ( .A(n2031), .B(n2032), .Z(\w0[4][115] ) );
  XNOR U2308 ( .A(n2033), .B(n1424), .Z(n2032) );
  XOR U2309 ( .A(n823), .B(n2029), .Z(n1424) );
  XOR U2310 ( .A(n1391), .B(n812), .Z(n2031) );
  XOR U2311 ( .A(n805), .B(n1390), .Z(n812) );
  XOR U2312 ( .A(key[625]), .B(\w0[4][113] ), .Z(n2001) );
  XNOR U2313 ( .A(n824), .B(n2034), .Z(\w0[4][113] ) );
  XNOR U2314 ( .A(n815), .B(n1435), .Z(n2034) );
  XOR U2315 ( .A(n808), .B(n1434), .Z(n824) );
  XOR U2316 ( .A(key[624]), .B(\w0[4][112] ), .Z(n1982) );
  XNOR U2317 ( .A(n1414), .B(n2035), .Z(\w0[4][112] ) );
  XNOR U2318 ( .A(n2036), .B(n810), .Z(n2035) );
  XOR U2319 ( .A(n2037), .B(n2038), .Z(out[15]) );
  XNOR U2320 ( .A(n4), .B(n2039), .Z(n2038) );
  XNOR U2321 ( .A(n3), .B(n2040), .Z(n2037) );
  XOR U2322 ( .A(key[527]), .B(n5), .Z(n2040) );
  XNOR U2323 ( .A(n2041), .B(n2042), .Z(out[14]) );
  XOR U2324 ( .A(key[526]), .B(n3), .Z(n2042) );
  XOR U2325 ( .A(n63), .B(n2043), .Z(n3) );
  IV U2326 ( .A(n2044), .Z(n63) );
  XOR U2327 ( .A(n2045), .B(n2046), .Z(out[13]) );
  XNOR U2328 ( .A(n2039), .B(n2047), .Z(n2046) );
  XNOR U2329 ( .A(n2048), .B(n61), .Z(n2047) );
  XNOR U2330 ( .A(n2049), .B(n2050), .Z(n2039) );
  XNOR U2331 ( .A(n2051), .B(n2052), .Z(n2050) );
  OR U2332 ( .A(n2053), .B(n2054), .Z(n2052) );
  XOR U2333 ( .A(n2055), .B(n2056), .Z(n2045) );
  XOR U2334 ( .A(key[525]), .B(n2057), .Z(n2056) );
  AND U2335 ( .A(n2058), .B(n2059), .Z(n2055) );
  XNOR U2336 ( .A(n2060), .B(n2061), .Z(out[12]) );
  XOR U2337 ( .A(key[524]), .B(n61), .Z(n2061) );
  XNOR U2338 ( .A(n2049), .B(n2062), .Z(n61) );
  XOR U2339 ( .A(n2063), .B(n2064), .Z(n2062) );
  ANDN U2340 ( .B(n2065), .A(n2066), .Z(n2063) );
  XNOR U2341 ( .A(n2067), .B(n2068), .Z(n2049) );
  XNOR U2342 ( .A(n2069), .B(n2070), .Z(n2068) );
  NAND U2343 ( .A(n2071), .B(n2072), .Z(n2070) );
  XOR U2344 ( .A(n2073), .B(n2074), .Z(out[127]) );
  XOR U2345 ( .A(n2075), .B(n2076), .Z(n2073) );
  XOR U2346 ( .A(key[639]), .B(n2077), .Z(n2076) );
  XNOR U2347 ( .A(n2078), .B(n2079), .Z(out[126]) );
  XNOR U2348 ( .A(key[638]), .B(n2080), .Z(n2079) );
  XOR U2349 ( .A(n2081), .B(n2082), .Z(out[125]) );
  XNOR U2350 ( .A(n2083), .B(n2084), .Z(n2082) );
  XOR U2351 ( .A(n2075), .B(n2085), .Z(n2084) );
  XNOR U2352 ( .A(n2087), .B(n2088), .Z(n2086) );
  NANDN U2353 ( .A(n2089), .B(n2090), .Z(n2088) );
  XOR U2354 ( .A(n2092), .B(n2093), .Z(n2081) );
  XOR U2355 ( .A(key[637]), .B(n2094), .Z(n2093) );
  ANDN U2356 ( .B(n2095), .A(n2096), .Z(n2092) );
  XNOR U2357 ( .A(n2097), .B(n2098), .Z(out[124]) );
  XNOR U2358 ( .A(key[636]), .B(n2099), .Z(n2098) );
  XOR U2359 ( .A(n2100), .B(n2101), .Z(out[123]) );
  XNOR U2360 ( .A(n2102), .B(n2078), .Z(n2101) );
  XNOR U2361 ( .A(n2103), .B(n2104), .Z(n2078) );
  XNOR U2362 ( .A(n2105), .B(n2094), .Z(n2104) );
  ANDN U2363 ( .B(n2106), .A(n2107), .Z(n2094) );
  NOR U2364 ( .A(n2108), .B(n2109), .Z(n2105) );
  XNOR U2365 ( .A(n2110), .B(n2111), .Z(n2100) );
  XOR U2366 ( .A(key[635]), .B(n2077), .Z(n2111) );
  XOR U2367 ( .A(key[634]), .B(n2097), .Z(out[122]) );
  XNOR U2368 ( .A(n2112), .B(n2113), .Z(n2097) );
  XOR U2369 ( .A(n2114), .B(n2074), .Z(out[121]) );
  XNOR U2370 ( .A(n2103), .B(n2115), .Z(n2102) );
  XNOR U2371 ( .A(n2116), .B(n2117), .Z(n2115) );
  NANDN U2372 ( .A(n2118), .B(n2090), .Z(n2117) );
  XNOR U2373 ( .A(n2085), .B(n2119), .Z(n2103) );
  XNOR U2374 ( .A(n2120), .B(n2121), .Z(n2119) );
  NANDN U2375 ( .A(n2122), .B(n2123), .Z(n2121) );
  XOR U2376 ( .A(n2113), .B(n2110), .Z(n2080) );
  XNOR U2377 ( .A(n2085), .B(n2124), .Z(n2110) );
  XNOR U2378 ( .A(n2116), .B(n2125), .Z(n2124) );
  NANDN U2379 ( .A(n2126), .B(n2127), .Z(n2125) );
  OR U2380 ( .A(n2128), .B(n2129), .Z(n2116) );
  XOR U2381 ( .A(n2130), .B(n2120), .Z(n2085) );
  NANDN U2382 ( .A(n2131), .B(n2132), .Z(n2120) );
  ANDN U2383 ( .B(n2133), .A(n2134), .Z(n2130) );
  XNOR U2384 ( .A(key[633]), .B(n2112), .Z(n2114) );
  IV U2385 ( .A(n2077), .Z(n2112) );
  XOR U2386 ( .A(n2135), .B(n2136), .Z(n2077) );
  XNOR U2387 ( .A(n2137), .B(n2138), .Z(n2136) );
  NAND U2388 ( .A(n2095), .B(n2139), .Z(n2138) );
  XNOR U2389 ( .A(n2083), .B(n2140), .Z(out[120]) );
  XOR U2390 ( .A(key[632]), .B(n2113), .Z(n2140) );
  XNOR U2391 ( .A(n2135), .B(n2141), .Z(n2113) );
  XOR U2392 ( .A(n2142), .B(n2087), .Z(n2141) );
  OR U2393 ( .A(n2143), .B(n2128), .Z(n2087) );
  XNOR U2394 ( .A(n2090), .B(n2127), .Z(n2128) );
  ANDN U2395 ( .B(n2144), .A(n2145), .Z(n2142) );
  IV U2396 ( .A(n2099), .Z(n2083) );
  XOR U2397 ( .A(n2091), .B(n2146), .Z(n2099) );
  XOR U2398 ( .A(n2147), .B(n2137), .Z(n2146) );
  XNOR U2399 ( .A(n2109), .B(n2095), .Z(n2106) );
  NOR U2400 ( .A(n2149), .B(n2109), .Z(n2147) );
  XNOR U2401 ( .A(n2135), .B(n2150), .Z(n2091) );
  XNOR U2402 ( .A(n2151), .B(n2152), .Z(n2150) );
  NANDN U2403 ( .A(n2122), .B(n2153), .Z(n2152) );
  XOR U2404 ( .A(n2154), .B(n2151), .Z(n2135) );
  OR U2405 ( .A(n2131), .B(n2155), .Z(n2151) );
  XOR U2406 ( .A(n2156), .B(n2122), .Z(n2131) );
  XNOR U2407 ( .A(n2127), .B(n2095), .Z(n2122) );
  XOR U2408 ( .A(n2157), .B(n2158), .Z(n2095) );
  NANDN U2409 ( .A(n2159), .B(n2160), .Z(n2158) );
  IV U2410 ( .A(n2145), .Z(n2127) );
  XNOR U2411 ( .A(n2161), .B(n2162), .Z(n2145) );
  NANDN U2412 ( .A(n2159), .B(n2163), .Z(n2162) );
  ANDN U2413 ( .B(n2156), .A(n2164), .Z(n2154) );
  IV U2414 ( .A(n2134), .Z(n2156) );
  XOR U2415 ( .A(n2109), .B(n2090), .Z(n2134) );
  XNOR U2416 ( .A(n2165), .B(n2161), .Z(n2090) );
  NANDN U2417 ( .A(n2166), .B(n2167), .Z(n2161) );
  XOR U2418 ( .A(n2163), .B(n2168), .Z(n2167) );
  ANDN U2419 ( .B(n2168), .A(n2169), .Z(n2165) );
  XOR U2420 ( .A(n2170), .B(n2157), .Z(n2109) );
  NANDN U2421 ( .A(n2166), .B(n2171), .Z(n2157) );
  XOR U2422 ( .A(n2172), .B(n2160), .Z(n2171) );
  XNOR U2423 ( .A(n2173), .B(n2174), .Z(n2159) );
  XOR U2424 ( .A(n2175), .B(n2176), .Z(n2174) );
  XNOR U2425 ( .A(n2177), .B(n2178), .Z(n2173) );
  XNOR U2426 ( .A(n2179), .B(n2180), .Z(n2178) );
  ANDN U2427 ( .B(n2172), .A(n2176), .Z(n2179) );
  ANDN U2428 ( .B(n2172), .A(n2169), .Z(n2170) );
  XNOR U2429 ( .A(n2175), .B(n2181), .Z(n2169) );
  XOR U2430 ( .A(n2182), .B(n2180), .Z(n2181) );
  NAND U2431 ( .A(n2183), .B(n2184), .Z(n2180) );
  XNOR U2432 ( .A(n2177), .B(n2160), .Z(n2184) );
  IV U2433 ( .A(n2172), .Z(n2177) );
  XNOR U2434 ( .A(n2163), .B(n2176), .Z(n2183) );
  IV U2435 ( .A(n2168), .Z(n2176) );
  XOR U2436 ( .A(n2185), .B(n2186), .Z(n2168) );
  XNOR U2437 ( .A(n2187), .B(n2188), .Z(n2186) );
  XNOR U2438 ( .A(n2189), .B(n2190), .Z(n2185) );
  NOR U2439 ( .A(n2108), .B(n2149), .Z(n2189) );
  AND U2440 ( .A(n2160), .B(n2163), .Z(n2182) );
  XNOR U2441 ( .A(n2160), .B(n2163), .Z(n2175) );
  XNOR U2442 ( .A(n2191), .B(n2192), .Z(n2163) );
  XNOR U2443 ( .A(n2193), .B(n2188), .Z(n2192) );
  XOR U2444 ( .A(n2194), .B(n2195), .Z(n2191) );
  XNOR U2445 ( .A(n2196), .B(n2190), .Z(n2195) );
  OR U2446 ( .A(n2107), .B(n2148), .Z(n2190) );
  XOR U2447 ( .A(n2149), .B(n2139), .Z(n2148) );
  XNOR U2448 ( .A(n2108), .B(n2096), .Z(n2107) );
  ANDN U2449 ( .B(n2139), .A(n2096), .Z(n2196) );
  XNOR U2450 ( .A(n2197), .B(n2198), .Z(n2160) );
  XNOR U2451 ( .A(n2188), .B(n2199), .Z(n2198) );
  XOR U2452 ( .A(n2118), .B(n2194), .Z(n2199) );
  XNOR U2453 ( .A(n2149), .B(n2200), .Z(n2188) );
  XNOR U2454 ( .A(n2201), .B(n2202), .Z(n2197) );
  XNOR U2455 ( .A(n2203), .B(n2204), .Z(n2202) );
  ANDN U2456 ( .B(n2144), .A(n2126), .Z(n2203) );
  XNOR U2457 ( .A(n2205), .B(n2206), .Z(n2172) );
  XNOR U2458 ( .A(n2193), .B(n2207), .Z(n2206) );
  XNOR U2459 ( .A(n2126), .B(n2187), .Z(n2207) );
  XOR U2460 ( .A(n2194), .B(n2208), .Z(n2187) );
  XNOR U2461 ( .A(n2209), .B(n2210), .Z(n2208) );
  NAND U2462 ( .A(n2153), .B(n2123), .Z(n2210) );
  XNOR U2463 ( .A(n2211), .B(n2209), .Z(n2194) );
  NANDN U2464 ( .A(n2155), .B(n2132), .Z(n2209) );
  XOR U2465 ( .A(n2133), .B(n2123), .Z(n2132) );
  XNOR U2466 ( .A(n2212), .B(n2096), .Z(n2123) );
  XOR U2467 ( .A(n2164), .B(n2153), .Z(n2155) );
  XOR U2468 ( .A(n2144), .B(n2139), .Z(n2153) );
  ANDN U2469 ( .B(n2133), .A(n2164), .Z(n2211) );
  XOR U2470 ( .A(n2201), .B(n2149), .Z(n2164) );
  XOR U2471 ( .A(n2213), .B(n2214), .Z(n2149) );
  XOR U2472 ( .A(n2215), .B(n2216), .Z(n2214) );
  XOR U2473 ( .A(n2217), .B(n2200), .Z(n2133) );
  XNOR U2474 ( .A(n2218), .B(n2219), .Z(n2096) );
  XNOR U2475 ( .A(n2220), .B(n2216), .Z(n2219) );
  XNOR U2476 ( .A(n2216), .B(n2218), .Z(n2139) );
  XNOR U2477 ( .A(n2144), .B(n2221), .Z(n2205) );
  XNOR U2478 ( .A(n2222), .B(n2204), .Z(n2221) );
  OR U2479 ( .A(n2129), .B(n2143), .Z(n2204) );
  XNOR U2480 ( .A(n2201), .B(n2144), .Z(n2143) );
  XOR U2481 ( .A(n2118), .B(n2212), .Z(n2129) );
  IV U2482 ( .A(n2126), .Z(n2212) );
  XOR U2483 ( .A(n2200), .B(n2223), .Z(n2126) );
  XNOR U2484 ( .A(n2220), .B(n2213), .Z(n2223) );
  XOR U2485 ( .A(key[634]), .B(\w0[4][122] ), .Z(n2213) );
  XOR U2486 ( .A(n2224), .B(n2225), .Z(\w0[4][122] ) );
  XNOR U2487 ( .A(n805), .B(n815), .Z(n2225) );
  XNOR U2488 ( .A(n2007), .B(n1392), .Z(n815) );
  IV U2489 ( .A(n1431), .Z(n2007) );
  XNOR U2490 ( .A(n2226), .B(n2227), .Z(n805) );
  XOR U2491 ( .A(n2228), .B(n2229), .Z(n2227) );
  XNOR U2492 ( .A(n2230), .B(n2231), .Z(n2226) );
  XOR U2493 ( .A(n2008), .B(n1425), .Z(n2224) );
  IV U2494 ( .A(n1430), .Z(n2008) );
  IV U2495 ( .A(n2108), .Z(n2200) );
  XNOR U2496 ( .A(n2218), .B(n2232), .Z(n2108) );
  XNOR U2497 ( .A(n2216), .B(n2233), .Z(n2232) );
  ANDN U2498 ( .B(n2217), .A(n2089), .Z(n2222) );
  IV U2499 ( .A(n2118), .Z(n2217) );
  XNOR U2500 ( .A(n2218), .B(n2234), .Z(n2118) );
  XNOR U2501 ( .A(n2216), .B(n2235), .Z(n2234) );
  XOR U2502 ( .A(n2089), .B(n2236), .Z(n2216) );
  XOR U2503 ( .A(key[638]), .B(\w0[4][126] ), .Z(n2236) );
  XNOR U2504 ( .A(n2015), .B(n2237), .Z(\w0[4][126] ) );
  XOR U2505 ( .A(n2238), .B(n2239), .Z(n1408) );
  XNOR U2506 ( .A(n2018), .B(n792), .Z(n819) );
  XOR U2507 ( .A(n2036), .B(n2025), .Z(n792) );
  XNOR U2508 ( .A(n2240), .B(n2241), .Z(n2025) );
  XNOR U2509 ( .A(n2242), .B(n2243), .Z(n2241) );
  XOR U2510 ( .A(n2230), .B(n2228), .Z(n2240) );
  IV U2511 ( .A(n2244), .Z(n2228) );
  XNOR U2512 ( .A(n1399), .B(n1407), .Z(n2018) );
  XNOR U2513 ( .A(n2245), .B(n2246), .Z(n1407) );
  XOR U2514 ( .A(n2247), .B(n1413), .Z(n2015) );
  IV U2515 ( .A(n2201), .Z(n2089) );
  XOR U2516 ( .A(key[637]), .B(\w0[4][125] ), .Z(n2218) );
  XOR U2517 ( .A(n2248), .B(n2249), .Z(\w0[4][125] ) );
  XNOR U2518 ( .A(n798), .B(n820), .Z(n2249) );
  XOR U2519 ( .A(n2231), .B(n2242), .Z(n820) );
  XNOR U2520 ( .A(n2251), .B(n2252), .Z(n2250) );
  ANDN U2521 ( .B(n2253), .A(n2254), .Z(n2251) );
  XNOR U2522 ( .A(n1405), .B(n2019), .Z(n798) );
  XNOR U2523 ( .A(n2256), .B(n2257), .Z(n2019) );
  XOR U2524 ( .A(n2258), .B(n2259), .Z(n2257) );
  XNOR U2525 ( .A(n2260), .B(n2261), .Z(n2256) );
  XOR U2526 ( .A(n2262), .B(n2263), .Z(n2261) );
  ANDN U2527 ( .B(n2264), .A(n2265), .Z(n2263) );
  XNOR U2528 ( .A(n1399), .B(n1418), .Z(n2248) );
  XNOR U2529 ( .A(n2266), .B(n2267), .Z(n1418) );
  XNOR U2530 ( .A(n2268), .B(n2269), .Z(n2267) );
  XNOR U2531 ( .A(n2270), .B(n2271), .Z(n2266) );
  XOR U2532 ( .A(n2272), .B(n2273), .Z(n2271) );
  ANDN U2533 ( .B(n2274), .A(n2275), .Z(n2273) );
  XOR U2534 ( .A(n2276), .B(n2277), .Z(n1399) );
  XOR U2535 ( .A(n2278), .B(n2279), .Z(n2144) );
  XNOR U2536 ( .A(n2235), .B(n2233), .Z(n2279) );
  XOR U2537 ( .A(key[639]), .B(\w0[4][127] ), .Z(n2233) );
  XNOR U2538 ( .A(n795), .B(n2280), .Z(\w0[4][127] ) );
  XNOR U2539 ( .A(n821), .B(n1402), .Z(n2280) );
  XOR U2540 ( .A(n2281), .B(n2282), .Z(n1402) );
  XOR U2541 ( .A(n2239), .B(n2269), .Z(n2282) );
  XNOR U2542 ( .A(n2283), .B(n2284), .Z(n2269) );
  XNOR U2543 ( .A(n2285), .B(n2286), .Z(n2284) );
  NANDN U2544 ( .A(n2287), .B(n2288), .Z(n2286) );
  XOR U2545 ( .A(n2289), .B(n2290), .Z(n2281) );
  XOR U2546 ( .A(n2036), .B(n2023), .Z(n821) );
  XNOR U2547 ( .A(n1413), .B(n2024), .Z(n795) );
  XNOR U2548 ( .A(n2291), .B(n2292), .Z(n2024) );
  XOR U2549 ( .A(n2246), .B(n2259), .Z(n2292) );
  XNOR U2550 ( .A(n2293), .B(n2294), .Z(n2259) );
  XNOR U2551 ( .A(n2295), .B(n2296), .Z(n2294) );
  NANDN U2552 ( .A(n2297), .B(n2298), .Z(n2296) );
  XOR U2553 ( .A(n2299), .B(n2300), .Z(n2291) );
  XNOR U2554 ( .A(n2301), .B(n2302), .Z(n1413) );
  XNOR U2555 ( .A(n2277), .B(n2303), .Z(n2302) );
  XOR U2556 ( .A(n2304), .B(n2305), .Z(n2301) );
  XOR U2557 ( .A(key[636]), .B(\w0[4][124] ), .Z(n2235) );
  XOR U2558 ( .A(n2306), .B(n2307), .Z(\w0[4][124] ) );
  XOR U2559 ( .A(n2028), .B(n783), .Z(n2307) );
  XOR U2560 ( .A(n1419), .B(n2029), .Z(n783) );
  XOR U2561 ( .A(n1431), .B(n2258), .Z(n2029) );
  XOR U2562 ( .A(n2299), .B(n2308), .Z(n1431) );
  IV U2563 ( .A(n2309), .Z(n2299) );
  XOR U2564 ( .A(n2247), .B(n1405), .Z(n2028) );
  XNOR U2565 ( .A(n2310), .B(n2311), .Z(n1405) );
  XOR U2566 ( .A(n2312), .B(n2303), .Z(n2311) );
  XNOR U2567 ( .A(n2313), .B(n2314), .Z(n2303) );
  XNOR U2568 ( .A(n2315), .B(n2316), .Z(n2314) );
  NANDN U2569 ( .A(n2317), .B(n2318), .Z(n2316) );
  XNOR U2570 ( .A(n2319), .B(n2320), .Z(n2310) );
  XOR U2571 ( .A(n2321), .B(n2322), .Z(n2320) );
  ANDN U2572 ( .B(n2323), .A(n2324), .Z(n2322) );
  XOR U2573 ( .A(n1426), .B(n786), .Z(n2306) );
  XOR U2574 ( .A(n2036), .B(n799), .Z(n786) );
  XNOR U2575 ( .A(n2325), .B(n2326), .Z(n799) );
  XNOR U2576 ( .A(n2327), .B(n2243), .Z(n2326) );
  XNOR U2577 ( .A(n2328), .B(n2329), .Z(n2243) );
  XNOR U2578 ( .A(n2330), .B(n2331), .Z(n2329) );
  NANDN U2579 ( .A(n2332), .B(n2333), .Z(n2331) );
  XNOR U2580 ( .A(n2334), .B(n2335), .Z(n2325) );
  XOR U2581 ( .A(n2252), .B(n2336), .Z(n2335) );
  ANDN U2582 ( .B(n2337), .A(n2338), .Z(n2336) );
  ANDN U2583 ( .B(n2339), .A(n2340), .Z(n2252) );
  XOR U2584 ( .A(n2270), .B(n1430), .Z(n1426) );
  XOR U2585 ( .A(n2289), .B(n2341), .Z(n1430) );
  XNOR U2586 ( .A(n2201), .B(n2215), .Z(n2278) );
  XOR U2587 ( .A(n2220), .B(n2342), .Z(n2215) );
  XOR U2588 ( .A(key[635]), .B(\w0[4][123] ), .Z(n2342) );
  XOR U2589 ( .A(n2343), .B(n2344), .Z(\w0[4][123] ) );
  XOR U2590 ( .A(n1390), .B(n2033), .Z(n2344) );
  XOR U2591 ( .A(n2023), .B(n1419), .Z(n2033) );
  XOR U2592 ( .A(n1392), .B(n2312), .Z(n1419) );
  IV U2593 ( .A(n2247), .Z(n2023) );
  XOR U2594 ( .A(n2345), .B(n2346), .Z(n1390) );
  XOR U2595 ( .A(n2290), .B(n2347), .Z(n2346) );
  IV U2596 ( .A(n2348), .Z(n2290) );
  XNOR U2597 ( .A(n2289), .B(n2238), .Z(n2345) );
  XNOR U2598 ( .A(n2350), .B(n2272), .Z(n2349) );
  ANDN U2599 ( .B(n2351), .A(n2352), .Z(n2272) );
  ANDN U2600 ( .B(n2353), .A(n2354), .Z(n2350) );
  XOR U2601 ( .A(n807), .B(n804), .Z(n2343) );
  IV U2602 ( .A(n2006), .Z(n804) );
  XOR U2603 ( .A(n1391), .B(n1425), .Z(n2006) );
  XOR U2604 ( .A(n2356), .B(n2357), .Z(n1425) );
  XNOR U2605 ( .A(n2358), .B(n2359), .Z(n2357) );
  XNOR U2606 ( .A(n2276), .B(n2360), .Z(n2356) );
  XNOR U2607 ( .A(n2362), .B(n2321), .Z(n2361) );
  ANDN U2608 ( .B(n2363), .A(n2364), .Z(n2321) );
  ANDN U2609 ( .B(n2365), .A(n2366), .Z(n2362) );
  XOR U2610 ( .A(n2368), .B(n2369), .Z(n1391) );
  XNOR U2611 ( .A(n2370), .B(n2371), .Z(n2369) );
  XNOR U2612 ( .A(n2245), .B(n2309), .Z(n2368) );
  XNOR U2613 ( .A(n2373), .B(n2262), .Z(n2372) );
  ANDN U2614 ( .B(n2374), .A(n2375), .Z(n2262) );
  ANDN U2615 ( .B(n2376), .A(n2377), .Z(n2373) );
  XOR U2616 ( .A(n2334), .B(n2379), .Z(n2036) );
  XOR U2617 ( .A(n2334), .B(n814), .Z(n785) );
  XNOR U2618 ( .A(n2328), .B(n2380), .Z(n2334) );
  XNOR U2619 ( .A(n2381), .B(n2382), .Z(n2380) );
  ANDN U2620 ( .B(n2383), .A(n2254), .Z(n2381) );
  IV U2621 ( .A(n2384), .Z(n2254) );
  XNOR U2622 ( .A(n2385), .B(n2386), .Z(n2328) );
  XNOR U2623 ( .A(n2387), .B(n2388), .Z(n2386) );
  NANDN U2624 ( .A(n2389), .B(n2390), .Z(n2388) );
  XOR U2625 ( .A(key[633]), .B(\w0[4][121] ), .Z(n2220) );
  XOR U2626 ( .A(n2391), .B(n2392), .Z(\w0[4][121] ) );
  XOR U2627 ( .A(n810), .B(n1434), .Z(n2392) );
  XNOR U2628 ( .A(n2239), .B(n2393), .Z(n1434) );
  XOR U2629 ( .A(n2289), .B(n2348), .Z(n2393) );
  XOR U2630 ( .A(n2355), .B(n2394), .Z(n2348) );
  XNOR U2631 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2632 ( .A(n2397), .B(n2288), .Z(n2396) );
  XNOR U2633 ( .A(n2268), .B(n2398), .Z(n2355) );
  XNOR U2634 ( .A(n2399), .B(n2400), .Z(n2398) );
  NANDN U2635 ( .A(n2401), .B(n2402), .Z(n2400) );
  XNOR U2636 ( .A(n2403), .B(n2404), .Z(n2289) );
  XOR U2637 ( .A(n2405), .B(n2406), .Z(n2404) );
  NANDN U2638 ( .A(n2407), .B(n2274), .Z(n2406) );
  XNOR U2639 ( .A(n2341), .B(n2347), .Z(n2239) );
  XOR U2640 ( .A(n2268), .B(n2408), .Z(n2347) );
  XNOR U2641 ( .A(n2395), .B(n2409), .Z(n2408) );
  NANDN U2642 ( .A(n2410), .B(n2411), .Z(n2409) );
  OR U2643 ( .A(n2412), .B(n2413), .Z(n2395) );
  XOR U2644 ( .A(n2414), .B(n2399), .Z(n2268) );
  NANDN U2645 ( .A(n2415), .B(n2416), .Z(n2399) );
  ANDN U2646 ( .B(n2417), .A(n2418), .Z(n2414) );
  IV U2647 ( .A(n2419), .Z(n2341) );
  XNOR U2648 ( .A(n1429), .B(n1435), .Z(n810) );
  XNOR U2649 ( .A(n2246), .B(n2420), .Z(n1435) );
  XNOR U2650 ( .A(n2309), .B(n2370), .Z(n2420) );
  IV U2651 ( .A(n2300), .Z(n2370) );
  XOR U2652 ( .A(n2378), .B(n2421), .Z(n2300) );
  XNOR U2653 ( .A(n2422), .B(n2423), .Z(n2421) );
  NAND U2654 ( .A(n2424), .B(n2298), .Z(n2423) );
  XNOR U2655 ( .A(n2260), .B(n2425), .Z(n2378) );
  XNOR U2656 ( .A(n2426), .B(n2427), .Z(n2425) );
  NANDN U2657 ( .A(n2428), .B(n2429), .Z(n2427) );
  XNOR U2658 ( .A(n2430), .B(n2431), .Z(n2309) );
  XNOR U2659 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2660 ( .A(n2434), .B(n2264), .Z(n2433) );
  XNOR U2661 ( .A(n2371), .B(n2308), .Z(n2246) );
  XNOR U2662 ( .A(n2260), .B(n2435), .Z(n2371) );
  XNOR U2663 ( .A(n2422), .B(n2436), .Z(n2435) );
  NANDN U2664 ( .A(n2437), .B(n2438), .Z(n2436) );
  OR U2665 ( .A(n2439), .B(n2440), .Z(n2422) );
  XOR U2666 ( .A(n2441), .B(n2426), .Z(n2260) );
  OR U2667 ( .A(n2442), .B(n2443), .Z(n2426) );
  ANDN U2668 ( .B(n2444), .A(n2445), .Z(n2441) );
  IV U2669 ( .A(n2446), .Z(n1429) );
  XOR U2670 ( .A(n2304), .B(n2447), .Z(n1392) );
  IV U2671 ( .A(n2360), .Z(n2304) );
  XOR U2672 ( .A(key[632]), .B(\w0[4][120] ), .Z(n2201) );
  XOR U2673 ( .A(n2448), .B(n2449), .Z(\w0[4][120] ) );
  XNOR U2674 ( .A(n2247), .B(n1414), .Z(n2449) );
  XOR U2675 ( .A(n1401), .B(n823), .Z(n1414) );
  XOR U2676 ( .A(n2308), .B(n2258), .Z(n823) );
  XOR U2677 ( .A(n2293), .B(n2450), .Z(n2258) );
  XOR U2678 ( .A(n2451), .B(n2432), .Z(n2450) );
  NANDN U2679 ( .A(n2452), .B(n2374), .Z(n2432) );
  XOR U2680 ( .A(n2376), .B(n2264), .Z(n2374) );
  AND U2681 ( .A(n2453), .B(n2376), .Z(n2451) );
  XNOR U2682 ( .A(n2430), .B(n2454), .Z(n2293) );
  XNOR U2683 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2684 ( .A(n2429), .B(n2457), .Z(n2456) );
  XOR U2685 ( .A(n2430), .B(n2458), .Z(n2308) );
  XOR U2686 ( .A(n2459), .B(n2295), .Z(n2458) );
  OR U2687 ( .A(n2439), .B(n2460), .Z(n2295) );
  XNOR U2688 ( .A(n2298), .B(n2438), .Z(n2439) );
  ANDN U2689 ( .B(n2438), .A(n2461), .Z(n2459) );
  XOR U2690 ( .A(n2462), .B(n2455), .Z(n2430) );
  NANDN U2691 ( .A(n2443), .B(n2463), .Z(n2455) );
  XNOR U2692 ( .A(n2444), .B(n2429), .Z(n2443) );
  XOR U2693 ( .A(n2438), .B(n2264), .Z(n2429) );
  XOR U2694 ( .A(n2464), .B(n2465), .Z(n2264) );
  NANDN U2695 ( .A(n2466), .B(n2467), .Z(n2465) );
  XOR U2696 ( .A(n2468), .B(n2469), .Z(n2438) );
  NANDN U2697 ( .A(n2466), .B(n2470), .Z(n2469) );
  AND U2698 ( .A(n2471), .B(n2444), .Z(n2462) );
  XOR U2699 ( .A(n2376), .B(n2298), .Z(n2444) );
  XNOR U2700 ( .A(n2472), .B(n2468), .Z(n2298) );
  NANDN U2701 ( .A(n2473), .B(n2474), .Z(n2468) );
  XOR U2702 ( .A(n2470), .B(n2475), .Z(n2474) );
  ANDN U2703 ( .B(n2475), .A(n2476), .Z(n2472) );
  XNOR U2704 ( .A(n2477), .B(n2464), .Z(n2376) );
  NANDN U2705 ( .A(n2473), .B(n2478), .Z(n2464) );
  XOR U2706 ( .A(n2479), .B(n2467), .Z(n2478) );
  XNOR U2707 ( .A(n2480), .B(n2481), .Z(n2466) );
  XOR U2708 ( .A(n2482), .B(n2483), .Z(n2481) );
  XNOR U2709 ( .A(n2484), .B(n2485), .Z(n2480) );
  XNOR U2710 ( .A(n2486), .B(n2487), .Z(n2485) );
  ANDN U2711 ( .B(n2479), .A(n2483), .Z(n2486) );
  ANDN U2712 ( .B(n2479), .A(n2476), .Z(n2477) );
  XNOR U2713 ( .A(n2482), .B(n2488), .Z(n2476) );
  XOR U2714 ( .A(n2489), .B(n2487), .Z(n2488) );
  NAND U2715 ( .A(n2490), .B(n2491), .Z(n2487) );
  XNOR U2716 ( .A(n2484), .B(n2467), .Z(n2491) );
  IV U2717 ( .A(n2479), .Z(n2484) );
  XNOR U2718 ( .A(n2470), .B(n2483), .Z(n2490) );
  IV U2719 ( .A(n2475), .Z(n2483) );
  XOR U2720 ( .A(n2492), .B(n2493), .Z(n2475) );
  XNOR U2721 ( .A(n2494), .B(n2495), .Z(n2493) );
  XNOR U2722 ( .A(n2496), .B(n2497), .Z(n2492) );
  ANDN U2723 ( .B(n2453), .A(n2377), .Z(n2496) );
  AND U2724 ( .A(n2467), .B(n2470), .Z(n2489) );
  XNOR U2725 ( .A(n2467), .B(n2470), .Z(n2482) );
  XNOR U2726 ( .A(n2498), .B(n2499), .Z(n2470) );
  XOR U2727 ( .A(n2500), .B(n2495), .Z(n2499) );
  XNOR U2728 ( .A(n2501), .B(n2502), .Z(n2498) );
  XNOR U2729 ( .A(n2503), .B(n2497), .Z(n2502) );
  OR U2730 ( .A(n2375), .B(n2452), .Z(n2497) );
  XNOR U2731 ( .A(n2504), .B(n2453), .Z(n2452) );
  XNOR U2732 ( .A(n2377), .B(n2265), .Z(n2375) );
  ANDN U2733 ( .B(n2505), .A(n2434), .Z(n2503) );
  XNOR U2734 ( .A(n2506), .B(n2507), .Z(n2467) );
  XNOR U2735 ( .A(n2495), .B(n2508), .Z(n2507) );
  XNOR U2736 ( .A(n2424), .B(n2500), .Z(n2508) );
  XNOR U2737 ( .A(n2377), .B(n2453), .Z(n2495) );
  XOR U2738 ( .A(n2297), .B(n2509), .Z(n2506) );
  XNOR U2739 ( .A(n2510), .B(n2511), .Z(n2509) );
  ANDN U2740 ( .B(n2512), .A(n2461), .Z(n2510) );
  XNOR U2741 ( .A(n2513), .B(n2514), .Z(n2479) );
  XNOR U2742 ( .A(n2494), .B(n2515), .Z(n2514) );
  XNOR U2743 ( .A(n2501), .B(n2516), .Z(n2515) );
  XNOR U2744 ( .A(n2265), .B(n2504), .Z(n2501) );
  XOR U2745 ( .A(n2500), .B(n2517), .Z(n2494) );
  XNOR U2746 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2747 ( .A(n2428), .B(n2457), .Z(n2519) );
  XNOR U2748 ( .A(n2520), .B(n2518), .Z(n2500) );
  NANDN U2749 ( .A(n2442), .B(n2463), .Z(n2518) );
  XOR U2750 ( .A(n2471), .B(n2457), .Z(n2463) );
  XNOR U2751 ( .A(n2434), .B(n2516), .Z(n2457) );
  IV U2752 ( .A(n2504), .Z(n2434) );
  XOR U2753 ( .A(n2521), .B(n2522), .Z(n2504) );
  XOR U2754 ( .A(n2523), .B(n2428), .Z(n2442) );
  XNOR U2755 ( .A(n2505), .B(n2512), .Z(n2428) );
  IV U2756 ( .A(n2265), .Z(n2505) );
  XOR U2757 ( .A(n2524), .B(n2525), .Z(n2265) );
  ANDN U2758 ( .B(n2471), .A(n2445), .Z(n2520) );
  IV U2759 ( .A(n2523), .Z(n2445) );
  XNOR U2760 ( .A(n2437), .B(n2526), .Z(n2513) );
  XNOR U2761 ( .A(n2527), .B(n2511), .Z(n2526) );
  OR U2762 ( .A(n2440), .B(n2460), .Z(n2511) );
  XNOR U2763 ( .A(n2297), .B(n2461), .Z(n2460) );
  IV U2764 ( .A(n2516), .Z(n2461) );
  XOR U2765 ( .A(n2528), .B(n2529), .Z(n2516) );
  XNOR U2766 ( .A(n2530), .B(n2531), .Z(n2529) );
  XNOR U2767 ( .A(n2532), .B(n2297), .Z(n2528) );
  XNOR U2768 ( .A(n2424), .B(n2512), .Z(n2440) );
  IV U2769 ( .A(n2437), .Z(n2512) );
  ANDN U2770 ( .B(n2424), .A(n2297), .Z(n2527) );
  XOR U2771 ( .A(n2530), .B(n2525), .Z(n2424) );
  XNOR U2772 ( .A(n2521), .B(n2533), .Z(n2525) );
  XOR U2773 ( .A(n2534), .B(n2535), .Z(n2530) );
  XOR U2774 ( .A(n2536), .B(n2537), .Z(n2535) );
  XNOR U2775 ( .A(n2538), .B(n2539), .Z(n2534) );
  XNOR U2776 ( .A(key[428]), .B(n2540), .Z(n2539) );
  XNOR U2777 ( .A(n2541), .B(n2542), .Z(n2437) );
  XOR U2778 ( .A(n2377), .B(n2524), .Z(n2542) );
  XOR U2779 ( .A(n2533), .B(n2543), .Z(n2377) );
  XOR U2780 ( .A(n2532), .B(n2521), .Z(n2543) );
  XNOR U2781 ( .A(n2544), .B(n2545), .Z(n2521) );
  XOR U2782 ( .A(n2546), .B(n2547), .Z(n2545) );
  XOR U2783 ( .A(n2548), .B(n2549), .Z(n2544) );
  XNOR U2784 ( .A(key[429]), .B(n2550), .Z(n2549) );
  XOR U2785 ( .A(n2551), .B(n2552), .Z(n2532) );
  XOR U2786 ( .A(n2553), .B(n2554), .Z(n2552) );
  XNOR U2787 ( .A(key[431]), .B(n2555), .Z(n2551) );
  IV U2788 ( .A(n2522), .Z(n2533) );
  XNOR U2789 ( .A(n2297), .B(n2453), .Z(n2471) );
  XNOR U2790 ( .A(n2531), .B(n2556), .Z(n2453) );
  XNOR U2791 ( .A(n2522), .B(n2541), .Z(n2556) );
  XOR U2792 ( .A(n2557), .B(n2558), .Z(n2541) );
  XNOR U2793 ( .A(n2559), .B(n2560), .Z(n2558) );
  XNOR U2794 ( .A(n2561), .B(n2562), .Z(n2557) );
  XOR U2795 ( .A(key[426]), .B(n2563), .Z(n2562) );
  XOR U2796 ( .A(n2564), .B(n2565), .Z(n2522) );
  XOR U2797 ( .A(n2297), .B(n2566), .Z(n2565) );
  XNOR U2798 ( .A(n2567), .B(n2568), .Z(n2564) );
  XNOR U2799 ( .A(key[430]), .B(n2569), .Z(n2568) );
  XOR U2800 ( .A(n2570), .B(n2571), .Z(n2531) );
  XOR U2801 ( .A(n2572), .B(n2573), .Z(n2571) );
  XOR U2802 ( .A(n2574), .B(n2524), .Z(n2573) );
  XNOR U2803 ( .A(n2575), .B(n2576), .Z(n2524) );
  XOR U2804 ( .A(n2577), .B(n2578), .Z(n2576) );
  XNOR U2805 ( .A(key[425]), .B(n2580), .Z(n2579) );
  XNOR U2806 ( .A(n2582), .B(n2583), .Z(n2570) );
  XNOR U2807 ( .A(key[427]), .B(n2584), .Z(n2583) );
  XNOR U2808 ( .A(n2585), .B(n2586), .Z(n2297) );
  XOR U2809 ( .A(n2587), .B(n2588), .Z(n2586) );
  XOR U2810 ( .A(n2589), .B(n2590), .Z(n2585) );
  XNOR U2811 ( .A(key[424]), .B(n2591), .Z(n2590) );
  XOR U2812 ( .A(n2270), .B(n2419), .Z(n1401) );
  XOR U2813 ( .A(n2403), .B(n2592), .Z(n2419) );
  XOR U2814 ( .A(n2593), .B(n2285), .Z(n2592) );
  OR U2815 ( .A(n2594), .B(n2412), .Z(n2285) );
  XNOR U2816 ( .A(n2288), .B(n2411), .Z(n2412) );
  ANDN U2817 ( .B(n2411), .A(n2595), .Z(n2593) );
  XNOR U2818 ( .A(n2283), .B(n2596), .Z(n2270) );
  XNOR U2819 ( .A(n2597), .B(n2405), .Z(n2596) );
  XOR U2820 ( .A(n2599), .B(n2274), .Z(n2351) );
  ANDN U2821 ( .B(n2600), .A(n2354), .Z(n2597) );
  IV U2822 ( .A(n2599), .Z(n2354) );
  XNOR U2823 ( .A(n2403), .B(n2601), .Z(n2283) );
  XNOR U2824 ( .A(n2602), .B(n2603), .Z(n2601) );
  NANDN U2825 ( .A(n2401), .B(n2604), .Z(n2603) );
  XOR U2826 ( .A(n2605), .B(n2602), .Z(n2403) );
  OR U2827 ( .A(n2415), .B(n2606), .Z(n2602) );
  XNOR U2828 ( .A(n2418), .B(n2401), .Z(n2415) );
  XNOR U2829 ( .A(n2411), .B(n2274), .Z(n2401) );
  XOR U2830 ( .A(n2607), .B(n2608), .Z(n2274) );
  NANDN U2831 ( .A(n2609), .B(n2610), .Z(n2608) );
  XOR U2832 ( .A(n2611), .B(n2612), .Z(n2411) );
  NANDN U2833 ( .A(n2609), .B(n2613), .Z(n2612) );
  NOR U2834 ( .A(n2418), .B(n2614), .Z(n2605) );
  XNOR U2835 ( .A(n2599), .B(n2288), .Z(n2418) );
  XNOR U2836 ( .A(n2615), .B(n2611), .Z(n2288) );
  NANDN U2837 ( .A(n2616), .B(n2617), .Z(n2611) );
  XOR U2838 ( .A(n2613), .B(n2618), .Z(n2617) );
  ANDN U2839 ( .B(n2618), .A(n2619), .Z(n2615) );
  XNOR U2840 ( .A(n2620), .B(n2607), .Z(n2599) );
  NANDN U2841 ( .A(n2616), .B(n2621), .Z(n2607) );
  XOR U2842 ( .A(n2622), .B(n2610), .Z(n2621) );
  XNOR U2843 ( .A(n2623), .B(n2624), .Z(n2609) );
  XOR U2844 ( .A(n2625), .B(n2626), .Z(n2624) );
  XNOR U2845 ( .A(n2627), .B(n2628), .Z(n2623) );
  XNOR U2846 ( .A(n2629), .B(n2630), .Z(n2628) );
  ANDN U2847 ( .B(n2622), .A(n2626), .Z(n2629) );
  ANDN U2848 ( .B(n2622), .A(n2619), .Z(n2620) );
  XNOR U2849 ( .A(n2625), .B(n2631), .Z(n2619) );
  XOR U2850 ( .A(n2632), .B(n2630), .Z(n2631) );
  NAND U2851 ( .A(n2633), .B(n2634), .Z(n2630) );
  XNOR U2852 ( .A(n2627), .B(n2610), .Z(n2634) );
  IV U2853 ( .A(n2622), .Z(n2627) );
  XNOR U2854 ( .A(n2613), .B(n2626), .Z(n2633) );
  IV U2855 ( .A(n2618), .Z(n2626) );
  XOR U2856 ( .A(n2635), .B(n2636), .Z(n2618) );
  XNOR U2857 ( .A(n2637), .B(n2638), .Z(n2636) );
  XNOR U2858 ( .A(n2639), .B(n2640), .Z(n2635) );
  ANDN U2859 ( .B(n2600), .A(n2641), .Z(n2639) );
  AND U2860 ( .A(n2610), .B(n2613), .Z(n2632) );
  XNOR U2861 ( .A(n2610), .B(n2613), .Z(n2625) );
  XNOR U2862 ( .A(n2642), .B(n2643), .Z(n2613) );
  XNOR U2863 ( .A(n2644), .B(n2638), .Z(n2643) );
  XOR U2864 ( .A(n2645), .B(n2646), .Z(n2642) );
  XNOR U2865 ( .A(n2647), .B(n2640), .Z(n2646) );
  OR U2866 ( .A(n2352), .B(n2598), .Z(n2640) );
  XNOR U2867 ( .A(n2600), .B(n2648), .Z(n2598) );
  XNOR U2868 ( .A(n2641), .B(n2275), .Z(n2352) );
  ANDN U2869 ( .B(n2649), .A(n2407), .Z(n2647) );
  XNOR U2870 ( .A(n2650), .B(n2651), .Z(n2610) );
  XNOR U2871 ( .A(n2638), .B(n2652), .Z(n2651) );
  XOR U2872 ( .A(n2397), .B(n2645), .Z(n2652) );
  XNOR U2873 ( .A(n2600), .B(n2641), .Z(n2638) );
  XOR U2874 ( .A(n2287), .B(n2653), .Z(n2650) );
  XNOR U2875 ( .A(n2654), .B(n2655), .Z(n2653) );
  ANDN U2876 ( .B(n2656), .A(n2595), .Z(n2654) );
  XNOR U2877 ( .A(n2657), .B(n2658), .Z(n2622) );
  XNOR U2878 ( .A(n2644), .B(n2659), .Z(n2658) );
  XNOR U2879 ( .A(n2410), .B(n2637), .Z(n2659) );
  XOR U2880 ( .A(n2645), .B(n2660), .Z(n2637) );
  XNOR U2881 ( .A(n2661), .B(n2662), .Z(n2660) );
  NAND U2882 ( .A(n2604), .B(n2402), .Z(n2662) );
  XNOR U2883 ( .A(n2663), .B(n2661), .Z(n2645) );
  NANDN U2884 ( .A(n2606), .B(n2416), .Z(n2661) );
  XOR U2885 ( .A(n2417), .B(n2402), .Z(n2416) );
  XNOR U2886 ( .A(n2656), .B(n2275), .Z(n2402) );
  XOR U2887 ( .A(n2614), .B(n2604), .Z(n2606) );
  XNOR U2888 ( .A(n2595), .B(n2648), .Z(n2604) );
  ANDN U2889 ( .B(n2417), .A(n2614), .Z(n2663) );
  XOR U2890 ( .A(n2287), .B(n2600), .Z(n2614) );
  XNOR U2891 ( .A(n2664), .B(n2665), .Z(n2600) );
  XNOR U2892 ( .A(n2666), .B(n2667), .Z(n2665) );
  XOR U2893 ( .A(n2648), .B(n2649), .Z(n2644) );
  IV U2894 ( .A(n2275), .Z(n2649) );
  XOR U2895 ( .A(n2668), .B(n2669), .Z(n2275) );
  XOR U2896 ( .A(n2670), .B(n2667), .Z(n2669) );
  IV U2897 ( .A(n2407), .Z(n2648) );
  XOR U2898 ( .A(n2667), .B(n2671), .Z(n2407) );
  XNOR U2899 ( .A(n2672), .B(n2673), .Z(n2657) );
  XNOR U2900 ( .A(n2674), .B(n2655), .Z(n2673) );
  OR U2901 ( .A(n2413), .B(n2594), .Z(n2655) );
  XNOR U2902 ( .A(n2287), .B(n2595), .Z(n2594) );
  IV U2903 ( .A(n2672), .Z(n2595) );
  XOR U2904 ( .A(n2397), .B(n2656), .Z(n2413) );
  IV U2905 ( .A(n2410), .Z(n2656) );
  XOR U2906 ( .A(n2353), .B(n2675), .Z(n2410) );
  XNOR U2907 ( .A(n2676), .B(n2664), .Z(n2675) );
  XOR U2908 ( .A(n2677), .B(n2678), .Z(n2664) );
  XOR U2909 ( .A(n2679), .B(n2680), .Z(n2678) );
  XOR U2910 ( .A(key[386]), .B(n2681), .Z(n2677) );
  IV U2911 ( .A(n2641), .Z(n2353) );
  XOR U2912 ( .A(n2668), .B(n2682), .Z(n2641) );
  XOR U2913 ( .A(n2667), .B(n2683), .Z(n2682) );
  NOR U2914 ( .A(n2397), .B(n2287), .Z(n2674) );
  XOR U2915 ( .A(n2668), .B(n2684), .Z(n2397) );
  XOR U2916 ( .A(n2667), .B(n2685), .Z(n2684) );
  XOR U2917 ( .A(n2686), .B(n2687), .Z(n2667) );
  XOR U2918 ( .A(n2287), .B(n2688), .Z(n2687) );
  XOR U2919 ( .A(n2689), .B(n2690), .Z(n2686) );
  XNOR U2920 ( .A(key[390]), .B(n2691), .Z(n2690) );
  IV U2921 ( .A(n2671), .Z(n2668) );
  XOR U2922 ( .A(n2692), .B(n2693), .Z(n2671) );
  XOR U2923 ( .A(n2694), .B(n2695), .Z(n2693) );
  XNOR U2924 ( .A(key[389]), .B(n2696), .Z(n2692) );
  XOR U2925 ( .A(n2697), .B(n2698), .Z(n2672) );
  XNOR U2926 ( .A(n2685), .B(n2683), .Z(n2698) );
  XNOR U2927 ( .A(n2699), .B(n2700), .Z(n2683) );
  XNOR U2928 ( .A(n2701), .B(n2702), .Z(n2700) );
  XNOR U2929 ( .A(key[391]), .B(n2703), .Z(n2699) );
  XNOR U2930 ( .A(n2704), .B(n2705), .Z(n2685) );
  XOR U2931 ( .A(n2706), .B(n2707), .Z(n2705) );
  XNOR U2932 ( .A(n2708), .B(n2709), .Z(n2704) );
  XNOR U2933 ( .A(key[388]), .B(n2710), .Z(n2709) );
  XNOR U2934 ( .A(n2287), .B(n2666), .Z(n2697) );
  XOR U2935 ( .A(n2711), .B(n2712), .Z(n2666) );
  XNOR U2936 ( .A(n2713), .B(n2714), .Z(n2712) );
  XOR U2937 ( .A(n2715), .B(n2676), .Z(n2714) );
  IV U2938 ( .A(n2670), .Z(n2676) );
  XNOR U2939 ( .A(n2716), .B(n2717), .Z(n2670) );
  XNOR U2940 ( .A(n2718), .B(n2719), .Z(n2717) );
  XNOR U2941 ( .A(key[385]), .B(n2720), .Z(n2716) );
  XOR U2942 ( .A(n2721), .B(n2722), .Z(n2711) );
  XNOR U2943 ( .A(key[387]), .B(n2723), .Z(n2722) );
  XNOR U2944 ( .A(n2724), .B(n2725), .Z(n2287) );
  XNOR U2945 ( .A(n2726), .B(n2727), .Z(n2725) );
  XNOR U2946 ( .A(n2447), .B(n2312), .Z(n2247) );
  XOR U2947 ( .A(n2313), .B(n2729), .Z(n2312) );
  XOR U2948 ( .A(n2730), .B(n2731), .Z(n2729) );
  AND U2949 ( .A(n2732), .B(n2365), .Z(n2730) );
  XNOR U2950 ( .A(n2733), .B(n2734), .Z(n2313) );
  XNOR U2951 ( .A(n2735), .B(n2736), .Z(n2734) );
  NAND U2952 ( .A(n2737), .B(n2738), .Z(n2736) );
  XOR U2953 ( .A(n2446), .B(n808), .Z(n2448) );
  XNOR U2954 ( .A(n2242), .B(n2739), .Z(n808) );
  XOR U2955 ( .A(n2230), .B(n2244), .Z(n2739) );
  XOR U2956 ( .A(n2255), .B(n2740), .Z(n2244) );
  XNOR U2957 ( .A(n2741), .B(n2742), .Z(n2740) );
  NANDN U2958 ( .A(n2743), .B(n2333), .Z(n2742) );
  XNOR U2959 ( .A(n2327), .B(n2744), .Z(n2255) );
  XNOR U2960 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2961 ( .A(n2389), .B(n2747), .Z(n2746) );
  XNOR U2962 ( .A(n2385), .B(n2748), .Z(n2230) );
  XOR U2963 ( .A(n2382), .B(n2749), .Z(n2748) );
  NANDN U2964 ( .A(n2750), .B(n2337), .Z(n2749) );
  XOR U2965 ( .A(n2384), .B(n2337), .Z(n2339) );
  XNOR U2966 ( .A(n2379), .B(n2229), .Z(n2242) );
  XOR U2967 ( .A(n2327), .B(n2752), .Z(n2229) );
  XNOR U2968 ( .A(n2741), .B(n2753), .Z(n2752) );
  NANDN U2969 ( .A(n2754), .B(n2755), .Z(n2753) );
  OR U2970 ( .A(n2756), .B(n2757), .Z(n2741) );
  XOR U2971 ( .A(n2758), .B(n2745), .Z(n2327) );
  NANDN U2972 ( .A(n2759), .B(n2760), .Z(n2745) );
  ANDN U2973 ( .B(n2761), .A(n2762), .Z(n2758) );
  XOR U2974 ( .A(n2385), .B(n2763), .Z(n2379) );
  XOR U2975 ( .A(n2764), .B(n2330), .Z(n2763) );
  OR U2976 ( .A(n2765), .B(n2756), .Z(n2330) );
  XNOR U2977 ( .A(n2333), .B(n2755), .Z(n2756) );
  ANDN U2978 ( .B(n2755), .A(n2766), .Z(n2764) );
  XOR U2979 ( .A(n2767), .B(n2387), .Z(n2385) );
  OR U2980 ( .A(n2759), .B(n2768), .Z(n2387) );
  XNOR U2981 ( .A(n2762), .B(n2389), .Z(n2759) );
  XNOR U2982 ( .A(n2755), .B(n2337), .Z(n2389) );
  XOR U2983 ( .A(n2769), .B(n2770), .Z(n2337) );
  NANDN U2984 ( .A(n2771), .B(n2772), .Z(n2770) );
  XOR U2985 ( .A(n2773), .B(n2774), .Z(n2755) );
  NANDN U2986 ( .A(n2771), .B(n2775), .Z(n2774) );
  NOR U2987 ( .A(n2762), .B(n2776), .Z(n2767) );
  XNOR U2988 ( .A(n2384), .B(n2333), .Z(n2762) );
  XNOR U2989 ( .A(n2777), .B(n2773), .Z(n2333) );
  NANDN U2990 ( .A(n2778), .B(n2779), .Z(n2773) );
  XOR U2991 ( .A(n2775), .B(n2780), .Z(n2779) );
  ANDN U2992 ( .B(n2780), .A(n2781), .Z(n2777) );
  XNOR U2993 ( .A(n2782), .B(n2769), .Z(n2384) );
  NANDN U2994 ( .A(n2778), .B(n2783), .Z(n2769) );
  XOR U2995 ( .A(n2784), .B(n2772), .Z(n2783) );
  XNOR U2996 ( .A(n2785), .B(n2786), .Z(n2771) );
  XOR U2997 ( .A(n2787), .B(n2788), .Z(n2786) );
  XNOR U2998 ( .A(n2789), .B(n2790), .Z(n2785) );
  XNOR U2999 ( .A(n2791), .B(n2792), .Z(n2790) );
  ANDN U3000 ( .B(n2784), .A(n2788), .Z(n2791) );
  ANDN U3001 ( .B(n2784), .A(n2781), .Z(n2782) );
  XNOR U3002 ( .A(n2787), .B(n2793), .Z(n2781) );
  XOR U3003 ( .A(n2794), .B(n2792), .Z(n2793) );
  NAND U3004 ( .A(n2795), .B(n2796), .Z(n2792) );
  XNOR U3005 ( .A(n2789), .B(n2772), .Z(n2796) );
  IV U3006 ( .A(n2784), .Z(n2789) );
  XNOR U3007 ( .A(n2775), .B(n2788), .Z(n2795) );
  IV U3008 ( .A(n2780), .Z(n2788) );
  XOR U3009 ( .A(n2797), .B(n2798), .Z(n2780) );
  XNOR U3010 ( .A(n2799), .B(n2800), .Z(n2798) );
  XNOR U3011 ( .A(n2801), .B(n2802), .Z(n2797) );
  ANDN U3012 ( .B(n2383), .A(n2803), .Z(n2801) );
  AND U3013 ( .A(n2772), .B(n2775), .Z(n2794) );
  XNOR U3014 ( .A(n2772), .B(n2775), .Z(n2787) );
  XNOR U3015 ( .A(n2804), .B(n2805), .Z(n2775) );
  XNOR U3016 ( .A(n2806), .B(n2800), .Z(n2805) );
  XOR U3017 ( .A(n2807), .B(n2808), .Z(n2804) );
  XNOR U3018 ( .A(n2809), .B(n2802), .Z(n2808) );
  OR U3019 ( .A(n2340), .B(n2751), .Z(n2802) );
  XNOR U3020 ( .A(n2383), .B(n2810), .Z(n2751) );
  XNOR U3021 ( .A(n2803), .B(n2338), .Z(n2340) );
  ANDN U3022 ( .B(n2811), .A(n2750), .Z(n2809) );
  XNOR U3023 ( .A(n2812), .B(n2813), .Z(n2772) );
  XNOR U3024 ( .A(n2800), .B(n2814), .Z(n2813) );
  XOR U3025 ( .A(n2743), .B(n2807), .Z(n2814) );
  XNOR U3026 ( .A(n2383), .B(n2803), .Z(n2800) );
  XOR U3027 ( .A(n2332), .B(n2815), .Z(n2812) );
  XNOR U3028 ( .A(n2816), .B(n2817), .Z(n2815) );
  ANDN U3029 ( .B(n2818), .A(n2766), .Z(n2816) );
  XNOR U3030 ( .A(n2819), .B(n2820), .Z(n2784) );
  XNOR U3031 ( .A(n2806), .B(n2821), .Z(n2820) );
  XNOR U3032 ( .A(n2754), .B(n2799), .Z(n2821) );
  XOR U3033 ( .A(n2807), .B(n2822), .Z(n2799) );
  XNOR U3034 ( .A(n2823), .B(n2824), .Z(n2822) );
  NAND U3035 ( .A(n2390), .B(n2747), .Z(n2824) );
  XNOR U3036 ( .A(n2825), .B(n2823), .Z(n2807) );
  NANDN U3037 ( .A(n2768), .B(n2760), .Z(n2823) );
  XOR U3038 ( .A(n2761), .B(n2747), .Z(n2760) );
  XNOR U3039 ( .A(n2818), .B(n2338), .Z(n2747) );
  XOR U3040 ( .A(n2776), .B(n2390), .Z(n2768) );
  XNOR U3041 ( .A(n2766), .B(n2810), .Z(n2390) );
  ANDN U3042 ( .B(n2761), .A(n2776), .Z(n2825) );
  XOR U3043 ( .A(n2332), .B(n2383), .Z(n2776) );
  XNOR U3044 ( .A(n2826), .B(n2827), .Z(n2383) );
  XNOR U3045 ( .A(n2828), .B(n2829), .Z(n2827) );
  XOR U3046 ( .A(n2810), .B(n2811), .Z(n2806) );
  IV U3047 ( .A(n2338), .Z(n2811) );
  XOR U3048 ( .A(n2830), .B(n2831), .Z(n2338) );
  XOR U3049 ( .A(n2832), .B(n2829), .Z(n2831) );
  IV U3050 ( .A(n2750), .Z(n2810) );
  XOR U3051 ( .A(n2829), .B(n2833), .Z(n2750) );
  XNOR U3052 ( .A(n2834), .B(n2835), .Z(n2819) );
  XNOR U3053 ( .A(n2836), .B(n2817), .Z(n2835) );
  OR U3054 ( .A(n2757), .B(n2765), .Z(n2817) );
  XNOR U3055 ( .A(n2332), .B(n2766), .Z(n2765) );
  IV U3056 ( .A(n2834), .Z(n2766) );
  XOR U3057 ( .A(n2743), .B(n2818), .Z(n2757) );
  IV U3058 ( .A(n2754), .Z(n2818) );
  XOR U3059 ( .A(n2253), .B(n2837), .Z(n2754) );
  XOR U3060 ( .A(n2838), .B(n2839), .Z(n2826) );
  XOR U3061 ( .A(n2840), .B(n2841), .Z(n2839) );
  XNOR U3062 ( .A(n2842), .B(n2843), .Z(n2838) );
  IV U3063 ( .A(n2803), .Z(n2253) );
  XOR U3064 ( .A(n2830), .B(n2845), .Z(n2803) );
  XOR U3065 ( .A(n2829), .B(n2846), .Z(n2845) );
  NOR U3066 ( .A(n2743), .B(n2332), .Z(n2836) );
  XOR U3067 ( .A(n2830), .B(n2847), .Z(n2743) );
  XOR U3068 ( .A(n2829), .B(n2848), .Z(n2847) );
  XOR U3069 ( .A(n2849), .B(n2850), .Z(n2829) );
  XNOR U3070 ( .A(n2332), .B(n2851), .Z(n2850) );
  XNOR U3071 ( .A(n2852), .B(n2853), .Z(n2849) );
  XNOR U3072 ( .A(key[510]), .B(n2854), .Z(n2853) );
  IV U3073 ( .A(n2833), .Z(n2830) );
  XOR U3074 ( .A(n2855), .B(n2856), .Z(n2833) );
  XOR U3075 ( .A(n2857), .B(n2858), .Z(n2856) );
  XNOR U3076 ( .A(n2859), .B(n2860), .Z(n2855) );
  XNOR U3077 ( .A(key[509]), .B(n2861), .Z(n2860) );
  XOR U3078 ( .A(n2862), .B(n2863), .Z(n2834) );
  XNOR U3079 ( .A(n2848), .B(n2846), .Z(n2863) );
  XNOR U3080 ( .A(n2864), .B(n2865), .Z(n2846) );
  XOR U3081 ( .A(n2866), .B(n2867), .Z(n2865) );
  XNOR U3082 ( .A(key[511]), .B(n2868), .Z(n2864) );
  XNOR U3083 ( .A(n2869), .B(n2870), .Z(n2848) );
  XOR U3084 ( .A(n2871), .B(n2872), .Z(n2870) );
  XNOR U3085 ( .A(n2873), .B(n2874), .Z(n2869) );
  XNOR U3086 ( .A(key[508]), .B(n2875), .Z(n2874) );
  XNOR U3087 ( .A(n2332), .B(n2828), .Z(n2862) );
  XOR U3088 ( .A(n2876), .B(n2877), .Z(n2828) );
  XNOR U3089 ( .A(n2878), .B(n2879), .Z(n2877) );
  XOR U3090 ( .A(n2880), .B(n2832), .Z(n2879) );
  XNOR U3091 ( .A(n2881), .B(n2882), .Z(n2832) );
  XOR U3092 ( .A(n2883), .B(n2884), .Z(n2882) );
  XNOR U3093 ( .A(n2885), .B(n2886), .Z(n2881) );
  XNOR U3094 ( .A(key[505]), .B(n2887), .Z(n2886) );
  XNOR U3095 ( .A(n2888), .B(n2889), .Z(n2876) );
  XNOR U3096 ( .A(key[507]), .B(n2890), .Z(n2889) );
  XNOR U3097 ( .A(n2891), .B(n2892), .Z(n2332) );
  XOR U3098 ( .A(n2893), .B(n2894), .Z(n2892) );
  XNOR U3099 ( .A(n2895), .B(n2896), .Z(n2891) );
  XNOR U3100 ( .A(key[504]), .B(n2897), .Z(n2896) );
  XNOR U3101 ( .A(n2360), .B(n2358), .Z(n2898) );
  IV U3102 ( .A(n2305), .Z(n2358) );
  XOR U3103 ( .A(n2367), .B(n2899), .Z(n2305) );
  XNOR U3104 ( .A(n2900), .B(n2901), .Z(n2899) );
  NAND U3105 ( .A(n2902), .B(n2318), .Z(n2901) );
  XNOR U3106 ( .A(n2319), .B(n2903), .Z(n2367) );
  XNOR U3107 ( .A(n2904), .B(n2905), .Z(n2903) );
  NANDN U3108 ( .A(n2906), .B(n2737), .Z(n2905) );
  XNOR U3109 ( .A(n2733), .B(n2907), .Z(n2360) );
  XNOR U3110 ( .A(n2731), .B(n2908), .Z(n2907) );
  NANDN U3111 ( .A(n2909), .B(n2323), .Z(n2908) );
  NANDN U3112 ( .A(n2910), .B(n2363), .Z(n2731) );
  XOR U3113 ( .A(n2365), .B(n2323), .Z(n2363) );
  XOR U3114 ( .A(n2359), .B(n2447), .Z(n2277) );
  XOR U3115 ( .A(n2733), .B(n2911), .Z(n2447) );
  XOR U3116 ( .A(n2912), .B(n2315), .Z(n2911) );
  OR U3117 ( .A(n2913), .B(n2914), .Z(n2315) );
  ANDN U3118 ( .B(n2915), .A(n2916), .Z(n2912) );
  XOR U3119 ( .A(n2917), .B(n2735), .Z(n2733) );
  NANDN U3120 ( .A(n2918), .B(n2919), .Z(n2735) );
  AND U3121 ( .A(n2920), .B(n2921), .Z(n2917) );
  XNOR U3122 ( .A(n2319), .B(n2922), .Z(n2359) );
  XNOR U3123 ( .A(n2900), .B(n2923), .Z(n2922) );
  NANDN U3124 ( .A(n2924), .B(n2915), .Z(n2923) );
  OR U3125 ( .A(n2913), .B(n2925), .Z(n2900) );
  XNOR U3126 ( .A(n2318), .B(n2915), .Z(n2913) );
  XOR U3127 ( .A(n2926), .B(n2904), .Z(n2319) );
  OR U3128 ( .A(n2927), .B(n2918), .Z(n2904) );
  XNOR U3129 ( .A(n2921), .B(n2737), .Z(n2918) );
  XOR U3130 ( .A(n2915), .B(n2323), .Z(n2737) );
  XOR U3131 ( .A(n2928), .B(n2929), .Z(n2323) );
  NANDN U3132 ( .A(n2930), .B(n2931), .Z(n2929) );
  XOR U3133 ( .A(n2932), .B(n2933), .Z(n2915) );
  NANDN U3134 ( .A(n2930), .B(n2934), .Z(n2933) );
  ANDN U3135 ( .B(n2921), .A(n2935), .Z(n2926) );
  XOR U3136 ( .A(n2365), .B(n2318), .Z(n2921) );
  XNOR U3137 ( .A(n2936), .B(n2932), .Z(n2318) );
  NANDN U3138 ( .A(n2937), .B(n2938), .Z(n2932) );
  XOR U3139 ( .A(n2934), .B(n2939), .Z(n2938) );
  ANDN U3140 ( .B(n2939), .A(n2940), .Z(n2936) );
  XNOR U3141 ( .A(n2941), .B(n2928), .Z(n2365) );
  NANDN U3142 ( .A(n2937), .B(n2942), .Z(n2928) );
  XOR U3143 ( .A(n2943), .B(n2931), .Z(n2942) );
  XNOR U3144 ( .A(n2944), .B(n2945), .Z(n2930) );
  XOR U3145 ( .A(n2946), .B(n2947), .Z(n2945) );
  XNOR U3146 ( .A(n2948), .B(n2949), .Z(n2944) );
  XNOR U3147 ( .A(n2950), .B(n2951), .Z(n2949) );
  ANDN U3148 ( .B(n2943), .A(n2947), .Z(n2950) );
  ANDN U3149 ( .B(n2943), .A(n2940), .Z(n2941) );
  XNOR U3150 ( .A(n2946), .B(n2952), .Z(n2940) );
  XOR U3151 ( .A(n2953), .B(n2951), .Z(n2952) );
  NAND U3152 ( .A(n2954), .B(n2955), .Z(n2951) );
  XNOR U3153 ( .A(n2948), .B(n2931), .Z(n2955) );
  IV U3154 ( .A(n2943), .Z(n2948) );
  XNOR U3155 ( .A(n2934), .B(n2947), .Z(n2954) );
  IV U3156 ( .A(n2939), .Z(n2947) );
  XOR U3157 ( .A(n2956), .B(n2957), .Z(n2939) );
  XNOR U3158 ( .A(n2958), .B(n2959), .Z(n2957) );
  XNOR U3159 ( .A(n2960), .B(n2961), .Z(n2956) );
  ANDN U3160 ( .B(n2732), .A(n2366), .Z(n2960) );
  AND U3161 ( .A(n2931), .B(n2934), .Z(n2953) );
  XNOR U3162 ( .A(n2931), .B(n2934), .Z(n2946) );
  XNOR U3163 ( .A(n2962), .B(n2963), .Z(n2934) );
  XOR U3164 ( .A(n2964), .B(n2959), .Z(n2963) );
  XNOR U3165 ( .A(n2965), .B(n2966), .Z(n2962) );
  XNOR U3166 ( .A(n2967), .B(n2961), .Z(n2966) );
  OR U3167 ( .A(n2364), .B(n2910), .Z(n2961) );
  XNOR U3168 ( .A(n2968), .B(n2732), .Z(n2910) );
  XNOR U3169 ( .A(n2366), .B(n2324), .Z(n2364) );
  ANDN U3170 ( .B(n2969), .A(n2909), .Z(n2967) );
  XNOR U3171 ( .A(n2970), .B(n2971), .Z(n2931) );
  XNOR U3172 ( .A(n2959), .B(n2972), .Z(n2971) );
  XNOR U3173 ( .A(n2902), .B(n2964), .Z(n2972) );
  XNOR U3174 ( .A(n2366), .B(n2732), .Z(n2959) );
  XOR U3175 ( .A(n2317), .B(n2973), .Z(n2970) );
  XNOR U3176 ( .A(n2974), .B(n2975), .Z(n2973) );
  ANDN U3177 ( .B(n2976), .A(n2916), .Z(n2974) );
  XNOR U3178 ( .A(n2977), .B(n2978), .Z(n2943) );
  XNOR U3179 ( .A(n2958), .B(n2979), .Z(n2978) );
  XNOR U3180 ( .A(n2965), .B(n2980), .Z(n2979) );
  XNOR U3181 ( .A(n2324), .B(n2968), .Z(n2965) );
  XOR U3182 ( .A(n2964), .B(n2981), .Z(n2958) );
  XNOR U3183 ( .A(n2982), .B(n2983), .Z(n2981) );
  NANDN U3184 ( .A(n2906), .B(n2738), .Z(n2983) );
  XNOR U3185 ( .A(n2984), .B(n2982), .Z(n2964) );
  NANDN U3186 ( .A(n2927), .B(n2919), .Z(n2982) );
  XOR U3187 ( .A(n2920), .B(n2738), .Z(n2919) );
  XNOR U3188 ( .A(n2909), .B(n2980), .Z(n2738) );
  IV U3189 ( .A(n2968), .Z(n2909) );
  XOR U3190 ( .A(n2985), .B(n2986), .Z(n2968) );
  XOR U3191 ( .A(n2987), .B(n2906), .Z(n2927) );
  XNOR U3192 ( .A(n2969), .B(n2976), .Z(n2906) );
  IV U3193 ( .A(n2324), .Z(n2969) );
  XOR U3194 ( .A(n2988), .B(n2989), .Z(n2324) );
  ANDN U3195 ( .B(n2920), .A(n2935), .Z(n2984) );
  IV U3196 ( .A(n2987), .Z(n2935) );
  XNOR U3197 ( .A(n2317), .B(n2732), .Z(n2920) );
  XNOR U3198 ( .A(n2990), .B(n2991), .Z(n2732) );
  XNOR U3199 ( .A(n2986), .B(n2992), .Z(n2991) );
  XNOR U3200 ( .A(n2924), .B(n2993), .Z(n2977) );
  XNOR U3201 ( .A(n2994), .B(n2975), .Z(n2993) );
  OR U3202 ( .A(n2925), .B(n2914), .Z(n2975) );
  XNOR U3203 ( .A(n2317), .B(n2916), .Z(n2914) );
  IV U3204 ( .A(n2980), .Z(n2916) );
  XOR U3205 ( .A(n2995), .B(n2996), .Z(n2980) );
  XNOR U3206 ( .A(n2997), .B(n2990), .Z(n2996) );
  XOR U3207 ( .A(n2998), .B(n2999), .Z(n2990) );
  XNOR U3208 ( .A(n3000), .B(n3001), .Z(n2999) );
  XOR U3209 ( .A(n3002), .B(n2988), .Z(n3001) );
  XNOR U3210 ( .A(n3003), .B(n3004), .Z(n2998) );
  XOR U3211 ( .A(key[467]), .B(n3005), .Z(n3004) );
  XNOR U3212 ( .A(n3006), .B(n2317), .Z(n2995) );
  XNOR U3213 ( .A(n2902), .B(n2976), .Z(n2925) );
  IV U3214 ( .A(n2924), .Z(n2976) );
  ANDN U3215 ( .B(n2902), .A(n2317), .Z(n2994) );
  XOR U3216 ( .A(n2997), .B(n2989), .Z(n2902) );
  XNOR U3217 ( .A(n2985), .B(n3007), .Z(n2989) );
  XOR U3218 ( .A(n3008), .B(n3009), .Z(n2997) );
  XOR U3219 ( .A(n3010), .B(n3011), .Z(n3009) );
  XNOR U3220 ( .A(n3012), .B(n3013), .Z(n3008) );
  XNOR U3221 ( .A(key[468]), .B(n3014), .Z(n3013) );
  XNOR U3222 ( .A(n2992), .B(n3015), .Z(n2924) );
  XOR U3223 ( .A(n2366), .B(n2988), .Z(n3015) );
  XNOR U3224 ( .A(n3016), .B(n3017), .Z(n2988) );
  XNOR U3225 ( .A(key[465]), .B(n3020), .Z(n3016) );
  XOR U3226 ( .A(n3007), .B(n3021), .Z(n2366) );
  XOR U3227 ( .A(n3006), .B(n2985), .Z(n3021) );
  XNOR U3228 ( .A(n3022), .B(n3023), .Z(n2985) );
  XNOR U3229 ( .A(n3024), .B(n3025), .Z(n3023) );
  XNOR U3230 ( .A(key[469]), .B(n3026), .Z(n3022) );
  XOR U3231 ( .A(n3027), .B(n3028), .Z(n3006) );
  XNOR U3232 ( .A(n3029), .B(n3030), .Z(n3028) );
  XNOR U3233 ( .A(key[471]), .B(n3031), .Z(n3027) );
  IV U3234 ( .A(n2986), .Z(n3007) );
  XOR U3235 ( .A(n3032), .B(n3033), .Z(n2986) );
  XOR U3236 ( .A(n2317), .B(n3034), .Z(n3033) );
  XNOR U3237 ( .A(n3035), .B(n3036), .Z(n2317) );
  XNOR U3238 ( .A(n3037), .B(n3038), .Z(n3036) );
  XNOR U3239 ( .A(key[464]), .B(n3039), .Z(n3035) );
  XOR U3240 ( .A(n3040), .B(n3041), .Z(n3032) );
  XNOR U3241 ( .A(key[470]), .B(n3042), .Z(n3041) );
  XOR U3242 ( .A(n3043), .B(n3044), .Z(n2992) );
  XOR U3243 ( .A(n3045), .B(n3046), .Z(n3044) );
  XNOR U3244 ( .A(key[466]), .B(n3047), .Z(n3043) );
  XOR U3245 ( .A(n3048), .B(n3049), .Z(out[11]) );
  XNOR U3246 ( .A(n4), .B(n2041), .Z(n3049) );
  XNOR U3247 ( .A(n3050), .B(n3051), .Z(n2041) );
  XNOR U3248 ( .A(n3052), .B(n2057), .Z(n3051) );
  ANDN U3249 ( .B(n3053), .A(n3054), .Z(n2057) );
  NOR U3250 ( .A(n2066), .B(n3055), .Z(n3052) );
  XNOR U3251 ( .A(n2043), .B(n3056), .Z(n3048) );
  XOR U3252 ( .A(key[523]), .B(n5), .Z(n3056) );
  XOR U3253 ( .A(n3050), .B(n3057), .Z(n5) );
  XNOR U3254 ( .A(n3058), .B(n3059), .Z(n3057) );
  NANDN U3255 ( .A(n2053), .B(n3060), .Z(n3059) );
  XNOR U3256 ( .A(n2048), .B(n3061), .Z(n3050) );
  XNOR U3257 ( .A(n3062), .B(n3063), .Z(n3061) );
  NAND U3258 ( .A(n3064), .B(n2071), .Z(n3063) );
  XNOR U3259 ( .A(n2048), .B(n3065), .Z(n2043) );
  XNOR U3260 ( .A(n3058), .B(n3066), .Z(n3065) );
  NANDN U3261 ( .A(n3067), .B(n3068), .Z(n3066) );
  OR U3262 ( .A(n3069), .B(n3070), .Z(n3058) );
  XOR U3263 ( .A(n3071), .B(n3062), .Z(n2048) );
  OR U3264 ( .A(n3072), .B(n3073), .Z(n3062) );
  ANDN U3265 ( .B(n3074), .A(n3075), .Z(n3071) );
  XOR U3266 ( .A(n3076), .B(n3077), .Z(out[119]) );
  XOR U3267 ( .A(n3078), .B(n3079), .Z(n3076) );
  XOR U3268 ( .A(key[631]), .B(n3080), .Z(n3079) );
  XNOR U3269 ( .A(n3081), .B(n3082), .Z(out[118]) );
  XNOR U3270 ( .A(key[630]), .B(n3083), .Z(n3082) );
  XOR U3271 ( .A(n3084), .B(n3085), .Z(out[117]) );
  XNOR U3272 ( .A(n3086), .B(n3087), .Z(n3085) );
  XOR U3273 ( .A(n3078), .B(n3088), .Z(n3087) );
  XNOR U3274 ( .A(n3090), .B(n3091), .Z(n3089) );
  NANDN U3275 ( .A(n3092), .B(n3093), .Z(n3091) );
  XOR U3276 ( .A(n3095), .B(n3096), .Z(n3084) );
  XOR U3277 ( .A(key[629]), .B(n3097), .Z(n3096) );
  ANDN U3278 ( .B(n3098), .A(n3099), .Z(n3095) );
  XNOR U3279 ( .A(n3100), .B(n3101), .Z(out[116]) );
  XNOR U3280 ( .A(key[628]), .B(n3102), .Z(n3101) );
  XOR U3281 ( .A(n3103), .B(n3104), .Z(out[115]) );
  XNOR U3282 ( .A(n3105), .B(n3081), .Z(n3104) );
  XNOR U3283 ( .A(n3106), .B(n3107), .Z(n3081) );
  XNOR U3284 ( .A(n3108), .B(n3097), .Z(n3107) );
  ANDN U3285 ( .B(n3109), .A(n3110), .Z(n3097) );
  NOR U3286 ( .A(n3111), .B(n3112), .Z(n3108) );
  XNOR U3287 ( .A(n3113), .B(n3114), .Z(n3103) );
  XOR U3288 ( .A(key[627]), .B(n3080), .Z(n3114) );
  XOR U3289 ( .A(key[626]), .B(n3100), .Z(out[114]) );
  XNOR U3290 ( .A(n3115), .B(n3116), .Z(n3100) );
  XOR U3291 ( .A(n3117), .B(n3077), .Z(out[113]) );
  XNOR U3292 ( .A(n3106), .B(n3118), .Z(n3105) );
  XNOR U3293 ( .A(n3119), .B(n3120), .Z(n3118) );
  NANDN U3294 ( .A(n3121), .B(n3093), .Z(n3120) );
  XNOR U3295 ( .A(n3088), .B(n3122), .Z(n3106) );
  XNOR U3296 ( .A(n3123), .B(n3124), .Z(n3122) );
  NANDN U3297 ( .A(n3125), .B(n3126), .Z(n3124) );
  XOR U3298 ( .A(n3116), .B(n3113), .Z(n3083) );
  XNOR U3299 ( .A(n3088), .B(n3127), .Z(n3113) );
  XNOR U3300 ( .A(n3119), .B(n3128), .Z(n3127) );
  NANDN U3301 ( .A(n3129), .B(n3130), .Z(n3128) );
  OR U3302 ( .A(n3131), .B(n3132), .Z(n3119) );
  XOR U3303 ( .A(n3133), .B(n3123), .Z(n3088) );
  NANDN U3304 ( .A(n3134), .B(n3135), .Z(n3123) );
  ANDN U3305 ( .B(n3136), .A(n3137), .Z(n3133) );
  XNOR U3306 ( .A(key[625]), .B(n3115), .Z(n3117) );
  IV U3307 ( .A(n3080), .Z(n3115) );
  XOR U3308 ( .A(n3138), .B(n3139), .Z(n3080) );
  XNOR U3309 ( .A(n3140), .B(n3141), .Z(n3139) );
  NANDN U3310 ( .A(n3142), .B(n3098), .Z(n3141) );
  XNOR U3311 ( .A(n3086), .B(n3143), .Z(out[112]) );
  XOR U3312 ( .A(key[624]), .B(n3116), .Z(n3143) );
  XNOR U3313 ( .A(n3138), .B(n3144), .Z(n3116) );
  XOR U3314 ( .A(n3145), .B(n3090), .Z(n3144) );
  OR U3315 ( .A(n3146), .B(n3131), .Z(n3090) );
  XNOR U3316 ( .A(n3093), .B(n3130), .Z(n3131) );
  ANDN U3317 ( .B(n3147), .A(n3148), .Z(n3145) );
  IV U3318 ( .A(n3102), .Z(n3086) );
  XOR U3319 ( .A(n3094), .B(n3149), .Z(n3102) );
  XOR U3320 ( .A(n3150), .B(n3140), .Z(n3149) );
  XNOR U3321 ( .A(n3112), .B(n3098), .Z(n3109) );
  NOR U3322 ( .A(n3152), .B(n3112), .Z(n3150) );
  XNOR U3323 ( .A(n3138), .B(n3153), .Z(n3094) );
  XNOR U3324 ( .A(n3154), .B(n3155), .Z(n3153) );
  NANDN U3325 ( .A(n3125), .B(n3156), .Z(n3155) );
  XOR U3326 ( .A(n3157), .B(n3154), .Z(n3138) );
  OR U3327 ( .A(n3134), .B(n3158), .Z(n3154) );
  XOR U3328 ( .A(n3159), .B(n3125), .Z(n3134) );
  XNOR U3329 ( .A(n3130), .B(n3098), .Z(n3125) );
  XOR U3330 ( .A(n3160), .B(n3161), .Z(n3098) );
  NANDN U3331 ( .A(n3162), .B(n3163), .Z(n3161) );
  IV U3332 ( .A(n3148), .Z(n3130) );
  XNOR U3333 ( .A(n3164), .B(n3165), .Z(n3148) );
  NANDN U3334 ( .A(n3162), .B(n3166), .Z(n3165) );
  ANDN U3335 ( .B(n3159), .A(n3167), .Z(n3157) );
  IV U3336 ( .A(n3137), .Z(n3159) );
  XOR U3337 ( .A(n3112), .B(n3093), .Z(n3137) );
  XNOR U3338 ( .A(n3168), .B(n3164), .Z(n3093) );
  NANDN U3339 ( .A(n3169), .B(n3170), .Z(n3164) );
  XOR U3340 ( .A(n3166), .B(n3171), .Z(n3170) );
  ANDN U3341 ( .B(n3171), .A(n3172), .Z(n3168) );
  XOR U3342 ( .A(n3173), .B(n3160), .Z(n3112) );
  NANDN U3343 ( .A(n3169), .B(n3174), .Z(n3160) );
  XOR U3344 ( .A(n3175), .B(n3163), .Z(n3174) );
  XNOR U3345 ( .A(n3176), .B(n3177), .Z(n3162) );
  XOR U3346 ( .A(n3178), .B(n3179), .Z(n3177) );
  XNOR U3347 ( .A(n3180), .B(n3181), .Z(n3176) );
  XNOR U3348 ( .A(n3182), .B(n3183), .Z(n3181) );
  ANDN U3349 ( .B(n3175), .A(n3179), .Z(n3182) );
  ANDN U3350 ( .B(n3175), .A(n3172), .Z(n3173) );
  XNOR U3351 ( .A(n3178), .B(n3184), .Z(n3172) );
  XOR U3352 ( .A(n3185), .B(n3183), .Z(n3184) );
  NAND U3353 ( .A(n3186), .B(n3187), .Z(n3183) );
  XNOR U3354 ( .A(n3180), .B(n3163), .Z(n3187) );
  IV U3355 ( .A(n3175), .Z(n3180) );
  XNOR U3356 ( .A(n3166), .B(n3179), .Z(n3186) );
  IV U3357 ( .A(n3171), .Z(n3179) );
  XOR U3358 ( .A(n3188), .B(n3189), .Z(n3171) );
  XNOR U3359 ( .A(n3190), .B(n3191), .Z(n3189) );
  XNOR U3360 ( .A(n3192), .B(n3193), .Z(n3188) );
  ANDN U3361 ( .B(n3194), .A(n3152), .Z(n3192) );
  AND U3362 ( .A(n3163), .B(n3166), .Z(n3185) );
  XNOR U3363 ( .A(n3163), .B(n3166), .Z(n3178) );
  XNOR U3364 ( .A(n3195), .B(n3196), .Z(n3166) );
  XNOR U3365 ( .A(n3197), .B(n3191), .Z(n3196) );
  XOR U3366 ( .A(n3198), .B(n3199), .Z(n3195) );
  XNOR U3367 ( .A(n3200), .B(n3193), .Z(n3199) );
  OR U3368 ( .A(n3110), .B(n3151), .Z(n3193) );
  XNOR U3369 ( .A(n3201), .B(n3202), .Z(n3151) );
  XNOR U3370 ( .A(n3111), .B(n3099), .Z(n3110) );
  ANDN U3371 ( .B(n3203), .A(n3142), .Z(n3200) );
  XNOR U3372 ( .A(n3204), .B(n3205), .Z(n3163) );
  XNOR U3373 ( .A(n3191), .B(n3206), .Z(n3205) );
  XOR U3374 ( .A(n3121), .B(n3198), .Z(n3206) );
  XNOR U3375 ( .A(n3201), .B(n3111), .Z(n3191) );
  XNOR U3376 ( .A(n3207), .B(n3208), .Z(n3204) );
  XNOR U3377 ( .A(n3209), .B(n3210), .Z(n3208) );
  ANDN U3378 ( .B(n3147), .A(n3129), .Z(n3209) );
  XNOR U3379 ( .A(n3211), .B(n3212), .Z(n3175) );
  XNOR U3380 ( .A(n3197), .B(n3213), .Z(n3212) );
  XNOR U3381 ( .A(n3129), .B(n3190), .Z(n3213) );
  XOR U3382 ( .A(n3198), .B(n3214), .Z(n3190) );
  XNOR U3383 ( .A(n3215), .B(n3216), .Z(n3214) );
  NAND U3384 ( .A(n3156), .B(n3126), .Z(n3216) );
  XNOR U3385 ( .A(n3217), .B(n3215), .Z(n3198) );
  NANDN U3386 ( .A(n3158), .B(n3135), .Z(n3215) );
  XOR U3387 ( .A(n3136), .B(n3126), .Z(n3135) );
  XNOR U3388 ( .A(n3218), .B(n3099), .Z(n3126) );
  XOR U3389 ( .A(n3167), .B(n3156), .Z(n3158) );
  XOR U3390 ( .A(n3147), .B(n3202), .Z(n3156) );
  ANDN U3391 ( .B(n3136), .A(n3167), .Z(n3217) );
  XNOR U3392 ( .A(n3207), .B(n3201), .Z(n3167) );
  IV U3393 ( .A(n3152), .Z(n3201) );
  XNOR U3394 ( .A(n3219), .B(n3220), .Z(n3152) );
  XOR U3395 ( .A(n3221), .B(n3222), .Z(n3220) );
  XOR U3396 ( .A(n3223), .B(n3194), .Z(n3136) );
  XOR U3397 ( .A(n3202), .B(n3203), .Z(n3197) );
  IV U3398 ( .A(n3099), .Z(n3203) );
  XOR U3399 ( .A(n3224), .B(n3225), .Z(n3099) );
  XNOR U3400 ( .A(n3226), .B(n3222), .Z(n3225) );
  IV U3401 ( .A(n3142), .Z(n3202) );
  XOR U3402 ( .A(n3222), .B(n3227), .Z(n3142) );
  XNOR U3403 ( .A(n3147), .B(n3228), .Z(n3211) );
  XNOR U3404 ( .A(n3229), .B(n3210), .Z(n3228) );
  OR U3405 ( .A(n3132), .B(n3146), .Z(n3210) );
  XNOR U3406 ( .A(n3207), .B(n3147), .Z(n3146) );
  XOR U3407 ( .A(n3121), .B(n3218), .Z(n3132) );
  IV U3408 ( .A(n3129), .Z(n3218) );
  XOR U3409 ( .A(n3194), .B(n3230), .Z(n3129) );
  XOR U3410 ( .A(n3226), .B(n3219), .Z(n3230) );
  XNOR U3411 ( .A(key[594]), .B(\w0[4][82] ), .Z(n3219) );
  XNOR U3412 ( .A(n1638), .B(n3231), .Z(\w0[4][82] ) );
  XOR U3413 ( .A(n3232), .B(n211), .Z(n3231) );
  XOR U3414 ( .A(n179), .B(n3233), .Z(n211) );
  IV U3415 ( .A(n3111), .Z(n3194) );
  XOR U3416 ( .A(n3224), .B(n3234), .Z(n3111) );
  XOR U3417 ( .A(n3222), .B(n3235), .Z(n3234) );
  ANDN U3418 ( .B(n3223), .A(n3092), .Z(n3229) );
  IV U3419 ( .A(n3121), .Z(n3223) );
  XOR U3420 ( .A(n3224), .B(n3236), .Z(n3121) );
  XOR U3421 ( .A(n3222), .B(n3237), .Z(n3236) );
  XOR U3422 ( .A(n3092), .B(n3238), .Z(n3222) );
  XOR U3423 ( .A(key[598]), .B(\w0[4][86] ), .Z(n3238) );
  XNOR U3424 ( .A(n3239), .B(n3240), .Z(\w0[4][86] ) );
  XNOR U3425 ( .A(n3241), .B(n185), .Z(n3240) );
  XOR U3426 ( .A(n1626), .B(n3242), .Z(n185) );
  IV U3427 ( .A(n3207), .Z(n3092) );
  IV U3428 ( .A(n3227), .Z(n3224) );
  XOR U3429 ( .A(key[597]), .B(\w0[4][85] ), .Z(n3227) );
  XNOR U3430 ( .A(n3243), .B(n3244), .Z(\w0[4][85] ) );
  XOR U3431 ( .A(n1612), .B(n1618), .Z(n3244) );
  XNOR U3432 ( .A(n193), .B(n3241), .Z(n1612) );
  XOR U3433 ( .A(n3245), .B(n3246), .Z(n3147) );
  XNOR U3434 ( .A(n3237), .B(n3235), .Z(n3246) );
  XNOR U3435 ( .A(key[599]), .B(\w0[4][87] ), .Z(n3235) );
  XNOR U3436 ( .A(n3247), .B(n3248), .Z(\w0[4][87] ) );
  XNOR U3437 ( .A(n224), .B(n3249), .Z(n3248) );
  XNOR U3438 ( .A(key[596]), .B(\w0[4][84] ), .Z(n3237) );
  XOR U3439 ( .A(n3250), .B(n3251), .Z(\w0[4][84] ) );
  XNOR U3440 ( .A(n3252), .B(n3253), .Z(n3251) );
  XOR U3441 ( .A(n206), .B(n1631), .Z(n3250) );
  XOR U3442 ( .A(n224), .B(n1617), .Z(n206) );
  IV U3443 ( .A(n3242), .Z(n224) );
  XNOR U3444 ( .A(n3207), .B(n3221), .Z(n3245) );
  XOR U3445 ( .A(n3226), .B(n3254), .Z(n3221) );
  XOR U3446 ( .A(key[595]), .B(\w0[4][83] ), .Z(n3254) );
  XOR U3447 ( .A(n3255), .B(n3256), .Z(\w0[4][83] ) );
  XOR U3448 ( .A(n1602), .B(n3257), .Z(n3256) );
  XOR U3449 ( .A(n213), .B(n3233), .Z(n3255) );
  IV U3450 ( .A(n3258), .Z(n3233) );
  XNOR U3451 ( .A(n3242), .B(n1632), .Z(n213) );
  XOR U3452 ( .A(key[593]), .B(\w0[4][81] ), .Z(n3226) );
  XNOR U3453 ( .A(n1640), .B(n3259), .Z(\w0[4][81] ) );
  XNOR U3454 ( .A(n176), .B(n3260), .Z(n3259) );
  IV U3455 ( .A(n1604), .Z(n176) );
  XNOR U3456 ( .A(n3232), .B(n218), .Z(n1604) );
  XOR U3457 ( .A(key[592]), .B(\w0[4][80] ), .Z(n3207) );
  XOR U3458 ( .A(n222), .B(n3261), .Z(\w0[4][80] ) );
  XNOR U3459 ( .A(n1623), .B(n217), .Z(n3261) );
  XNOR U3460 ( .A(n3260), .B(n225), .Z(n217) );
  IV U3461 ( .A(n1633), .Z(n1623) );
  XOR U3462 ( .A(n3262), .B(n3263), .Z(out[111]) );
  XOR U3463 ( .A(n3264), .B(n3265), .Z(n3262) );
  XOR U3464 ( .A(key[623]), .B(n3266), .Z(n3265) );
  XNOR U3465 ( .A(n3267), .B(n3268), .Z(out[110]) );
  XNOR U3466 ( .A(key[622]), .B(n3269), .Z(n3268) );
  XOR U3467 ( .A(key[522]), .B(n2060), .Z(out[10]) );
  XNOR U3468 ( .A(n2044), .B(n4), .Z(n2060) );
  XNOR U3469 ( .A(n2067), .B(n3270), .Z(n4) );
  XNOR U3470 ( .A(n2064), .B(n3271), .Z(n3270) );
  NANDN U3471 ( .A(n3272), .B(n2059), .Z(n3271) );
  XNOR U3472 ( .A(n2066), .B(n2059), .Z(n3053) );
  XNOR U3473 ( .A(n2067), .B(n3274), .Z(n2044) );
  XOR U3474 ( .A(n3275), .B(n2051), .Z(n3274) );
  OR U3475 ( .A(n3069), .B(n3276), .Z(n2051) );
  XNOR U3476 ( .A(n2053), .B(n3067), .Z(n3069) );
  NOR U3477 ( .A(n3277), .B(n3067), .Z(n3275) );
  XOR U3478 ( .A(n3278), .B(n2069), .Z(n2067) );
  NANDN U3479 ( .A(n3073), .B(n3279), .Z(n2069) );
  XNOR U3480 ( .A(n3074), .B(n2071), .Z(n3073) );
  XNOR U3481 ( .A(n3067), .B(n2059), .Z(n2071) );
  XOR U3482 ( .A(n3280), .B(n3281), .Z(n2059) );
  NANDN U3483 ( .A(n3282), .B(n3283), .Z(n3281) );
  XNOR U3484 ( .A(n3284), .B(n3285), .Z(n3067) );
  OR U3485 ( .A(n3282), .B(n3286), .Z(n3285) );
  AND U3486 ( .A(n3074), .B(n3287), .Z(n3278) );
  XOR U3487 ( .A(n2053), .B(n2066), .Z(n3074) );
  XOR U3488 ( .A(n3288), .B(n3280), .Z(n2066) );
  NANDN U3489 ( .A(n3289), .B(n3290), .Z(n3280) );
  ANDN U3490 ( .B(n3291), .A(n3292), .Z(n3288) );
  NANDN U3491 ( .A(n3289), .B(n3294), .Z(n3284) );
  XOR U3492 ( .A(n3295), .B(n3282), .Z(n3289) );
  XNOR U3493 ( .A(n3296), .B(n3297), .Z(n3282) );
  XOR U3494 ( .A(n3298), .B(n3291), .Z(n3297) );
  XNOR U3495 ( .A(n3299), .B(n3300), .Z(n3296) );
  XNOR U3496 ( .A(n3301), .B(n3302), .Z(n3300) );
  ANDN U3497 ( .B(n3291), .A(n3303), .Z(n3301) );
  IV U3498 ( .A(n3304), .Z(n3291) );
  ANDN U3499 ( .B(n3295), .A(n3303), .Z(n3293) );
  IV U3500 ( .A(n3299), .Z(n3303) );
  IV U3501 ( .A(n3292), .Z(n3295) );
  XNOR U3502 ( .A(n3298), .B(n3305), .Z(n3292) );
  XOR U3503 ( .A(n3306), .B(n3302), .Z(n3305) );
  NAND U3504 ( .A(n3294), .B(n3290), .Z(n3302) );
  XNOR U3505 ( .A(n3283), .B(n3304), .Z(n3290) );
  XOR U3506 ( .A(n3307), .B(n3308), .Z(n3304) );
  XOR U3507 ( .A(n3309), .B(n3310), .Z(n3308) );
  XOR U3508 ( .A(n3311), .B(n3312), .Z(n3310) );
  XOR U3509 ( .A(n3068), .B(n3313), .Z(n3307) );
  XNOR U3510 ( .A(n3314), .B(n3315), .Z(n3313) );
  ANDN U3511 ( .B(n3060), .A(n2054), .Z(n3314) );
  XNOR U3512 ( .A(n3299), .B(n3286), .Z(n3294) );
  XOR U3513 ( .A(n3316), .B(n3317), .Z(n3299) );
  XNOR U3514 ( .A(n3318), .B(n3312), .Z(n3317) );
  XOR U3515 ( .A(n3319), .B(n3320), .Z(n3312) );
  XNOR U3516 ( .A(n3321), .B(n3322), .Z(n3320) );
  NAND U3517 ( .A(n2072), .B(n3064), .Z(n3322) );
  XNOR U3518 ( .A(n3323), .B(n3324), .Z(n3316) );
  ANDN U3519 ( .B(n2065), .A(n3055), .Z(n3323) );
  ANDN U3520 ( .B(n3283), .A(n3286), .Z(n3306) );
  XOR U3521 ( .A(n3286), .B(n3283), .Z(n3298) );
  XNOR U3522 ( .A(n3325), .B(n3326), .Z(n3283) );
  XNOR U3523 ( .A(n3319), .B(n3327), .Z(n3326) );
  XNOR U3524 ( .A(n3060), .B(n3318), .Z(n3327) );
  XOR U3525 ( .A(n2054), .B(n3328), .Z(n3325) );
  XNOR U3526 ( .A(n3329), .B(n3315), .Z(n3328) );
  OR U3527 ( .A(n3070), .B(n3276), .Z(n3315) );
  XNOR U3528 ( .A(n3330), .B(n3311), .Z(n3276) );
  XNOR U3529 ( .A(n3060), .B(n3068), .Z(n3070) );
  ANDN U3530 ( .B(n3068), .A(n3277), .Z(n3329) );
  IV U3531 ( .A(n3311), .Z(n3277) );
  XOR U3532 ( .A(n3331), .B(n3332), .Z(n3286) );
  XOR U3533 ( .A(n3319), .B(n3309), .Z(n3332) );
  XOR U3534 ( .A(n2058), .B(n3272), .Z(n3309) );
  XOR U3535 ( .A(n3333), .B(n3321), .Z(n3319) );
  NANDN U3536 ( .A(n3072), .B(n3279), .Z(n3321) );
  XOR U3537 ( .A(n3287), .B(n2072), .Z(n3279) );
  XNOR U3538 ( .A(n3272), .B(n3311), .Z(n2072) );
  XOR U3539 ( .A(n3334), .B(n3335), .Z(n3311) );
  XNOR U3540 ( .A(n3336), .B(n3337), .Z(n3335) );
  XOR U3541 ( .A(n3330), .B(n3338), .Z(n3334) );
  XOR U3542 ( .A(n3075), .B(n3064), .Z(n3072) );
  XOR U3543 ( .A(n2058), .B(n3068), .Z(n3064) );
  XOR U3544 ( .A(n3339), .B(n3340), .Z(n3068) );
  XNOR U3545 ( .A(n3055), .B(n3341), .Z(n3340) );
  ANDN U3546 ( .B(n3287), .A(n3075), .Z(n3333) );
  XOR U3547 ( .A(n3055), .B(n3060), .Z(n3075) );
  XOR U3548 ( .A(n3336), .B(n3342), .Z(n3060) );
  XOR U3549 ( .A(key[588]), .B(\w0[4][76] ), .Z(n3336) );
  XOR U3550 ( .A(n3343), .B(n3344), .Z(\w0[4][76] ) );
  XOR U3551 ( .A(n3253), .B(n1630), .Z(n3344) );
  XNOR U3552 ( .A(n194), .B(n1621), .Z(n1630) );
  XOR U3553 ( .A(n203), .B(n1629), .Z(n3253) );
  XNOR U3554 ( .A(n3345), .B(n219), .Z(n1629) );
  XNOR U3555 ( .A(n1632), .B(n3252), .Z(n3343) );
  XNOR U3556 ( .A(n1618), .B(n3346), .Z(n3252) );
  XNOR U3557 ( .A(n3347), .B(n3348), .Z(n1618) );
  XNOR U3558 ( .A(n3349), .B(n3350), .Z(n3348) );
  XOR U3559 ( .A(n3351), .B(n3352), .Z(n3347) );
  XNOR U3560 ( .A(n3353), .B(n3354), .Z(n3352) );
  ANDN U3561 ( .B(n3355), .A(n3356), .Z(n3354) );
  XOR U3562 ( .A(n3357), .B(n218), .Z(n1632) );
  XOR U3563 ( .A(n3330), .B(n2065), .Z(n3287) );
  XOR U3564 ( .A(n3318), .B(n3358), .Z(n3331) );
  XNOR U3565 ( .A(n3359), .B(n3324), .Z(n3358) );
  OR U3566 ( .A(n3273), .B(n3054), .Z(n3324) );
  XOR U3567 ( .A(n3055), .B(n2058), .Z(n3054) );
  XNOR U3568 ( .A(n2065), .B(n3342), .Z(n3273) );
  ANDN U3569 ( .B(n2058), .A(n3272), .Z(n3359) );
  IV U3570 ( .A(n3342), .Z(n3272) );
  XOR U3571 ( .A(n3341), .B(n3342), .Z(n2058) );
  XOR U3572 ( .A(n3055), .B(n2065), .Z(n3318) );
  XNOR U3573 ( .A(n3337), .B(n3360), .Z(n2065) );
  XNOR U3574 ( .A(n3361), .B(n3339), .Z(n3360) );
  XOR U3575 ( .A(key[586]), .B(\w0[4][74] ), .Z(n3339) );
  XOR U3576 ( .A(n3362), .B(n3363), .Z(\w0[4][74] ) );
  XOR U3577 ( .A(n3258), .B(n1638), .Z(n3363) );
  XOR U3578 ( .A(n178), .B(n219), .Z(n1638) );
  XNOR U3579 ( .A(n3364), .B(n3365), .Z(n219) );
  XNOR U3580 ( .A(n3366), .B(n3367), .Z(n3258) );
  XOR U3581 ( .A(n3368), .B(n3369), .Z(n3367) );
  XOR U3582 ( .A(n3370), .B(n3371), .Z(n3366) );
  XNOR U3583 ( .A(n218), .B(n210), .Z(n3362) );
  XOR U3584 ( .A(n3372), .B(n3373), .Z(n218) );
  XNOR U3585 ( .A(n3341), .B(n3374), .Z(n3337) );
  XOR U3586 ( .A(key[587]), .B(\w0[4][75] ), .Z(n3374) );
  XOR U3587 ( .A(n3375), .B(n3376), .Z(\w0[4][75] ) );
  XOR U3588 ( .A(n3257), .B(n1637), .Z(n3376) );
  XNOR U3589 ( .A(n203), .B(n1621), .Z(n1637) );
  XOR U3590 ( .A(n3377), .B(n3378), .Z(n203) );
  XNOR U3591 ( .A(n1631), .B(n1642), .Z(n3257) );
  XNOR U3592 ( .A(n3350), .B(n3232), .Z(n1631) );
  XNOR U3593 ( .A(n179), .B(n1602), .Z(n3375) );
  XNOR U3594 ( .A(n210), .B(n177), .Z(n1602) );
  XNOR U3595 ( .A(n3379), .B(n3380), .Z(n177) );
  XOR U3596 ( .A(n3381), .B(n3382), .Z(n3380) );
  XOR U3597 ( .A(n3365), .B(n3383), .Z(n3379) );
  XOR U3598 ( .A(n3384), .B(n3385), .Z(n210) );
  XOR U3599 ( .A(n3388), .B(n3389), .Z(n3384) );
  XOR U3600 ( .A(n3390), .B(n3391), .Z(n179) );
  XOR U3601 ( .A(n3392), .B(n3393), .Z(n3391) );
  XOR U3602 ( .A(n3372), .B(n3394), .Z(n3390) );
  XOR U3603 ( .A(key[585]), .B(\w0[4][73] ), .Z(n3341) );
  XOR U3604 ( .A(n3395), .B(n3396), .Z(\w0[4][73] ) );
  XOR U3605 ( .A(n225), .B(n1640), .Z(n3396) );
  XNOR U3606 ( .A(n216), .B(n223), .Z(n1640) );
  XNOR U3607 ( .A(n3397), .B(n3398), .Z(n223) );
  XNOR U3608 ( .A(n3365), .B(n3383), .Z(n3398) );
  XOR U3609 ( .A(n3399), .B(n3400), .Z(n225) );
  XNOR U3610 ( .A(n3372), .B(n3394), .Z(n3400) );
  XNOR U3611 ( .A(n3378), .B(n3232), .Z(n3395) );
  XOR U3612 ( .A(n3370), .B(n3401), .Z(n3232) );
  IV U3613 ( .A(n178), .Z(n3378) );
  XNOR U3614 ( .A(n3338), .B(n3342), .Z(n3055) );
  XNOR U3615 ( .A(n3403), .B(n3361), .Z(n3342) );
  XOR U3616 ( .A(n2054), .B(n3404), .Z(n3361) );
  XOR U3617 ( .A(key[590]), .B(\w0[4][78] ), .Z(n3404) );
  XNOR U3618 ( .A(n1610), .B(n3405), .Z(\w0[4][78] ) );
  XNOR U3619 ( .A(n193), .B(n3239), .Z(n3405) );
  XOR U3620 ( .A(n3249), .B(n1614), .Z(n3239) );
  XOR U3621 ( .A(n188), .B(n192), .Z(n1614) );
  XOR U3622 ( .A(n3406), .B(n3382), .Z(n192) );
  XNOR U3623 ( .A(n3407), .B(n3408), .Z(n3382) );
  XNOR U3624 ( .A(n3409), .B(n3410), .Z(n3408) );
  ANDN U3625 ( .B(n3411), .A(n3412), .Z(n3409) );
  XNOR U3626 ( .A(n1625), .B(n1642), .Z(n3249) );
  XOR U3627 ( .A(n3413), .B(n3414), .Z(n1625) );
  XOR U3628 ( .A(n3415), .B(n3368), .Z(n3414) );
  XNOR U3629 ( .A(n3417), .B(n3418), .Z(n3416) );
  OR U3630 ( .A(n3419), .B(n3420), .Z(n3418) );
  XOR U3631 ( .A(n3399), .B(n3393), .Z(n193) );
  XNOR U3632 ( .A(n3422), .B(n3423), .Z(n3393) );
  XNOR U3633 ( .A(n3424), .B(n3425), .Z(n3423) );
  ANDN U3634 ( .B(n3426), .A(n3427), .Z(n3424) );
  XNOR U3635 ( .A(n199), .B(n3428), .Z(n1610) );
  IV U3636 ( .A(n3330), .Z(n2054) );
  XOR U3637 ( .A(key[584]), .B(\w0[4][72] ), .Z(n3330) );
  XOR U3638 ( .A(n3429), .B(n3430), .Z(\w0[4][72] ) );
  XNOR U3639 ( .A(n3260), .B(n3428), .Z(n3430) );
  IV U3640 ( .A(n1621), .Z(n3428) );
  XOR U3641 ( .A(n3368), .B(n3431), .Z(n3260) );
  XOR U3642 ( .A(n3370), .B(n3415), .Z(n3431) );
  XOR U3643 ( .A(n3432), .B(n3433), .Z(n3370) );
  XOR U3644 ( .A(n3434), .B(n3435), .Z(n3433) );
  ANDN U3645 ( .B(n3436), .A(n3356), .Z(n3434) );
  XOR U3646 ( .A(n3437), .B(n3438), .Z(n3368) );
  XOR U3647 ( .A(n3439), .B(n3440), .Z(n3438) );
  NOR U3648 ( .A(n3441), .B(n3419), .Z(n3439) );
  XOR U3649 ( .A(n197), .B(n216), .Z(n3429) );
  XOR U3650 ( .A(n3387), .B(n3442), .Z(n216) );
  XOR U3651 ( .A(n3443), .B(n3389), .Z(n3442) );
  XOR U3652 ( .A(n1633), .B(n3242), .Z(n197) );
  XOR U3653 ( .A(n3373), .B(n3357), .Z(n3242) );
  XOR U3654 ( .A(key[589]), .B(\w0[4][77] ), .Z(n3403) );
  XOR U3655 ( .A(n3444), .B(n3445), .Z(\w0[4][77] ) );
  XOR U3656 ( .A(n1617), .B(n3243), .Z(n3445) );
  XOR U3657 ( .A(n194), .B(n1616), .Z(n3243) );
  XNOR U3658 ( .A(n3446), .B(n3447), .Z(n1616) );
  XNOR U3659 ( .A(n3448), .B(n3449), .Z(n3447) );
  XNOR U3660 ( .A(n3345), .B(n3450), .Z(n3446) );
  XOR U3661 ( .A(n3410), .B(n3451), .Z(n3450) );
  ANDN U3662 ( .B(n3452), .A(n3453), .Z(n3451) );
  ANDN U3663 ( .B(n3454), .A(n3455), .Z(n3410) );
  XNOR U3664 ( .A(n3456), .B(n3457), .Z(n3345) );
  XNOR U3665 ( .A(n3458), .B(n3459), .Z(n3457) );
  ANDN U3666 ( .B(n3460), .A(n3412), .Z(n3458) );
  IV U3667 ( .A(n3461), .Z(n3412) );
  XOR U3668 ( .A(n3462), .B(n3463), .Z(n194) );
  XNOR U3669 ( .A(n3464), .B(n3377), .Z(n3463) );
  XNOR U3670 ( .A(n3465), .B(n3466), .Z(n3462) );
  XNOR U3671 ( .A(n3467), .B(n3468), .Z(n3466) );
  ANDN U3672 ( .B(n3469), .A(n3470), .Z(n3467) );
  XNOR U3673 ( .A(n3471), .B(n3472), .Z(n1617) );
  XOR U3674 ( .A(n3473), .B(n3357), .Z(n3472) );
  XOR U3675 ( .A(n3474), .B(n3475), .Z(n3357) );
  XNOR U3676 ( .A(n3476), .B(n3477), .Z(n3475) );
  ANDN U3677 ( .B(n3478), .A(n3427), .Z(n3476) );
  IV U3678 ( .A(n3479), .Z(n3427) );
  XNOR U3679 ( .A(n3480), .B(n3481), .Z(n3471) );
  XOR U3680 ( .A(n3425), .B(n3482), .Z(n3481) );
  ANDN U3681 ( .B(n3483), .A(n3484), .Z(n3482) );
  ANDN U3682 ( .B(n3485), .A(n3486), .Z(n3425) );
  XNOR U3683 ( .A(n3241), .B(n188), .Z(n3444) );
  XOR U3684 ( .A(n3386), .B(n3443), .Z(n188) );
  XNOR U3685 ( .A(n3487), .B(n3488), .Z(n3386) );
  XNOR U3686 ( .A(n3468), .B(n3489), .Z(n3488) );
  OR U3687 ( .A(n3490), .B(n3491), .Z(n3489) );
  NANDN U3688 ( .A(n3492), .B(n3493), .Z(n3468) );
  XNOR U3689 ( .A(n3369), .B(n3415), .Z(n3241) );
  XOR U3690 ( .A(n3371), .B(n3401), .Z(n3415) );
  XOR U3691 ( .A(n3349), .B(n3494), .Z(n3371) );
  XNOR U3692 ( .A(n3440), .B(n3495), .Z(n3494) );
  NANDN U3693 ( .A(n3496), .B(n3497), .Z(n3495) );
  OR U3694 ( .A(n3498), .B(n3499), .Z(n3440) );
  XNOR U3695 ( .A(n3437), .B(n3500), .Z(n3369) );
  XOR U3696 ( .A(n3501), .B(n3353), .Z(n3500) );
  OR U3697 ( .A(n3502), .B(n3503), .Z(n3353) );
  ANDN U3698 ( .B(n3504), .A(n3505), .Z(n3501) );
  XNOR U3699 ( .A(n3349), .B(n3506), .Z(n3437) );
  XNOR U3700 ( .A(n3507), .B(n3508), .Z(n3506) );
  NAND U3701 ( .A(n3509), .B(n3510), .Z(n3508) );
  XOR U3702 ( .A(n3511), .B(n3507), .Z(n3349) );
  NANDN U3703 ( .A(n3512), .B(n3513), .Z(n3507) );
  ANDN U3704 ( .B(n3514), .A(n3515), .Z(n3511) );
  XOR U3705 ( .A(key[591]), .B(\w0[4][79] ), .Z(n3338) );
  XNOR U3706 ( .A(n3247), .B(n3516), .Z(\w0[4][79] ) );
  XOR U3707 ( .A(n1626), .B(n222), .Z(n3516) );
  XOR U3708 ( .A(n1621), .B(n3346), .Z(n222) );
  IV U3709 ( .A(n1642), .Z(n3346) );
  XNOR U3710 ( .A(n3401), .B(n3350), .Z(n1642) );
  XNOR U3711 ( .A(n3421), .B(n3517), .Z(n3350) );
  XNOR U3712 ( .A(n3435), .B(n3518), .Z(n3517) );
  NANDN U3713 ( .A(n3519), .B(n3504), .Z(n3518) );
  OR U3714 ( .A(n3520), .B(n3502), .Z(n3435) );
  XNOR U3715 ( .A(n3504), .B(n3521), .Z(n3502) );
  XNOR U3716 ( .A(n3432), .B(n3522), .Z(n3421) );
  XNOR U3717 ( .A(n3523), .B(n3524), .Z(n3522) );
  NAND U3718 ( .A(n3510), .B(n3525), .Z(n3524) );
  XNOR U3719 ( .A(n3432), .B(n3526), .Z(n3401) );
  XOR U3720 ( .A(n3527), .B(n3417), .Z(n3526) );
  OR U3721 ( .A(n3528), .B(n3498), .Z(n3417) );
  XNOR U3722 ( .A(n3419), .B(n3496), .Z(n3498) );
  NOR U3723 ( .A(n3529), .B(n3496), .Z(n3527) );
  XOR U3724 ( .A(n3530), .B(n3523), .Z(n3432) );
  OR U3725 ( .A(n3512), .B(n3531), .Z(n3523) );
  XNOR U3726 ( .A(n3532), .B(n3510), .Z(n3512) );
  XOR U3727 ( .A(n3496), .B(n3356), .Z(n3510) );
  IV U3728 ( .A(n3521), .Z(n3356) );
  XOR U3729 ( .A(n3533), .B(n3534), .Z(n3521) );
  NANDN U3730 ( .A(n3535), .B(n3536), .Z(n3534) );
  XNOR U3731 ( .A(n3537), .B(n3538), .Z(n3496) );
  OR U3732 ( .A(n3535), .B(n3539), .Z(n3538) );
  ANDN U3733 ( .B(n3532), .A(n3540), .Z(n3530) );
  IV U3734 ( .A(n3515), .Z(n3532) );
  XOR U3735 ( .A(n3419), .B(n3504), .Z(n3515) );
  XOR U3736 ( .A(n3533), .B(n3541), .Z(n3504) );
  NANDN U3737 ( .A(n3542), .B(n3543), .Z(n3541) );
  NANDN U3738 ( .A(n3544), .B(n3545), .Z(n3533) );
  OR U3739 ( .A(n3547), .B(n3544), .Z(n3537) );
  XOR U3740 ( .A(n3548), .B(n3535), .Z(n3544) );
  XNOR U3741 ( .A(n3549), .B(n3550), .Z(n3535) );
  XOR U3742 ( .A(n3551), .B(n3543), .Z(n3550) );
  XNOR U3743 ( .A(n3552), .B(n3553), .Z(n3549) );
  XNOR U3744 ( .A(n3554), .B(n3555), .Z(n3553) );
  ANDN U3745 ( .B(n3543), .A(n3556), .Z(n3554) );
  IV U3746 ( .A(n3557), .Z(n3543) );
  ANDN U3747 ( .B(n3548), .A(n3556), .Z(n3546) );
  IV U3748 ( .A(n3542), .Z(n3548) );
  XNOR U3749 ( .A(n3551), .B(n3558), .Z(n3542) );
  XNOR U3750 ( .A(n3555), .B(n3559), .Z(n3558) );
  NANDN U3751 ( .A(n3539), .B(n3536), .Z(n3559) );
  NANDN U3752 ( .A(n3547), .B(n3545), .Z(n3555) );
  XNOR U3753 ( .A(n3536), .B(n3557), .Z(n3545) );
  XOR U3754 ( .A(n3560), .B(n3561), .Z(n3557) );
  XOR U3755 ( .A(n3562), .B(n3563), .Z(n3561) );
  XNOR U3756 ( .A(n3497), .B(n3564), .Z(n3563) );
  XNOR U3757 ( .A(n3565), .B(n3566), .Z(n3560) );
  XNOR U3758 ( .A(n3567), .B(n3568), .Z(n3566) );
  ANDN U3759 ( .B(n3569), .A(n3420), .Z(n3567) );
  XNOR U3760 ( .A(n3556), .B(n3539), .Z(n3547) );
  IV U3761 ( .A(n3552), .Z(n3556) );
  XOR U3762 ( .A(n3570), .B(n3571), .Z(n3552) );
  XNOR U3763 ( .A(n3572), .B(n3564), .Z(n3571) );
  XOR U3764 ( .A(n3573), .B(n3574), .Z(n3564) );
  XNOR U3765 ( .A(n3575), .B(n3576), .Z(n3574) );
  NAND U3766 ( .A(n3525), .B(n3509), .Z(n3576) );
  XNOR U3767 ( .A(n3577), .B(n3578), .Z(n3570) );
  ANDN U3768 ( .B(n3579), .A(n3519), .Z(n3577) );
  XOR U3769 ( .A(n3539), .B(n3536), .Z(n3551) );
  XNOR U3770 ( .A(n3580), .B(n3581), .Z(n3536) );
  XNOR U3771 ( .A(n3573), .B(n3582), .Z(n3581) );
  XOR U3772 ( .A(n3572), .B(n3441), .Z(n3582) );
  XOR U3773 ( .A(n3420), .B(n3583), .Z(n3580) );
  XNOR U3774 ( .A(n3584), .B(n3568), .Z(n3583) );
  OR U3775 ( .A(n3499), .B(n3528), .Z(n3568) );
  XNOR U3776 ( .A(n3420), .B(n3529), .Z(n3528) );
  XOR U3777 ( .A(n3441), .B(n3497), .Z(n3499) );
  ANDN U3778 ( .B(n3497), .A(n3529), .Z(n3584) );
  XOR U3779 ( .A(n3585), .B(n3586), .Z(n3539) );
  XOR U3780 ( .A(n3573), .B(n3562), .Z(n3586) );
  XNOR U3781 ( .A(n3436), .B(n3355), .Z(n3562) );
  XOR U3782 ( .A(n3587), .B(n3575), .Z(n3573) );
  NANDN U3783 ( .A(n3531), .B(n3513), .Z(n3575) );
  XOR U3784 ( .A(n3514), .B(n3509), .Z(n3513) );
  XOR U3785 ( .A(n3355), .B(n3497), .Z(n3509) );
  XNOR U3786 ( .A(n3579), .B(n3588), .Z(n3497) );
  XOR U3787 ( .A(n3589), .B(n3590), .Z(n3588) );
  XOR U3788 ( .A(n3540), .B(n3525), .Z(n3531) );
  XNOR U3789 ( .A(n3529), .B(n3436), .Z(n3525) );
  IV U3790 ( .A(n3565), .Z(n3529) );
  XOR U3791 ( .A(n3591), .B(n3592), .Z(n3565) );
  XOR U3792 ( .A(n3593), .B(n3594), .Z(n3592) );
  XNOR U3793 ( .A(n3420), .B(n3595), .Z(n3591) );
  ANDN U3794 ( .B(n3514), .A(n3540), .Z(n3587) );
  XNOR U3795 ( .A(n3420), .B(n3519), .Z(n3540) );
  XOR U3796 ( .A(n3579), .B(n3569), .Z(n3514) );
  IV U3797 ( .A(n3441), .Z(n3569) );
  XOR U3798 ( .A(n3596), .B(n3597), .Z(n3441) );
  XOR U3799 ( .A(n3598), .B(n3594), .Z(n3597) );
  XNOR U3800 ( .A(n3599), .B(n3600), .Z(n3594) );
  XOR U3801 ( .A(n2707), .B(n3601), .Z(n3600) );
  XNOR U3802 ( .A(n3602), .B(n3603), .Z(n2707) );
  XNOR U3803 ( .A(key[396]), .B(n3604), .Z(n3599) );
  XOR U3804 ( .A(n3572), .B(n3605), .Z(n3585) );
  XNOR U3805 ( .A(n3606), .B(n3578), .Z(n3605) );
  OR U3806 ( .A(n3503), .B(n3520), .Z(n3578) );
  XNOR U3807 ( .A(n3607), .B(n3436), .Z(n3520) );
  XNOR U3808 ( .A(n3579), .B(n3355), .Z(n3503) );
  IV U3809 ( .A(n3505), .Z(n3579) );
  AND U3810 ( .A(n3355), .B(n3436), .Z(n3606) );
  XOR U3811 ( .A(n3598), .B(n3596), .Z(n3436) );
  XNOR U3812 ( .A(n3596), .B(n3608), .Z(n3355) );
  XNOR U3813 ( .A(n3609), .B(n3598), .Z(n3608) );
  XNOR U3814 ( .A(n3519), .B(n3505), .Z(n3572) );
  XOR U3815 ( .A(n3596), .B(n3610), .Z(n3505) );
  XNOR U3816 ( .A(n3598), .B(n3593), .Z(n3610) );
  XOR U3817 ( .A(n3611), .B(n3612), .Z(n3593) );
  XOR U3818 ( .A(n3613), .B(n3614), .Z(n3612) );
  XNOR U3819 ( .A(key[399]), .B(n3615), .Z(n3611) );
  XNOR U3820 ( .A(n3616), .B(n3617), .Z(n3596) );
  XNOR U3821 ( .A(n3618), .B(n3619), .Z(n3617) );
  XNOR U3822 ( .A(n3620), .B(n3621), .Z(n3616) );
  XOR U3823 ( .A(key[397]), .B(n3622), .Z(n3621) );
  IV U3824 ( .A(n3607), .Z(n3519) );
  XNOR U3825 ( .A(n3590), .B(n3623), .Z(n3607) );
  XOR U3826 ( .A(n3624), .B(n3625), .Z(n3598) );
  XNOR U3827 ( .A(n3420), .B(n3626), .Z(n3625) );
  XNOR U3828 ( .A(n3627), .B(n3628), .Z(n3420) );
  XNOR U3829 ( .A(n3629), .B(n2726), .Z(n3628) );
  XNOR U3830 ( .A(n3630), .B(n3631), .Z(n3627) );
  XOR U3831 ( .A(key[392]), .B(n3602), .Z(n3631) );
  XNOR U3832 ( .A(n2688), .B(n3632), .Z(n3624) );
  XNOR U3833 ( .A(key[398]), .B(n3633), .Z(n3632) );
  XNOR U3834 ( .A(n3602), .B(n3634), .Z(n2688) );
  XOR U3835 ( .A(n3635), .B(n3636), .Z(n3595) );
  XNOR U3836 ( .A(n3637), .B(n3638), .Z(n3636) );
  XOR U3837 ( .A(n2680), .B(n3609), .Z(n3638) );
  IV U3838 ( .A(n3589), .Z(n3609) );
  XNOR U3839 ( .A(n3639), .B(n3640), .Z(n3589) );
  XOR U3840 ( .A(n3641), .B(n2727), .Z(n3640) );
  XOR U3841 ( .A(n3642), .B(n3643), .Z(n3639) );
  XOR U3842 ( .A(key[393]), .B(n3644), .Z(n3643) );
  XNOR U3843 ( .A(n2713), .B(n3645), .Z(n3635) );
  XNOR U3844 ( .A(key[395]), .B(n3646), .Z(n3645) );
  XOR U3845 ( .A(n2703), .B(n3647), .Z(n2713) );
  IV U3846 ( .A(n3602), .Z(n2703) );
  XOR U3847 ( .A(n3648), .B(n3649), .Z(n3590) );
  XNOR U3848 ( .A(n3650), .B(n2719), .Z(n3649) );
  XOR U3849 ( .A(n3651), .B(n3652), .Z(n3648) );
  XNOR U3850 ( .A(key[394]), .B(n3653), .Z(n3652) );
  XOR U3851 ( .A(n3402), .B(n3377), .Z(n1621) );
  XNOR U3852 ( .A(n3654), .B(n3655), .Z(n3377) );
  XOR U3853 ( .A(n3656), .B(n3657), .Z(n3655) );
  NOR U3854 ( .A(n3658), .B(n3490), .Z(n3656) );
  XOR U3855 ( .A(n3659), .B(n3660), .Z(n1626) );
  XOR U3856 ( .A(n3394), .B(n3399), .Z(n3660) );
  XOR U3857 ( .A(n3373), .B(n3392), .Z(n3399) );
  XNOR U3858 ( .A(n3473), .B(n3661), .Z(n3392) );
  XNOR U3859 ( .A(n3662), .B(n3663), .Z(n3661) );
  NANDN U3860 ( .A(n3664), .B(n3665), .Z(n3663) );
  XOR U3861 ( .A(n3666), .B(n3667), .Z(n3373) );
  XOR U3862 ( .A(n3668), .B(n3669), .Z(n3667) );
  ANDN U3863 ( .B(n3665), .A(n3670), .Z(n3668) );
  XNOR U3864 ( .A(n3422), .B(n3671), .Z(n3394) );
  XNOR U3865 ( .A(n3662), .B(n3672), .Z(n3671) );
  NANDN U3866 ( .A(n3673), .B(n3674), .Z(n3672) );
  OR U3867 ( .A(n3675), .B(n3676), .Z(n3662) );
  XOR U3868 ( .A(n3473), .B(n3677), .Z(n3422) );
  XNOR U3869 ( .A(n3678), .B(n3679), .Z(n3677) );
  NANDN U3870 ( .A(n3680), .B(n3681), .Z(n3679) );
  XOR U3871 ( .A(n3682), .B(n3678), .Z(n3473) );
  NANDN U3872 ( .A(n3683), .B(n3684), .Z(n3678) );
  ANDN U3873 ( .B(n3685), .A(n3686), .Z(n3682) );
  XOR U3874 ( .A(n3666), .B(n3687), .Z(n3372) );
  XOR U3875 ( .A(n3477), .B(n3688), .Z(n3687) );
  NANDN U3876 ( .A(n3689), .B(n3483), .Z(n3688) );
  XOR U3877 ( .A(n3479), .B(n3483), .Z(n3485) );
  XNOR U3878 ( .A(n3474), .B(n3691), .Z(n3480) );
  XNOR U3879 ( .A(n3669), .B(n3692), .Z(n3691) );
  NANDN U3880 ( .A(n3693), .B(n3674), .Z(n3692) );
  OR U3881 ( .A(n3694), .B(n3675), .Z(n3669) );
  XNOR U3882 ( .A(n3674), .B(n3665), .Z(n3675) );
  XNOR U3883 ( .A(n3666), .B(n3695), .Z(n3474) );
  XNOR U3884 ( .A(n3696), .B(n3697), .Z(n3695) );
  NANDN U3885 ( .A(n3680), .B(n3698), .Z(n3697) );
  XOR U3886 ( .A(n3699), .B(n3696), .Z(n3666) );
  OR U3887 ( .A(n3683), .B(n3700), .Z(n3696) );
  XNOR U3888 ( .A(n3686), .B(n3680), .Z(n3683) );
  XNOR U3889 ( .A(n3665), .B(n3483), .Z(n3680) );
  XOR U3890 ( .A(n3701), .B(n3702), .Z(n3483) );
  NANDN U3891 ( .A(n3703), .B(n3704), .Z(n3702) );
  XOR U3892 ( .A(n3705), .B(n3706), .Z(n3665) );
  NANDN U3893 ( .A(n3703), .B(n3707), .Z(n3706) );
  NOR U3894 ( .A(n3686), .B(n3708), .Z(n3699) );
  XNOR U3895 ( .A(n3479), .B(n3674), .Z(n3686) );
  XNOR U3896 ( .A(n3709), .B(n3705), .Z(n3674) );
  NANDN U3897 ( .A(n3710), .B(n3711), .Z(n3705) );
  XOR U3898 ( .A(n3707), .B(n3712), .Z(n3711) );
  ANDN U3899 ( .B(n3712), .A(n3713), .Z(n3709) );
  XNOR U3900 ( .A(n3714), .B(n3701), .Z(n3479) );
  NANDN U3901 ( .A(n3710), .B(n3715), .Z(n3701) );
  XOR U3902 ( .A(n3716), .B(n3704), .Z(n3715) );
  XNOR U3903 ( .A(n3717), .B(n3718), .Z(n3703) );
  XOR U3904 ( .A(n3719), .B(n3720), .Z(n3718) );
  XNOR U3905 ( .A(n3721), .B(n3722), .Z(n3717) );
  XNOR U3906 ( .A(n3723), .B(n3724), .Z(n3722) );
  ANDN U3907 ( .B(n3716), .A(n3720), .Z(n3723) );
  ANDN U3908 ( .B(n3716), .A(n3713), .Z(n3714) );
  XNOR U3909 ( .A(n3719), .B(n3725), .Z(n3713) );
  XOR U3910 ( .A(n3726), .B(n3724), .Z(n3725) );
  NAND U3911 ( .A(n3727), .B(n3728), .Z(n3724) );
  XNOR U3912 ( .A(n3721), .B(n3704), .Z(n3728) );
  IV U3913 ( .A(n3716), .Z(n3721) );
  XNOR U3914 ( .A(n3707), .B(n3720), .Z(n3727) );
  IV U3915 ( .A(n3712), .Z(n3720) );
  XOR U3916 ( .A(n3729), .B(n3730), .Z(n3712) );
  XNOR U3917 ( .A(n3731), .B(n3732), .Z(n3730) );
  XNOR U3918 ( .A(n3733), .B(n3734), .Z(n3729) );
  ANDN U3919 ( .B(n3478), .A(n3735), .Z(n3733) );
  AND U3920 ( .A(n3704), .B(n3707), .Z(n3726) );
  XNOR U3921 ( .A(n3704), .B(n3707), .Z(n3719) );
  XNOR U3922 ( .A(n3736), .B(n3737), .Z(n3707) );
  XNOR U3923 ( .A(n3738), .B(n3732), .Z(n3737) );
  XOR U3924 ( .A(n3739), .B(n3740), .Z(n3736) );
  XNOR U3925 ( .A(n3741), .B(n3734), .Z(n3740) );
  OR U3926 ( .A(n3486), .B(n3690), .Z(n3734) );
  XNOR U3927 ( .A(n3478), .B(n3742), .Z(n3690) );
  XNOR U3928 ( .A(n3735), .B(n3484), .Z(n3486) );
  ANDN U3929 ( .B(n3743), .A(n3689), .Z(n3741) );
  XNOR U3930 ( .A(n3744), .B(n3745), .Z(n3704) );
  XNOR U3931 ( .A(n3732), .B(n3746), .Z(n3745) );
  XOR U3932 ( .A(n3673), .B(n3739), .Z(n3746) );
  XNOR U3933 ( .A(n3478), .B(n3735), .Z(n3732) );
  XOR U3934 ( .A(n3693), .B(n3747), .Z(n3744) );
  XNOR U3935 ( .A(n3748), .B(n3749), .Z(n3747) );
  ANDN U3936 ( .B(n3750), .A(n3670), .Z(n3748) );
  XNOR U3937 ( .A(n3751), .B(n3752), .Z(n3716) );
  XNOR U3938 ( .A(n3738), .B(n3753), .Z(n3752) );
  XNOR U3939 ( .A(n3664), .B(n3731), .Z(n3753) );
  XOR U3940 ( .A(n3739), .B(n3754), .Z(n3731) );
  XNOR U3941 ( .A(n3755), .B(n3756), .Z(n3754) );
  NAND U3942 ( .A(n3698), .B(n3681), .Z(n3756) );
  XNOR U3943 ( .A(n3757), .B(n3755), .Z(n3739) );
  NANDN U3944 ( .A(n3700), .B(n3684), .Z(n3755) );
  XOR U3945 ( .A(n3685), .B(n3681), .Z(n3684) );
  XNOR U3946 ( .A(n3750), .B(n3484), .Z(n3681) );
  XOR U3947 ( .A(n3708), .B(n3698), .Z(n3700) );
  XNOR U3948 ( .A(n3670), .B(n3742), .Z(n3698) );
  ANDN U3949 ( .B(n3685), .A(n3708), .Z(n3757) );
  XOR U3950 ( .A(n3693), .B(n3478), .Z(n3708) );
  XNOR U3951 ( .A(n3758), .B(n3759), .Z(n3478) );
  XNOR U3952 ( .A(n3760), .B(n3761), .Z(n3759) );
  XOR U3953 ( .A(n3742), .B(n3743), .Z(n3738) );
  IV U3954 ( .A(n3484), .Z(n3743) );
  XOR U3955 ( .A(n3762), .B(n3763), .Z(n3484) );
  XOR U3956 ( .A(n3764), .B(n3761), .Z(n3763) );
  IV U3957 ( .A(n3689), .Z(n3742) );
  XOR U3958 ( .A(n3761), .B(n3765), .Z(n3689) );
  XNOR U3959 ( .A(n3766), .B(n3767), .Z(n3751) );
  XNOR U3960 ( .A(n3768), .B(n3749), .Z(n3767) );
  OR U3961 ( .A(n3676), .B(n3694), .Z(n3749) );
  XNOR U3962 ( .A(n3693), .B(n3670), .Z(n3694) );
  IV U3963 ( .A(n3766), .Z(n3670) );
  XOR U3964 ( .A(n3673), .B(n3750), .Z(n3676) );
  IV U3965 ( .A(n3664), .Z(n3750) );
  XOR U3966 ( .A(n3426), .B(n3769), .Z(n3664) );
  XNOR U3967 ( .A(n3770), .B(n3758), .Z(n3769) );
  XOR U3968 ( .A(n3771), .B(n3772), .Z(n3758) );
  XOR U3969 ( .A(n3773), .B(n2578), .Z(n3772) );
  XOR U3970 ( .A(key[434]), .B(n2563), .Z(n3771) );
  IV U3971 ( .A(n3735), .Z(n3426) );
  XOR U3972 ( .A(n3762), .B(n3774), .Z(n3735) );
  XOR U3973 ( .A(n3761), .B(n3775), .Z(n3774) );
  NOR U3974 ( .A(n3673), .B(n3693), .Z(n3768) );
  XOR U3975 ( .A(n3762), .B(n3776), .Z(n3673) );
  XOR U3976 ( .A(n3761), .B(n3777), .Z(n3776) );
  XOR U3977 ( .A(n3778), .B(n3779), .Z(n3761) );
  XOR U3978 ( .A(n3693), .B(n3780), .Z(n3779) );
  XNOR U3979 ( .A(n2566), .B(n3781), .Z(n3778) );
  XNOR U3980 ( .A(key[438]), .B(n2550), .Z(n3781) );
  XOR U3981 ( .A(n3782), .B(n3783), .Z(n2566) );
  IV U3982 ( .A(n3765), .Z(n3762) );
  XOR U3983 ( .A(n3784), .B(n3785), .Z(n3765) );
  XNOR U3984 ( .A(n3786), .B(n2547), .Z(n3785) );
  XOR U3985 ( .A(n3787), .B(n3788), .Z(n2547) );
  XNOR U3986 ( .A(key[437]), .B(n3789), .Z(n3784) );
  XOR U3987 ( .A(n3790), .B(n3791), .Z(n3766) );
  XNOR U3988 ( .A(n3777), .B(n3775), .Z(n3791) );
  XNOR U3989 ( .A(n3792), .B(n3793), .Z(n3775) );
  XOR U3990 ( .A(n2553), .B(n3783), .Z(n3793) );
  XNOR U3991 ( .A(n3794), .B(n3795), .Z(n3783) );
  XOR U3992 ( .A(n3796), .B(n3797), .Z(n2553) );
  XNOR U3993 ( .A(key[439]), .B(n3798), .Z(n3792) );
  XNOR U3994 ( .A(n3799), .B(n3800), .Z(n3777) );
  XNOR U3995 ( .A(n2537), .B(n3801), .Z(n3800) );
  XNOR U3996 ( .A(n3802), .B(n3803), .Z(n2537) );
  XNOR U3997 ( .A(n2536), .B(n3804), .Z(n3799) );
  XOR U3998 ( .A(key[436]), .B(n3805), .Z(n3804) );
  XNOR U3999 ( .A(n3806), .B(n3786), .Z(n2536) );
  XNOR U4000 ( .A(n3693), .B(n3760), .Z(n3790) );
  XOR U4001 ( .A(n3807), .B(n3808), .Z(n3760) );
  XNOR U4002 ( .A(n3809), .B(n3810), .Z(n3808) );
  XOR U4003 ( .A(n2572), .B(n3770), .Z(n3810) );
  IV U4004 ( .A(n3764), .Z(n3770) );
  XNOR U4005 ( .A(n3811), .B(n3812), .Z(n3764) );
  XOR U4006 ( .A(n2588), .B(n3813), .Z(n3812) );
  XOR U4007 ( .A(key[433]), .B(n3814), .Z(n3811) );
  XNOR U4008 ( .A(n3794), .B(n3805), .Z(n2572) );
  XOR U4009 ( .A(n3815), .B(n3816), .Z(n3807) );
  XNOR U4010 ( .A(key[435]), .B(n2561), .Z(n3816) );
  XNOR U4011 ( .A(n3817), .B(n3818), .Z(n3693) );
  XNOR U4012 ( .A(n3819), .B(n2554), .Z(n3818) );
  XOR U4013 ( .A(key[432]), .B(n3820), .Z(n3817) );
  XOR U4014 ( .A(n199), .B(n1624), .Z(n3247) );
  XNOR U4015 ( .A(n3821), .B(n3822), .Z(n1624) );
  XOR U4016 ( .A(n3383), .B(n3397), .Z(n3822) );
  IV U4017 ( .A(n3406), .Z(n3397) );
  XOR U4018 ( .A(n3364), .B(n3381), .Z(n3406) );
  XNOR U4019 ( .A(n3449), .B(n3823), .Z(n3381) );
  XNOR U4020 ( .A(n3824), .B(n3825), .Z(n3823) );
  NANDN U4021 ( .A(n3826), .B(n3827), .Z(n3825) );
  XNOR U4022 ( .A(n3828), .B(n3829), .Z(n3364) );
  XOR U4023 ( .A(n3830), .B(n3831), .Z(n3829) );
  ANDN U4024 ( .B(n3827), .A(n3832), .Z(n3830) );
  XNOR U4025 ( .A(n3407), .B(n3833), .Z(n3383) );
  XNOR U4026 ( .A(n3824), .B(n3834), .Z(n3833) );
  NANDN U4027 ( .A(n3835), .B(n3836), .Z(n3834) );
  OR U4028 ( .A(n3837), .B(n3838), .Z(n3824) );
  XOR U4029 ( .A(n3449), .B(n3839), .Z(n3407) );
  XNOR U4030 ( .A(n3840), .B(n3841), .Z(n3839) );
  NANDN U4031 ( .A(n3842), .B(n3843), .Z(n3841) );
  XOR U4032 ( .A(n3844), .B(n3840), .Z(n3449) );
  NANDN U4033 ( .A(n3845), .B(n3846), .Z(n3840) );
  ANDN U4034 ( .B(n3847), .A(n3848), .Z(n3844) );
  XNOR U4035 ( .A(n3448), .B(n3365), .Z(n3821) );
  XOR U4036 ( .A(n3828), .B(n3849), .Z(n3365) );
  XOR U4037 ( .A(n3459), .B(n3850), .Z(n3849) );
  NANDN U4038 ( .A(n3851), .B(n3452), .Z(n3850) );
  XOR U4039 ( .A(n3461), .B(n3452), .Z(n3454) );
  XNOR U4040 ( .A(n3456), .B(n3853), .Z(n3448) );
  XNOR U4041 ( .A(n3831), .B(n3854), .Z(n3853) );
  NANDN U4042 ( .A(n3855), .B(n3836), .Z(n3854) );
  OR U4043 ( .A(n3856), .B(n3837), .Z(n3831) );
  XNOR U4044 ( .A(n3836), .B(n3827), .Z(n3837) );
  XNOR U4045 ( .A(n3828), .B(n3857), .Z(n3456) );
  XNOR U4046 ( .A(n3858), .B(n3859), .Z(n3857) );
  NANDN U4047 ( .A(n3842), .B(n3860), .Z(n3859) );
  XOR U4048 ( .A(n3861), .B(n3858), .Z(n3828) );
  OR U4049 ( .A(n3845), .B(n3862), .Z(n3858) );
  XNOR U4050 ( .A(n3848), .B(n3842), .Z(n3845) );
  XNOR U4051 ( .A(n3827), .B(n3452), .Z(n3842) );
  XOR U4052 ( .A(n3863), .B(n3864), .Z(n3452) );
  NANDN U4053 ( .A(n3865), .B(n3866), .Z(n3864) );
  XOR U4054 ( .A(n3867), .B(n3868), .Z(n3827) );
  NANDN U4055 ( .A(n3865), .B(n3869), .Z(n3868) );
  NOR U4056 ( .A(n3848), .B(n3870), .Z(n3861) );
  XNOR U4057 ( .A(n3461), .B(n3836), .Z(n3848) );
  XNOR U4058 ( .A(n3871), .B(n3867), .Z(n3836) );
  NANDN U4059 ( .A(n3872), .B(n3873), .Z(n3867) );
  XOR U4060 ( .A(n3869), .B(n3874), .Z(n3873) );
  ANDN U4061 ( .B(n3874), .A(n3875), .Z(n3871) );
  XNOR U4062 ( .A(n3876), .B(n3863), .Z(n3461) );
  NANDN U4063 ( .A(n3872), .B(n3877), .Z(n3863) );
  XOR U4064 ( .A(n3878), .B(n3866), .Z(n3877) );
  XNOR U4065 ( .A(n3879), .B(n3880), .Z(n3865) );
  XOR U4066 ( .A(n3881), .B(n3882), .Z(n3880) );
  XNOR U4067 ( .A(n3883), .B(n3884), .Z(n3879) );
  XNOR U4068 ( .A(n3885), .B(n3886), .Z(n3884) );
  ANDN U4069 ( .B(n3878), .A(n3882), .Z(n3885) );
  ANDN U4070 ( .B(n3878), .A(n3875), .Z(n3876) );
  XNOR U4071 ( .A(n3881), .B(n3887), .Z(n3875) );
  XOR U4072 ( .A(n3888), .B(n3886), .Z(n3887) );
  NAND U4073 ( .A(n3889), .B(n3890), .Z(n3886) );
  XNOR U4074 ( .A(n3883), .B(n3866), .Z(n3890) );
  IV U4075 ( .A(n3878), .Z(n3883) );
  XNOR U4076 ( .A(n3869), .B(n3882), .Z(n3889) );
  IV U4077 ( .A(n3874), .Z(n3882) );
  XOR U4078 ( .A(n3891), .B(n3892), .Z(n3874) );
  XNOR U4079 ( .A(n3893), .B(n3894), .Z(n3892) );
  XNOR U4080 ( .A(n3895), .B(n3896), .Z(n3891) );
  ANDN U4081 ( .B(n3460), .A(n3897), .Z(n3895) );
  AND U4082 ( .A(n3866), .B(n3869), .Z(n3888) );
  XNOR U4083 ( .A(n3866), .B(n3869), .Z(n3881) );
  XNOR U4084 ( .A(n3898), .B(n3899), .Z(n3869) );
  XNOR U4085 ( .A(n3900), .B(n3894), .Z(n3899) );
  XOR U4086 ( .A(n3901), .B(n3902), .Z(n3898) );
  XNOR U4087 ( .A(n3903), .B(n3896), .Z(n3902) );
  OR U4088 ( .A(n3455), .B(n3852), .Z(n3896) );
  XNOR U4089 ( .A(n3460), .B(n3904), .Z(n3852) );
  XNOR U4090 ( .A(n3897), .B(n3453), .Z(n3455) );
  ANDN U4091 ( .B(n3905), .A(n3851), .Z(n3903) );
  XNOR U4092 ( .A(n3906), .B(n3907), .Z(n3866) );
  XNOR U4093 ( .A(n3894), .B(n3908), .Z(n3907) );
  XOR U4094 ( .A(n3835), .B(n3901), .Z(n3908) );
  XNOR U4095 ( .A(n3460), .B(n3897), .Z(n3894) );
  XOR U4096 ( .A(n3855), .B(n3909), .Z(n3906) );
  XNOR U4097 ( .A(n3910), .B(n3911), .Z(n3909) );
  ANDN U4098 ( .B(n3912), .A(n3832), .Z(n3910) );
  XNOR U4099 ( .A(n3913), .B(n3914), .Z(n3878) );
  XNOR U4100 ( .A(n3900), .B(n3915), .Z(n3914) );
  XNOR U4101 ( .A(n3826), .B(n3893), .Z(n3915) );
  XOR U4102 ( .A(n3901), .B(n3916), .Z(n3893) );
  XNOR U4103 ( .A(n3917), .B(n3918), .Z(n3916) );
  NAND U4104 ( .A(n3860), .B(n3843), .Z(n3918) );
  XNOR U4105 ( .A(n3919), .B(n3917), .Z(n3901) );
  NANDN U4106 ( .A(n3862), .B(n3846), .Z(n3917) );
  XOR U4107 ( .A(n3847), .B(n3843), .Z(n3846) );
  XNOR U4108 ( .A(n3912), .B(n3453), .Z(n3843) );
  XOR U4109 ( .A(n3870), .B(n3860), .Z(n3862) );
  XNOR U4110 ( .A(n3832), .B(n3904), .Z(n3860) );
  ANDN U4111 ( .B(n3847), .A(n3870), .Z(n3919) );
  XOR U4112 ( .A(n3855), .B(n3460), .Z(n3870) );
  XNOR U4113 ( .A(n3920), .B(n3921), .Z(n3460) );
  XNOR U4114 ( .A(n3922), .B(n3923), .Z(n3921) );
  XOR U4115 ( .A(n3904), .B(n3905), .Z(n3900) );
  IV U4116 ( .A(n3453), .Z(n3905) );
  XOR U4117 ( .A(n3924), .B(n3925), .Z(n3453) );
  XOR U4118 ( .A(n3926), .B(n3923), .Z(n3925) );
  IV U4119 ( .A(n3851), .Z(n3904) );
  XOR U4120 ( .A(n3923), .B(n3927), .Z(n3851) );
  XNOR U4121 ( .A(n3928), .B(n3929), .Z(n3913) );
  XNOR U4122 ( .A(n3930), .B(n3911), .Z(n3929) );
  OR U4123 ( .A(n3838), .B(n3856), .Z(n3911) );
  XNOR U4124 ( .A(n3855), .B(n3832), .Z(n3856) );
  IV U4125 ( .A(n3928), .Z(n3832) );
  XOR U4126 ( .A(n3835), .B(n3912), .Z(n3838) );
  IV U4127 ( .A(n3826), .Z(n3912) );
  XOR U4128 ( .A(n3411), .B(n3931), .Z(n3826) );
  XNOR U4129 ( .A(n3932), .B(n3920), .Z(n3931) );
  XOR U4130 ( .A(n3933), .B(n3934), .Z(n3920) );
  XOR U4131 ( .A(n3935), .B(n3019), .Z(n3934) );
  XOR U4132 ( .A(n3936), .B(n3937), .Z(n3933) );
  XNOR U4133 ( .A(key[474]), .B(n3938), .Z(n3937) );
  IV U4134 ( .A(n3897), .Z(n3411) );
  XOR U4135 ( .A(n3924), .B(n3939), .Z(n3897) );
  XOR U4136 ( .A(n3923), .B(n3940), .Z(n3939) );
  NOR U4137 ( .A(n3835), .B(n3855), .Z(n3930) );
  XOR U4138 ( .A(n3924), .B(n3941), .Z(n3835) );
  XOR U4139 ( .A(n3923), .B(n3942), .Z(n3941) );
  XOR U4140 ( .A(n3943), .B(n3944), .Z(n3923) );
  XNOR U4141 ( .A(n3855), .B(n3945), .Z(n3944) );
  XNOR U4142 ( .A(n3034), .B(n3946), .Z(n3943) );
  XNOR U4143 ( .A(key[478]), .B(n3947), .Z(n3946) );
  XNOR U4144 ( .A(n3948), .B(n3949), .Z(n3034) );
  IV U4145 ( .A(n3927), .Z(n3924) );
  XOR U4146 ( .A(n3950), .B(n3951), .Z(n3927) );
  XNOR U4147 ( .A(n3952), .B(n3953), .Z(n3951) );
  XNOR U4148 ( .A(n3954), .B(n3955), .Z(n3950) );
  XNOR U4149 ( .A(key[477]), .B(n3956), .Z(n3955) );
  XOR U4150 ( .A(n3957), .B(n3958), .Z(n3928) );
  XNOR U4151 ( .A(n3942), .B(n3940), .Z(n3958) );
  XNOR U4152 ( .A(n3959), .B(n3960), .Z(n3940) );
  XNOR U4153 ( .A(n3961), .B(n3962), .Z(n3960) );
  XNOR U4154 ( .A(key[479]), .B(n3963), .Z(n3959) );
  XNOR U4155 ( .A(n3964), .B(n3965), .Z(n3942) );
  XNOR U4156 ( .A(n3011), .B(n3966), .Z(n3964) );
  XNOR U4157 ( .A(key[476]), .B(n3967), .Z(n3966) );
  XNOR U4158 ( .A(n3948), .B(n3968), .Z(n3011) );
  XNOR U4159 ( .A(n3855), .B(n3922), .Z(n3957) );
  XOR U4160 ( .A(n3969), .B(n3970), .Z(n3922) );
  XNOR U4161 ( .A(n3971), .B(n3972), .Z(n3970) );
  XNOR U4162 ( .A(n3000), .B(n3932), .Z(n3972) );
  IV U4163 ( .A(n3926), .Z(n3932) );
  XNOR U4164 ( .A(n3973), .B(n3974), .Z(n3926) );
  XNOR U4165 ( .A(n3975), .B(n3038), .Z(n3974) );
  XOR U4166 ( .A(n3976), .B(n3977), .Z(n3973) );
  XNOR U4167 ( .A(key[473]), .B(n3978), .Z(n3977) );
  XNOR U4168 ( .A(n3031), .B(n3979), .Z(n3000) );
  XNOR U4169 ( .A(n3046), .B(n3980), .Z(n3969) );
  XNOR U4170 ( .A(key[475]), .B(n3981), .Z(n3980) );
  IV U4171 ( .A(n3982), .Z(n3046) );
  XNOR U4172 ( .A(n3983), .B(n3984), .Z(n3855) );
  XNOR U4173 ( .A(n3985), .B(n3037), .Z(n3984) );
  XNOR U4174 ( .A(n3986), .B(n3987), .Z(n3983) );
  XOR U4175 ( .A(key[472]), .B(n3948), .Z(n3987) );
  XOR U4176 ( .A(n3988), .B(n3989), .Z(n199) );
  XNOR U4177 ( .A(n3389), .B(n3387), .Z(n3989) );
  XOR U4178 ( .A(n3990), .B(n3991), .Z(n3387) );
  XNOR U4179 ( .A(n3657), .B(n3992), .Z(n3991) );
  NAND U4180 ( .A(n3993), .B(n3469), .Z(n3992) );
  NANDN U4181 ( .A(n3994), .B(n3493), .Z(n3657) );
  XNOR U4182 ( .A(n3490), .B(n3469), .Z(n3493) );
  XOR U4183 ( .A(n3487), .B(n3995), .Z(n3389) );
  XNOR U4184 ( .A(n3996), .B(n3997), .Z(n3995) );
  OR U4185 ( .A(n3998), .B(n3999), .Z(n3997) );
  XNOR U4186 ( .A(n3465), .B(n4000), .Z(n3487) );
  XNOR U4187 ( .A(n4001), .B(n4002), .Z(n4000) );
  NANDN U4188 ( .A(n4003), .B(n4004), .Z(n4002) );
  XOR U4189 ( .A(n3443), .B(n3464), .Z(n3988) );
  XNOR U4190 ( .A(n3654), .B(n4005), .Z(n3464) );
  XNOR U4191 ( .A(n4006), .B(n4007), .Z(n4005) );
  OR U4192 ( .A(n3998), .B(n4008), .Z(n4007) );
  XNOR U4193 ( .A(n3990), .B(n4009), .Z(n3654) );
  XNOR U4194 ( .A(n4010), .B(n4011), .Z(n4009) );
  NANDN U4195 ( .A(n4003), .B(n4012), .Z(n4011) );
  XOR U4196 ( .A(n3402), .B(n3388), .Z(n3443) );
  XOR U4197 ( .A(n3465), .B(n4013), .Z(n3388) );
  XOR U4198 ( .A(n4014), .B(n3996), .Z(n4013) );
  OR U4199 ( .A(n4015), .B(n4016), .Z(n3996) );
  AND U4200 ( .A(n4017), .B(n4018), .Z(n4014) );
  XOR U4201 ( .A(n4019), .B(n4001), .Z(n3465) );
  NANDN U4202 ( .A(n4020), .B(n4021), .Z(n4001) );
  AND U4203 ( .A(n4022), .B(n4023), .Z(n4019) );
  XNOR U4204 ( .A(n3990), .B(n4024), .Z(n3402) );
  XOR U4205 ( .A(n4025), .B(n4006), .Z(n4024) );
  OR U4206 ( .A(n4026), .B(n4015), .Z(n4006) );
  XOR U4207 ( .A(n3998), .B(n4018), .Z(n4015) );
  ANDN U4208 ( .B(n4018), .A(n4027), .Z(n4025) );
  XOR U4209 ( .A(n4028), .B(n4010), .Z(n3990) );
  OR U4210 ( .A(n4020), .B(n4029), .Z(n4010) );
  XOR U4211 ( .A(n4022), .B(n4003), .Z(n4020) );
  XNOR U4212 ( .A(n4018), .B(n3469), .Z(n4003) );
  XOR U4213 ( .A(n4030), .B(n4031), .Z(n3469) );
  NANDN U4214 ( .A(n4032), .B(n4033), .Z(n4031) );
  XOR U4215 ( .A(n4034), .B(n4035), .Z(n4018) );
  OR U4216 ( .A(n4032), .B(n4036), .Z(n4035) );
  ANDN U4217 ( .B(n4022), .A(n4037), .Z(n4028) );
  XOR U4218 ( .A(n3998), .B(n3490), .Z(n4022) );
  XOR U4219 ( .A(n4038), .B(n4030), .Z(n3490) );
  NANDN U4220 ( .A(n4039), .B(n4040), .Z(n4030) );
  ANDN U4221 ( .B(n4041), .A(n4042), .Z(n4038) );
  NANDN U4222 ( .A(n4039), .B(n4044), .Z(n4034) );
  XOR U4223 ( .A(n4045), .B(n4032), .Z(n4039) );
  XNOR U4224 ( .A(n4046), .B(n4047), .Z(n4032) );
  XOR U4225 ( .A(n4048), .B(n4041), .Z(n4047) );
  XNOR U4226 ( .A(n4049), .B(n4050), .Z(n4046) );
  XNOR U4227 ( .A(n4051), .B(n4052), .Z(n4050) );
  ANDN U4228 ( .B(n4041), .A(n4053), .Z(n4051) );
  IV U4229 ( .A(n4054), .Z(n4041) );
  ANDN U4230 ( .B(n4045), .A(n4053), .Z(n4043) );
  IV U4231 ( .A(n4049), .Z(n4053) );
  IV U4232 ( .A(n4042), .Z(n4045) );
  XNOR U4233 ( .A(n4048), .B(n4055), .Z(n4042) );
  XOR U4234 ( .A(n4056), .B(n4052), .Z(n4055) );
  NAND U4235 ( .A(n4044), .B(n4040), .Z(n4052) );
  XNOR U4236 ( .A(n4033), .B(n4054), .Z(n4040) );
  XOR U4237 ( .A(n4057), .B(n4058), .Z(n4054) );
  XOR U4238 ( .A(n4059), .B(n4060), .Z(n4058) );
  XNOR U4239 ( .A(n4017), .B(n4061), .Z(n4060) );
  XNOR U4240 ( .A(n4062), .B(n4063), .Z(n4057) );
  XNOR U4241 ( .A(n4064), .B(n4065), .Z(n4063) );
  ANDN U4242 ( .B(n4066), .A(n4008), .Z(n4064) );
  XNOR U4243 ( .A(n4049), .B(n4036), .Z(n4044) );
  XOR U4244 ( .A(n4067), .B(n4068), .Z(n4049) );
  XNOR U4245 ( .A(n4069), .B(n4061), .Z(n4068) );
  XOR U4246 ( .A(n4070), .B(n4071), .Z(n4061) );
  XNOR U4247 ( .A(n4072), .B(n4073), .Z(n4071) );
  NAND U4248 ( .A(n4012), .B(n4004), .Z(n4073) );
  XNOR U4249 ( .A(n4074), .B(n4075), .Z(n4067) );
  ANDN U4250 ( .B(n4076), .A(n3658), .Z(n4074) );
  ANDN U4251 ( .B(n4033), .A(n4036), .Z(n4056) );
  XOR U4252 ( .A(n4036), .B(n4033), .Z(n4048) );
  XNOR U4253 ( .A(n4077), .B(n4078), .Z(n4033) );
  XNOR U4254 ( .A(n4070), .B(n4079), .Z(n4078) );
  XOR U4255 ( .A(n4069), .B(n3999), .Z(n4079) );
  XOR U4256 ( .A(n4008), .B(n4080), .Z(n4077) );
  XNOR U4257 ( .A(n4081), .B(n4065), .Z(n4080) );
  OR U4258 ( .A(n4016), .B(n4026), .Z(n4065) );
  XNOR U4259 ( .A(n4008), .B(n4027), .Z(n4026) );
  XOR U4260 ( .A(n3999), .B(n4017), .Z(n4016) );
  ANDN U4261 ( .B(n4017), .A(n4027), .Z(n4081) );
  XOR U4262 ( .A(n4082), .B(n4083), .Z(n4036) );
  XOR U4263 ( .A(n4070), .B(n4059), .Z(n4083) );
  XOR U4264 ( .A(n3993), .B(n3470), .Z(n4059) );
  XOR U4265 ( .A(n4084), .B(n4072), .Z(n4070) );
  NANDN U4266 ( .A(n4029), .B(n4021), .Z(n4072) );
  XOR U4267 ( .A(n4023), .B(n4004), .Z(n4021) );
  XNOR U4268 ( .A(n4076), .B(n4085), .Z(n4017) );
  XOR U4269 ( .A(n4086), .B(n4087), .Z(n4085) );
  XOR U4270 ( .A(n4037), .B(n4012), .Z(n4029) );
  XNOR U4271 ( .A(n4027), .B(n3993), .Z(n4012) );
  IV U4272 ( .A(n4062), .Z(n4027) );
  XOR U4273 ( .A(n4088), .B(n4089), .Z(n4062) );
  XOR U4274 ( .A(n4090), .B(n4091), .Z(n4089) );
  XNOR U4275 ( .A(n4008), .B(n4092), .Z(n4088) );
  ANDN U4276 ( .B(n4023), .A(n4037), .Z(n4084) );
  XNOR U4277 ( .A(n4008), .B(n3658), .Z(n4037) );
  XOR U4278 ( .A(n4076), .B(n4066), .Z(n4023) );
  IV U4279 ( .A(n3999), .Z(n4066) );
  XOR U4280 ( .A(n4093), .B(n4094), .Z(n3999) );
  XOR U4281 ( .A(n4095), .B(n4091), .Z(n4094) );
  XNOR U4282 ( .A(n4096), .B(n4097), .Z(n4091) );
  XNOR U4283 ( .A(n2872), .B(n4098), .Z(n4097) );
  XNOR U4284 ( .A(n4099), .B(n4100), .Z(n2872) );
  XNOR U4285 ( .A(n2871), .B(n4101), .Z(n4096) );
  XOR U4286 ( .A(key[484]), .B(n4102), .Z(n4101) );
  XOR U4287 ( .A(n4103), .B(n4104), .Z(n2871) );
  IV U4288 ( .A(n3491), .Z(n4076) );
  XOR U4289 ( .A(n4069), .B(n4105), .Z(n4082) );
  XNOR U4290 ( .A(n4106), .B(n4075), .Z(n4105) );
  OR U4291 ( .A(n3492), .B(n3994), .Z(n4075) );
  XNOR U4292 ( .A(n4107), .B(n3993), .Z(n3994) );
  XNOR U4293 ( .A(n3491), .B(n3470), .Z(n3492) );
  ANDN U4294 ( .B(n3993), .A(n3470), .Z(n4106) );
  XOR U4295 ( .A(n4093), .B(n4108), .Z(n3470) );
  XNOR U4296 ( .A(n4109), .B(n4095), .Z(n4108) );
  XOR U4297 ( .A(n4095), .B(n4093), .Z(n3993) );
  XNOR U4298 ( .A(n3658), .B(n3491), .Z(n4069) );
  XOR U4299 ( .A(n4093), .B(n4110), .Z(n3491) );
  XNOR U4300 ( .A(n4095), .B(n4090), .Z(n4110) );
  XOR U4301 ( .A(n4111), .B(n4112), .Z(n4090) );
  XOR U4302 ( .A(n4113), .B(n2866), .Z(n4112) );
  XNOR U4303 ( .A(n4114), .B(n4115), .Z(n2866) );
  XNOR U4304 ( .A(key[487]), .B(n4116), .Z(n4111) );
  XNOR U4305 ( .A(n4117), .B(n4118), .Z(n4093) );
  XNOR U4306 ( .A(n4104), .B(n2858), .Z(n4118) );
  XOR U4307 ( .A(n4119), .B(n4120), .Z(n2858) );
  XNOR U4308 ( .A(key[485]), .B(n4121), .Z(n4117) );
  IV U4309 ( .A(n4107), .Z(n3658) );
  XNOR U4310 ( .A(n4086), .B(n4092), .Z(n4122) );
  XOR U4311 ( .A(n4123), .B(n4124), .Z(n4092) );
  XNOR U4312 ( .A(n4125), .B(n4126), .Z(n4124) );
  XOR U4313 ( .A(n2878), .B(n4087), .Z(n4126) );
  IV U4314 ( .A(n4109), .Z(n4087) );
  XOR U4315 ( .A(n4127), .B(n4128), .Z(n4109) );
  XOR U4316 ( .A(n2893), .B(n4129), .Z(n4128) );
  XNOR U4317 ( .A(key[481]), .B(n2887), .Z(n4127) );
  XNOR U4318 ( .A(n4130), .B(n4102), .Z(n2878) );
  XOR U4319 ( .A(n4131), .B(n4132), .Z(n4123) );
  XNOR U4320 ( .A(key[483]), .B(n2842), .Z(n4132) );
  XOR U4321 ( .A(n4133), .B(n4134), .Z(n4086) );
  XOR U4322 ( .A(n4135), .B(n2884), .Z(n4134) );
  XOR U4323 ( .A(key[482]), .B(n2844), .Z(n4133) );
  XOR U4324 ( .A(n4136), .B(n4137), .Z(n4095) );
  XNOR U4325 ( .A(n4008), .B(n4138), .Z(n4137) );
  XNOR U4326 ( .A(n4139), .B(n4140), .Z(n4008) );
  XNOR U4327 ( .A(n4141), .B(n2867), .Z(n4140) );
  XNOR U4328 ( .A(key[480]), .B(n4142), .Z(n4139) );
  XOR U4329 ( .A(n2851), .B(n4143), .Z(n4136) );
  XNOR U4330 ( .A(key[486]), .B(n2861), .Z(n4143) );
  XNOR U4331 ( .A(n4144), .B(n4113), .Z(n2851) );
  XNOR U4332 ( .A(n4130), .B(n4145), .Z(n4113) );
  XOR U4333 ( .A(n4146), .B(n4147), .Z(out[109]) );
  XNOR U4334 ( .A(n4148), .B(n4149), .Z(n4147) );
  XOR U4335 ( .A(n3264), .B(n4150), .Z(n4149) );
  XNOR U4336 ( .A(n4152), .B(n4153), .Z(n4151) );
  NANDN U4337 ( .A(n4154), .B(n4155), .Z(n4153) );
  XOR U4338 ( .A(n4157), .B(n4158), .Z(n4146) );
  XOR U4339 ( .A(key[621]), .B(n4159), .Z(n4158) );
  ANDN U4340 ( .B(n4160), .A(n4161), .Z(n4157) );
  XNOR U4341 ( .A(n4162), .B(n4163), .Z(out[108]) );
  XNOR U4342 ( .A(key[620]), .B(n4164), .Z(n4163) );
  XOR U4343 ( .A(n4165), .B(n4166), .Z(out[107]) );
  XNOR U4344 ( .A(n4167), .B(n3267), .Z(n4166) );
  XNOR U4345 ( .A(n4168), .B(n4169), .Z(n3267) );
  XNOR U4346 ( .A(n4170), .B(n4159), .Z(n4169) );
  ANDN U4347 ( .B(n4171), .A(n4172), .Z(n4159) );
  NOR U4348 ( .A(n4173), .B(n4174), .Z(n4170) );
  XNOR U4349 ( .A(n4175), .B(n4176), .Z(n4165) );
  XOR U4350 ( .A(key[619]), .B(n3266), .Z(n4176) );
  XOR U4351 ( .A(key[618]), .B(n4162), .Z(out[106]) );
  XNOR U4352 ( .A(n4177), .B(n4178), .Z(n4162) );
  XOR U4353 ( .A(n4179), .B(n3263), .Z(out[105]) );
  XNOR U4354 ( .A(n4168), .B(n4180), .Z(n4167) );
  XNOR U4355 ( .A(n4181), .B(n4182), .Z(n4180) );
  NANDN U4356 ( .A(n4183), .B(n4155), .Z(n4182) );
  XNOR U4357 ( .A(n4150), .B(n4184), .Z(n4168) );
  XNOR U4358 ( .A(n4185), .B(n4186), .Z(n4184) );
  NANDN U4359 ( .A(n4187), .B(n4188), .Z(n4186) );
  XOR U4360 ( .A(n4178), .B(n4175), .Z(n3269) );
  XNOR U4361 ( .A(n4150), .B(n4189), .Z(n4175) );
  XNOR U4362 ( .A(n4181), .B(n4190), .Z(n4189) );
  NANDN U4363 ( .A(n4191), .B(n4192), .Z(n4190) );
  OR U4364 ( .A(n4193), .B(n4194), .Z(n4181) );
  XOR U4365 ( .A(n4195), .B(n4185), .Z(n4150) );
  NANDN U4366 ( .A(n4196), .B(n4197), .Z(n4185) );
  ANDN U4367 ( .B(n4198), .A(n4199), .Z(n4195) );
  XNOR U4368 ( .A(key[617]), .B(n4177), .Z(n4179) );
  IV U4369 ( .A(n3266), .Z(n4177) );
  XOR U4370 ( .A(n4200), .B(n4201), .Z(n3266) );
  XNOR U4371 ( .A(n4202), .B(n4203), .Z(n4201) );
  NANDN U4372 ( .A(n4204), .B(n4160), .Z(n4203) );
  XNOR U4373 ( .A(n4148), .B(n4205), .Z(out[104]) );
  XOR U4374 ( .A(key[616]), .B(n4178), .Z(n4205) );
  XNOR U4375 ( .A(n4200), .B(n4206), .Z(n4178) );
  XOR U4376 ( .A(n4207), .B(n4152), .Z(n4206) );
  OR U4377 ( .A(n4208), .B(n4193), .Z(n4152) );
  XNOR U4378 ( .A(n4155), .B(n4192), .Z(n4193) );
  ANDN U4379 ( .B(n4209), .A(n4210), .Z(n4207) );
  IV U4380 ( .A(n4164), .Z(n4148) );
  XOR U4381 ( .A(n4156), .B(n4211), .Z(n4164) );
  XOR U4382 ( .A(n4212), .B(n4202), .Z(n4211) );
  XNOR U4383 ( .A(n4174), .B(n4160), .Z(n4171) );
  NOR U4384 ( .A(n4214), .B(n4174), .Z(n4212) );
  XNOR U4385 ( .A(n4200), .B(n4215), .Z(n4156) );
  XNOR U4386 ( .A(n4216), .B(n4217), .Z(n4215) );
  NANDN U4387 ( .A(n4187), .B(n4218), .Z(n4217) );
  XOR U4388 ( .A(n4219), .B(n4216), .Z(n4200) );
  OR U4389 ( .A(n4196), .B(n4220), .Z(n4216) );
  XOR U4390 ( .A(n4221), .B(n4187), .Z(n4196) );
  XNOR U4391 ( .A(n4192), .B(n4160), .Z(n4187) );
  XOR U4392 ( .A(n4222), .B(n4223), .Z(n4160) );
  NANDN U4393 ( .A(n4224), .B(n4225), .Z(n4223) );
  IV U4394 ( .A(n4210), .Z(n4192) );
  XNOR U4395 ( .A(n4226), .B(n4227), .Z(n4210) );
  NANDN U4396 ( .A(n4224), .B(n4228), .Z(n4227) );
  ANDN U4397 ( .B(n4221), .A(n4229), .Z(n4219) );
  IV U4398 ( .A(n4199), .Z(n4221) );
  XOR U4399 ( .A(n4174), .B(n4155), .Z(n4199) );
  XNOR U4400 ( .A(n4230), .B(n4226), .Z(n4155) );
  NANDN U4401 ( .A(n4231), .B(n4232), .Z(n4226) );
  XOR U4402 ( .A(n4228), .B(n4233), .Z(n4232) );
  ANDN U4403 ( .B(n4233), .A(n4234), .Z(n4230) );
  XOR U4404 ( .A(n4235), .B(n4222), .Z(n4174) );
  NANDN U4405 ( .A(n4231), .B(n4236), .Z(n4222) );
  XOR U4406 ( .A(n4237), .B(n4225), .Z(n4236) );
  XNOR U4407 ( .A(n4238), .B(n4239), .Z(n4224) );
  XOR U4408 ( .A(n4240), .B(n4241), .Z(n4239) );
  XNOR U4409 ( .A(n4242), .B(n4243), .Z(n4238) );
  XNOR U4410 ( .A(n4244), .B(n4245), .Z(n4243) );
  ANDN U4411 ( .B(n4237), .A(n4241), .Z(n4244) );
  ANDN U4412 ( .B(n4237), .A(n4234), .Z(n4235) );
  XNOR U4413 ( .A(n4240), .B(n4246), .Z(n4234) );
  XOR U4414 ( .A(n4247), .B(n4245), .Z(n4246) );
  NAND U4415 ( .A(n4248), .B(n4249), .Z(n4245) );
  XNOR U4416 ( .A(n4242), .B(n4225), .Z(n4249) );
  IV U4417 ( .A(n4237), .Z(n4242) );
  XNOR U4418 ( .A(n4228), .B(n4241), .Z(n4248) );
  IV U4419 ( .A(n4233), .Z(n4241) );
  XOR U4420 ( .A(n4250), .B(n4251), .Z(n4233) );
  XNOR U4421 ( .A(n4252), .B(n4253), .Z(n4251) );
  XNOR U4422 ( .A(n4254), .B(n4255), .Z(n4250) );
  ANDN U4423 ( .B(n4256), .A(n4214), .Z(n4254) );
  AND U4424 ( .A(n4225), .B(n4228), .Z(n4247) );
  XNOR U4425 ( .A(n4225), .B(n4228), .Z(n4240) );
  XNOR U4426 ( .A(n4257), .B(n4258), .Z(n4228) );
  XNOR U4427 ( .A(n4259), .B(n4253), .Z(n4258) );
  XOR U4428 ( .A(n4260), .B(n4261), .Z(n4257) );
  XNOR U4429 ( .A(n4262), .B(n4255), .Z(n4261) );
  OR U4430 ( .A(n4172), .B(n4213), .Z(n4255) );
  XNOR U4431 ( .A(n4263), .B(n4264), .Z(n4213) );
  XNOR U4432 ( .A(n4173), .B(n4161), .Z(n4172) );
  ANDN U4433 ( .B(n4265), .A(n4204), .Z(n4262) );
  XNOR U4434 ( .A(n4266), .B(n4267), .Z(n4225) );
  XNOR U4435 ( .A(n4253), .B(n4268), .Z(n4267) );
  XOR U4436 ( .A(n4183), .B(n4260), .Z(n4268) );
  XNOR U4437 ( .A(n4263), .B(n4173), .Z(n4253) );
  XNOR U4438 ( .A(n4269), .B(n4270), .Z(n4266) );
  XNOR U4439 ( .A(n4271), .B(n4272), .Z(n4270) );
  ANDN U4440 ( .B(n4209), .A(n4191), .Z(n4271) );
  XNOR U4441 ( .A(n4273), .B(n4274), .Z(n4237) );
  XNOR U4442 ( .A(n4259), .B(n4275), .Z(n4274) );
  XNOR U4443 ( .A(n4191), .B(n4252), .Z(n4275) );
  XOR U4444 ( .A(n4260), .B(n4276), .Z(n4252) );
  XNOR U4445 ( .A(n4277), .B(n4278), .Z(n4276) );
  NAND U4446 ( .A(n4218), .B(n4188), .Z(n4278) );
  XNOR U4447 ( .A(n4279), .B(n4277), .Z(n4260) );
  NANDN U4448 ( .A(n4220), .B(n4197), .Z(n4277) );
  XOR U4449 ( .A(n4198), .B(n4188), .Z(n4197) );
  XNOR U4450 ( .A(n4280), .B(n4161), .Z(n4188) );
  XOR U4451 ( .A(n4229), .B(n4218), .Z(n4220) );
  XOR U4452 ( .A(n4209), .B(n4264), .Z(n4218) );
  ANDN U4453 ( .B(n4198), .A(n4229), .Z(n4279) );
  XNOR U4454 ( .A(n4269), .B(n4263), .Z(n4229) );
  IV U4455 ( .A(n4214), .Z(n4263) );
  XNOR U4456 ( .A(n4281), .B(n4282), .Z(n4214) );
  XOR U4457 ( .A(n4283), .B(n4284), .Z(n4282) );
  XOR U4458 ( .A(n4285), .B(n4256), .Z(n4198) );
  XOR U4459 ( .A(n4264), .B(n4265), .Z(n4259) );
  IV U4460 ( .A(n4161), .Z(n4265) );
  XOR U4461 ( .A(n4286), .B(n4287), .Z(n4161) );
  XNOR U4462 ( .A(n4288), .B(n4284), .Z(n4287) );
  IV U4463 ( .A(n4204), .Z(n4264) );
  XOR U4464 ( .A(n4284), .B(n4289), .Z(n4204) );
  XNOR U4465 ( .A(n4209), .B(n4290), .Z(n4273) );
  XNOR U4466 ( .A(n4291), .B(n4272), .Z(n4290) );
  OR U4467 ( .A(n4194), .B(n4208), .Z(n4272) );
  XNOR U4468 ( .A(n4269), .B(n4209), .Z(n4208) );
  XOR U4469 ( .A(n4183), .B(n4280), .Z(n4194) );
  IV U4470 ( .A(n4191), .Z(n4280) );
  XOR U4471 ( .A(n4256), .B(n4292), .Z(n4191) );
  XOR U4472 ( .A(n4288), .B(n4281), .Z(n4292) );
  XNOR U4473 ( .A(key[554]), .B(\w0[4][42] ), .Z(n4281) );
  XOR U4474 ( .A(n4293), .B(n4294), .Z(\w0[4][42] ) );
  XOR U4475 ( .A(n1029), .B(n377), .Z(n4294) );
  XNOR U4476 ( .A(n1036), .B(n412), .Z(n4293) );
  IV U4477 ( .A(n4173), .Z(n4256) );
  XOR U4478 ( .A(n4286), .B(n4295), .Z(n4173) );
  XNOR U4479 ( .A(n4284), .B(n4296), .Z(n4295) );
  ANDN U4480 ( .B(n4285), .A(n4154), .Z(n4291) );
  IV U4481 ( .A(n4183), .Z(n4285) );
  XOR U4482 ( .A(n4286), .B(n4297), .Z(n4183) );
  XOR U4483 ( .A(n4284), .B(n4298), .Z(n4297) );
  XOR U4484 ( .A(n4154), .B(n4299), .Z(n4284) );
  XOR U4485 ( .A(key[558]), .B(\w0[4][46] ), .Z(n4299) );
  XNOR U4486 ( .A(n4300), .B(n4301), .Z(\w0[4][46] ) );
  XNOR U4487 ( .A(n1011), .B(n386), .Z(n4301) );
  XOR U4488 ( .A(n399), .B(n4302), .Z(n386) );
  XNOR U4489 ( .A(n4303), .B(n4304), .Z(n399) );
  IV U4490 ( .A(n4269), .Z(n4154) );
  IV U4491 ( .A(n4289), .Z(n4286) );
  XOR U4492 ( .A(key[557]), .B(\w0[4][45] ), .Z(n4289) );
  XOR U4493 ( .A(n4305), .B(n4306), .Z(\w0[4][45] ) );
  XOR U4494 ( .A(n1024), .B(n390), .Z(n4306) );
  XOR U4495 ( .A(n1009), .B(n4307), .Z(n390) );
  XNOR U4496 ( .A(n4308), .B(n1005), .Z(n4305) );
  IV U4497 ( .A(n4309), .Z(n1005) );
  XOR U4498 ( .A(n4310), .B(n4311), .Z(n4209) );
  XOR U4499 ( .A(n4298), .B(n4296), .Z(n4311) );
  XOR U4500 ( .A(key[559]), .B(\w0[4][47] ), .Z(n4296) );
  XNOR U4501 ( .A(n396), .B(n4312), .Z(\w0[4][47] ) );
  XOR U4502 ( .A(n1006), .B(n417), .Z(n4312) );
  XOR U4503 ( .A(n4313), .B(n4314), .Z(n417) );
  XOR U4504 ( .A(n1017), .B(n4315), .Z(n396) );
  XNOR U4505 ( .A(key[556]), .B(\w0[4][44] ), .Z(n4298) );
  XOR U4506 ( .A(n4316), .B(n4317), .Z(\w0[4][44] ) );
  XOR U4507 ( .A(n403), .B(n4318), .Z(n4317) );
  XOR U4508 ( .A(n1021), .B(n4319), .Z(n403) );
  XOR U4509 ( .A(n1031), .B(n402), .Z(n4316) );
  XNOR U4510 ( .A(n393), .B(n4314), .Z(n402) );
  XNOR U4511 ( .A(n4269), .B(n4283), .Z(n4310) );
  XOR U4512 ( .A(n4288), .B(n4320), .Z(n4283) );
  XOR U4513 ( .A(key[555]), .B(\w0[4][43] ), .Z(n4320) );
  XOR U4514 ( .A(n4321), .B(n4322), .Z(\w0[4][43] ) );
  XOR U4515 ( .A(n410), .B(n4323), .Z(n4322) );
  XOR U4516 ( .A(n405), .B(n4314), .Z(n410) );
  IV U4517 ( .A(n4304), .Z(n4314) );
  XOR U4518 ( .A(n997), .B(n409), .Z(n4321) );
  IV U4519 ( .A(n4324), .Z(n409) );
  XOR U4520 ( .A(key[553]), .B(\w0[4][41] ), .Z(n4288) );
  XOR U4521 ( .A(n4325), .B(n4326), .Z(\w0[4][41] ) );
  XNOR U4522 ( .A(n1040), .B(n413), .Z(n4326) );
  XOR U4523 ( .A(n4327), .B(n379), .Z(n4325) );
  XOR U4524 ( .A(key[552]), .B(\w0[4][40] ), .Z(n4269) );
  XOR U4525 ( .A(n4328), .B(n4329), .Z(\w0[4][40] ) );
  XNOR U4526 ( .A(n416), .B(n4313), .Z(n4329) );
  XOR U4527 ( .A(n1015), .B(n1034), .Z(n4328) );
  XOR U4528 ( .A(n4330), .B(n4331), .Z(out[103]) );
  XNOR U4529 ( .A(n16), .B(n4332), .Z(n4331) );
  IV U4530 ( .A(n4333), .Z(n16) );
  XNOR U4531 ( .A(n8), .B(n4334), .Z(n4330) );
  XNOR U4532 ( .A(key[615]), .B(n12), .Z(n4334) );
  XNOR U4533 ( .A(n4335), .B(n4336), .Z(n8) );
  XNOR U4534 ( .A(n4337), .B(n4338), .Z(n4336) );
  NANDN U4535 ( .A(n4339), .B(n4340), .Z(n4338) );
  XOR U4536 ( .A(n4333), .B(n4341), .Z(out[102]) );
  XNOR U4537 ( .A(key[614]), .B(n10), .Z(n4341) );
  XNOR U4538 ( .A(n4343), .B(n4344), .Z(n4342) );
  OR U4539 ( .A(n4345), .B(n4346), .Z(n4344) );
  XNOR U4540 ( .A(n4347), .B(n4348), .Z(n4335) );
  XNOR U4541 ( .A(n4349), .B(n4350), .Z(n4348) );
  NAND U4542 ( .A(n4351), .B(n4352), .Z(n4350) );
  XNOR U4543 ( .A(n9), .B(n19), .Z(n4333) );
  XNOR U4544 ( .A(n4347), .B(n4353), .Z(n9) );
  XNOR U4545 ( .A(n4337), .B(n4354), .Z(n4353) );
  NANDN U4546 ( .A(n4355), .B(n4356), .Z(n4354) );
  OR U4547 ( .A(n4357), .B(n4358), .Z(n4337) );
  XOR U4548 ( .A(n4359), .B(n4360), .Z(out[101]) );
  XNOR U4549 ( .A(n4332), .B(n4361), .Z(n4360) );
  XOR U4550 ( .A(n4347), .B(n17), .Z(n4361) );
  XOR U4551 ( .A(n4362), .B(n4349), .Z(n4347) );
  NANDN U4552 ( .A(n4363), .B(n4364), .Z(n4349) );
  ANDN U4553 ( .B(n4365), .A(n4366), .Z(n4362) );
  XNOR U4554 ( .A(n4367), .B(n4368), .Z(n4332) );
  XNOR U4555 ( .A(n4369), .B(n4370), .Z(n4368) );
  NANDN U4556 ( .A(n4371), .B(n4340), .Z(n4370) );
  XOR U4557 ( .A(n4372), .B(n4373), .Z(n4359) );
  XNOR U4558 ( .A(key[613]), .B(n4343), .Z(n4373) );
  NANDN U4559 ( .A(n4374), .B(n4375), .Z(n4343) );
  ANDN U4560 ( .B(n4376), .A(n4377), .Z(n4372) );
  XOR U4561 ( .A(n17), .B(n4378), .Z(out[100]) );
  XNOR U4562 ( .A(key[612]), .B(n13), .Z(n4378) );
  XOR U4563 ( .A(n4379), .B(n4380), .Z(n19) );
  XOR U4564 ( .A(n4381), .B(n4369), .Z(n4380) );
  OR U4565 ( .A(n4357), .B(n4382), .Z(n4369) );
  XNOR U4566 ( .A(n4340), .B(n4356), .Z(n4357) );
  ANDN U4567 ( .B(n4383), .A(n4384), .Z(n4381) );
  XNOR U4568 ( .A(n4379), .B(n4385), .Z(n12) );
  XNOR U4569 ( .A(n4386), .B(n4387), .Z(n4385) );
  NAND U4570 ( .A(n4376), .B(n4388), .Z(n4387) );
  XOR U4571 ( .A(n4367), .B(n4389), .Z(n17) );
  XOR U4572 ( .A(n4390), .B(n4386), .Z(n4389) );
  NANDN U4573 ( .A(n4391), .B(n4375), .Z(n4386) );
  XNOR U4574 ( .A(n4345), .B(n4376), .Z(n4375) );
  NOR U4575 ( .A(n4392), .B(n4345), .Z(n4390) );
  XNOR U4576 ( .A(n4379), .B(n4393), .Z(n4367) );
  XNOR U4577 ( .A(n4394), .B(n4395), .Z(n4393) );
  NAND U4578 ( .A(n4352), .B(n4396), .Z(n4395) );
  XOR U4579 ( .A(n4397), .B(n4394), .Z(n4379) );
  OR U4580 ( .A(n4363), .B(n4398), .Z(n4394) );
  XOR U4581 ( .A(n4366), .B(n4352), .Z(n4363) );
  XOR U4582 ( .A(n4356), .B(n4376), .Z(n4352) );
  XOR U4583 ( .A(n4399), .B(n4400), .Z(n4376) );
  NANDN U4584 ( .A(n4401), .B(n4402), .Z(n4400) );
  IV U4585 ( .A(n4384), .Z(n4356) );
  XNOR U4586 ( .A(n4403), .B(n4404), .Z(n4384) );
  NANDN U4587 ( .A(n4401), .B(n4405), .Z(n4404) );
  NOR U4588 ( .A(n4366), .B(n4406), .Z(n4397) );
  XOR U4589 ( .A(n4345), .B(n4340), .Z(n4366) );
  XNOR U4590 ( .A(n4407), .B(n4403), .Z(n4340) );
  NANDN U4591 ( .A(n4408), .B(n4409), .Z(n4403) );
  XOR U4592 ( .A(n4405), .B(n4410), .Z(n4409) );
  ANDN U4593 ( .B(n4410), .A(n4411), .Z(n4407) );
  XOR U4594 ( .A(n4412), .B(n4399), .Z(n4345) );
  NANDN U4595 ( .A(n4408), .B(n4413), .Z(n4399) );
  XOR U4596 ( .A(n4414), .B(n4402), .Z(n4413) );
  XNOR U4597 ( .A(n4415), .B(n4416), .Z(n4401) );
  XOR U4598 ( .A(n4417), .B(n4418), .Z(n4416) );
  XNOR U4599 ( .A(n4419), .B(n4420), .Z(n4415) );
  XNOR U4600 ( .A(n4421), .B(n4422), .Z(n4420) );
  ANDN U4601 ( .B(n4414), .A(n4418), .Z(n4421) );
  ANDN U4602 ( .B(n4414), .A(n4411), .Z(n4412) );
  XNOR U4603 ( .A(n4417), .B(n4423), .Z(n4411) );
  XOR U4604 ( .A(n4424), .B(n4422), .Z(n4423) );
  NAND U4605 ( .A(n4425), .B(n4426), .Z(n4422) );
  XNOR U4606 ( .A(n4419), .B(n4402), .Z(n4426) );
  IV U4607 ( .A(n4414), .Z(n4419) );
  XNOR U4608 ( .A(n4405), .B(n4418), .Z(n4425) );
  IV U4609 ( .A(n4410), .Z(n4418) );
  XOR U4610 ( .A(n4427), .B(n4428), .Z(n4410) );
  XNOR U4611 ( .A(n4429), .B(n4430), .Z(n4428) );
  XNOR U4612 ( .A(n4431), .B(n4432), .Z(n4427) );
  ANDN U4613 ( .B(n4433), .A(n4392), .Z(n4431) );
  AND U4614 ( .A(n4402), .B(n4405), .Z(n4424) );
  XNOR U4615 ( .A(n4402), .B(n4405), .Z(n4417) );
  XNOR U4616 ( .A(n4434), .B(n4435), .Z(n4405) );
  XOR U4617 ( .A(n4436), .B(n4430), .Z(n4435) );
  XNOR U4618 ( .A(n4437), .B(n4438), .Z(n4434) );
  XNOR U4619 ( .A(n4439), .B(n4432), .Z(n4438) );
  OR U4620 ( .A(n4374), .B(n4391), .Z(n4432) );
  XNOR U4621 ( .A(n4440), .B(n4388), .Z(n4391) );
  XNOR U4622 ( .A(n4377), .B(n4346), .Z(n4374) );
  ANDN U4623 ( .B(n4388), .A(n4377), .Z(n4439) );
  XNOR U4624 ( .A(n4441), .B(n4442), .Z(n4402) );
  XNOR U4625 ( .A(n4430), .B(n4443), .Z(n4442) );
  XOR U4626 ( .A(n4339), .B(n4436), .Z(n4443) );
  XNOR U4627 ( .A(n4440), .B(n4346), .Z(n4430) );
  XNOR U4628 ( .A(n4444), .B(n4445), .Z(n4441) );
  XNOR U4629 ( .A(n4446), .B(n4447), .Z(n4445) );
  ANDN U4630 ( .B(n4383), .A(n4355), .Z(n4446) );
  XNOR U4631 ( .A(n4448), .B(n4449), .Z(n4414) );
  XNOR U4632 ( .A(n4429), .B(n4450), .Z(n4449) );
  XNOR U4633 ( .A(n4437), .B(n4355), .Z(n4450) );
  XOR U4634 ( .A(n4388), .B(n4451), .Z(n4437) );
  XOR U4635 ( .A(n4436), .B(n4452), .Z(n4429) );
  XNOR U4636 ( .A(n4453), .B(n4454), .Z(n4452) );
  NAND U4637 ( .A(n4396), .B(n4351), .Z(n4454) );
  XNOR U4638 ( .A(n4455), .B(n4453), .Z(n4436) );
  NANDN U4639 ( .A(n4398), .B(n4364), .Z(n4453) );
  XOR U4640 ( .A(n4365), .B(n4351), .Z(n4364) );
  XNOR U4641 ( .A(n4451), .B(n4355), .Z(n4351) );
  IV U4642 ( .A(n4377), .Z(n4451) );
  XOR U4643 ( .A(n4456), .B(n4457), .Z(n4377) );
  XOR U4644 ( .A(n4458), .B(n4459), .Z(n4457) );
  XOR U4645 ( .A(n4406), .B(n4396), .Z(n4398) );
  XOR U4646 ( .A(n4388), .B(n4383), .Z(n4396) );
  ANDN U4647 ( .B(n4365), .A(n4406), .Z(n4455) );
  XNOR U4648 ( .A(n4444), .B(n4440), .Z(n4406) );
  IV U4649 ( .A(n4392), .Z(n4440) );
  XOR U4650 ( .A(n4460), .B(n4461), .Z(n4392) );
  XOR U4651 ( .A(n4462), .B(n4458), .Z(n4461) );
  XOR U4652 ( .A(n4463), .B(n4433), .Z(n4365) );
  XNOR U4653 ( .A(n4383), .B(n4464), .Z(n4448) );
  XNOR U4654 ( .A(n4465), .B(n4447), .Z(n4464) );
  OR U4655 ( .A(n4358), .B(n4382), .Z(n4447) );
  XNOR U4656 ( .A(n4444), .B(n4383), .Z(n4382) );
  XNOR U4657 ( .A(n4339), .B(n4355), .Z(n4358) );
  XOR U4658 ( .A(n4433), .B(n4466), .Z(n4355) );
  XNOR U4659 ( .A(n4462), .B(n4459), .Z(n4466) );
  XOR U4660 ( .A(key[514]), .B(\w0[4][2] ), .Z(n4462) );
  XOR U4661 ( .A(n612), .B(n4467), .Z(\w0[4][2] ) );
  XNOR U4662 ( .A(n1824), .B(n1232), .Z(n4467) );
  XNOR U4663 ( .A(n4468), .B(n626), .Z(n1232) );
  IV U4664 ( .A(n1231), .Z(n612) );
  XNOR U4665 ( .A(n1797), .B(n624), .Z(n1231) );
  XOR U4666 ( .A(n4469), .B(n4470), .Z(n624) );
  XNOR U4667 ( .A(n4471), .B(n4472), .Z(n4470) );
  XNOR U4668 ( .A(n4473), .B(n4474), .Z(n4469) );
  IV U4669 ( .A(n4346), .Z(n4433) );
  XNOR U4670 ( .A(n4475), .B(n4388), .Z(n4346) );
  IV U4671 ( .A(n4463), .Z(n4339) );
  ANDN U4672 ( .B(n4463), .A(n4371), .Z(n4465) );
  XOR U4673 ( .A(n4476), .B(n4388), .Z(n4463) );
  XNOR U4674 ( .A(n4458), .B(n4456), .Z(n4388) );
  XNOR U4675 ( .A(key[517]), .B(\w0[4][5] ), .Z(n4456) );
  XNOR U4676 ( .A(n1209), .B(n4477), .Z(\w0[4][5] ) );
  XNOR U4677 ( .A(n1204), .B(n1808), .Z(n4477) );
  XNOR U4678 ( .A(n1208), .B(n593), .Z(n1808) );
  XNOR U4679 ( .A(n4478), .B(n4479), .Z(n593) );
  XNOR U4680 ( .A(n4480), .B(n4481), .Z(n4479) );
  XNOR U4681 ( .A(n4482), .B(n4483), .Z(n4478) );
  XOR U4682 ( .A(n4484), .B(n4485), .Z(n4483) );
  ANDN U4683 ( .B(n4486), .A(n4487), .Z(n4485) );
  IV U4684 ( .A(n1225), .Z(n1208) );
  XOR U4685 ( .A(n4488), .B(n4489), .Z(n1225) );
  XNOR U4686 ( .A(n4490), .B(n4491), .Z(n4489) );
  XNOR U4687 ( .A(n4492), .B(n4493), .Z(n4488) );
  XNOR U4688 ( .A(n4494), .B(n4495), .Z(n4493) );
  ANDN U4689 ( .B(n4496), .A(n4497), .Z(n4495) );
  XOR U4690 ( .A(n1809), .B(n596), .Z(n1204) );
  XOR U4691 ( .A(n4498), .B(n4472), .Z(n596) );
  XNOR U4692 ( .A(n4499), .B(n4500), .Z(n4472) );
  XNOR U4693 ( .A(n4501), .B(n4502), .Z(n4500) );
  ANDN U4694 ( .B(n4503), .A(n4504), .Z(n4501) );
  XNOR U4695 ( .A(n4371), .B(n4505), .Z(n4458) );
  XOR U4696 ( .A(key[518]), .B(\w0[4][6] ), .Z(n4505) );
  XNOR U4697 ( .A(n1809), .B(n4506), .Z(\w0[4][6] ) );
  XOR U4698 ( .A(n601), .B(n1804), .Z(n4506) );
  XOR U4699 ( .A(n4507), .B(n1207), .Z(n1804) );
  XNOR U4700 ( .A(n602), .B(n595), .Z(n1207) );
  XNOR U4701 ( .A(n4508), .B(n4509), .Z(n595) );
  XOR U4702 ( .A(n4510), .B(n4511), .Z(n602) );
  XOR U4703 ( .A(n605), .B(n1218), .Z(n601) );
  XOR U4704 ( .A(n4512), .B(n4513), .Z(n1218) );
  XNOR U4705 ( .A(n4498), .B(n4514), .Z(n4513) );
  XOR U4706 ( .A(n4515), .B(n4474), .Z(n4512) );
  XOR U4707 ( .A(n4516), .B(n4517), .Z(n1809) );
  IV U4708 ( .A(n4444), .Z(n4371) );
  XOR U4709 ( .A(n4518), .B(n4519), .Z(n4383) );
  XNOR U4710 ( .A(n4476), .B(n4475), .Z(n4519) );
  XOR U4711 ( .A(key[519]), .B(\w0[4][7] ), .Z(n4475) );
  XNOR U4712 ( .A(n4507), .B(n4520), .Z(\w0[4][7] ) );
  XNOR U4713 ( .A(n605), .B(n1813), .Z(n4520) );
  XNOR U4714 ( .A(n589), .B(n1215), .Z(n1813) );
  XOR U4715 ( .A(n4521), .B(n4522), .Z(n1215) );
  XNOR U4716 ( .A(n4523), .B(n4490), .Z(n4522) );
  XNOR U4717 ( .A(n4524), .B(n4525), .Z(n4490) );
  XNOR U4718 ( .A(n4526), .B(n4527), .Z(n4525) );
  NANDN U4719 ( .A(n4528), .B(n4529), .Z(n4527) );
  XNOR U4720 ( .A(n4530), .B(n4508), .Z(n4521) );
  XNOR U4721 ( .A(n4531), .B(n4532), .Z(n589) );
  XNOR U4722 ( .A(n4510), .B(n4481), .Z(n4532) );
  XNOR U4723 ( .A(n4533), .B(n4534), .Z(n4481) );
  XNOR U4724 ( .A(n4535), .B(n4536), .Z(n4534) );
  OR U4725 ( .A(n4537), .B(n4538), .Z(n4536) );
  XOR U4726 ( .A(n1235), .B(n1217), .Z(n4507) );
  XOR U4727 ( .A(n4539), .B(n4540), .Z(n1217) );
  XNOR U4728 ( .A(n4516), .B(n4541), .Z(n4540) );
  XOR U4729 ( .A(key[516]), .B(\w0[4][4] ), .Z(n4476) );
  XOR U4730 ( .A(n4542), .B(n4543), .Z(\w0[4][4] ) );
  XOR U4731 ( .A(n4544), .B(n1817), .Z(n4543) );
  XOR U4732 ( .A(n1220), .B(n581), .Z(n1817) );
  XNOR U4733 ( .A(n4480), .B(n626), .Z(n581) );
  XOR U4734 ( .A(n4545), .B(n4546), .Z(n626) );
  XNOR U4735 ( .A(n621), .B(n4491), .Z(n1220) );
  IV U4736 ( .A(n4468), .Z(n621) );
  XOR U4737 ( .A(n4547), .B(n4548), .Z(n4468) );
  XOR U4738 ( .A(n580), .B(n1816), .Z(n4542) );
  XNOR U4739 ( .A(n4549), .B(n1209), .Z(n1816) );
  XOR U4740 ( .A(n4550), .B(n4551), .Z(n1209) );
  XNOR U4741 ( .A(n4552), .B(n4541), .Z(n4551) );
  XNOR U4742 ( .A(n4553), .B(n4554), .Z(n4541) );
  XNOR U4743 ( .A(n4555), .B(n4556), .Z(n4554) );
  OR U4744 ( .A(n4557), .B(n4558), .Z(n4556) );
  XNOR U4745 ( .A(n4559), .B(n4560), .Z(n4550) );
  XOR U4746 ( .A(n4561), .B(n4562), .Z(n4560) );
  ANDN U4747 ( .B(n4563), .A(n4564), .Z(n4562) );
  XNOR U4748 ( .A(n605), .B(n1210), .Z(n580) );
  XNOR U4749 ( .A(n4565), .B(n4566), .Z(n1210) );
  XOR U4750 ( .A(n4567), .B(n4514), .Z(n4566) );
  XNOR U4751 ( .A(n4568), .B(n4569), .Z(n4514) );
  XNOR U4752 ( .A(n4570), .B(n4571), .Z(n4569) );
  OR U4753 ( .A(n4572), .B(n4573), .Z(n4571) );
  XNOR U4754 ( .A(n4574), .B(n4575), .Z(n4565) );
  XOR U4755 ( .A(n4502), .B(n4576), .Z(n4575) );
  ANDN U4756 ( .B(n4577), .A(n4578), .Z(n4576) );
  ANDN U4757 ( .B(n4579), .A(n4580), .Z(n4502) );
  XOR U4758 ( .A(n4444), .B(n4460), .Z(n4518) );
  XNOR U4759 ( .A(n4459), .B(n4581), .Z(n4460) );
  XOR U4760 ( .A(key[515]), .B(\w0[4][3] ), .Z(n4581) );
  XOR U4761 ( .A(n4582), .B(n4583), .Z(\w0[4][3] ) );
  XNOR U4762 ( .A(n1797), .B(n1196), .Z(n4583) );
  XNOR U4763 ( .A(n615), .B(n627), .Z(n1196) );
  XOR U4764 ( .A(n4584), .B(n4585), .Z(n627) );
  XNOR U4765 ( .A(n4586), .B(n4509), .Z(n4585) );
  XNOR U4766 ( .A(n4587), .B(n4588), .Z(n4509) );
  XOR U4767 ( .A(n4589), .B(n4494), .Z(n4588) );
  OR U4768 ( .A(n4590), .B(n4591), .Z(n4494) );
  NOR U4769 ( .A(n4592), .B(n4593), .Z(n4589) );
  XNOR U4770 ( .A(n4547), .B(n4594), .Z(n4584) );
  IV U4771 ( .A(n4530), .Z(n4547) );
  XOR U4772 ( .A(n4531), .B(n4595), .Z(n615) );
  XOR U4773 ( .A(n4596), .B(n4511), .Z(n4595) );
  XOR U4774 ( .A(n4597), .B(n4598), .Z(n4511) );
  XNOR U4775 ( .A(n4599), .B(n4484), .Z(n4598) );
  ANDN U4776 ( .B(n4600), .A(n4601), .Z(n4484) );
  ANDN U4777 ( .B(n4602), .A(n4603), .Z(n4599) );
  XNOR U4778 ( .A(n4604), .B(n4605), .Z(n4531) );
  XOR U4779 ( .A(n4539), .B(n4606), .Z(n1797) );
  XOR U4780 ( .A(n4607), .B(n4517), .Z(n4606) );
  XOR U4781 ( .A(n4608), .B(n4609), .Z(n4517) );
  XNOR U4782 ( .A(n4610), .B(n4561), .Z(n4609) );
  ANDN U4783 ( .B(n4611), .A(n4612), .Z(n4561) );
  ANDN U4784 ( .B(n4613), .A(n4614), .Z(n4610) );
  XNOR U4785 ( .A(n4615), .B(n4616), .Z(n4539) );
  XNOR U4786 ( .A(n614), .B(n1821), .Z(n4582) );
  XNOR U4787 ( .A(n4549), .B(n4544), .Z(n1821) );
  IV U4788 ( .A(n1226), .Z(n4544) );
  XNOR U4789 ( .A(n4552), .B(n1824), .Z(n1226) );
  XOR U4790 ( .A(n605), .B(n1224), .Z(n614) );
  XOR U4791 ( .A(n619), .B(n4567), .Z(n1224) );
  XOR U4792 ( .A(n4617), .B(n4567), .Z(n605) );
  XOR U4793 ( .A(n4568), .B(n4618), .Z(n4567) );
  XOR U4794 ( .A(n4619), .B(n4620), .Z(n4618) );
  ANDN U4795 ( .B(n4503), .A(n4621), .Z(n4619) );
  XNOR U4796 ( .A(n4622), .B(n4623), .Z(n4568) );
  XNOR U4797 ( .A(n4624), .B(n4625), .Z(n4623) );
  NAND U4798 ( .A(n4626), .B(n4627), .Z(n4625) );
  XOR U4799 ( .A(key[513]), .B(\w0[4][1] ), .Z(n4459) );
  XNOR U4800 ( .A(n625), .B(n4628), .Z(\w0[4][1] ) );
  XOR U4801 ( .A(n4629), .B(n1236), .Z(n4628) );
  XOR U4802 ( .A(n618), .B(n606), .Z(n1236) );
  XNOR U4803 ( .A(n4586), .B(n4630), .Z(n606) );
  XOR U4804 ( .A(n4530), .B(n4508), .Z(n4630) );
  XOR U4805 ( .A(n4548), .B(n4594), .Z(n4508) );
  XNOR U4806 ( .A(n4492), .B(n4631), .Z(n4594) );
  XNOR U4807 ( .A(n4632), .B(n4633), .Z(n4631) );
  NANDN U4808 ( .A(n4634), .B(n4635), .Z(n4633) );
  XNOR U4809 ( .A(n4636), .B(n4637), .Z(n4530) );
  XNOR U4810 ( .A(n4638), .B(n4639), .Z(n4637) );
  NAND U4811 ( .A(n4496), .B(n4640), .Z(n4639) );
  IV U4812 ( .A(n4523), .Z(n4586) );
  XOR U4813 ( .A(n4587), .B(n4641), .Z(n4523) );
  XNOR U4814 ( .A(n4632), .B(n4642), .Z(n4641) );
  NANDN U4815 ( .A(n4643), .B(n4529), .Z(n4642) );
  OR U4816 ( .A(n4644), .B(n4645), .Z(n4632) );
  XOR U4817 ( .A(n4492), .B(n4646), .Z(n4587) );
  XNOR U4818 ( .A(n4647), .B(n4648), .Z(n4646) );
  NAND U4819 ( .A(n4649), .B(n4650), .Z(n4648) );
  XOR U4820 ( .A(n4651), .B(n4647), .Z(n4492) );
  NANDN U4821 ( .A(n4652), .B(n4653), .Z(n4647) );
  ANDN U4822 ( .B(n4654), .A(n4655), .Z(n4651) );
  XNOR U4823 ( .A(n4510), .B(n4656), .Z(n618) );
  XOR U4824 ( .A(n4604), .B(n4605), .Z(n4656) );
  XOR U4825 ( .A(n4597), .B(n4657), .Z(n4605) );
  XNOR U4826 ( .A(n4658), .B(n4659), .Z(n4657) );
  OR U4827 ( .A(n4537), .B(n4660), .Z(n4659) );
  XNOR U4828 ( .A(n4482), .B(n4661), .Z(n4597) );
  XNOR U4829 ( .A(n4662), .B(n4663), .Z(n4661) );
  NAND U4830 ( .A(n4664), .B(n4665), .Z(n4663) );
  IV U4831 ( .A(n4545), .Z(n4604) );
  XOR U4832 ( .A(n4666), .B(n4667), .Z(n4545) );
  XNOR U4833 ( .A(n4668), .B(n4669), .Z(n4667) );
  NAND U4834 ( .A(n4670), .B(n4486), .Z(n4669) );
  XOR U4835 ( .A(n4546), .B(n4596), .Z(n4510) );
  XNOR U4836 ( .A(n4482), .B(n4671), .Z(n4596) );
  XNOR U4837 ( .A(n4658), .B(n4672), .Z(n4671) );
  NANDN U4838 ( .A(n4673), .B(n4674), .Z(n4672) );
  OR U4839 ( .A(n4675), .B(n4676), .Z(n4658) );
  XOR U4840 ( .A(n4677), .B(n4662), .Z(n4482) );
  NANDN U4841 ( .A(n4678), .B(n4679), .Z(n4662) );
  ANDN U4842 ( .B(n4680), .A(n4681), .Z(n4677) );
  XNOR U4843 ( .A(n619), .B(n1824), .Z(n625) );
  XOR U4844 ( .A(n4682), .B(n4683), .Z(n1824) );
  XOR U4845 ( .A(n4515), .B(n4617), .Z(n619) );
  XOR U4846 ( .A(key[512]), .B(\w0[4][0] ), .Z(n4444) );
  XOR U4847 ( .A(n1216), .B(n4684), .Z(\w0[4][0] ) );
  XNOR U4848 ( .A(n620), .B(n608), .Z(n4684) );
  XNOR U4849 ( .A(n1214), .B(n1235), .Z(n608) );
  IV U4850 ( .A(n4549), .Z(n1235) );
  XOR U4851 ( .A(n4683), .B(n4552), .Z(n4549) );
  XNOR U4852 ( .A(n4553), .B(n4685), .Z(n4552) );
  XOR U4853 ( .A(n4686), .B(n4687), .Z(n4685) );
  ANDN U4854 ( .B(n4613), .A(n4688), .Z(n4686) );
  XNOR U4855 ( .A(n4689), .B(n4690), .Z(n4553) );
  XNOR U4856 ( .A(n4691), .B(n4692), .Z(n4690) );
  NAND U4857 ( .A(n4693), .B(n4694), .Z(n4692) );
  IV U4858 ( .A(n1805), .Z(n1214) );
  XOR U4859 ( .A(n4546), .B(n4480), .Z(n1805) );
  XNOR U4860 ( .A(n4533), .B(n4695), .Z(n4480) );
  XOR U4861 ( .A(n4696), .B(n4668), .Z(n4695) );
  XOR U4862 ( .A(n4602), .B(n4486), .Z(n4600) );
  ANDN U4863 ( .B(n4602), .A(n4698), .Z(n4696) );
  XNOR U4864 ( .A(n4666), .B(n4699), .Z(n4533) );
  XNOR U4865 ( .A(n4700), .B(n4701), .Z(n4699) );
  NAND U4866 ( .A(n4665), .B(n4702), .Z(n4701) );
  XOR U4867 ( .A(n4666), .B(n4703), .Z(n4546) );
  XOR U4868 ( .A(n4704), .B(n4535), .Z(n4703) );
  OR U4869 ( .A(n4705), .B(n4675), .Z(n4535) );
  XNOR U4870 ( .A(n4537), .B(n4673), .Z(n4675) );
  NOR U4871 ( .A(n4706), .B(n4673), .Z(n4704) );
  XOR U4872 ( .A(n4707), .B(n4700), .Z(n4666) );
  OR U4873 ( .A(n4678), .B(n4708), .Z(n4700) );
  XNOR U4874 ( .A(n4709), .B(n4665), .Z(n4678) );
  XNOR U4875 ( .A(n4673), .B(n4486), .Z(n4665) );
  XOR U4876 ( .A(n4710), .B(n4711), .Z(n4486) );
  NANDN U4877 ( .A(n4712), .B(n4713), .Z(n4711) );
  XNOR U4878 ( .A(n4714), .B(n4715), .Z(n4673) );
  OR U4879 ( .A(n4712), .B(n4716), .Z(n4715) );
  ANDN U4880 ( .B(n4709), .A(n4717), .Z(n4707) );
  IV U4881 ( .A(n4681), .Z(n4709) );
  XOR U4882 ( .A(n4537), .B(n4602), .Z(n4681) );
  XNOR U4883 ( .A(n4718), .B(n4710), .Z(n4602) );
  NANDN U4884 ( .A(n4719), .B(n4720), .Z(n4710) );
  ANDN U4885 ( .B(n4721), .A(n4722), .Z(n4718) );
  NANDN U4886 ( .A(n4719), .B(n4724), .Z(n4714) );
  XOR U4887 ( .A(n4725), .B(n4712), .Z(n4719) );
  XNOR U4888 ( .A(n4726), .B(n4727), .Z(n4712) );
  XOR U4889 ( .A(n4728), .B(n4721), .Z(n4727) );
  XNOR U4890 ( .A(n4729), .B(n4730), .Z(n4726) );
  XNOR U4891 ( .A(n4731), .B(n4732), .Z(n4730) );
  ANDN U4892 ( .B(n4721), .A(n4733), .Z(n4731) );
  IV U4893 ( .A(n4734), .Z(n4721) );
  ANDN U4894 ( .B(n4725), .A(n4733), .Z(n4723) );
  IV U4895 ( .A(n4729), .Z(n4733) );
  IV U4896 ( .A(n4722), .Z(n4725) );
  XNOR U4897 ( .A(n4728), .B(n4735), .Z(n4722) );
  XOR U4898 ( .A(n4736), .B(n4732), .Z(n4735) );
  NAND U4899 ( .A(n4724), .B(n4720), .Z(n4732) );
  XNOR U4900 ( .A(n4713), .B(n4734), .Z(n4720) );
  XOR U4901 ( .A(n4737), .B(n4738), .Z(n4734) );
  XOR U4902 ( .A(n4739), .B(n4740), .Z(n4738) );
  XNOR U4903 ( .A(n4674), .B(n4741), .Z(n4740) );
  XNOR U4904 ( .A(n4742), .B(n4743), .Z(n4737) );
  XNOR U4905 ( .A(n4744), .B(n4745), .Z(n4743) );
  ANDN U4906 ( .B(n4746), .A(n4538), .Z(n4744) );
  XNOR U4907 ( .A(n4729), .B(n4716), .Z(n4724) );
  XOR U4908 ( .A(n4747), .B(n4748), .Z(n4729) );
  XNOR U4909 ( .A(n4749), .B(n4741), .Z(n4748) );
  XOR U4910 ( .A(n4750), .B(n4751), .Z(n4741) );
  XNOR U4911 ( .A(n4752), .B(n4753), .Z(n4751) );
  NAND U4912 ( .A(n4702), .B(n4664), .Z(n4753) );
  XNOR U4913 ( .A(n4754), .B(n4755), .Z(n4747) );
  ANDN U4914 ( .B(n4756), .A(n4698), .Z(n4754) );
  ANDN U4915 ( .B(n4713), .A(n4716), .Z(n4736) );
  XOR U4916 ( .A(n4716), .B(n4713), .Z(n4728) );
  XNOR U4917 ( .A(n4757), .B(n4758), .Z(n4713) );
  XNOR U4918 ( .A(n4750), .B(n4759), .Z(n4758) );
  XOR U4919 ( .A(n4749), .B(n4660), .Z(n4759) );
  XOR U4920 ( .A(n4538), .B(n4760), .Z(n4757) );
  XNOR U4921 ( .A(n4761), .B(n4745), .Z(n4760) );
  OR U4922 ( .A(n4676), .B(n4705), .Z(n4745) );
  XNOR U4923 ( .A(n4538), .B(n4706), .Z(n4705) );
  XOR U4924 ( .A(n4660), .B(n4674), .Z(n4676) );
  ANDN U4925 ( .B(n4674), .A(n4706), .Z(n4761) );
  XOR U4926 ( .A(n4762), .B(n4763), .Z(n4716) );
  XOR U4927 ( .A(n4750), .B(n4739), .Z(n4763) );
  XOR U4928 ( .A(n4670), .B(n4487), .Z(n4739) );
  XOR U4929 ( .A(n4764), .B(n4752), .Z(n4750) );
  NANDN U4930 ( .A(n4708), .B(n4679), .Z(n4752) );
  XOR U4931 ( .A(n4680), .B(n4664), .Z(n4679) );
  XNOR U4932 ( .A(n4756), .B(n4765), .Z(n4674) );
  XNOR U4933 ( .A(n4766), .B(n4767), .Z(n4765) );
  XOR U4934 ( .A(n4717), .B(n4702), .Z(n4708) );
  XNOR U4935 ( .A(n4706), .B(n4670), .Z(n4702) );
  IV U4936 ( .A(n4742), .Z(n4706) );
  XOR U4937 ( .A(n4768), .B(n4769), .Z(n4742) );
  XOR U4938 ( .A(n4770), .B(n4771), .Z(n4769) );
  XNOR U4939 ( .A(n4538), .B(n4772), .Z(n4768) );
  ANDN U4940 ( .B(n4680), .A(n4717), .Z(n4764) );
  XNOR U4941 ( .A(n4538), .B(n4698), .Z(n4717) );
  XOR U4942 ( .A(n4756), .B(n4746), .Z(n4680) );
  IV U4943 ( .A(n4660), .Z(n4746) );
  XOR U4944 ( .A(n4773), .B(n4774), .Z(n4660) );
  XOR U4945 ( .A(n4775), .B(n4771), .Z(n4774) );
  XNOR U4946 ( .A(n4776), .B(n4777), .Z(n4771) );
  XNOR U4947 ( .A(n4778), .B(n2873), .Z(n4777) );
  XOR U4948 ( .A(n2894), .B(n4120), .Z(n2873) );
  XNOR U4949 ( .A(n4779), .B(n4780), .Z(n4776) );
  XNOR U4950 ( .A(key[500]), .B(n4099), .Z(n4780) );
  IV U4951 ( .A(n4603), .Z(n4756) );
  XOR U4952 ( .A(n4749), .B(n4781), .Z(n4762) );
  XNOR U4953 ( .A(n4782), .B(n4755), .Z(n4781) );
  OR U4954 ( .A(n4601), .B(n4697), .Z(n4755) );
  XNOR U4955 ( .A(n4783), .B(n4670), .Z(n4697) );
  XNOR U4956 ( .A(n4603), .B(n4487), .Z(n4601) );
  ANDN U4957 ( .B(n4670), .A(n4487), .Z(n4782) );
  XOR U4958 ( .A(n4773), .B(n4784), .Z(n4487) );
  XOR U4959 ( .A(n4766), .B(n4785), .Z(n4784) );
  XOR U4960 ( .A(n4775), .B(n4773), .Z(n4670) );
  XNOR U4961 ( .A(n4698), .B(n4603), .Z(n4749) );
  XOR U4962 ( .A(n4773), .B(n4786), .Z(n4603) );
  XNOR U4963 ( .A(n4775), .B(n4770), .Z(n4786) );
  XOR U4964 ( .A(n4787), .B(n4788), .Z(n4770) );
  XNOR U4965 ( .A(n4789), .B(n4790), .Z(n4788) );
  XNOR U4966 ( .A(key[503]), .B(n2894), .Z(n4787) );
  XNOR U4967 ( .A(n4791), .B(n4792), .Z(n4773) );
  XOR U4968 ( .A(n4793), .B(n4144), .Z(n4792) );
  XOR U4969 ( .A(n4794), .B(n4795), .Z(n4144) );
  XOR U4970 ( .A(key[501]), .B(n4119), .Z(n4791) );
  IV U4971 ( .A(n4783), .Z(n4698) );
  XNOR U4972 ( .A(n4767), .B(n4796), .Z(n4783) );
  XOR U4973 ( .A(n4772), .B(n4785), .Z(n4796) );
  IV U4974 ( .A(n4775), .Z(n4785) );
  XOR U4975 ( .A(n4797), .B(n4798), .Z(n4775) );
  XOR U4976 ( .A(n4794), .B(n2852), .Z(n4798) );
  XOR U4977 ( .A(n2894), .B(n4115), .Z(n2852) );
  XNOR U4978 ( .A(n4799), .B(n4800), .Z(n4797) );
  XOR U4979 ( .A(key[502]), .B(n4538), .Z(n4800) );
  XNOR U4980 ( .A(n4801), .B(n4802), .Z(n4538) );
  XOR U4981 ( .A(n2887), .B(n4803), .Z(n4802) );
  XOR U4982 ( .A(n4804), .B(n4805), .Z(n2887) );
  XNOR U4983 ( .A(key[496]), .B(n4103), .Z(n4801) );
  XOR U4984 ( .A(n4806), .B(n4807), .Z(n4772) );
  XNOR U4985 ( .A(n4135), .B(n4808), .Z(n4807) );
  XNOR U4986 ( .A(n4766), .B(n2890), .Z(n4808) );
  XOR U4987 ( .A(n2894), .B(n4100), .Z(n2890) );
  XOR U4988 ( .A(n4809), .B(n4810), .Z(n4766) );
  XOR U4989 ( .A(n4141), .B(n2844), .Z(n4810) );
  XOR U4990 ( .A(n4811), .B(n4812), .Z(n2844) );
  XNOR U4991 ( .A(key[497]), .B(n4804), .Z(n4809) );
  IV U4992 ( .A(n4813), .Z(n4135) );
  XNOR U4993 ( .A(n4814), .B(n4815), .Z(n4806) );
  XNOR U4994 ( .A(key[499]), .B(n4816), .Z(n4815) );
  XOR U4995 ( .A(n4817), .B(n4818), .Z(n4767) );
  XNOR U4996 ( .A(n4129), .B(n2880), .Z(n4818) );
  IV U4997 ( .A(n4131), .Z(n2880) );
  XNOR U4998 ( .A(n4814), .B(n2841), .Z(n4131) );
  XOR U4999 ( .A(key[498]), .B(n4811), .Z(n4817) );
  XNOR U5000 ( .A(n4629), .B(n607), .Z(n620) );
  XOR U5001 ( .A(n4498), .B(n4819), .Z(n607) );
  XOR U5002 ( .A(n4473), .B(n4474), .Z(n4819) );
  XOR U5003 ( .A(n4499), .B(n4820), .Z(n4474) );
  XNOR U5004 ( .A(n4821), .B(n4822), .Z(n4820) );
  NANDN U5005 ( .A(n4572), .B(n4823), .Z(n4822) );
  XNOR U5006 ( .A(n4574), .B(n4824), .Z(n4499) );
  XNOR U5007 ( .A(n4825), .B(n4826), .Z(n4824) );
  NAND U5008 ( .A(n4827), .B(n4626), .Z(n4826) );
  IV U5009 ( .A(n4515), .Z(n4473) );
  XOR U5010 ( .A(n4622), .B(n4828), .Z(n4515) );
  XNOR U5011 ( .A(n4620), .B(n4829), .Z(n4828) );
  NAND U5012 ( .A(n4830), .B(n4577), .Z(n4829) );
  XOR U5013 ( .A(n4503), .B(n4577), .Z(n4579) );
  XOR U5014 ( .A(n4471), .B(n4617), .Z(n4498) );
  XOR U5015 ( .A(n4622), .B(n4832), .Z(n4617) );
  XOR U5016 ( .A(n4833), .B(n4570), .Z(n4832) );
  OR U5017 ( .A(n4834), .B(n4835), .Z(n4570) );
  NOR U5018 ( .A(n4836), .B(n4837), .Z(n4833) );
  XOR U5019 ( .A(n4838), .B(n4624), .Z(n4622) );
  OR U5020 ( .A(n4839), .B(n4840), .Z(n4624) );
  ANDN U5021 ( .B(n4841), .A(n4842), .Z(n4838) );
  XNOR U5022 ( .A(n4574), .B(n4843), .Z(n4471) );
  XNOR U5023 ( .A(n4821), .B(n4844), .Z(n4843) );
  NANDN U5024 ( .A(n4837), .B(n4845), .Z(n4844) );
  OR U5025 ( .A(n4834), .B(n4846), .Z(n4821) );
  XNOR U5026 ( .A(n4572), .B(n4837), .Z(n4834) );
  XOR U5027 ( .A(n4847), .B(n4825), .Z(n4574) );
  NANDN U5028 ( .A(n4839), .B(n4848), .Z(n4825) );
  XOR U5029 ( .A(n4842), .B(n4626), .Z(n4839) );
  XNOR U5030 ( .A(n4837), .B(n4577), .Z(n4626) );
  XOR U5031 ( .A(n4849), .B(n4850), .Z(n4577) );
  NANDN U5032 ( .A(n4851), .B(n4852), .Z(n4850) );
  XNOR U5033 ( .A(n4853), .B(n4854), .Z(n4837) );
  OR U5034 ( .A(n4851), .B(n4855), .Z(n4854) );
  ANDN U5035 ( .B(n4856), .A(n4842), .Z(n4847) );
  XOR U5036 ( .A(n4572), .B(n4503), .Z(n4842) );
  XNOR U5037 ( .A(n4857), .B(n4849), .Z(n4503) );
  NANDN U5038 ( .A(n4858), .B(n4859), .Z(n4849) );
  ANDN U5039 ( .B(n4860), .A(n4861), .Z(n4857) );
  NANDN U5040 ( .A(n4858), .B(n4863), .Z(n4853) );
  XOR U5041 ( .A(n4864), .B(n4851), .Z(n4858) );
  XNOR U5042 ( .A(n4865), .B(n4866), .Z(n4851) );
  XOR U5043 ( .A(n4867), .B(n4860), .Z(n4866) );
  XNOR U5044 ( .A(n4868), .B(n4869), .Z(n4865) );
  XNOR U5045 ( .A(n4870), .B(n4871), .Z(n4869) );
  ANDN U5046 ( .B(n4860), .A(n4872), .Z(n4870) );
  IV U5047 ( .A(n4873), .Z(n4860) );
  ANDN U5048 ( .B(n4864), .A(n4872), .Z(n4862) );
  IV U5049 ( .A(n4868), .Z(n4872) );
  IV U5050 ( .A(n4861), .Z(n4864) );
  XNOR U5051 ( .A(n4867), .B(n4874), .Z(n4861) );
  XOR U5052 ( .A(n4875), .B(n4871), .Z(n4874) );
  NAND U5053 ( .A(n4863), .B(n4859), .Z(n4871) );
  XNOR U5054 ( .A(n4852), .B(n4873), .Z(n4859) );
  XOR U5055 ( .A(n4876), .B(n4877), .Z(n4873) );
  XOR U5056 ( .A(n4878), .B(n4879), .Z(n4877) );
  XNOR U5057 ( .A(n4845), .B(n4880), .Z(n4879) );
  XNOR U5058 ( .A(n4881), .B(n4882), .Z(n4876) );
  XNOR U5059 ( .A(n4883), .B(n4884), .Z(n4882) );
  ANDN U5060 ( .B(n4823), .A(n4573), .Z(n4883) );
  XNOR U5061 ( .A(n4868), .B(n4855), .Z(n4863) );
  XOR U5062 ( .A(n4885), .B(n4886), .Z(n4868) );
  XNOR U5063 ( .A(n4887), .B(n4880), .Z(n4886) );
  XOR U5064 ( .A(n4888), .B(n4889), .Z(n4880) );
  XNOR U5065 ( .A(n4890), .B(n4891), .Z(n4889) );
  NAND U5066 ( .A(n4627), .B(n4827), .Z(n4891) );
  XNOR U5067 ( .A(n4892), .B(n4893), .Z(n4885) );
  ANDN U5068 ( .B(n4894), .A(n4621), .Z(n4892) );
  ANDN U5069 ( .B(n4852), .A(n4855), .Z(n4875) );
  XOR U5070 ( .A(n4855), .B(n4852), .Z(n4867) );
  XNOR U5071 ( .A(n4895), .B(n4896), .Z(n4852) );
  XNOR U5072 ( .A(n4888), .B(n4897), .Z(n4896) );
  XNOR U5073 ( .A(n4887), .B(n4823), .Z(n4897) );
  XNOR U5074 ( .A(n4898), .B(n4899), .Z(n4895) );
  XNOR U5075 ( .A(n4900), .B(n4884), .Z(n4899) );
  OR U5076 ( .A(n4846), .B(n4835), .Z(n4884) );
  XNOR U5077 ( .A(n4898), .B(n4881), .Z(n4835) );
  XNOR U5078 ( .A(n4823), .B(n4845), .Z(n4846) );
  ANDN U5079 ( .B(n4845), .A(n4836), .Z(n4900) );
  XOR U5080 ( .A(n4901), .B(n4902), .Z(n4855) );
  XOR U5081 ( .A(n4888), .B(n4878), .Z(n4902) );
  XOR U5082 ( .A(n4830), .B(n4578), .Z(n4878) );
  XOR U5083 ( .A(n4903), .B(n4890), .Z(n4888) );
  NANDN U5084 ( .A(n4840), .B(n4848), .Z(n4890) );
  XOR U5085 ( .A(n4856), .B(n4827), .Z(n4848) );
  XNOR U5086 ( .A(n4894), .B(n4904), .Z(n4845) );
  XNOR U5087 ( .A(n4905), .B(n4906), .Z(n4904) );
  XNOR U5088 ( .A(n4841), .B(n4627), .Z(n4840) );
  XNOR U5089 ( .A(n4836), .B(n4830), .Z(n4627) );
  IV U5090 ( .A(n4881), .Z(n4836) );
  XOR U5091 ( .A(n4907), .B(n4908), .Z(n4881) );
  XOR U5092 ( .A(n4909), .B(n4910), .Z(n4908) );
  XOR U5093 ( .A(n4898), .B(n4911), .Z(n4907) );
  AND U5094 ( .A(n4856), .B(n4841), .Z(n4903) );
  XOR U5095 ( .A(n4573), .B(n4621), .Z(n4841) );
  IV U5096 ( .A(n4898), .Z(n4573) );
  XOR U5097 ( .A(n4887), .B(n4912), .Z(n4901) );
  XNOR U5098 ( .A(n4913), .B(n4893), .Z(n4912) );
  OR U5099 ( .A(n4580), .B(n4831), .Z(n4893) );
  XNOR U5100 ( .A(n4914), .B(n4830), .Z(n4831) );
  XNOR U5101 ( .A(n4504), .B(n4578), .Z(n4580) );
  ANDN U5102 ( .B(n4830), .A(n4578), .Z(n4913) );
  XOR U5103 ( .A(n4915), .B(n4916), .Z(n4578) );
  XOR U5104 ( .A(n4905), .B(n4917), .Z(n4916) );
  XOR U5105 ( .A(n4918), .B(n4915), .Z(n4830) );
  XNOR U5106 ( .A(n4621), .B(n4504), .Z(n4887) );
  IV U5107 ( .A(n4914), .Z(n4621) );
  XNOR U5108 ( .A(n4906), .B(n4919), .Z(n4914) );
  XOR U5109 ( .A(n4911), .B(n4917), .Z(n4919) );
  IV U5110 ( .A(n4918), .Z(n4917) );
  XOR U5111 ( .A(n4920), .B(n4921), .Z(n4911) );
  XNOR U5112 ( .A(n3773), .B(n4922), .Z(n4921) );
  XOR U5113 ( .A(n4905), .B(n4923), .Z(n4922) );
  XOR U5114 ( .A(n4924), .B(n4925), .Z(n4905) );
  XOR U5115 ( .A(n2581), .B(n4926), .Z(n2563) );
  XNOR U5116 ( .A(key[417]), .B(n4927), .Z(n4924) );
  IV U5117 ( .A(n4928), .Z(n3773) );
  XNOR U5118 ( .A(n4929), .B(n4930), .Z(n4920) );
  XNOR U5119 ( .A(key[419]), .B(n2584), .Z(n4930) );
  XOR U5120 ( .A(n4931), .B(n3802), .Z(n2584) );
  XOR U5121 ( .A(n4932), .B(n4933), .Z(n4906) );
  XNOR U5122 ( .A(n2574), .B(n3813), .Z(n4933) );
  IV U5123 ( .A(n3815), .Z(n2574) );
  XOR U5124 ( .A(n4929), .B(n2559), .Z(n3815) );
  XOR U5125 ( .A(key[418]), .B(n4926), .Z(n4932) );
  XOR U5126 ( .A(n4894), .B(n4823), .Z(n4856) );
  XNOR U5127 ( .A(n4915), .B(n4934), .Z(n4823) );
  XOR U5128 ( .A(n4918), .B(n4910), .Z(n4934) );
  XNOR U5129 ( .A(n4935), .B(n4936), .Z(n4910) );
  XNOR U5130 ( .A(n4937), .B(n4938), .Z(n4936) );
  XNOR U5131 ( .A(n2540), .B(n4939), .Z(n4935) );
  XOR U5132 ( .A(key[420]), .B(n3803), .Z(n4939) );
  XOR U5133 ( .A(n4931), .B(n3787), .Z(n2540) );
  IV U5134 ( .A(n4504), .Z(n4894) );
  XOR U5135 ( .A(n4915), .B(n4940), .Z(n4504) );
  XNOR U5136 ( .A(n4918), .B(n4909), .Z(n4940) );
  XOR U5137 ( .A(n4941), .B(n4942), .Z(n4909) );
  XNOR U5138 ( .A(n4943), .B(n4944), .Z(n4942) );
  XNOR U5139 ( .A(key[423]), .B(n2587), .Z(n4941) );
  XOR U5140 ( .A(n4945), .B(n4946), .Z(n4918) );
  XNOR U5141 ( .A(n4947), .B(n4948), .Z(n4946) );
  XNOR U5142 ( .A(n2569), .B(n4949), .Z(n4945) );
  XNOR U5143 ( .A(key[422]), .B(n4898), .Z(n4949) );
  XOR U5144 ( .A(n4950), .B(n4951), .Z(n4898) );
  XOR U5145 ( .A(n3794), .B(n2589), .Z(n4951) );
  IV U5146 ( .A(n3806), .Z(n3794) );
  XNOR U5147 ( .A(key[416]), .B(n2580), .Z(n4950) );
  IV U5148 ( .A(n3814), .Z(n2580) );
  XOR U5149 ( .A(n4927), .B(n2591), .Z(n3814) );
  XOR U5150 ( .A(n4931), .B(n3796), .Z(n2569) );
  IV U5151 ( .A(n2587), .Z(n4931) );
  XNOR U5152 ( .A(n4952), .B(n4953), .Z(n4915) );
  XNOR U5153 ( .A(n4954), .B(n3782), .Z(n4953) );
  XOR U5154 ( .A(n4948), .B(n4955), .Z(n3782) );
  XNOR U5155 ( .A(key[421]), .B(n3788), .Z(n4952) );
  IV U5156 ( .A(n1827), .Z(n4629) );
  XNOR U5157 ( .A(n4516), .B(n4956), .Z(n1827) );
  XOR U5158 ( .A(n4615), .B(n4616), .Z(n4956) );
  XOR U5159 ( .A(n4608), .B(n4957), .Z(n4616) );
  XNOR U5160 ( .A(n4958), .B(n4959), .Z(n4957) );
  OR U5161 ( .A(n4557), .B(n4960), .Z(n4959) );
  XNOR U5162 ( .A(n4559), .B(n4961), .Z(n4608) );
  XNOR U5163 ( .A(n4962), .B(n4963), .Z(n4961) );
  NAND U5164 ( .A(n4964), .B(n4693), .Z(n4963) );
  IV U5165 ( .A(n4682), .Z(n4615) );
  XOR U5166 ( .A(n4689), .B(n4965), .Z(n4682) );
  XNOR U5167 ( .A(n4687), .B(n4966), .Z(n4965) );
  NAND U5168 ( .A(n4967), .B(n4563), .Z(n4966) );
  XOR U5169 ( .A(n4613), .B(n4563), .Z(n4611) );
  XOR U5170 ( .A(n4683), .B(n4607), .Z(n4516) );
  XNOR U5171 ( .A(n4559), .B(n4969), .Z(n4607) );
  XNOR U5172 ( .A(n4958), .B(n4970), .Z(n4969) );
  NANDN U5173 ( .A(n4971), .B(n4972), .Z(n4970) );
  OR U5174 ( .A(n4973), .B(n4974), .Z(n4958) );
  XOR U5175 ( .A(n4975), .B(n4962), .Z(n4559) );
  NANDN U5176 ( .A(n4976), .B(n4977), .Z(n4962) );
  ANDN U5177 ( .B(n4978), .A(n4979), .Z(n4975) );
  XOR U5178 ( .A(n4689), .B(n4980), .Z(n4683) );
  XOR U5179 ( .A(n4981), .B(n4555), .Z(n4980) );
  OR U5180 ( .A(n4982), .B(n4973), .Z(n4555) );
  XNOR U5181 ( .A(n4557), .B(n4971), .Z(n4973) );
  NOR U5182 ( .A(n4983), .B(n4971), .Z(n4981) );
  XOR U5183 ( .A(n4984), .B(n4691), .Z(n4689) );
  OR U5184 ( .A(n4976), .B(n4985), .Z(n4691) );
  XNOR U5185 ( .A(n4986), .B(n4693), .Z(n4976) );
  XNOR U5186 ( .A(n4971), .B(n4563), .Z(n4693) );
  XOR U5187 ( .A(n4987), .B(n4988), .Z(n4563) );
  NANDN U5188 ( .A(n4989), .B(n4990), .Z(n4988) );
  XNOR U5189 ( .A(n4991), .B(n4992), .Z(n4971) );
  OR U5190 ( .A(n4989), .B(n4993), .Z(n4992) );
  ANDN U5191 ( .B(n4986), .A(n4994), .Z(n4984) );
  IV U5192 ( .A(n4979), .Z(n4986) );
  XOR U5193 ( .A(n4557), .B(n4613), .Z(n4979) );
  XNOR U5194 ( .A(n4995), .B(n4987), .Z(n4613) );
  NANDN U5195 ( .A(n4996), .B(n4997), .Z(n4987) );
  ANDN U5196 ( .B(n4998), .A(n4999), .Z(n4995) );
  NANDN U5197 ( .A(n4996), .B(n5001), .Z(n4991) );
  XOR U5198 ( .A(n5002), .B(n4989), .Z(n4996) );
  XNOR U5199 ( .A(n5003), .B(n5004), .Z(n4989) );
  XOR U5200 ( .A(n5005), .B(n4998), .Z(n5004) );
  XNOR U5201 ( .A(n5006), .B(n5007), .Z(n5003) );
  XNOR U5202 ( .A(n5008), .B(n5009), .Z(n5007) );
  ANDN U5203 ( .B(n4998), .A(n5010), .Z(n5008) );
  IV U5204 ( .A(n5011), .Z(n4998) );
  ANDN U5205 ( .B(n5002), .A(n5010), .Z(n5000) );
  IV U5206 ( .A(n5006), .Z(n5010) );
  IV U5207 ( .A(n4999), .Z(n5002) );
  XNOR U5208 ( .A(n5005), .B(n5012), .Z(n4999) );
  XOR U5209 ( .A(n5013), .B(n5009), .Z(n5012) );
  NAND U5210 ( .A(n5001), .B(n4997), .Z(n5009) );
  XNOR U5211 ( .A(n4990), .B(n5011), .Z(n4997) );
  XOR U5212 ( .A(n5014), .B(n5015), .Z(n5011) );
  XOR U5213 ( .A(n5016), .B(n5017), .Z(n5015) );
  XNOR U5214 ( .A(n4972), .B(n5018), .Z(n5017) );
  XNOR U5215 ( .A(n5019), .B(n5020), .Z(n5014) );
  XNOR U5216 ( .A(n5021), .B(n5022), .Z(n5020) );
  ANDN U5217 ( .B(n5023), .A(n4558), .Z(n5021) );
  XNOR U5218 ( .A(n5006), .B(n4993), .Z(n5001) );
  XOR U5219 ( .A(n5024), .B(n5025), .Z(n5006) );
  XNOR U5220 ( .A(n5026), .B(n5018), .Z(n5025) );
  XOR U5221 ( .A(n5027), .B(n5028), .Z(n5018) );
  XNOR U5222 ( .A(n5029), .B(n5030), .Z(n5028) );
  NAND U5223 ( .A(n4694), .B(n4964), .Z(n5030) );
  XNOR U5224 ( .A(n5031), .B(n5032), .Z(n5024) );
  ANDN U5225 ( .B(n5033), .A(n4688), .Z(n5031) );
  ANDN U5226 ( .B(n4990), .A(n4993), .Z(n5013) );
  XOR U5227 ( .A(n4993), .B(n4990), .Z(n5005) );
  XNOR U5228 ( .A(n5034), .B(n5035), .Z(n4990) );
  XNOR U5229 ( .A(n5027), .B(n5036), .Z(n5035) );
  XOR U5230 ( .A(n5026), .B(n4960), .Z(n5036) );
  XOR U5231 ( .A(n4558), .B(n5037), .Z(n5034) );
  XNOR U5232 ( .A(n5038), .B(n5022), .Z(n5037) );
  OR U5233 ( .A(n4974), .B(n4982), .Z(n5022) );
  XNOR U5234 ( .A(n4558), .B(n4983), .Z(n4982) );
  XOR U5235 ( .A(n4960), .B(n4972), .Z(n4974) );
  ANDN U5236 ( .B(n4972), .A(n4983), .Z(n5038) );
  XOR U5237 ( .A(n5039), .B(n5040), .Z(n4993) );
  XOR U5238 ( .A(n5027), .B(n5016), .Z(n5040) );
  XOR U5239 ( .A(n4967), .B(n4564), .Z(n5016) );
  XOR U5240 ( .A(n5041), .B(n5029), .Z(n5027) );
  NANDN U5241 ( .A(n4985), .B(n4977), .Z(n5029) );
  XOR U5242 ( .A(n4978), .B(n4964), .Z(n4977) );
  XNOR U5243 ( .A(n5033), .B(n5042), .Z(n4972) );
  XNOR U5244 ( .A(n5043), .B(n5044), .Z(n5042) );
  XOR U5245 ( .A(n4994), .B(n4694), .Z(n4985) );
  XNOR U5246 ( .A(n4983), .B(n4967), .Z(n4694) );
  IV U5247 ( .A(n5019), .Z(n4983) );
  XOR U5248 ( .A(n5045), .B(n5046), .Z(n5019) );
  XOR U5249 ( .A(n5047), .B(n5048), .Z(n5046) );
  XNOR U5250 ( .A(n4558), .B(n5049), .Z(n5045) );
  ANDN U5251 ( .B(n4978), .A(n4994), .Z(n5041) );
  XNOR U5252 ( .A(n4558), .B(n4688), .Z(n4994) );
  XOR U5253 ( .A(n5033), .B(n5023), .Z(n4978) );
  IV U5254 ( .A(n4960), .Z(n5023) );
  XOR U5255 ( .A(n5050), .B(n5051), .Z(n4960) );
  XOR U5256 ( .A(n5052), .B(n5048), .Z(n5051) );
  XNOR U5257 ( .A(n5053), .B(n5054), .Z(n5048) );
  XNOR U5258 ( .A(n3647), .B(n2706), .Z(n5054) );
  XOR U5259 ( .A(n3604), .B(n5055), .Z(n2706) );
  XNOR U5260 ( .A(n5056), .B(n5057), .Z(n5053) );
  XNOR U5261 ( .A(key[412]), .B(n2708), .Z(n5057) );
  XOR U5262 ( .A(n5058), .B(n2696), .Z(n2708) );
  IV U5263 ( .A(n4614), .Z(n5033) );
  XOR U5264 ( .A(n5026), .B(n5059), .Z(n5039) );
  XNOR U5265 ( .A(n5060), .B(n5032), .Z(n5059) );
  OR U5266 ( .A(n4612), .B(n4968), .Z(n5032) );
  XNOR U5267 ( .A(n5061), .B(n4967), .Z(n4968) );
  XNOR U5268 ( .A(n4614), .B(n4564), .Z(n4612) );
  ANDN U5269 ( .B(n4967), .A(n4564), .Z(n5060) );
  XOR U5270 ( .A(n5050), .B(n5062), .Z(n4564) );
  XOR U5271 ( .A(n5043), .B(n5063), .Z(n5062) );
  XOR U5272 ( .A(n5052), .B(n5050), .Z(n4967) );
  XNOR U5273 ( .A(n4688), .B(n4614), .Z(n5026) );
  XOR U5274 ( .A(n5050), .B(n5064), .Z(n4614) );
  XNOR U5275 ( .A(n5052), .B(n5047), .Z(n5064) );
  XOR U5276 ( .A(n5065), .B(n5066), .Z(n5047) );
  XNOR U5277 ( .A(n2726), .B(n3634), .Z(n5066) );
  XOR U5278 ( .A(n5067), .B(n5058), .Z(n2726) );
  XNOR U5279 ( .A(key[415]), .B(n2702), .Z(n5065) );
  XOR U5280 ( .A(n3613), .B(n5068), .Z(n2702) );
  XNOR U5281 ( .A(n5069), .B(n5070), .Z(n5050) );
  XNOR U5282 ( .A(n2689), .B(n3603), .Z(n5070) );
  XNOR U5283 ( .A(n2694), .B(n5071), .Z(n5069) );
  XNOR U5284 ( .A(key[413]), .B(n3633), .Z(n5071) );
  XNOR U5285 ( .A(n3618), .B(n5072), .Z(n2694) );
  IV U5286 ( .A(n5061), .Z(n4688) );
  XNOR U5287 ( .A(n5044), .B(n5073), .Z(n5061) );
  XOR U5288 ( .A(n5049), .B(n5063), .Z(n5073) );
  IV U5289 ( .A(n5052), .Z(n5063) );
  XOR U5290 ( .A(n5074), .B(n5075), .Z(n5052) );
  XNOR U5291 ( .A(n5076), .B(n2701), .Z(n2691) );
  XOR U5292 ( .A(n5058), .B(n5077), .Z(n2701) );
  XNOR U5293 ( .A(n5078), .B(n5079), .Z(n5074) );
  XOR U5294 ( .A(key[414]), .B(n4558), .Z(n5079) );
  XNOR U5295 ( .A(n5080), .B(n5081), .Z(n4558) );
  XOR U5296 ( .A(n3644), .B(n2720), .Z(n5081) );
  XNOR U5297 ( .A(n3615), .B(n5082), .Z(n5080) );
  XOR U5298 ( .A(n5083), .B(n5084), .Z(n5049) );
  XOR U5299 ( .A(n2721), .B(n5085), .Z(n5084) );
  XOR U5300 ( .A(n5086), .B(n5087), .Z(n5043) );
  XOR U5301 ( .A(n2718), .B(n3629), .Z(n5087) );
  XNOR U5302 ( .A(n3653), .B(n5088), .Z(n5086) );
  XNOR U5303 ( .A(n5089), .B(n5090), .Z(n5083) );
  XNOR U5304 ( .A(key[411]), .B(n2723), .Z(n5090) );
  XOR U5305 ( .A(n5058), .B(n2710), .Z(n2723) );
  IV U5306 ( .A(n5091), .Z(n5058) );
  XOR U5307 ( .A(n5092), .B(n5093), .Z(n5044) );
  XOR U5308 ( .A(n2715), .B(n3641), .Z(n5093) );
  XNOR U5309 ( .A(n2679), .B(n5094), .Z(n5092) );
  XNOR U5310 ( .A(key[410]), .B(n3646), .Z(n5094) );
  XOR U5311 ( .A(n4548), .B(n4491), .Z(n1216) );
  XNOR U5312 ( .A(n4524), .B(n5095), .Z(n4491) );
  XOR U5313 ( .A(n5096), .B(n4638), .Z(n5095) );
  OR U5314 ( .A(n5097), .B(n4590), .Z(n4638) );
  XOR U5315 ( .A(n4593), .B(n4496), .Z(n4590) );
  NOR U5316 ( .A(n5098), .B(n4593), .Z(n5096) );
  XNOR U5317 ( .A(n4636), .B(n5099), .Z(n4524) );
  XNOR U5318 ( .A(n5100), .B(n5101), .Z(n5099) );
  NAND U5319 ( .A(n4650), .B(n5102), .Z(n5101) );
  XNOR U5320 ( .A(n4636), .B(n5103), .Z(n4548) );
  XOR U5321 ( .A(n5104), .B(n4526), .Z(n5103) );
  OR U5322 ( .A(n5105), .B(n4644), .Z(n4526) );
  XNOR U5323 ( .A(n4529), .B(n4635), .Z(n4644) );
  ANDN U5324 ( .B(n4635), .A(n5106), .Z(n5104) );
  XOR U5325 ( .A(n5107), .B(n5100), .Z(n4636) );
  OR U5326 ( .A(n4652), .B(n5108), .Z(n5100) );
  XNOR U5327 ( .A(n5109), .B(n4650), .Z(n4652) );
  XOR U5328 ( .A(n4496), .B(n4635), .Z(n4650) );
  XOR U5329 ( .A(n5110), .B(n5111), .Z(n4635) );
  NANDN U5330 ( .A(n5112), .B(n5113), .Z(n5111) );
  XOR U5331 ( .A(n5114), .B(n5115), .Z(n4496) );
  NANDN U5332 ( .A(n5112), .B(n5116), .Z(n5115) );
  ANDN U5333 ( .B(n5109), .A(n5117), .Z(n5107) );
  IV U5334 ( .A(n4655), .Z(n5109) );
  XOR U5335 ( .A(n4593), .B(n4529), .Z(n4655) );
  XNOR U5336 ( .A(n5118), .B(n5110), .Z(n4529) );
  NANDN U5337 ( .A(n5119), .B(n5120), .Z(n5110) );
  XOR U5338 ( .A(n5113), .B(n5121), .Z(n5120) );
  ANDN U5339 ( .B(n5121), .A(n5122), .Z(n5118) );
  NANDN U5340 ( .A(n5119), .B(n5124), .Z(n5114) );
  XOR U5341 ( .A(n5125), .B(n5116), .Z(n5124) );
  XNOR U5342 ( .A(n5126), .B(n5127), .Z(n5112) );
  XOR U5343 ( .A(n5128), .B(n5129), .Z(n5127) );
  XNOR U5344 ( .A(n5130), .B(n5131), .Z(n5126) );
  XNOR U5345 ( .A(n5132), .B(n5133), .Z(n5131) );
  ANDN U5346 ( .B(n5125), .A(n5129), .Z(n5132) );
  ANDN U5347 ( .B(n5125), .A(n5122), .Z(n5123) );
  XNOR U5348 ( .A(n5128), .B(n5134), .Z(n5122) );
  XOR U5349 ( .A(n5135), .B(n5133), .Z(n5134) );
  NAND U5350 ( .A(n5136), .B(n5137), .Z(n5133) );
  XNOR U5351 ( .A(n5130), .B(n5116), .Z(n5137) );
  IV U5352 ( .A(n5125), .Z(n5130) );
  XNOR U5353 ( .A(n5113), .B(n5129), .Z(n5136) );
  IV U5354 ( .A(n5121), .Z(n5129) );
  XOR U5355 ( .A(n5138), .B(n5139), .Z(n5121) );
  XNOR U5356 ( .A(n5140), .B(n5141), .Z(n5139) );
  XNOR U5357 ( .A(n5142), .B(n5143), .Z(n5138) );
  ANDN U5358 ( .B(n5144), .A(n5098), .Z(n5142) );
  AND U5359 ( .A(n5116), .B(n5113), .Z(n5135) );
  XNOR U5360 ( .A(n5116), .B(n5113), .Z(n5128) );
  XNOR U5361 ( .A(n5145), .B(n5146), .Z(n5113) );
  XOR U5362 ( .A(n5147), .B(n5141), .Z(n5146) );
  XNOR U5363 ( .A(n5148), .B(n5149), .Z(n5145) );
  XNOR U5364 ( .A(n5150), .B(n5143), .Z(n5149) );
  OR U5365 ( .A(n4591), .B(n5097), .Z(n5143) );
  XNOR U5366 ( .A(n5151), .B(n4640), .Z(n5097) );
  XNOR U5367 ( .A(n4497), .B(n4592), .Z(n4591) );
  ANDN U5368 ( .B(n4640), .A(n4497), .Z(n5150) );
  XNOR U5369 ( .A(n5152), .B(n5153), .Z(n5116) );
  XNOR U5370 ( .A(n5141), .B(n5154), .Z(n5153) );
  XOR U5371 ( .A(n4643), .B(n5147), .Z(n5154) );
  XNOR U5372 ( .A(n5151), .B(n4592), .Z(n5141) );
  XOR U5373 ( .A(n4528), .B(n5155), .Z(n5152) );
  XNOR U5374 ( .A(n5156), .B(n5157), .Z(n5155) );
  XNOR U5375 ( .A(n5158), .B(n5159), .Z(n5125) );
  XNOR U5376 ( .A(n5140), .B(n5160), .Z(n5159) );
  XNOR U5377 ( .A(n5148), .B(n4634), .Z(n5160) );
  XOR U5378 ( .A(n4640), .B(n5161), .Z(n5148) );
  XOR U5379 ( .A(n5147), .B(n5162), .Z(n5140) );
  XNOR U5380 ( .A(n5163), .B(n5164), .Z(n5162) );
  NAND U5381 ( .A(n5102), .B(n4649), .Z(n5164) );
  XNOR U5382 ( .A(n5165), .B(n5163), .Z(n5147) );
  NANDN U5383 ( .A(n5108), .B(n4653), .Z(n5163) );
  XOR U5384 ( .A(n4654), .B(n4649), .Z(n4653) );
  XNOR U5385 ( .A(n5161), .B(n4634), .Z(n4649) );
  IV U5386 ( .A(n4497), .Z(n5161) );
  XOR U5387 ( .A(n5166), .B(n5167), .Z(n4497) );
  XOR U5388 ( .A(n5168), .B(n5169), .Z(n5167) );
  XOR U5389 ( .A(n5117), .B(n5102), .Z(n5108) );
  XOR U5390 ( .A(n4640), .B(n5170), .Z(n5102) );
  ANDN U5391 ( .B(n4654), .A(n5117), .Z(n5165) );
  XOR U5392 ( .A(n4528), .B(n5151), .Z(n5117) );
  IV U5393 ( .A(n5098), .Z(n5151) );
  XOR U5394 ( .A(n5171), .B(n5172), .Z(n5098) );
  XOR U5395 ( .A(n5173), .B(n5168), .Z(n5172) );
  XOR U5396 ( .A(n5174), .B(n5144), .Z(n4654) );
  XNOR U5397 ( .A(n5170), .B(n5175), .Z(n5158) );
  XNOR U5398 ( .A(n5176), .B(n5157), .Z(n5175) );
  OR U5399 ( .A(n4645), .B(n5105), .Z(n5157) );
  XNOR U5400 ( .A(n4528), .B(n5106), .Z(n5105) );
  IV U5401 ( .A(n5170), .Z(n5106) );
  XNOR U5402 ( .A(n4643), .B(n4634), .Z(n4645) );
  XOR U5403 ( .A(n5144), .B(n5177), .Z(n4634) );
  XNOR U5404 ( .A(n5173), .B(n5169), .Z(n5177) );
  XOR U5405 ( .A(n5178), .B(n5179), .Z(n5173) );
  XOR U5406 ( .A(n3047), .B(n3005), .Z(n5179) );
  IV U5407 ( .A(n5180), .Z(n3047) );
  XNOR U5408 ( .A(n5181), .B(n5182), .Z(n5178) );
  XNOR U5409 ( .A(key[458]), .B(n3981), .Z(n5182) );
  IV U5410 ( .A(n4592), .Z(n5144) );
  XNOR U5411 ( .A(n5183), .B(n4640), .Z(n4592) );
  NOR U5412 ( .A(n4643), .B(n4528), .Z(n5176) );
  IV U5413 ( .A(n5174), .Z(n4643) );
  XOR U5414 ( .A(n5184), .B(n4640), .Z(n5174) );
  XNOR U5415 ( .A(n5168), .B(n5166), .Z(n4640) );
  XNOR U5416 ( .A(n5185), .B(n5186), .Z(n5166) );
  XNOR U5417 ( .A(n3040), .B(n3968), .Z(n5186) );
  XNOR U5418 ( .A(n3026), .B(n5187), .Z(n5185) );
  XNOR U5419 ( .A(key[461]), .B(n3947), .Z(n5187) );
  XNOR U5420 ( .A(n5189), .B(n5190), .Z(n5168) );
  XNOR U5421 ( .A(n3956), .B(n3042), .Z(n5190) );
  XNOR U5422 ( .A(n5191), .B(n3029), .Z(n3042) );
  XOR U5423 ( .A(n5192), .B(n5193), .Z(n3029) );
  XNOR U5424 ( .A(n5194), .B(n5195), .Z(n5189) );
  XOR U5425 ( .A(key[462]), .B(n4528), .Z(n5195) );
  XOR U5426 ( .A(n5196), .B(n5197), .Z(n5170) );
  XNOR U5427 ( .A(n5184), .B(n5183), .Z(n5197) );
  XOR U5428 ( .A(n5198), .B(n5199), .Z(n5183) );
  XNOR U5429 ( .A(n3037), .B(n3949), .Z(n5199) );
  XOR U5430 ( .A(n5200), .B(n5192), .Z(n3037) );
  XNOR U5431 ( .A(key[463]), .B(n3030), .Z(n5198) );
  XNOR U5432 ( .A(n3961), .B(n5201), .Z(n3030) );
  XOR U5433 ( .A(n5202), .B(n5203), .Z(n5184) );
  XOR U5434 ( .A(n3979), .B(n3010), .Z(n5203) );
  XOR U5435 ( .A(n3967), .B(n5204), .Z(n3010) );
  XNOR U5436 ( .A(n5205), .B(n5206), .Z(n5202) );
  XNOR U5437 ( .A(key[460]), .B(n3012), .Z(n5206) );
  XNOR U5438 ( .A(n5207), .B(n3024), .Z(n3012) );
  XNOR U5439 ( .A(n4528), .B(n5171), .Z(n5196) );
  XOR U5440 ( .A(n5208), .B(n5209), .Z(n5171) );
  XNOR U5441 ( .A(n3002), .B(n5210), .Z(n5209) );
  XOR U5442 ( .A(n3936), .B(n3003), .Z(n5210) );
  XOR U5443 ( .A(n5192), .B(n3014), .Z(n3003) );
  IV U5444 ( .A(n5211), .Z(n3002) );
  XNOR U5445 ( .A(n5169), .B(n5212), .Z(n5208) );
  XNOR U5446 ( .A(key[459]), .B(n5213), .Z(n5212) );
  XOR U5447 ( .A(n5214), .B(n5215), .Z(n5169) );
  XNOR U5448 ( .A(n3045), .B(n3985), .Z(n5215) );
  XNOR U5449 ( .A(n3018), .B(n5216), .Z(n5214) );
  XNOR U5450 ( .A(key[457]), .B(n3938), .Z(n5216) );
  IV U5451 ( .A(n5217), .Z(n3938) );
  XNOR U5452 ( .A(n5218), .B(n5219), .Z(n4528) );
  XOR U5453 ( .A(n5200), .B(n3020), .Z(n5219) );
  XNOR U5454 ( .A(n3978), .B(n5220), .Z(n5218) );
  XNOR U5455 ( .A(key[456]), .B(n3963), .Z(n5220) );
  XNOR U5456 ( .A(n854), .B(n5221), .Z(out[0]) );
  XOR U5457 ( .A(key[512]), .B(n1651), .Z(n5221) );
  XNOR U5458 ( .A(n1876), .B(n5222), .Z(n1651) );
  XOR U5459 ( .A(n5223), .B(n858), .Z(n5222) );
  OR U5460 ( .A(n5224), .B(n1869), .Z(n858) );
  XNOR U5461 ( .A(n861), .B(n1868), .Z(n1869) );
  ANDN U5462 ( .B(n5225), .A(n5226), .Z(n5223) );
  IV U5463 ( .A(n1084), .Z(n854) );
  XOR U5464 ( .A(n862), .B(n5227), .Z(n1084) );
  XOR U5465 ( .A(n5228), .B(n1878), .Z(n5227) );
  XNOR U5466 ( .A(n1445), .B(n866), .Z(n1442) );
  NOR U5467 ( .A(n5230), .B(n1445), .Z(n5228) );
  XNOR U5468 ( .A(n1876), .B(n5231), .Z(n862) );
  XNOR U5469 ( .A(n5232), .B(n5233), .Z(n5231) );
  NANDN U5470 ( .A(n1863), .B(n5234), .Z(n5233) );
  XOR U5471 ( .A(n5235), .B(n5232), .Z(n1876) );
  OR U5472 ( .A(n1872), .B(n5236), .Z(n5232) );
  XOR U5473 ( .A(n5237), .B(n1863), .Z(n1872) );
  XNOR U5474 ( .A(n1868), .B(n866), .Z(n1863) );
  XOR U5475 ( .A(n5238), .B(n5239), .Z(n866) );
  NANDN U5476 ( .A(n5240), .B(n5241), .Z(n5239) );
  IV U5477 ( .A(n5226), .Z(n1868) );
  XNOR U5478 ( .A(n5242), .B(n5243), .Z(n5226) );
  NANDN U5479 ( .A(n5240), .B(n5244), .Z(n5243) );
  ANDN U5480 ( .B(n5237), .A(n5245), .Z(n5235) );
  IV U5481 ( .A(n1875), .Z(n5237) );
  XOR U5482 ( .A(n1445), .B(n861), .Z(n1875) );
  XNOR U5483 ( .A(n5246), .B(n5242), .Z(n861) );
  NANDN U5484 ( .A(n5247), .B(n5248), .Z(n5242) );
  XOR U5485 ( .A(n5244), .B(n5249), .Z(n5248) );
  ANDN U5486 ( .B(n5249), .A(n5250), .Z(n5246) );
  XOR U5487 ( .A(n5251), .B(n5238), .Z(n1445) );
  NANDN U5488 ( .A(n5247), .B(n5252), .Z(n5238) );
  XOR U5489 ( .A(n5253), .B(n5241), .Z(n5252) );
  XNOR U5490 ( .A(n5254), .B(n5255), .Z(n5240) );
  XOR U5491 ( .A(n5256), .B(n5257), .Z(n5255) );
  XNOR U5492 ( .A(n5258), .B(n5259), .Z(n5254) );
  XNOR U5493 ( .A(n5260), .B(n5261), .Z(n5259) );
  ANDN U5494 ( .B(n5253), .A(n5257), .Z(n5260) );
  ANDN U5495 ( .B(n5253), .A(n5250), .Z(n5251) );
  XNOR U5496 ( .A(n5256), .B(n5262), .Z(n5250) );
  XOR U5497 ( .A(n5263), .B(n5261), .Z(n5262) );
  NAND U5498 ( .A(n5264), .B(n5265), .Z(n5261) );
  XNOR U5499 ( .A(n5258), .B(n5241), .Z(n5265) );
  IV U5500 ( .A(n5253), .Z(n5258) );
  XNOR U5501 ( .A(n5244), .B(n5257), .Z(n5264) );
  IV U5502 ( .A(n5249), .Z(n5257) );
  XOR U5503 ( .A(n5266), .B(n5267), .Z(n5249) );
  XNOR U5504 ( .A(n5268), .B(n5269), .Z(n5267) );
  XNOR U5505 ( .A(n5270), .B(n5271), .Z(n5266) );
  ANDN U5506 ( .B(n5272), .A(n5230), .Z(n5270) );
  AND U5507 ( .A(n5241), .B(n5244), .Z(n5263) );
  XNOR U5508 ( .A(n5241), .B(n5244), .Z(n5256) );
  XNOR U5509 ( .A(n5273), .B(n5274), .Z(n5244) );
  XNOR U5510 ( .A(n5275), .B(n5269), .Z(n5274) );
  XOR U5511 ( .A(n5276), .B(n5277), .Z(n5273) );
  XNOR U5512 ( .A(n5278), .B(n5271), .Z(n5277) );
  OR U5513 ( .A(n1443), .B(n5229), .Z(n5271) );
  XNOR U5514 ( .A(n5279), .B(n1880), .Z(n5229) );
  XNOR U5515 ( .A(n1444), .B(n867), .Z(n1443) );
  ANDN U5516 ( .B(n1880), .A(n867), .Z(n5278) );
  XNOR U5517 ( .A(n5280), .B(n5281), .Z(n5241) );
  XNOR U5518 ( .A(n5269), .B(n5282), .Z(n5281) );
  XOR U5519 ( .A(n1859), .B(n5276), .Z(n5282) );
  XNOR U5520 ( .A(n5279), .B(n1444), .Z(n5269) );
  XNOR U5521 ( .A(n5283), .B(n5284), .Z(n5280) );
  XNOR U5522 ( .A(n5285), .B(n5286), .Z(n5284) );
  ANDN U5523 ( .B(n5225), .A(n1867), .Z(n5285) );
  XNOR U5524 ( .A(n5287), .B(n5288), .Z(n5253) );
  XNOR U5525 ( .A(n5275), .B(n5289), .Z(n5288) );
  XNOR U5526 ( .A(n1867), .B(n5268), .Z(n5289) );
  XOR U5527 ( .A(n5276), .B(n5290), .Z(n5268) );
  XNOR U5528 ( .A(n5291), .B(n5292), .Z(n5290) );
  NAND U5529 ( .A(n5234), .B(n1864), .Z(n5292) );
  XNOR U5530 ( .A(n5293), .B(n5291), .Z(n5276) );
  NANDN U5531 ( .A(n5236), .B(n1873), .Z(n5291) );
  XOR U5532 ( .A(n1874), .B(n1864), .Z(n1873) );
  XNOR U5533 ( .A(n5294), .B(n867), .Z(n1864) );
  XOR U5534 ( .A(n5245), .B(n5234), .Z(n5236) );
  XOR U5535 ( .A(n5225), .B(n1880), .Z(n5234) );
  ANDN U5536 ( .B(n1874), .A(n5245), .Z(n5293) );
  XNOR U5537 ( .A(n5283), .B(n5279), .Z(n5245) );
  IV U5538 ( .A(n5230), .Z(n5279) );
  XNOR U5539 ( .A(n5295), .B(n5296), .Z(n5230) );
  XOR U5540 ( .A(n5297), .B(n5298), .Z(n5296) );
  XOR U5541 ( .A(n5299), .B(n5272), .Z(n1874) );
  XNOR U5542 ( .A(n5300), .B(n5301), .Z(n867) );
  XNOR U5543 ( .A(n5302), .B(n5298), .Z(n5301) );
  XNOR U5544 ( .A(n5298), .B(n5300), .Z(n1880) );
  XNOR U5545 ( .A(n5225), .B(n5303), .Z(n5287) );
  XNOR U5546 ( .A(n5304), .B(n5286), .Z(n5303) );
  OR U5547 ( .A(n1870), .B(n5224), .Z(n5286) );
  XNOR U5548 ( .A(n5283), .B(n5225), .Z(n5224) );
  XOR U5549 ( .A(n1859), .B(n5294), .Z(n1870) );
  IV U5550 ( .A(n1867), .Z(n5294) );
  XOR U5551 ( .A(n5272), .B(n5305), .Z(n1867) );
  XOR U5552 ( .A(n5302), .B(n5295), .Z(n5305) );
  XNOR U5553 ( .A(key[546]), .B(\w0[4][34] ), .Z(n5295) );
  XOR U5554 ( .A(n4324), .B(n5306), .Z(\w0[4][34] ) );
  XNOR U5555 ( .A(n1035), .B(n995), .Z(n5306) );
  XOR U5556 ( .A(n1036), .B(n379), .Z(n995) );
  XOR U5557 ( .A(n1029), .B(n994), .Z(n4324) );
  XNOR U5558 ( .A(n5307), .B(n5308), .Z(n1029) );
  XNOR U5559 ( .A(n5309), .B(n5310), .Z(n5308) );
  XNOR U5560 ( .A(n5311), .B(n5312), .Z(n5307) );
  IV U5561 ( .A(n1444), .Z(n5272) );
  XNOR U5562 ( .A(n5300), .B(n5313), .Z(n1444) );
  XNOR U5563 ( .A(n5298), .B(n5314), .Z(n5313) );
  ANDN U5564 ( .B(n5299), .A(n860), .Z(n5304) );
  IV U5565 ( .A(n1859), .Z(n5299) );
  XNOR U5566 ( .A(n5300), .B(n5315), .Z(n1859) );
  XNOR U5567 ( .A(n5298), .B(n5316), .Z(n5315) );
  XOR U5568 ( .A(n860), .B(n5317), .Z(n5298) );
  XOR U5569 ( .A(key[550]), .B(\w0[4][38] ), .Z(n5317) );
  XNOR U5570 ( .A(n4300), .B(n5318), .Z(\w0[4][38] ) );
  XOR U5571 ( .A(n1004), .B(n1010), .Z(n5318) );
  XNOR U5572 ( .A(n392), .B(n5319), .Z(n1004) );
  XOR U5573 ( .A(n1011), .B(n4308), .Z(n392) );
  IV U5574 ( .A(n388), .Z(n4308) );
  XOR U5575 ( .A(n5320), .B(n5321), .Z(n388) );
  XOR U5576 ( .A(n5322), .B(n5323), .Z(n1011) );
  XNOR U5577 ( .A(n1017), .B(n5324), .Z(n4300) );
  XOR U5578 ( .A(n5325), .B(n5326), .Z(n1017) );
  XNOR U5579 ( .A(n5327), .B(n5309), .Z(n5326) );
  IV U5580 ( .A(n5283), .Z(n860) );
  XOR U5581 ( .A(key[549]), .B(\w0[4][37] ), .Z(n5300) );
  XOR U5582 ( .A(n4302), .B(n5329), .Z(\w0[4][37] ) );
  XOR U5583 ( .A(n1012), .B(n4307), .Z(n5329) );
  XNOR U5584 ( .A(n1024), .B(n393), .Z(n1012) );
  XNOR U5585 ( .A(n5330), .B(n5331), .Z(n393) );
  XNOR U5586 ( .A(n5332), .B(n5333), .Z(n5331) );
  XOR U5587 ( .A(n5334), .B(n5335), .Z(n5330) );
  XOR U5588 ( .A(n5336), .B(n5337), .Z(n5335) );
  ANDN U5589 ( .B(n5338), .A(n5339), .Z(n5337) );
  XNOR U5590 ( .A(n5340), .B(n5341), .Z(n1024) );
  XOR U5591 ( .A(n5342), .B(n5343), .Z(n5341) );
  XNOR U5592 ( .A(n5344), .B(n5345), .Z(n5340) );
  XOR U5593 ( .A(n5346), .B(n5347), .Z(n5345) );
  ANDN U5594 ( .B(n5348), .A(n5349), .Z(n5347) );
  XOR U5595 ( .A(n4309), .B(n1010), .Z(n4302) );
  XOR U5596 ( .A(n5350), .B(n5351), .Z(n1010) );
  XOR U5597 ( .A(n5327), .B(n5310), .Z(n4309) );
  XOR U5598 ( .A(n5352), .B(n5353), .Z(n5310) );
  XNOR U5599 ( .A(n5354), .B(n5355), .Z(n5353) );
  NOR U5600 ( .A(n5356), .B(n5357), .Z(n5354) );
  XOR U5601 ( .A(n5358), .B(n5359), .Z(n5225) );
  XNOR U5602 ( .A(n5316), .B(n5314), .Z(n5359) );
  XOR U5603 ( .A(key[551]), .B(\w0[4][39] ), .Z(n5314) );
  XNOR U5604 ( .A(n5324), .B(n5360), .Z(\w0[4][39] ) );
  XNOR U5605 ( .A(n1018), .B(n5319), .Z(n5360) );
  XNOR U5606 ( .A(n419), .B(n4315), .Z(n5319) );
  XNOR U5607 ( .A(n5361), .B(n5362), .Z(n4315) );
  XNOR U5608 ( .A(n5364), .B(n5365), .Z(n5361) );
  IV U5609 ( .A(n5366), .Z(n419) );
  XNOR U5610 ( .A(n1006), .B(n4303), .Z(n1018) );
  XOR U5611 ( .A(n5367), .B(n5368), .Z(n4303) );
  XOR U5612 ( .A(n5369), .B(n5320), .Z(n5368) );
  XNOR U5613 ( .A(n5372), .B(n5373), .Z(n5371) );
  NANDN U5614 ( .A(n5374), .B(n5375), .Z(n5373) );
  XOR U5615 ( .A(n5377), .B(n5378), .Z(n1006) );
  XOR U5616 ( .A(n5379), .B(n5322), .Z(n5378) );
  XNOR U5617 ( .A(n5381), .B(n5382), .Z(n5344) );
  XNOR U5618 ( .A(n5383), .B(n5384), .Z(n5382) );
  NANDN U5619 ( .A(n5385), .B(n5386), .Z(n5384) );
  XOR U5620 ( .A(key[548]), .B(\w0[4][36] ), .Z(n5316) );
  XOR U5621 ( .A(n5387), .B(n5388), .Z(\w0[4][36] ) );
  XNOR U5622 ( .A(n4319), .B(n4318), .Z(n5388) );
  XNOR U5623 ( .A(n1009), .B(n4313), .Z(n4318) );
  XOR U5624 ( .A(n5389), .B(n5390), .Z(n1009) );
  XNOR U5625 ( .A(n5391), .B(n5392), .Z(n5390) );
  XOR U5626 ( .A(n5328), .B(n5393), .Z(n5389) );
  XOR U5627 ( .A(n5355), .B(n5394), .Z(n5393) );
  ANDN U5628 ( .B(n5395), .A(n5396), .Z(n5394) );
  ANDN U5629 ( .B(n5397), .A(n5398), .Z(n5355) );
  XNOR U5630 ( .A(n5400), .B(n5401), .Z(n5399) );
  NANDN U5631 ( .A(n5402), .B(n5403), .Z(n5401) );
  XOR U5632 ( .A(n1023), .B(n1022), .Z(n5387) );
  XOR U5633 ( .A(n5333), .B(n379), .Z(n405) );
  XOR U5634 ( .A(n5370), .B(n5405), .Z(n379) );
  XNOR U5635 ( .A(n5343), .B(n1036), .Z(n1031) );
  XNOR U5636 ( .A(n5380), .B(n5406), .Z(n1036) );
  XOR U5637 ( .A(n5366), .B(n4307), .Z(n1023) );
  XNOR U5638 ( .A(n5407), .B(n5408), .Z(n4307) );
  XNOR U5639 ( .A(n5364), .B(n5409), .Z(n5408) );
  XNOR U5640 ( .A(n5410), .B(n5411), .Z(n5364) );
  XNOR U5641 ( .A(n5412), .B(n5413), .Z(n5411) );
  NANDN U5642 ( .A(n5414), .B(n5415), .Z(n5413) );
  XNOR U5643 ( .A(n5416), .B(n5417), .Z(n5407) );
  XOR U5644 ( .A(n5418), .B(n5419), .Z(n5417) );
  ANDN U5645 ( .B(n5420), .A(n5421), .Z(n5419) );
  XNOR U5646 ( .A(n5283), .B(n5297), .Z(n5358) );
  XOR U5647 ( .A(n5302), .B(n5422), .Z(n5297) );
  XOR U5648 ( .A(key[547]), .B(\w0[4][35] ), .Z(n5422) );
  XOR U5649 ( .A(n5423), .B(n5424), .Z(\w0[4][35] ) );
  XNOR U5650 ( .A(n994), .B(n4323), .Z(n5424) );
  XNOR U5651 ( .A(n1021), .B(n4313), .Z(n4323) );
  IV U5652 ( .A(n5324), .Z(n4313) );
  XOR U5653 ( .A(n5425), .B(n5392), .Z(n5324) );
  XOR U5654 ( .A(n5392), .B(n4327), .Z(n1021) );
  IV U5655 ( .A(n996), .Z(n4327) );
  XNOR U5656 ( .A(n5404), .B(n5426), .Z(n5392) );
  XOR U5657 ( .A(n5427), .B(n5428), .Z(n5426) );
  NOR U5658 ( .A(n5429), .B(n5357), .Z(n5427) );
  XNOR U5659 ( .A(n5430), .B(n5431), .Z(n5404) );
  XNOR U5660 ( .A(n5432), .B(n5433), .Z(n5431) );
  NANDN U5661 ( .A(n5434), .B(n5435), .Z(n5433) );
  XNOR U5662 ( .A(n5436), .B(n5437), .Z(n994) );
  XNOR U5663 ( .A(n5363), .B(n5351), .Z(n5437) );
  XOR U5664 ( .A(n5438), .B(n5439), .Z(n5351) );
  XNOR U5665 ( .A(n5440), .B(n5418), .Z(n5439) );
  ANDN U5666 ( .B(n5441), .A(n5442), .Z(n5418) );
  ANDN U5667 ( .B(n5443), .A(n5444), .Z(n5440) );
  XNOR U5668 ( .A(n5365), .B(n5445), .Z(n5436) );
  XOR U5669 ( .A(n1030), .B(n1028), .Z(n5423) );
  IV U5670 ( .A(n380), .Z(n1028) );
  XOR U5671 ( .A(n997), .B(n412), .Z(n380) );
  XOR U5672 ( .A(n5446), .B(n5447), .Z(n412) );
  XOR U5673 ( .A(n5448), .B(n5321), .Z(n5447) );
  XNOR U5674 ( .A(n5449), .B(n5450), .Z(n5321) );
  XNOR U5675 ( .A(n5451), .B(n5336), .Z(n5450) );
  ANDN U5676 ( .B(n5452), .A(n5453), .Z(n5336) );
  NOR U5677 ( .A(n5454), .B(n5455), .Z(n5451) );
  XOR U5678 ( .A(n5370), .B(n5369), .Z(n5446) );
  XOR U5679 ( .A(n5456), .B(n5457), .Z(n997) );
  XOR U5680 ( .A(n5458), .B(n5323), .Z(n5457) );
  XNOR U5681 ( .A(n5459), .B(n5460), .Z(n5323) );
  XNOR U5682 ( .A(n5461), .B(n5346), .Z(n5460) );
  ANDN U5683 ( .B(n5462), .A(n5463), .Z(n5346) );
  ANDN U5684 ( .B(n5464), .A(n5465), .Z(n5461) );
  XOR U5685 ( .A(n5380), .B(n5379), .Z(n5456) );
  XOR U5686 ( .A(n5366), .B(n4319), .Z(n1030) );
  XNOR U5687 ( .A(n5416), .B(n1035), .Z(n4319) );
  XOR U5688 ( .A(key[545]), .B(\w0[4][33] ), .Z(n5302) );
  XNOR U5689 ( .A(n377), .B(n5466), .Z(\w0[4][33] ) );
  XOR U5690 ( .A(n420), .B(n1039), .Z(n5466) );
  XNOR U5691 ( .A(n1040), .B(n416), .Z(n420) );
  XOR U5692 ( .A(n5320), .B(n5467), .Z(n416) );
  XNOR U5693 ( .A(n5370), .B(n5369), .Z(n5467) );
  XNOR U5694 ( .A(n5449), .B(n5468), .Z(n5369) );
  XNOR U5695 ( .A(n5469), .B(n5470), .Z(n5468) );
  NANDN U5696 ( .A(n5471), .B(n5375), .Z(n5470) );
  XOR U5697 ( .A(n5332), .B(n5472), .Z(n5449) );
  XNOR U5698 ( .A(n5473), .B(n5474), .Z(n5472) );
  NANDN U5699 ( .A(n5475), .B(n5476), .Z(n5474) );
  XOR U5700 ( .A(n5477), .B(n5478), .Z(n5370) );
  XNOR U5701 ( .A(n5479), .B(n5480), .Z(n5478) );
  NANDN U5702 ( .A(n5481), .B(n5338), .Z(n5480) );
  XOR U5703 ( .A(n5405), .B(n5448), .Z(n5320) );
  XNOR U5704 ( .A(n5332), .B(n5482), .Z(n5448) );
  XNOR U5705 ( .A(n5469), .B(n5483), .Z(n5482) );
  NANDN U5706 ( .A(n5484), .B(n5485), .Z(n5483) );
  OR U5707 ( .A(n5486), .B(n5487), .Z(n5469) );
  XOR U5708 ( .A(n5488), .B(n5473), .Z(n5332) );
  NANDN U5709 ( .A(n5489), .B(n5490), .Z(n5473) );
  ANDN U5710 ( .B(n5491), .A(n5492), .Z(n5488) );
  XNOR U5711 ( .A(n5322), .B(n5493), .Z(n1040) );
  XNOR U5712 ( .A(n5380), .B(n5379), .Z(n5493) );
  XNOR U5713 ( .A(n5459), .B(n5494), .Z(n5379) );
  XNOR U5714 ( .A(n5495), .B(n5496), .Z(n5494) );
  NANDN U5715 ( .A(n5497), .B(n5386), .Z(n5496) );
  XOR U5716 ( .A(n5342), .B(n5498), .Z(n5459) );
  XNOR U5717 ( .A(n5499), .B(n5500), .Z(n5498) );
  NANDN U5718 ( .A(n5501), .B(n5502), .Z(n5500) );
  XOR U5719 ( .A(n5503), .B(n5504), .Z(n5380) );
  XOR U5720 ( .A(n5505), .B(n5506), .Z(n5504) );
  NANDN U5721 ( .A(n5507), .B(n5348), .Z(n5506) );
  XOR U5722 ( .A(n5508), .B(n5458), .Z(n5322) );
  XNOR U5723 ( .A(n5342), .B(n5509), .Z(n5458) );
  XNOR U5724 ( .A(n5495), .B(n5510), .Z(n5509) );
  NANDN U5725 ( .A(n5511), .B(n5512), .Z(n5510) );
  OR U5726 ( .A(n5513), .B(n5514), .Z(n5495) );
  XOR U5727 ( .A(n5515), .B(n5499), .Z(n5342) );
  NANDN U5728 ( .A(n5516), .B(n5517), .Z(n5499) );
  ANDN U5729 ( .B(n5518), .A(n5519), .Z(n5515) );
  XOR U5730 ( .A(n996), .B(n1035), .Z(n377) );
  XNOR U5731 ( .A(n5520), .B(n5365), .Z(n1035) );
  XNOR U5732 ( .A(n5311), .B(n5425), .Z(n996) );
  XOR U5733 ( .A(key[544]), .B(\w0[4][32] ), .Z(n5283) );
  XNOR U5734 ( .A(n413), .B(n5521), .Z(\w0[4][32] ) );
  XNOR U5735 ( .A(n1015), .B(n4304), .Z(n5521) );
  XOR U5736 ( .A(n5405), .B(n5333), .Z(n4304) );
  XNOR U5737 ( .A(n5376), .B(n5522), .Z(n5333) );
  XOR U5738 ( .A(n5523), .B(n5479), .Z(n5522) );
  XNOR U5739 ( .A(n5455), .B(n5338), .Z(n5452) );
  NOR U5740 ( .A(n5525), .B(n5455), .Z(n5523) );
  XNOR U5741 ( .A(n5477), .B(n5526), .Z(n5376) );
  XNOR U5742 ( .A(n5527), .B(n5528), .Z(n5526) );
  NANDN U5743 ( .A(n5475), .B(n5529), .Z(n5528) );
  XOR U5744 ( .A(n5477), .B(n5530), .Z(n5405) );
  XOR U5745 ( .A(n5531), .B(n5372), .Z(n5530) );
  OR U5746 ( .A(n5532), .B(n5486), .Z(n5372) );
  XNOR U5747 ( .A(n5375), .B(n5485), .Z(n5486) );
  ANDN U5748 ( .B(n5533), .A(n5534), .Z(n5531) );
  XOR U5749 ( .A(n5535), .B(n5527), .Z(n5477) );
  OR U5750 ( .A(n5489), .B(n5536), .Z(n5527) );
  XOR U5751 ( .A(n5537), .B(n5475), .Z(n5489) );
  XNOR U5752 ( .A(n5485), .B(n5338), .Z(n5475) );
  XOR U5753 ( .A(n5538), .B(n5539), .Z(n5338) );
  NANDN U5754 ( .A(n5540), .B(n5541), .Z(n5539) );
  IV U5755 ( .A(n5534), .Z(n5485) );
  XNOR U5756 ( .A(n5542), .B(n5543), .Z(n5534) );
  NANDN U5757 ( .A(n5540), .B(n5544), .Z(n5543) );
  ANDN U5758 ( .B(n5537), .A(n5545), .Z(n5535) );
  IV U5759 ( .A(n5492), .Z(n5537) );
  XOR U5760 ( .A(n5455), .B(n5375), .Z(n5492) );
  XNOR U5761 ( .A(n5546), .B(n5542), .Z(n5375) );
  NANDN U5762 ( .A(n5547), .B(n5548), .Z(n5542) );
  XOR U5763 ( .A(n5544), .B(n5549), .Z(n5548) );
  ANDN U5764 ( .B(n5549), .A(n5550), .Z(n5546) );
  XOR U5765 ( .A(n5551), .B(n5538), .Z(n5455) );
  NANDN U5766 ( .A(n5547), .B(n5552), .Z(n5538) );
  XOR U5767 ( .A(n5553), .B(n5541), .Z(n5552) );
  XNOR U5768 ( .A(n5554), .B(n5555), .Z(n5540) );
  XOR U5769 ( .A(n5556), .B(n5557), .Z(n5555) );
  XNOR U5770 ( .A(n5558), .B(n5559), .Z(n5554) );
  XNOR U5771 ( .A(n5560), .B(n5561), .Z(n5559) );
  ANDN U5772 ( .B(n5553), .A(n5557), .Z(n5560) );
  ANDN U5773 ( .B(n5553), .A(n5550), .Z(n5551) );
  XNOR U5774 ( .A(n5556), .B(n5562), .Z(n5550) );
  XOR U5775 ( .A(n5563), .B(n5561), .Z(n5562) );
  NAND U5776 ( .A(n5564), .B(n5565), .Z(n5561) );
  XNOR U5777 ( .A(n5558), .B(n5541), .Z(n5565) );
  IV U5778 ( .A(n5553), .Z(n5558) );
  XNOR U5779 ( .A(n5544), .B(n5557), .Z(n5564) );
  IV U5780 ( .A(n5549), .Z(n5557) );
  XOR U5781 ( .A(n5566), .B(n5567), .Z(n5549) );
  XNOR U5782 ( .A(n5568), .B(n5569), .Z(n5567) );
  XNOR U5783 ( .A(n5570), .B(n5571), .Z(n5566) );
  NOR U5784 ( .A(n5454), .B(n5525), .Z(n5570) );
  AND U5785 ( .A(n5541), .B(n5544), .Z(n5563) );
  XNOR U5786 ( .A(n5541), .B(n5544), .Z(n5556) );
  XNOR U5787 ( .A(n5572), .B(n5573), .Z(n5544) );
  XNOR U5788 ( .A(n5574), .B(n5569), .Z(n5573) );
  XOR U5789 ( .A(n5575), .B(n5576), .Z(n5572) );
  XNOR U5790 ( .A(n5577), .B(n5571), .Z(n5576) );
  OR U5791 ( .A(n5453), .B(n5524), .Z(n5571) );
  XNOR U5792 ( .A(n5525), .B(n5481), .Z(n5524) );
  XNOR U5793 ( .A(n5454), .B(n5339), .Z(n5453) );
  ANDN U5794 ( .B(n5578), .A(n5481), .Z(n5577) );
  XNOR U5795 ( .A(n5579), .B(n5580), .Z(n5541) );
  XNOR U5796 ( .A(n5569), .B(n5581), .Z(n5580) );
  XOR U5797 ( .A(n5471), .B(n5575), .Z(n5581) );
  XNOR U5798 ( .A(n5525), .B(n5582), .Z(n5569) );
  XNOR U5799 ( .A(n5583), .B(n5584), .Z(n5579) );
  XNOR U5800 ( .A(n5585), .B(n5586), .Z(n5584) );
  ANDN U5801 ( .B(n5533), .A(n5484), .Z(n5585) );
  XNOR U5802 ( .A(n5587), .B(n5588), .Z(n5553) );
  XNOR U5803 ( .A(n5574), .B(n5589), .Z(n5588) );
  XNOR U5804 ( .A(n5484), .B(n5568), .Z(n5589) );
  XOR U5805 ( .A(n5575), .B(n5590), .Z(n5568) );
  XNOR U5806 ( .A(n5591), .B(n5592), .Z(n5590) );
  NAND U5807 ( .A(n5529), .B(n5476), .Z(n5592) );
  XNOR U5808 ( .A(n5593), .B(n5591), .Z(n5575) );
  NANDN U5809 ( .A(n5536), .B(n5490), .Z(n5591) );
  XOR U5810 ( .A(n5491), .B(n5476), .Z(n5490) );
  XNOR U5811 ( .A(n5594), .B(n5339), .Z(n5476) );
  XOR U5812 ( .A(n5545), .B(n5529), .Z(n5536) );
  XOR U5813 ( .A(n5533), .B(n5595), .Z(n5529) );
  ANDN U5814 ( .B(n5491), .A(n5545), .Z(n5593) );
  XOR U5815 ( .A(n5583), .B(n5525), .Z(n5545) );
  XOR U5816 ( .A(n5596), .B(n5597), .Z(n5525) );
  XNOR U5817 ( .A(n5598), .B(n5599), .Z(n5597) );
  XOR U5818 ( .A(n5600), .B(n5582), .Z(n5491) );
  XOR U5819 ( .A(n5595), .B(n5578), .Z(n5574) );
  IV U5820 ( .A(n5339), .Z(n5578) );
  XOR U5821 ( .A(n5601), .B(n5602), .Z(n5339) );
  XNOR U5822 ( .A(n5603), .B(n5599), .Z(n5602) );
  IV U5823 ( .A(n5481), .Z(n5595) );
  XOR U5824 ( .A(n5599), .B(n5604), .Z(n5481) );
  XNOR U5825 ( .A(n5533), .B(n5605), .Z(n5587) );
  XNOR U5826 ( .A(n5606), .B(n5586), .Z(n5605) );
  OR U5827 ( .A(n5487), .B(n5532), .Z(n5586) );
  XNOR U5828 ( .A(n5583), .B(n5533), .Z(n5532) );
  XOR U5829 ( .A(n5471), .B(n5594), .Z(n5487) );
  IV U5830 ( .A(n5484), .Z(n5594) );
  XOR U5831 ( .A(n5582), .B(n5607), .Z(n5484) );
  XNOR U5832 ( .A(n5603), .B(n5596), .Z(n5607) );
  XOR U5833 ( .A(n5608), .B(n5609), .Z(n5596) );
  XNOR U5834 ( .A(n2888), .B(n4129), .Z(n5609) );
  XNOR U5835 ( .A(n2840), .B(n5610), .Z(n4129) );
  XOR U5836 ( .A(n4812), .B(n5611), .Z(n5608) );
  XNOR U5837 ( .A(key[490]), .B(n4814), .Z(n5611) );
  XOR U5838 ( .A(n5612), .B(n5613), .Z(n4814) );
  XNOR U5839 ( .A(n5614), .B(n5615), .Z(n5613) );
  XNOR U5840 ( .A(n5616), .B(n5617), .Z(n5612) );
  IV U5841 ( .A(n2883), .Z(n4812) );
  IV U5842 ( .A(n5454), .Z(n5582) );
  XOR U5843 ( .A(n5601), .B(n5618), .Z(n5454) );
  XOR U5844 ( .A(n5599), .B(n5619), .Z(n5618) );
  ANDN U5845 ( .B(n5600), .A(n5374), .Z(n5606) );
  IV U5846 ( .A(n5471), .Z(n5600) );
  XOR U5847 ( .A(n5601), .B(n5620), .Z(n5471) );
  XOR U5848 ( .A(n5599), .B(n5621), .Z(n5620) );
  XOR U5849 ( .A(n5622), .B(n5623), .Z(n5599) );
  XNOR U5850 ( .A(n4138), .B(n5374), .Z(n5623) );
  IV U5851 ( .A(n5583), .Z(n5374) );
  XOR U5852 ( .A(n5624), .B(n5625), .Z(n4138) );
  XOR U5853 ( .A(n4795), .B(n5626), .Z(n5622) );
  XNOR U5854 ( .A(key[494]), .B(n4799), .Z(n5626) );
  XNOR U5855 ( .A(n4121), .B(n4789), .Z(n4799) );
  XNOR U5856 ( .A(n4142), .B(n4114), .Z(n4789) );
  XOR U5857 ( .A(n5627), .B(n5628), .Z(n4114) );
  XNOR U5858 ( .A(n5629), .B(n5630), .Z(n5628) );
  XOR U5859 ( .A(n5631), .B(n5617), .Z(n5627) );
  XNOR U5860 ( .A(n2854), .B(n2861), .Z(n4121) );
  XOR U5861 ( .A(n5632), .B(n5633), .Z(n2861) );
  IV U5862 ( .A(n2857), .Z(n4795) );
  XNOR U5863 ( .A(n5634), .B(n5635), .Z(n2857) );
  IV U5864 ( .A(n5604), .Z(n5601) );
  XOR U5865 ( .A(n5636), .B(n5637), .Z(n5604) );
  XOR U5866 ( .A(n4120), .B(n4793), .Z(n5637) );
  XNOR U5867 ( .A(n4104), .B(n5638), .Z(n4793) );
  XNOR U5868 ( .A(n5639), .B(n5640), .Z(n4104) );
  XNOR U5869 ( .A(n5641), .B(n5642), .Z(n5640) );
  XNOR U5870 ( .A(n5643), .B(n5644), .Z(n5639) );
  XOR U5871 ( .A(n5645), .B(n5646), .Z(n5644) );
  ANDN U5872 ( .B(n5647), .A(n5648), .Z(n5646) );
  XNOR U5873 ( .A(n5649), .B(n5650), .Z(n4120) );
  XOR U5874 ( .A(n5651), .B(n5652), .Z(n5650) );
  XNOR U5875 ( .A(n5653), .B(n5654), .Z(n5649) );
  XOR U5876 ( .A(n5655), .B(n5656), .Z(n5654) );
  ANDN U5877 ( .B(n5657), .A(n5658), .Z(n5656) );
  XOR U5878 ( .A(n4794), .B(n5659), .Z(n5636) );
  XNOR U5879 ( .A(key[493]), .B(n2854), .Z(n5659) );
  XOR U5880 ( .A(n5660), .B(n5661), .Z(n2854) );
  XOR U5881 ( .A(n5629), .B(n5615), .Z(n4794) );
  XNOR U5882 ( .A(n5662), .B(n5663), .Z(n5615) );
  XNOR U5883 ( .A(n5664), .B(n5665), .Z(n5663) );
  NOR U5884 ( .A(n5666), .B(n5667), .Z(n5664) );
  XOR U5885 ( .A(n5668), .B(n5669), .Z(n5533) );
  XNOR U5886 ( .A(n5621), .B(n5619), .Z(n5669) );
  XNOR U5887 ( .A(n5670), .B(n5671), .Z(n5619) );
  XOR U5888 ( .A(n4115), .B(n4790), .Z(n5671) );
  XNOR U5889 ( .A(n5625), .B(n4145), .Z(n4790) );
  XNOR U5890 ( .A(n5672), .B(n5673), .Z(n4145) );
  XOR U5891 ( .A(n5674), .B(n5642), .Z(n5673) );
  XNOR U5892 ( .A(n5675), .B(n5676), .Z(n5642) );
  XNOR U5893 ( .A(n5677), .B(n5678), .Z(n5676) );
  NANDN U5894 ( .A(n5679), .B(n5680), .Z(n5678) );
  XOR U5895 ( .A(n5681), .B(n5632), .Z(n5672) );
  IV U5896 ( .A(n2868), .Z(n5625) );
  XOR U5897 ( .A(n5682), .B(n5683), .Z(n2868) );
  XOR U5898 ( .A(n5684), .B(n5685), .Z(n5683) );
  XOR U5899 ( .A(n5686), .B(n5660), .Z(n5682) );
  XNOR U5900 ( .A(n5687), .B(n5688), .Z(n4115) );
  XNOR U5901 ( .A(n5634), .B(n5652), .Z(n5688) );
  XNOR U5902 ( .A(n5689), .B(n5690), .Z(n5652) );
  XNOR U5903 ( .A(n5691), .B(n5692), .Z(n5690) );
  OR U5904 ( .A(n5693), .B(n5694), .Z(n5692) );
  XOR U5905 ( .A(n5695), .B(n5696), .Z(n5687) );
  XOR U5906 ( .A(key[495]), .B(n4803), .Z(n5670) );
  IV U5907 ( .A(n2895), .Z(n4803) );
  XOR U5908 ( .A(n4142), .B(n5624), .Z(n2895) );
  XNOR U5909 ( .A(n5697), .B(n5698), .Z(n5621) );
  XOR U5910 ( .A(n4778), .B(n4098), .Z(n5698) );
  XOR U5911 ( .A(n5624), .B(n5638), .Z(n4098) );
  IV U5912 ( .A(n2859), .Z(n5638) );
  XOR U5913 ( .A(n5699), .B(n5700), .Z(n2859) );
  XNOR U5914 ( .A(n5701), .B(n5685), .Z(n5700) );
  XNOR U5915 ( .A(n5702), .B(n5703), .Z(n5685) );
  XNOR U5916 ( .A(n5704), .B(n5705), .Z(n5703) );
  NANDN U5917 ( .A(n5706), .B(n5707), .Z(n5705) );
  XNOR U5918 ( .A(n5708), .B(n5709), .Z(n5699) );
  XOR U5919 ( .A(n5710), .B(n5711), .Z(n5709) );
  ANDN U5920 ( .B(n5712), .A(n5713), .Z(n5711) );
  XOR U5921 ( .A(n2875), .B(n4102), .Z(n4778) );
  XNOR U5922 ( .A(n5643), .B(n2884), .Z(n4102) );
  IV U5923 ( .A(n5610), .Z(n2884) );
  XNOR U5924 ( .A(n5714), .B(n5674), .Z(n5610) );
  XNOR U5925 ( .A(n4779), .B(n5715), .Z(n5697) );
  XOR U5926 ( .A(key[492]), .B(n4100), .Z(n5715) );
  XNOR U5927 ( .A(n2883), .B(n5651), .Z(n4100) );
  XOR U5928 ( .A(n5695), .B(n5716), .Z(n2883) );
  IV U5929 ( .A(n5717), .Z(n5695) );
  XOR U5930 ( .A(n4142), .B(n4119), .Z(n4779) );
  XNOR U5931 ( .A(n5718), .B(n5719), .Z(n4119) );
  XNOR U5932 ( .A(n5720), .B(n5630), .Z(n5719) );
  XNOR U5933 ( .A(n5721), .B(n5722), .Z(n5630) );
  XNOR U5934 ( .A(n5723), .B(n5724), .Z(n5722) );
  OR U5935 ( .A(n5725), .B(n5726), .Z(n5724) );
  XNOR U5936 ( .A(n5727), .B(n5728), .Z(n5718) );
  XOR U5937 ( .A(n5665), .B(n5729), .Z(n5728) );
  ANDN U5938 ( .B(n5730), .A(n5731), .Z(n5729) );
  ANDN U5939 ( .B(n5732), .A(n5733), .Z(n5665) );
  XOR U5940 ( .A(n5583), .B(n5598), .Z(n5668) );
  XOR U5941 ( .A(n5734), .B(n5735), .Z(n5598) );
  XNOR U5942 ( .A(n5603), .B(n5736), .Z(n5735) );
  XOR U5943 ( .A(n2841), .B(n4125), .Z(n5736) );
  XNOR U5944 ( .A(n4116), .B(n2875), .Z(n4125) );
  XNOR U5945 ( .A(n5708), .B(n2840), .Z(n2875) );
  IV U5946 ( .A(n5624), .Z(n4116) );
  XNOR U5947 ( .A(n5737), .B(n5738), .Z(n2841) );
  XOR U5948 ( .A(n5739), .B(n5635), .Z(n5738) );
  XNOR U5949 ( .A(n5740), .B(n5741), .Z(n5635) );
  XNOR U5950 ( .A(n5742), .B(n5655), .Z(n5741) );
  ANDN U5951 ( .B(n5743), .A(n5744), .Z(n5655) );
  NOR U5952 ( .A(n5745), .B(n5746), .Z(n5742) );
  XNOR U5953 ( .A(n5717), .B(n5696), .Z(n5737) );
  XOR U5954 ( .A(n5747), .B(n5748), .Z(n5603) );
  XNOR U5955 ( .A(n4141), .B(n2840), .Z(n5748) );
  XNOR U5956 ( .A(n5749), .B(n5684), .Z(n2840) );
  XNOR U5957 ( .A(n5750), .B(n2893), .Z(n4141) );
  XNOR U5958 ( .A(n5674), .B(n5751), .Z(n2893) );
  XOR U5959 ( .A(n5714), .B(n5752), .Z(n5632) );
  IV U5960 ( .A(n5753), .Z(n5714) );
  XOR U5961 ( .A(n4811), .B(n5754), .Z(n5747) );
  XOR U5962 ( .A(key[489]), .B(n4805), .Z(n5754) );
  IV U5963 ( .A(n2897), .Z(n4805) );
  XNOR U5964 ( .A(n5634), .B(n5755), .Z(n2897) );
  XOR U5965 ( .A(n5717), .B(n5696), .Z(n5755) );
  XNOR U5966 ( .A(n5757), .B(n5758), .Z(n5756) );
  NANDN U5967 ( .A(n5693), .B(n5759), .Z(n5758) );
  XNOR U5968 ( .A(n5653), .B(n5760), .Z(n5740) );
  XNOR U5969 ( .A(n5761), .B(n5762), .Z(n5760) );
  NAND U5970 ( .A(n5763), .B(n5764), .Z(n5762) );
  XNOR U5971 ( .A(n5765), .B(n5766), .Z(n5717) );
  XNOR U5972 ( .A(n5767), .B(n5768), .Z(n5766) );
  NAND U5973 ( .A(n5769), .B(n5657), .Z(n5768) );
  XOR U5974 ( .A(n5716), .B(n5739), .Z(n5634) );
  XOR U5975 ( .A(n5653), .B(n5770), .Z(n5739) );
  XNOR U5976 ( .A(n5757), .B(n5771), .Z(n5770) );
  NANDN U5977 ( .A(n5772), .B(n5773), .Z(n5771) );
  OR U5978 ( .A(n5774), .B(n5775), .Z(n5757) );
  XOR U5979 ( .A(n5776), .B(n5761), .Z(n5653) );
  NANDN U5980 ( .A(n5777), .B(n5778), .Z(n5761) );
  AND U5981 ( .A(n5779), .B(n5780), .Z(n5776) );
  XOR U5982 ( .A(n4813), .B(n5781), .Z(n5734) );
  XNOR U5983 ( .A(key[491]), .B(n4816), .Z(n5781) );
  XOR U5984 ( .A(n5720), .B(n4811), .Z(n4099) );
  XOR U5985 ( .A(n5631), .B(n5782), .Z(n4811) );
  IV U5986 ( .A(n5616), .Z(n5631) );
  XOR U5987 ( .A(n5782), .B(n5720), .Z(n4142) );
  XNOR U5988 ( .A(n5721), .B(n5783), .Z(n5720) );
  XOR U5989 ( .A(n5784), .B(n5785), .Z(n5783) );
  NOR U5990 ( .A(n5786), .B(n5667), .Z(n5784) );
  XNOR U5991 ( .A(n5787), .B(n5788), .Z(n5721) );
  XNOR U5992 ( .A(n5789), .B(n5790), .Z(n5788) );
  NAND U5993 ( .A(n5791), .B(n5792), .Z(n5790) );
  IV U5994 ( .A(n5793), .Z(n5782) );
  XOR U5995 ( .A(n2888), .B(n2842), .Z(n4813) );
  XOR U5996 ( .A(n5794), .B(n5795), .Z(n2842) );
  XNOR U5997 ( .A(n5796), .B(n5797), .Z(n5633) );
  XNOR U5998 ( .A(n5798), .B(n5645), .Z(n5797) );
  ANDN U5999 ( .B(n5799), .A(n5800), .Z(n5645) );
  NOR U6000 ( .A(n5801), .B(n5802), .Z(n5798) );
  XOR U6001 ( .A(n5803), .B(n5804), .Z(n5674) );
  XNOR U6002 ( .A(n5805), .B(n5806), .Z(n5804) );
  NANDN U6003 ( .A(n5807), .B(n5647), .Z(n5806) );
  XOR U6004 ( .A(n5681), .B(n5752), .Z(n5794) );
  XOR U6005 ( .A(n5641), .B(n5808), .Z(n5752) );
  XNOR U6006 ( .A(n5809), .B(n5810), .Z(n5808) );
  NANDN U6007 ( .A(n5811), .B(n5812), .Z(n5810) );
  XNOR U6008 ( .A(n5809), .B(n5814), .Z(n5813) );
  NANDN U6009 ( .A(n5815), .B(n5680), .Z(n5814) );
  OR U6010 ( .A(n5816), .B(n5817), .Z(n5809) );
  XNOR U6011 ( .A(n5641), .B(n5818), .Z(n5796) );
  XNOR U6012 ( .A(n5819), .B(n5820), .Z(n5818) );
  NAND U6013 ( .A(n5821), .B(n5822), .Z(n5820) );
  XOR U6014 ( .A(n5823), .B(n5819), .Z(n5641) );
  NANDN U6015 ( .A(n5824), .B(n5825), .Z(n5819) );
  ANDN U6016 ( .B(n5826), .A(n5827), .Z(n5823) );
  XOR U6017 ( .A(n5828), .B(n5829), .Z(n2888) );
  XNOR U6018 ( .A(n5830), .B(n5831), .Z(n5661) );
  XNOR U6019 ( .A(n5832), .B(n5710), .Z(n5831) );
  ANDN U6020 ( .B(n5833), .A(n5834), .Z(n5710) );
  NOR U6021 ( .A(n5835), .B(n5836), .Z(n5832) );
  XOR U6022 ( .A(n5686), .B(n5837), .Z(n5828) );
  XOR U6023 ( .A(n5838), .B(n5839), .Z(n5583) );
  XOR U6024 ( .A(n5750), .B(n2867), .Z(n5839) );
  XNOR U6025 ( .A(n4103), .B(n2894), .Z(n2867) );
  XOR U6026 ( .A(n5716), .B(n5651), .Z(n2894) );
  XOR U6027 ( .A(n5689), .B(n5840), .Z(n5651) );
  XOR U6028 ( .A(n5841), .B(n5767), .Z(n5840) );
  XNOR U6029 ( .A(n5746), .B(n5657), .Z(n5743) );
  NOR U6030 ( .A(n5843), .B(n5746), .Z(n5841) );
  XNOR U6031 ( .A(n5765), .B(n5844), .Z(n5689) );
  XNOR U6032 ( .A(n5845), .B(n5846), .Z(n5844) );
  NAND U6033 ( .A(n5764), .B(n5847), .Z(n5846) );
  XNOR U6034 ( .A(n5765), .B(n5848), .Z(n5716) );
  XOR U6035 ( .A(n5849), .B(n5691), .Z(n5848) );
  OR U6036 ( .A(n5774), .B(n5850), .Z(n5691) );
  XNOR U6037 ( .A(n5693), .B(n5772), .Z(n5774) );
  NOR U6038 ( .A(n5851), .B(n5772), .Z(n5849) );
  XOR U6039 ( .A(n5852), .B(n5845), .Z(n5765) );
  OR U6040 ( .A(n5777), .B(n5853), .Z(n5845) );
  XNOR U6041 ( .A(n5779), .B(n5764), .Z(n5777) );
  XNOR U6042 ( .A(n5772), .B(n5657), .Z(n5764) );
  XOR U6043 ( .A(n5854), .B(n5855), .Z(n5657) );
  NANDN U6044 ( .A(n5856), .B(n5857), .Z(n5855) );
  XNOR U6045 ( .A(n5858), .B(n5859), .Z(n5772) );
  OR U6046 ( .A(n5856), .B(n5860), .Z(n5859) );
  ANDN U6047 ( .B(n5779), .A(n5861), .Z(n5852) );
  XOR U6048 ( .A(n5693), .B(n5746), .Z(n5779) );
  XOR U6049 ( .A(n5862), .B(n5854), .Z(n5746) );
  NANDN U6050 ( .A(n5863), .B(n5864), .Z(n5854) );
  ANDN U6051 ( .B(n5865), .A(n5866), .Z(n5862) );
  NANDN U6052 ( .A(n5863), .B(n5868), .Z(n5858) );
  XOR U6053 ( .A(n5869), .B(n5856), .Z(n5863) );
  XNOR U6054 ( .A(n5870), .B(n5871), .Z(n5856) );
  XOR U6055 ( .A(n5872), .B(n5865), .Z(n5871) );
  XNOR U6056 ( .A(n5873), .B(n5874), .Z(n5870) );
  XNOR U6057 ( .A(n5875), .B(n5876), .Z(n5874) );
  ANDN U6058 ( .B(n5865), .A(n5877), .Z(n5875) );
  IV U6059 ( .A(n5878), .Z(n5865) );
  ANDN U6060 ( .B(n5869), .A(n5877), .Z(n5867) );
  IV U6061 ( .A(n5873), .Z(n5877) );
  IV U6062 ( .A(n5866), .Z(n5869) );
  XNOR U6063 ( .A(n5872), .B(n5879), .Z(n5866) );
  XOR U6064 ( .A(n5880), .B(n5876), .Z(n5879) );
  NAND U6065 ( .A(n5868), .B(n5864), .Z(n5876) );
  XNOR U6066 ( .A(n5857), .B(n5878), .Z(n5864) );
  XOR U6067 ( .A(n5881), .B(n5882), .Z(n5878) );
  XOR U6068 ( .A(n5883), .B(n5884), .Z(n5882) );
  XNOR U6069 ( .A(n5773), .B(n5885), .Z(n5884) );
  XNOR U6070 ( .A(n5886), .B(n5887), .Z(n5881) );
  XNOR U6071 ( .A(n5888), .B(n5889), .Z(n5887) );
  ANDN U6072 ( .B(n5759), .A(n5694), .Z(n5888) );
  XNOR U6073 ( .A(n5873), .B(n5860), .Z(n5868) );
  XOR U6074 ( .A(n5890), .B(n5891), .Z(n5873) );
  XNOR U6075 ( .A(n5892), .B(n5885), .Z(n5891) );
  XOR U6076 ( .A(n5893), .B(n5894), .Z(n5885) );
  XNOR U6077 ( .A(n5895), .B(n5896), .Z(n5894) );
  NAND U6078 ( .A(n5847), .B(n5763), .Z(n5896) );
  XNOR U6079 ( .A(n5897), .B(n5898), .Z(n5890) );
  ANDN U6080 ( .B(n5899), .A(n5843), .Z(n5897) );
  ANDN U6081 ( .B(n5857), .A(n5860), .Z(n5880) );
  XOR U6082 ( .A(n5860), .B(n5857), .Z(n5872) );
  XNOR U6083 ( .A(n5900), .B(n5901), .Z(n5857) );
  XNOR U6084 ( .A(n5893), .B(n5902), .Z(n5901) );
  XNOR U6085 ( .A(n5892), .B(n5759), .Z(n5902) );
  XNOR U6086 ( .A(n5903), .B(n5904), .Z(n5900) );
  XNOR U6087 ( .A(n5905), .B(n5889), .Z(n5904) );
  OR U6088 ( .A(n5775), .B(n5850), .Z(n5889) );
  XNOR U6089 ( .A(n5903), .B(n5886), .Z(n5850) );
  XNOR U6090 ( .A(n5759), .B(n5773), .Z(n5775) );
  ANDN U6091 ( .B(n5773), .A(n5851), .Z(n5905) );
  XOR U6092 ( .A(n5906), .B(n5907), .Z(n5860) );
  XOR U6093 ( .A(n5893), .B(n5883), .Z(n5907) );
  XOR U6094 ( .A(n5769), .B(n5658), .Z(n5883) );
  XOR U6095 ( .A(n5908), .B(n5895), .Z(n5893) );
  NANDN U6096 ( .A(n5853), .B(n5778), .Z(n5895) );
  XOR U6097 ( .A(n5780), .B(n5763), .Z(n5778) );
  XNOR U6098 ( .A(n5899), .B(n5909), .Z(n5773) );
  XNOR U6099 ( .A(n5910), .B(n5911), .Z(n5909) );
  XOR U6100 ( .A(n5861), .B(n5847), .Z(n5853) );
  XNOR U6101 ( .A(n5851), .B(n5769), .Z(n5847) );
  IV U6102 ( .A(n5886), .Z(n5851) );
  XOR U6103 ( .A(n5912), .B(n5913), .Z(n5886) );
  XOR U6104 ( .A(n5914), .B(n5915), .Z(n5913) );
  XOR U6105 ( .A(n5903), .B(n5916), .Z(n5912) );
  ANDN U6106 ( .B(n5780), .A(n5861), .Z(n5908) );
  XNOR U6107 ( .A(n5903), .B(n5917), .Z(n5861) );
  XOR U6108 ( .A(n5899), .B(n5759), .Z(n5780) );
  XNOR U6109 ( .A(n5918), .B(n5919), .Z(n5759) );
  XOR U6110 ( .A(n5920), .B(n5915), .Z(n5919) );
  XNOR U6111 ( .A(n5921), .B(n5922), .Z(n5915) );
  XNOR U6112 ( .A(n5923), .B(n5924), .Z(n5922) );
  XNOR U6113 ( .A(n5925), .B(n5926), .Z(n5921) );
  XNOR U6114 ( .A(key[340]), .B(n5927), .Z(n5926) );
  IV U6115 ( .A(n5745), .Z(n5899) );
  XOR U6116 ( .A(n5892), .B(n5928), .Z(n5906) );
  XNOR U6117 ( .A(n5929), .B(n5898), .Z(n5928) );
  OR U6118 ( .A(n5744), .B(n5842), .Z(n5898) );
  XNOR U6119 ( .A(n5917), .B(n5769), .Z(n5842) );
  XNOR U6120 ( .A(n5745), .B(n5658), .Z(n5744) );
  ANDN U6121 ( .B(n5769), .A(n5658), .Z(n5929) );
  XOR U6122 ( .A(n5918), .B(n5930), .Z(n5658) );
  XOR U6123 ( .A(n5910), .B(n5931), .Z(n5930) );
  XOR U6124 ( .A(n5920), .B(n5918), .Z(n5769) );
  XNOR U6125 ( .A(n5843), .B(n5745), .Z(n5892) );
  XOR U6126 ( .A(n5918), .B(n5932), .Z(n5745) );
  XNOR U6127 ( .A(n5920), .B(n5914), .Z(n5932) );
  XOR U6128 ( .A(n5933), .B(n5934), .Z(n5914) );
  XNOR U6129 ( .A(n5935), .B(n5936), .Z(n5934) );
  XOR U6130 ( .A(key[343]), .B(n5937), .Z(n5933) );
  XNOR U6131 ( .A(n5938), .B(n5939), .Z(n5918) );
  XNOR U6132 ( .A(n5940), .B(n5941), .Z(n5939) );
  XNOR U6133 ( .A(key[341]), .B(n5942), .Z(n5938) );
  IV U6134 ( .A(n5917), .Z(n5843) );
  XNOR U6135 ( .A(n5911), .B(n5943), .Z(n5917) );
  XOR U6136 ( .A(n5916), .B(n5931), .Z(n5943) );
  IV U6137 ( .A(n5920), .Z(n5931) );
  XOR U6138 ( .A(n5944), .B(n5945), .Z(n5920) );
  XOR U6139 ( .A(n5946), .B(n5694), .Z(n5945) );
  IV U6140 ( .A(n5903), .Z(n5694) );
  XOR U6141 ( .A(n5947), .B(n5948), .Z(n5903) );
  XNOR U6142 ( .A(n5949), .B(n5950), .Z(n5948) );
  XNOR U6143 ( .A(key[336]), .B(n5951), .Z(n5947) );
  XOR U6144 ( .A(n5952), .B(n5953), .Z(n5944) );
  XNOR U6145 ( .A(key[342]), .B(n5954), .Z(n5953) );
  XOR U6146 ( .A(n5955), .B(n5956), .Z(n5916) );
  XNOR U6147 ( .A(n5910), .B(n5957), .Z(n5956) );
  XOR U6148 ( .A(n5958), .B(n5959), .Z(n5957) );
  XOR U6149 ( .A(n5960), .B(n5961), .Z(n5910) );
  XNOR U6150 ( .A(n5962), .B(n5963), .Z(n5961) );
  XOR U6151 ( .A(key[337]), .B(n5964), .Z(n5960) );
  XOR U6152 ( .A(n5965), .B(n5966), .Z(n5955) );
  XNOR U6153 ( .A(key[339]), .B(n5967), .Z(n5966) );
  XOR U6154 ( .A(n5968), .B(n5969), .Z(n5911) );
  XNOR U6155 ( .A(n5970), .B(n5971), .Z(n5969) );
  XOR U6156 ( .A(key[338]), .B(n5972), .Z(n5968) );
  IV U6157 ( .A(n4130), .Z(n4103) );
  XOR U6158 ( .A(n5643), .B(n5753), .Z(n4130) );
  XNOR U6159 ( .A(n5803), .B(n5973), .Z(n5753) );
  XOR U6160 ( .A(n5974), .B(n5677), .Z(n5973) );
  OR U6161 ( .A(n5975), .B(n5816), .Z(n5677) );
  XNOR U6162 ( .A(n5680), .B(n5812), .Z(n5816) );
  ANDN U6163 ( .B(n5976), .A(n5977), .Z(n5974) );
  XNOR U6164 ( .A(n5675), .B(n5978), .Z(n5643) );
  XOR U6165 ( .A(n5979), .B(n5805), .Z(n5978) );
  XNOR U6166 ( .A(n5802), .B(n5647), .Z(n5799) );
  NOR U6167 ( .A(n5981), .B(n5802), .Z(n5979) );
  XNOR U6168 ( .A(n5803), .B(n5982), .Z(n5675) );
  XNOR U6169 ( .A(n5983), .B(n5984), .Z(n5982) );
  NAND U6170 ( .A(n5822), .B(n5985), .Z(n5984) );
  XOR U6171 ( .A(n5986), .B(n5983), .Z(n5803) );
  OR U6172 ( .A(n5824), .B(n5987), .Z(n5983) );
  XNOR U6173 ( .A(n5988), .B(n5822), .Z(n5824) );
  XOR U6174 ( .A(n5812), .B(n5647), .Z(n5822) );
  XOR U6175 ( .A(n5989), .B(n5990), .Z(n5647) );
  NANDN U6176 ( .A(n5991), .B(n5992), .Z(n5990) );
  IV U6177 ( .A(n5977), .Z(n5812) );
  XNOR U6178 ( .A(n5993), .B(n5994), .Z(n5977) );
  NANDN U6179 ( .A(n5991), .B(n5995), .Z(n5994) );
  ANDN U6180 ( .B(n5988), .A(n5996), .Z(n5986) );
  IV U6181 ( .A(n5827), .Z(n5988) );
  XOR U6182 ( .A(n5802), .B(n5680), .Z(n5827) );
  XNOR U6183 ( .A(n5997), .B(n5993), .Z(n5680) );
  NANDN U6184 ( .A(n5998), .B(n5999), .Z(n5993) );
  XOR U6185 ( .A(n5995), .B(n6000), .Z(n5999) );
  ANDN U6186 ( .B(n6000), .A(n6001), .Z(n5997) );
  XOR U6187 ( .A(n6002), .B(n5989), .Z(n5802) );
  NANDN U6188 ( .A(n5998), .B(n6003), .Z(n5989) );
  XOR U6189 ( .A(n6004), .B(n5992), .Z(n6003) );
  XNOR U6190 ( .A(n6005), .B(n6006), .Z(n5991) );
  XOR U6191 ( .A(n6007), .B(n6008), .Z(n6006) );
  XNOR U6192 ( .A(n6009), .B(n6010), .Z(n6005) );
  XNOR U6193 ( .A(n6011), .B(n6012), .Z(n6010) );
  ANDN U6194 ( .B(n6004), .A(n6008), .Z(n6011) );
  ANDN U6195 ( .B(n6004), .A(n6001), .Z(n6002) );
  XNOR U6196 ( .A(n6007), .B(n6013), .Z(n6001) );
  XOR U6197 ( .A(n6014), .B(n6012), .Z(n6013) );
  NAND U6198 ( .A(n6015), .B(n6016), .Z(n6012) );
  XNOR U6199 ( .A(n6009), .B(n5992), .Z(n6016) );
  IV U6200 ( .A(n6004), .Z(n6009) );
  XNOR U6201 ( .A(n5995), .B(n6008), .Z(n6015) );
  IV U6202 ( .A(n6000), .Z(n6008) );
  XOR U6203 ( .A(n6017), .B(n6018), .Z(n6000) );
  XNOR U6204 ( .A(n6019), .B(n6020), .Z(n6018) );
  XNOR U6205 ( .A(n6021), .B(n6022), .Z(n6017) );
  NOR U6206 ( .A(n5801), .B(n5981), .Z(n6021) );
  AND U6207 ( .A(n5992), .B(n5995), .Z(n6014) );
  XNOR U6208 ( .A(n5992), .B(n5995), .Z(n6007) );
  XNOR U6209 ( .A(n6023), .B(n6024), .Z(n5995) );
  XNOR U6210 ( .A(n6025), .B(n6020), .Z(n6024) );
  XOR U6211 ( .A(n6026), .B(n6027), .Z(n6023) );
  XNOR U6212 ( .A(n6028), .B(n6022), .Z(n6027) );
  OR U6213 ( .A(n5800), .B(n5980), .Z(n6022) );
  XNOR U6214 ( .A(n5981), .B(n5807), .Z(n5980) );
  XNOR U6215 ( .A(n5801), .B(n5648), .Z(n5800) );
  ANDN U6216 ( .B(n6029), .A(n5807), .Z(n6028) );
  XNOR U6217 ( .A(n6030), .B(n6031), .Z(n5992) );
  XNOR U6218 ( .A(n6020), .B(n6032), .Z(n6031) );
  XOR U6219 ( .A(n5815), .B(n6026), .Z(n6032) );
  XNOR U6220 ( .A(n5981), .B(n6033), .Z(n6020) );
  XNOR U6221 ( .A(n6034), .B(n6035), .Z(n6030) );
  XNOR U6222 ( .A(n6036), .B(n6037), .Z(n6035) );
  ANDN U6223 ( .B(n5976), .A(n5811), .Z(n6036) );
  XNOR U6224 ( .A(n6038), .B(n6039), .Z(n6004) );
  XNOR U6225 ( .A(n6025), .B(n6040), .Z(n6039) );
  XNOR U6226 ( .A(n5811), .B(n6019), .Z(n6040) );
  XOR U6227 ( .A(n6026), .B(n6041), .Z(n6019) );
  XNOR U6228 ( .A(n6042), .B(n6043), .Z(n6041) );
  NAND U6229 ( .A(n5985), .B(n5821), .Z(n6043) );
  XNOR U6230 ( .A(n6044), .B(n6042), .Z(n6026) );
  NANDN U6231 ( .A(n5987), .B(n5825), .Z(n6042) );
  XOR U6232 ( .A(n5826), .B(n5821), .Z(n5825) );
  XNOR U6233 ( .A(n6045), .B(n5648), .Z(n5821) );
  XOR U6234 ( .A(n5996), .B(n5985), .Z(n5987) );
  XOR U6235 ( .A(n5976), .B(n6046), .Z(n5985) );
  ANDN U6236 ( .B(n5826), .A(n5996), .Z(n6044) );
  XOR U6237 ( .A(n6034), .B(n5981), .Z(n5996) );
  XOR U6238 ( .A(n6047), .B(n6048), .Z(n5981) );
  XNOR U6239 ( .A(n6049), .B(n6050), .Z(n6048) );
  XOR U6240 ( .A(n6051), .B(n6033), .Z(n5826) );
  XOR U6241 ( .A(n6046), .B(n6029), .Z(n6025) );
  IV U6242 ( .A(n5648), .Z(n6029) );
  XOR U6243 ( .A(n6052), .B(n6053), .Z(n5648) );
  XNOR U6244 ( .A(n6054), .B(n6050), .Z(n6053) );
  IV U6245 ( .A(n5807), .Z(n6046) );
  XOR U6246 ( .A(n6050), .B(n6055), .Z(n5807) );
  XNOR U6247 ( .A(n5976), .B(n6056), .Z(n6038) );
  XNOR U6248 ( .A(n6057), .B(n6037), .Z(n6056) );
  OR U6249 ( .A(n5817), .B(n5975), .Z(n6037) );
  XNOR U6250 ( .A(n6034), .B(n5976), .Z(n5975) );
  XOR U6251 ( .A(n5815), .B(n6045), .Z(n5817) );
  IV U6252 ( .A(n5811), .Z(n6045) );
  XOR U6253 ( .A(n6033), .B(n6058), .Z(n5811) );
  XNOR U6254 ( .A(n6054), .B(n6047), .Z(n6058) );
  XOR U6255 ( .A(n6059), .B(n6060), .Z(n6047) );
  XOR U6256 ( .A(n6061), .B(n6062), .Z(n6060) );
  XNOR U6257 ( .A(n6063), .B(n6064), .Z(n6059) );
  XOR U6258 ( .A(key[378]), .B(n6065), .Z(n6064) );
  IV U6259 ( .A(n5801), .Z(n6033) );
  XOR U6260 ( .A(n6052), .B(n6066), .Z(n5801) );
  XOR U6261 ( .A(n6050), .B(n6067), .Z(n6066) );
  ANDN U6262 ( .B(n6051), .A(n5679), .Z(n6057) );
  IV U6263 ( .A(n5815), .Z(n6051) );
  XOR U6264 ( .A(n6052), .B(n6068), .Z(n5815) );
  XOR U6265 ( .A(n6050), .B(n6069), .Z(n6068) );
  XOR U6266 ( .A(n6070), .B(n6071), .Z(n6050) );
  XNOR U6267 ( .A(n6072), .B(n5679), .Z(n6071) );
  IV U6268 ( .A(n6034), .Z(n5679) );
  XNOR U6269 ( .A(n6073), .B(n6074), .Z(n6070) );
  XOR U6270 ( .A(key[382]), .B(n6075), .Z(n6074) );
  IV U6271 ( .A(n6055), .Z(n6052) );
  XOR U6272 ( .A(n6076), .B(n6077), .Z(n6055) );
  XOR U6273 ( .A(n6078), .B(n6079), .Z(n6077) );
  XOR U6274 ( .A(n6080), .B(n6081), .Z(n6076) );
  XNOR U6275 ( .A(key[381]), .B(n6082), .Z(n6081) );
  XOR U6276 ( .A(n6083), .B(n6084), .Z(n5976) );
  XNOR U6277 ( .A(n6069), .B(n6067), .Z(n6084) );
  XNOR U6278 ( .A(n6085), .B(n6086), .Z(n6067) );
  XOR U6279 ( .A(n6087), .B(n6088), .Z(n6086) );
  XNOR U6280 ( .A(key[383]), .B(n6089), .Z(n6085) );
  XNOR U6281 ( .A(n6090), .B(n6091), .Z(n6069) );
  XOR U6282 ( .A(n6092), .B(n6093), .Z(n6090) );
  XOR U6283 ( .A(key[380]), .B(n6094), .Z(n6093) );
  XOR U6284 ( .A(n6034), .B(n6049), .Z(n6083) );
  XOR U6285 ( .A(n6095), .B(n6096), .Z(n6049) );
  XNOR U6286 ( .A(n6054), .B(n6097), .Z(n6096) );
  XOR U6287 ( .A(n6098), .B(n6099), .Z(n6097) );
  XOR U6288 ( .A(n6100), .B(n6101), .Z(n6054) );
  XNOR U6289 ( .A(n6102), .B(n6103), .Z(n6101) );
  XOR U6290 ( .A(n6104), .B(n6105), .Z(n6100) );
  XNOR U6291 ( .A(key[377]), .B(n6106), .Z(n6105) );
  XNOR U6292 ( .A(n6107), .B(n6108), .Z(n6095) );
  XOR U6293 ( .A(key[379]), .B(n6109), .Z(n6108) );
  XOR U6294 ( .A(n6110), .B(n6111), .Z(n6034) );
  XOR U6295 ( .A(n6112), .B(n6113), .Z(n6111) );
  XOR U6296 ( .A(n6114), .B(n6115), .Z(n6110) );
  XOR U6297 ( .A(key[376]), .B(n6116), .Z(n6115) );
  IV U6298 ( .A(n2885), .Z(n5750) );
  XOR U6299 ( .A(n5684), .B(n6117), .Z(n2885) );
  XOR U6300 ( .A(n5749), .B(n5837), .Z(n5660) );
  XOR U6301 ( .A(n5701), .B(n6118), .Z(n5837) );
  XNOR U6302 ( .A(n6119), .B(n6120), .Z(n6118) );
  NANDN U6303 ( .A(n6121), .B(n6122), .Z(n6120) );
  IV U6304 ( .A(n6123), .Z(n5749) );
  XNOR U6305 ( .A(n6119), .B(n6125), .Z(n6124) );
  NANDN U6306 ( .A(n6126), .B(n5707), .Z(n6125) );
  OR U6307 ( .A(n6127), .B(n6128), .Z(n6119) );
  XNOR U6308 ( .A(n5701), .B(n6129), .Z(n5830) );
  XNOR U6309 ( .A(n6130), .B(n6131), .Z(n6129) );
  NAND U6310 ( .A(n6132), .B(n6133), .Z(n6131) );
  XOR U6311 ( .A(n6134), .B(n6130), .Z(n5701) );
  NANDN U6312 ( .A(n6135), .B(n6136), .Z(n6130) );
  ANDN U6313 ( .B(n6137), .A(n6138), .Z(n6134) );
  XOR U6314 ( .A(n6139), .B(n6140), .Z(n5684) );
  XNOR U6315 ( .A(n6141), .B(n6142), .Z(n6140) );
  NANDN U6316 ( .A(n6143), .B(n5712), .Z(n6142) );
  XOR U6317 ( .A(n5624), .B(n6144), .Z(n5838) );
  XNOR U6318 ( .A(key[488]), .B(n4804), .Z(n6144) );
  XNOR U6319 ( .A(n5629), .B(n6145), .Z(n4804) );
  XOR U6320 ( .A(n5616), .B(n5617), .Z(n6145) );
  XNOR U6321 ( .A(n6147), .B(n6148), .Z(n6146) );
  NANDN U6322 ( .A(n5725), .B(n6149), .Z(n6148) );
  XNOR U6323 ( .A(n5727), .B(n6150), .Z(n5662) );
  XNOR U6324 ( .A(n6151), .B(n6152), .Z(n6150) );
  NAND U6325 ( .A(n6153), .B(n5791), .Z(n6152) );
  XNOR U6326 ( .A(n5787), .B(n6154), .Z(n5616) );
  XNOR U6327 ( .A(n5785), .B(n6155), .Z(n6154) );
  NAND U6328 ( .A(n6156), .B(n5730), .Z(n6155) );
  XNOR U6329 ( .A(n5667), .B(n5730), .Z(n5732) );
  XNOR U6330 ( .A(n5614), .B(n5793), .Z(n5629) );
  XNOR U6331 ( .A(n5787), .B(n6158), .Z(n5793) );
  XOR U6332 ( .A(n6159), .B(n5723), .Z(n6158) );
  OR U6333 ( .A(n6160), .B(n6161), .Z(n5723) );
  NOR U6334 ( .A(n6162), .B(n6163), .Z(n6159) );
  XOR U6335 ( .A(n6164), .B(n5789), .Z(n5787) );
  OR U6336 ( .A(n6165), .B(n6166), .Z(n5789) );
  ANDN U6337 ( .B(n6167), .A(n6168), .Z(n6164) );
  XNOR U6338 ( .A(n5727), .B(n6169), .Z(n5614) );
  XNOR U6339 ( .A(n6147), .B(n6170), .Z(n6169) );
  NANDN U6340 ( .A(n6163), .B(n6171), .Z(n6170) );
  OR U6341 ( .A(n6161), .B(n6172), .Z(n6147) );
  XNOR U6342 ( .A(n5725), .B(n6163), .Z(n6161) );
  XOR U6343 ( .A(n6173), .B(n6151), .Z(n5727) );
  NANDN U6344 ( .A(n6165), .B(n6174), .Z(n6151) );
  XNOR U6345 ( .A(n6167), .B(n5791), .Z(n6165) );
  XNOR U6346 ( .A(n6163), .B(n5730), .Z(n5791) );
  XOR U6347 ( .A(n6175), .B(n6176), .Z(n5730) );
  NANDN U6348 ( .A(n6177), .B(n6178), .Z(n6176) );
  XNOR U6349 ( .A(n6179), .B(n6180), .Z(n6163) );
  OR U6350 ( .A(n6177), .B(n6181), .Z(n6180) );
  AND U6351 ( .A(n6167), .B(n6182), .Z(n6173) );
  XOR U6352 ( .A(n5725), .B(n5667), .Z(n6167) );
  XOR U6353 ( .A(n6183), .B(n6175), .Z(n5667) );
  NANDN U6354 ( .A(n6184), .B(n6185), .Z(n6175) );
  ANDN U6355 ( .B(n6186), .A(n6187), .Z(n6183) );
  NANDN U6356 ( .A(n6184), .B(n6189), .Z(n6179) );
  XOR U6357 ( .A(n6190), .B(n6177), .Z(n6184) );
  XNOR U6358 ( .A(n6191), .B(n6192), .Z(n6177) );
  XOR U6359 ( .A(n6193), .B(n6186), .Z(n6192) );
  XNOR U6360 ( .A(n6194), .B(n6195), .Z(n6191) );
  XNOR U6361 ( .A(n6196), .B(n6197), .Z(n6195) );
  ANDN U6362 ( .B(n6186), .A(n6198), .Z(n6196) );
  IV U6363 ( .A(n6199), .Z(n6186) );
  ANDN U6364 ( .B(n6190), .A(n6198), .Z(n6188) );
  IV U6365 ( .A(n6194), .Z(n6198) );
  IV U6366 ( .A(n6187), .Z(n6190) );
  XNOR U6367 ( .A(n6193), .B(n6200), .Z(n6187) );
  XOR U6368 ( .A(n6201), .B(n6197), .Z(n6200) );
  NAND U6369 ( .A(n6189), .B(n6185), .Z(n6197) );
  XNOR U6370 ( .A(n6178), .B(n6199), .Z(n6185) );
  XOR U6371 ( .A(n6202), .B(n6203), .Z(n6199) );
  XOR U6372 ( .A(n6204), .B(n6205), .Z(n6203) );
  XNOR U6373 ( .A(n6171), .B(n6206), .Z(n6205) );
  XNOR U6374 ( .A(n6207), .B(n6208), .Z(n6202) );
  XNOR U6375 ( .A(n6209), .B(n6210), .Z(n6208) );
  ANDN U6376 ( .B(n6149), .A(n5726), .Z(n6209) );
  XNOR U6377 ( .A(n6194), .B(n6181), .Z(n6189) );
  XOR U6378 ( .A(n6211), .B(n6212), .Z(n6194) );
  XNOR U6379 ( .A(n6213), .B(n6206), .Z(n6212) );
  XOR U6380 ( .A(n6214), .B(n6215), .Z(n6206) );
  XNOR U6381 ( .A(n6216), .B(n6217), .Z(n6215) );
  NAND U6382 ( .A(n5792), .B(n6153), .Z(n6217) );
  XNOR U6383 ( .A(n6218), .B(n6219), .Z(n6211) );
  ANDN U6384 ( .B(n6220), .A(n5786), .Z(n6218) );
  ANDN U6385 ( .B(n6178), .A(n6181), .Z(n6201) );
  XOR U6386 ( .A(n6181), .B(n6178), .Z(n6193) );
  XNOR U6387 ( .A(n6221), .B(n6222), .Z(n6178) );
  XNOR U6388 ( .A(n6214), .B(n6223), .Z(n6222) );
  XNOR U6389 ( .A(n6213), .B(n6149), .Z(n6223) );
  XNOR U6390 ( .A(n6224), .B(n6225), .Z(n6221) );
  XNOR U6391 ( .A(n6226), .B(n6210), .Z(n6225) );
  OR U6392 ( .A(n6172), .B(n6160), .Z(n6210) );
  XNOR U6393 ( .A(n6224), .B(n6207), .Z(n6160) );
  XNOR U6394 ( .A(n6149), .B(n6171), .Z(n6172) );
  ANDN U6395 ( .B(n6171), .A(n6162), .Z(n6226) );
  XOR U6396 ( .A(n6227), .B(n6228), .Z(n6181) );
  XOR U6397 ( .A(n6214), .B(n6204), .Z(n6228) );
  XOR U6398 ( .A(n6156), .B(n5731), .Z(n6204) );
  XOR U6399 ( .A(n6229), .B(n6216), .Z(n6214) );
  NANDN U6400 ( .A(n6166), .B(n6174), .Z(n6216) );
  XOR U6401 ( .A(n6182), .B(n6153), .Z(n6174) );
  XNOR U6402 ( .A(n6220), .B(n6230), .Z(n6171) );
  XNOR U6403 ( .A(n6231), .B(n6232), .Z(n6230) );
  XOR U6404 ( .A(n6168), .B(n5792), .Z(n6166) );
  XNOR U6405 ( .A(n6162), .B(n6156), .Z(n5792) );
  IV U6406 ( .A(n6207), .Z(n6162) );
  XOR U6407 ( .A(n6233), .B(n6234), .Z(n6207) );
  XOR U6408 ( .A(n6235), .B(n6236), .Z(n6234) );
  XOR U6409 ( .A(n6224), .B(n6237), .Z(n6233) );
  ANDN U6410 ( .B(n6182), .A(n6168), .Z(n6229) );
  XNOR U6411 ( .A(n6224), .B(n6238), .Z(n6168) );
  XOR U6412 ( .A(n6220), .B(n6149), .Z(n6182) );
  XNOR U6413 ( .A(n6239), .B(n6240), .Z(n6149) );
  XOR U6414 ( .A(n6241), .B(n6236), .Z(n6240) );
  XNOR U6415 ( .A(n6242), .B(n6243), .Z(n6236) );
  XOR U6416 ( .A(n6244), .B(n6245), .Z(n6242) );
  XNOR U6417 ( .A(key[300]), .B(n6246), .Z(n6245) );
  IV U6418 ( .A(n5666), .Z(n6220) );
  XOR U6419 ( .A(n6213), .B(n6247), .Z(n6227) );
  XNOR U6420 ( .A(n6248), .B(n6219), .Z(n6247) );
  OR U6421 ( .A(n5733), .B(n6157), .Z(n6219) );
  XNOR U6422 ( .A(n6238), .B(n6156), .Z(n6157) );
  XNOR U6423 ( .A(n5666), .B(n5731), .Z(n5733) );
  ANDN U6424 ( .B(n6156), .A(n5731), .Z(n6248) );
  XOR U6425 ( .A(n6239), .B(n6249), .Z(n5731) );
  XOR U6426 ( .A(n6231), .B(n6250), .Z(n6249) );
  XOR U6427 ( .A(n6241), .B(n6239), .Z(n6156) );
  XNOR U6428 ( .A(n5786), .B(n5666), .Z(n6213) );
  XOR U6429 ( .A(n6239), .B(n6251), .Z(n5666) );
  XNOR U6430 ( .A(n6241), .B(n6235), .Z(n6251) );
  XOR U6431 ( .A(n6252), .B(n6253), .Z(n6235) );
  XNOR U6432 ( .A(n6254), .B(n6255), .Z(n6253) );
  XNOR U6433 ( .A(key[303]), .B(n6256), .Z(n6252) );
  XNOR U6434 ( .A(n6257), .B(n6258), .Z(n6239) );
  XNOR U6435 ( .A(n6259), .B(n6260), .Z(n6258) );
  XOR U6436 ( .A(n6261), .B(n6262), .Z(n6257) );
  XNOR U6437 ( .A(key[301]), .B(n6263), .Z(n6262) );
  IV U6438 ( .A(n6238), .Z(n5786) );
  XNOR U6439 ( .A(n6232), .B(n6264), .Z(n6238) );
  XOR U6440 ( .A(n6237), .B(n6250), .Z(n6264) );
  IV U6441 ( .A(n6241), .Z(n6250) );
  XOR U6442 ( .A(n6265), .B(n6266), .Z(n6241) );
  XNOR U6443 ( .A(n6267), .B(n5726), .Z(n6266) );
  IV U6444 ( .A(n6224), .Z(n5726) );
  XOR U6445 ( .A(n6268), .B(n6269), .Z(n6224) );
  XOR U6446 ( .A(n6270), .B(n6271), .Z(n6269) );
  XOR U6447 ( .A(n6272), .B(n6273), .Z(n6268) );
  XOR U6448 ( .A(key[296]), .B(n6274), .Z(n6273) );
  XOR U6449 ( .A(n6275), .B(n6276), .Z(n6265) );
  XNOR U6450 ( .A(key[302]), .B(n6277), .Z(n6276) );
  XOR U6451 ( .A(n6278), .B(n6279), .Z(n6237) );
  XNOR U6452 ( .A(n6231), .B(n6280), .Z(n6279) );
  XOR U6453 ( .A(n6281), .B(n6282), .Z(n6280) );
  XOR U6454 ( .A(n6283), .B(n6284), .Z(n6231) );
  XNOR U6455 ( .A(n6285), .B(n6286), .Z(n6284) );
  XOR U6456 ( .A(n6287), .B(n6288), .Z(n6283) );
  XNOR U6457 ( .A(key[297]), .B(n6289), .Z(n6288) );
  XNOR U6458 ( .A(n6290), .B(n6291), .Z(n6278) );
  XNOR U6459 ( .A(key[299]), .B(n6292), .Z(n6291) );
  XOR U6460 ( .A(n6293), .B(n6294), .Z(n6232) );
  XOR U6461 ( .A(n6295), .B(n6296), .Z(n6294) );
  XNOR U6462 ( .A(n6297), .B(n6298), .Z(n6293) );
  XOR U6463 ( .A(key[298]), .B(n6299), .Z(n6298) );
  XOR U6464 ( .A(n5708), .B(n6123), .Z(n5624) );
  XNOR U6465 ( .A(n6139), .B(n6300), .Z(n6123) );
  XOR U6466 ( .A(n6301), .B(n5704), .Z(n6300) );
  OR U6467 ( .A(n6302), .B(n6127), .Z(n5704) );
  XNOR U6468 ( .A(n5707), .B(n6122), .Z(n6127) );
  ANDN U6469 ( .B(n6303), .A(n6304), .Z(n6301) );
  XNOR U6470 ( .A(n5702), .B(n6305), .Z(n5708) );
  XOR U6471 ( .A(n6306), .B(n6141), .Z(n6305) );
  XNOR U6472 ( .A(n5836), .B(n5712), .Z(n5833) );
  NOR U6473 ( .A(n6308), .B(n5836), .Z(n6306) );
  XNOR U6474 ( .A(n6139), .B(n6309), .Z(n5702) );
  XNOR U6475 ( .A(n6310), .B(n6311), .Z(n6309) );
  NAND U6476 ( .A(n6133), .B(n6312), .Z(n6311) );
  XOR U6477 ( .A(n6313), .B(n6310), .Z(n6139) );
  OR U6478 ( .A(n6135), .B(n6314), .Z(n6310) );
  XNOR U6479 ( .A(n6315), .B(n6133), .Z(n6135) );
  XOR U6480 ( .A(n6122), .B(n5712), .Z(n6133) );
  XOR U6481 ( .A(n6316), .B(n6317), .Z(n5712) );
  NANDN U6482 ( .A(n6318), .B(n6319), .Z(n6317) );
  IV U6483 ( .A(n6304), .Z(n6122) );
  XNOR U6484 ( .A(n6320), .B(n6321), .Z(n6304) );
  NANDN U6485 ( .A(n6318), .B(n6322), .Z(n6321) );
  ANDN U6486 ( .B(n6315), .A(n6323), .Z(n6313) );
  IV U6487 ( .A(n6138), .Z(n6315) );
  XOR U6488 ( .A(n5836), .B(n5707), .Z(n6138) );
  XNOR U6489 ( .A(n6324), .B(n6320), .Z(n5707) );
  NANDN U6490 ( .A(n6325), .B(n6326), .Z(n6320) );
  XOR U6491 ( .A(n6322), .B(n6327), .Z(n6326) );
  ANDN U6492 ( .B(n6327), .A(n6328), .Z(n6324) );
  XOR U6493 ( .A(n6329), .B(n6316), .Z(n5836) );
  NANDN U6494 ( .A(n6325), .B(n6330), .Z(n6316) );
  XOR U6495 ( .A(n6331), .B(n6319), .Z(n6330) );
  XNOR U6496 ( .A(n6332), .B(n6333), .Z(n6318) );
  XOR U6497 ( .A(n6334), .B(n6335), .Z(n6333) );
  XNOR U6498 ( .A(n6336), .B(n6337), .Z(n6332) );
  XNOR U6499 ( .A(n6338), .B(n6339), .Z(n6337) );
  ANDN U6500 ( .B(n6331), .A(n6335), .Z(n6338) );
  ANDN U6501 ( .B(n6331), .A(n6328), .Z(n6329) );
  XNOR U6502 ( .A(n6334), .B(n6340), .Z(n6328) );
  XOR U6503 ( .A(n6341), .B(n6339), .Z(n6340) );
  NAND U6504 ( .A(n6342), .B(n6343), .Z(n6339) );
  XNOR U6505 ( .A(n6336), .B(n6319), .Z(n6343) );
  IV U6506 ( .A(n6331), .Z(n6336) );
  XNOR U6507 ( .A(n6322), .B(n6335), .Z(n6342) );
  IV U6508 ( .A(n6327), .Z(n6335) );
  XOR U6509 ( .A(n6344), .B(n6345), .Z(n6327) );
  XNOR U6510 ( .A(n6346), .B(n6347), .Z(n6345) );
  XNOR U6511 ( .A(n6348), .B(n6349), .Z(n6344) );
  NOR U6512 ( .A(n5835), .B(n6308), .Z(n6348) );
  AND U6513 ( .A(n6319), .B(n6322), .Z(n6341) );
  XNOR U6514 ( .A(n6319), .B(n6322), .Z(n6334) );
  XNOR U6515 ( .A(n6350), .B(n6351), .Z(n6322) );
  XNOR U6516 ( .A(n6352), .B(n6347), .Z(n6351) );
  XOR U6517 ( .A(n6353), .B(n6354), .Z(n6350) );
  XNOR U6518 ( .A(n6355), .B(n6349), .Z(n6354) );
  OR U6519 ( .A(n5834), .B(n6307), .Z(n6349) );
  XNOR U6520 ( .A(n6308), .B(n6143), .Z(n6307) );
  XNOR U6521 ( .A(n5835), .B(n5713), .Z(n5834) );
  ANDN U6522 ( .B(n6356), .A(n6143), .Z(n6355) );
  XNOR U6523 ( .A(n6357), .B(n6358), .Z(n6319) );
  XNOR U6524 ( .A(n6347), .B(n6359), .Z(n6358) );
  XOR U6525 ( .A(n6126), .B(n6353), .Z(n6359) );
  XNOR U6526 ( .A(n6308), .B(n6360), .Z(n6347) );
  XNOR U6527 ( .A(n6361), .B(n6362), .Z(n6357) );
  XNOR U6528 ( .A(n6363), .B(n6364), .Z(n6362) );
  ANDN U6529 ( .B(n6303), .A(n6121), .Z(n6363) );
  XNOR U6530 ( .A(n6365), .B(n6366), .Z(n6331) );
  XNOR U6531 ( .A(n6352), .B(n6367), .Z(n6366) );
  XNOR U6532 ( .A(n6121), .B(n6346), .Z(n6367) );
  XOR U6533 ( .A(n6353), .B(n6368), .Z(n6346) );
  XNOR U6534 ( .A(n6369), .B(n6370), .Z(n6368) );
  NAND U6535 ( .A(n6312), .B(n6132), .Z(n6370) );
  XNOR U6536 ( .A(n6371), .B(n6369), .Z(n6353) );
  NANDN U6537 ( .A(n6314), .B(n6136), .Z(n6369) );
  XOR U6538 ( .A(n6137), .B(n6132), .Z(n6136) );
  XNOR U6539 ( .A(n6372), .B(n5713), .Z(n6132) );
  XOR U6540 ( .A(n6323), .B(n6312), .Z(n6314) );
  XOR U6541 ( .A(n6303), .B(n6373), .Z(n6312) );
  ANDN U6542 ( .B(n6137), .A(n6323), .Z(n6371) );
  XOR U6543 ( .A(n6361), .B(n6308), .Z(n6323) );
  XOR U6544 ( .A(n6374), .B(n6375), .Z(n6308) );
  XNOR U6545 ( .A(n6376), .B(n6377), .Z(n6375) );
  XOR U6546 ( .A(n6378), .B(n6360), .Z(n6137) );
  XOR U6547 ( .A(n6373), .B(n6356), .Z(n6352) );
  IV U6548 ( .A(n5713), .Z(n6356) );
  XOR U6549 ( .A(n6379), .B(n6380), .Z(n5713) );
  XNOR U6550 ( .A(n6381), .B(n6377), .Z(n6380) );
  IV U6551 ( .A(n6143), .Z(n6373) );
  XOR U6552 ( .A(n6377), .B(n6382), .Z(n6143) );
  XNOR U6553 ( .A(n6303), .B(n6383), .Z(n6365) );
  XNOR U6554 ( .A(n6384), .B(n6364), .Z(n6383) );
  OR U6555 ( .A(n6128), .B(n6302), .Z(n6364) );
  XNOR U6556 ( .A(n6361), .B(n6303), .Z(n6302) );
  XOR U6557 ( .A(n6126), .B(n6372), .Z(n6128) );
  IV U6558 ( .A(n6121), .Z(n6372) );
  XOR U6559 ( .A(n6360), .B(n6385), .Z(n6121) );
  XNOR U6560 ( .A(n6381), .B(n6374), .Z(n6385) );
  XOR U6561 ( .A(n6386), .B(n6387), .Z(n6374) );
  XOR U6562 ( .A(n6388), .B(n6389), .Z(n6387) );
  XOR U6563 ( .A(key[258]), .B(n6390), .Z(n6386) );
  IV U6564 ( .A(n5835), .Z(n6360) );
  XOR U6565 ( .A(n6379), .B(n6391), .Z(n5835) );
  XOR U6566 ( .A(n6377), .B(n6392), .Z(n6391) );
  ANDN U6567 ( .B(n6378), .A(n5706), .Z(n6384) );
  IV U6568 ( .A(n6126), .Z(n6378) );
  XOR U6569 ( .A(n6379), .B(n6393), .Z(n6126) );
  XOR U6570 ( .A(n6377), .B(n6394), .Z(n6393) );
  XOR U6571 ( .A(n6395), .B(n6396), .Z(n6377) );
  XOR U6572 ( .A(n6397), .B(n5706), .Z(n6396) );
  IV U6573 ( .A(n6361), .Z(n5706) );
  XOR U6574 ( .A(n6398), .B(n6399), .Z(n6395) );
  XNOR U6575 ( .A(key[262]), .B(n6400), .Z(n6399) );
  IV U6576 ( .A(n6382), .Z(n6379) );
  XOR U6577 ( .A(n6401), .B(n6402), .Z(n6382) );
  XOR U6578 ( .A(n6403), .B(n6404), .Z(n6402) );
  XNOR U6579 ( .A(key[261]), .B(n6405), .Z(n6401) );
  XOR U6580 ( .A(n6406), .B(n6407), .Z(n6303) );
  XNOR U6581 ( .A(n6394), .B(n6392), .Z(n6407) );
  XNOR U6582 ( .A(n6408), .B(n6409), .Z(n6392) );
  XNOR U6583 ( .A(n6410), .B(n6411), .Z(n6409) );
  XOR U6584 ( .A(key[263]), .B(n6412), .Z(n6408) );
  XNOR U6585 ( .A(n6413), .B(n6414), .Z(n6394) );
  XNOR U6586 ( .A(n6415), .B(n6416), .Z(n6414) );
  XNOR U6587 ( .A(n6417), .B(n6418), .Z(n6413) );
  XNOR U6588 ( .A(key[260]), .B(n6419), .Z(n6418) );
  XOR U6589 ( .A(n6361), .B(n6376), .Z(n6406) );
  XOR U6590 ( .A(n6420), .B(n6421), .Z(n6376) );
  XNOR U6591 ( .A(n6381), .B(n6422), .Z(n6421) );
  XOR U6592 ( .A(n6423), .B(n6424), .Z(n6422) );
  XOR U6593 ( .A(n6425), .B(n6426), .Z(n6381) );
  XOR U6594 ( .A(n6427), .B(n6428), .Z(n6426) );
  XNOR U6595 ( .A(key[257]), .B(n6429), .Z(n6425) );
  XOR U6596 ( .A(n6430), .B(n6431), .Z(n6420) );
  XNOR U6597 ( .A(key[259]), .B(n6432), .Z(n6431) );
  XOR U6598 ( .A(n6433), .B(n6434), .Z(n6361) );
  XNOR U6599 ( .A(n6435), .B(n6436), .Z(n6434) );
  XOR U6600 ( .A(key[256]), .B(n6437), .Z(n6433) );
  XOR U6601 ( .A(n5366), .B(n398), .Z(n1015) );
  XOR U6602 ( .A(n5508), .B(n5343), .Z(n398) );
  XOR U6603 ( .A(n5381), .B(n6438), .Z(n5343) );
  XNOR U6604 ( .A(n6439), .B(n5505), .Z(n6438) );
  XOR U6605 ( .A(n6441), .B(n5348), .Z(n5462) );
  ANDN U6606 ( .B(n6442), .A(n5465), .Z(n6439) );
  IV U6607 ( .A(n6441), .Z(n5465) );
  XNOR U6608 ( .A(n5503), .B(n6443), .Z(n5381) );
  XNOR U6609 ( .A(n6444), .B(n6445), .Z(n6443) );
  NANDN U6610 ( .A(n5501), .B(n6446), .Z(n6445) );
  IV U6611 ( .A(n5406), .Z(n5508) );
  XNOR U6612 ( .A(n5503), .B(n6447), .Z(n5406) );
  XOR U6613 ( .A(n6448), .B(n5383), .Z(n6447) );
  OR U6614 ( .A(n6449), .B(n5513), .Z(n5383) );
  XNOR U6615 ( .A(n5386), .B(n5512), .Z(n5513) );
  ANDN U6616 ( .B(n6450), .A(n6451), .Z(n6448) );
  XOR U6617 ( .A(n6452), .B(n6444), .Z(n5503) );
  OR U6618 ( .A(n5516), .B(n6453), .Z(n6444) );
  XNOR U6619 ( .A(n5519), .B(n5501), .Z(n5516) );
  XNOR U6620 ( .A(n5512), .B(n5348), .Z(n5501) );
  XOR U6621 ( .A(n6454), .B(n6455), .Z(n5348) );
  NANDN U6622 ( .A(n6456), .B(n6457), .Z(n6455) );
  IV U6623 ( .A(n6451), .Z(n5512) );
  XNOR U6624 ( .A(n6458), .B(n6459), .Z(n6451) );
  NANDN U6625 ( .A(n6456), .B(n6460), .Z(n6459) );
  NOR U6626 ( .A(n5519), .B(n6461), .Z(n6452) );
  XNOR U6627 ( .A(n6441), .B(n5386), .Z(n5519) );
  XNOR U6628 ( .A(n6462), .B(n6458), .Z(n5386) );
  NANDN U6629 ( .A(n6463), .B(n6464), .Z(n6458) );
  XOR U6630 ( .A(n6460), .B(n6465), .Z(n6464) );
  ANDN U6631 ( .B(n6465), .A(n6466), .Z(n6462) );
  XNOR U6632 ( .A(n6467), .B(n6454), .Z(n6441) );
  NANDN U6633 ( .A(n6463), .B(n6468), .Z(n6454) );
  XOR U6634 ( .A(n6469), .B(n6457), .Z(n6468) );
  XNOR U6635 ( .A(n6470), .B(n6471), .Z(n6456) );
  XOR U6636 ( .A(n6472), .B(n6473), .Z(n6471) );
  XNOR U6637 ( .A(n6474), .B(n6475), .Z(n6470) );
  XNOR U6638 ( .A(n6476), .B(n6477), .Z(n6475) );
  ANDN U6639 ( .B(n6469), .A(n6473), .Z(n6476) );
  ANDN U6640 ( .B(n6469), .A(n6466), .Z(n6467) );
  XNOR U6641 ( .A(n6472), .B(n6478), .Z(n6466) );
  XOR U6642 ( .A(n6479), .B(n6477), .Z(n6478) );
  NAND U6643 ( .A(n6480), .B(n6481), .Z(n6477) );
  XNOR U6644 ( .A(n6474), .B(n6457), .Z(n6481) );
  IV U6645 ( .A(n6469), .Z(n6474) );
  XNOR U6646 ( .A(n6460), .B(n6473), .Z(n6480) );
  IV U6647 ( .A(n6465), .Z(n6473) );
  XOR U6648 ( .A(n6482), .B(n6483), .Z(n6465) );
  XNOR U6649 ( .A(n6484), .B(n6485), .Z(n6483) );
  XNOR U6650 ( .A(n6486), .B(n6487), .Z(n6482) );
  ANDN U6651 ( .B(n6442), .A(n6488), .Z(n6486) );
  AND U6652 ( .A(n6457), .B(n6460), .Z(n6479) );
  XNOR U6653 ( .A(n6457), .B(n6460), .Z(n6472) );
  XNOR U6654 ( .A(n6489), .B(n6490), .Z(n6460) );
  XNOR U6655 ( .A(n6491), .B(n6485), .Z(n6490) );
  XOR U6656 ( .A(n6492), .B(n6493), .Z(n6489) );
  XNOR U6657 ( .A(n6494), .B(n6487), .Z(n6493) );
  OR U6658 ( .A(n5463), .B(n6440), .Z(n6487) );
  XNOR U6659 ( .A(n6442), .B(n6495), .Z(n6440) );
  XNOR U6660 ( .A(n6488), .B(n5349), .Z(n5463) );
  ANDN U6661 ( .B(n6496), .A(n5507), .Z(n6494) );
  XNOR U6662 ( .A(n6497), .B(n6498), .Z(n6457) );
  XNOR U6663 ( .A(n6485), .B(n6499), .Z(n6498) );
  XOR U6664 ( .A(n5497), .B(n6492), .Z(n6499) );
  XNOR U6665 ( .A(n6442), .B(n6488), .Z(n6485) );
  XNOR U6666 ( .A(n6500), .B(n6501), .Z(n6497) );
  XNOR U6667 ( .A(n6502), .B(n6503), .Z(n6501) );
  ANDN U6668 ( .B(n6450), .A(n5511), .Z(n6502) );
  XNOR U6669 ( .A(n6504), .B(n6505), .Z(n6469) );
  XNOR U6670 ( .A(n6491), .B(n6506), .Z(n6505) );
  XNOR U6671 ( .A(n5511), .B(n6484), .Z(n6506) );
  XOR U6672 ( .A(n6492), .B(n6507), .Z(n6484) );
  XNOR U6673 ( .A(n6508), .B(n6509), .Z(n6507) );
  NAND U6674 ( .A(n6446), .B(n5502), .Z(n6509) );
  XNOR U6675 ( .A(n6510), .B(n6508), .Z(n6492) );
  NANDN U6676 ( .A(n6453), .B(n5517), .Z(n6508) );
  XOR U6677 ( .A(n5518), .B(n5502), .Z(n5517) );
  XNOR U6678 ( .A(n6511), .B(n5349), .Z(n5502) );
  XOR U6679 ( .A(n6461), .B(n6446), .Z(n6453) );
  XOR U6680 ( .A(n6450), .B(n6495), .Z(n6446) );
  ANDN U6681 ( .B(n5518), .A(n6461), .Z(n6510) );
  XNOR U6682 ( .A(n6500), .B(n6442), .Z(n6461) );
  XNOR U6683 ( .A(n6512), .B(n6513), .Z(n6442) );
  XNOR U6684 ( .A(n6514), .B(n6515), .Z(n6513) );
  XOR U6685 ( .A(n6516), .B(n5464), .Z(n5518) );
  XOR U6686 ( .A(n6495), .B(n6496), .Z(n6491) );
  IV U6687 ( .A(n5349), .Z(n6496) );
  XOR U6688 ( .A(n6517), .B(n6518), .Z(n5349) );
  XNOR U6689 ( .A(n6519), .B(n6515), .Z(n6518) );
  IV U6690 ( .A(n5507), .Z(n6495) );
  XOR U6691 ( .A(n6515), .B(n6520), .Z(n5507) );
  XNOR U6692 ( .A(n6450), .B(n6521), .Z(n6504) );
  XNOR U6693 ( .A(n6522), .B(n6503), .Z(n6521) );
  OR U6694 ( .A(n5514), .B(n6449), .Z(n6503) );
  XNOR U6695 ( .A(n6500), .B(n6450), .Z(n6449) );
  XOR U6696 ( .A(n5497), .B(n6511), .Z(n5514) );
  IV U6697 ( .A(n5511), .Z(n6511) );
  XOR U6698 ( .A(n5464), .B(n6523), .Z(n5511) );
  XNOR U6699 ( .A(n6519), .B(n6512), .Z(n6523) );
  XOR U6700 ( .A(n6524), .B(n6525), .Z(n6512) );
  XOR U6701 ( .A(n3642), .B(n2719), .Z(n6525) );
  XOR U6702 ( .A(n2681), .B(n3641), .Z(n2719) );
  XOR U6703 ( .A(key[402]), .B(n2721), .Z(n6524) );
  XOR U6704 ( .A(n3646), .B(n3650), .Z(n2721) );
  XOR U6705 ( .A(n6526), .B(n6527), .Z(n3646) );
  XOR U6706 ( .A(n6528), .B(n6529), .Z(n6527) );
  XNOR U6707 ( .A(n6530), .B(n6531), .Z(n6526) );
  IV U6708 ( .A(n6488), .Z(n5464) );
  XOR U6709 ( .A(n6517), .B(n6532), .Z(n6488) );
  XOR U6710 ( .A(n6515), .B(n6533), .Z(n6532) );
  ANDN U6711 ( .B(n6516), .A(n5385), .Z(n6522) );
  IV U6712 ( .A(n5497), .Z(n6516) );
  XOR U6713 ( .A(n6517), .B(n6534), .Z(n5497) );
  XOR U6714 ( .A(n6515), .B(n6535), .Z(n6534) );
  XOR U6715 ( .A(n6536), .B(n6537), .Z(n6515) );
  XNOR U6716 ( .A(n3626), .B(n5385), .Z(n6537) );
  IV U6717 ( .A(n6500), .Z(n5385) );
  XNOR U6718 ( .A(n2695), .B(n6538), .Z(n3626) );
  XOR U6719 ( .A(n3622), .B(n2689), .Z(n2695) );
  XNOR U6720 ( .A(n6539), .B(n6540), .Z(n2689) );
  XOR U6721 ( .A(n6541), .B(n6542), .Z(n3622) );
  XNOR U6722 ( .A(n3620), .B(n6543), .Z(n6536) );
  XNOR U6723 ( .A(key[406]), .B(n5078), .Z(n6543) );
  XOR U6724 ( .A(n5067), .B(n3613), .Z(n5078) );
  XOR U6725 ( .A(n6544), .B(n6545), .Z(n3613) );
  XOR U6726 ( .A(n6546), .B(n6547), .Z(n6545) );
  XOR U6727 ( .A(n6548), .B(n6531), .Z(n6544) );
  IV U6728 ( .A(n6520), .Z(n6517) );
  XOR U6729 ( .A(n6549), .B(n6550), .Z(n6520) );
  XNOR U6730 ( .A(n5072), .B(n3619), .Z(n6550) );
  XNOR U6731 ( .A(n2696), .B(n3603), .Z(n3619) );
  XNOR U6732 ( .A(n6551), .B(n6552), .Z(n3603) );
  XNOR U6733 ( .A(n6553), .B(n6554), .Z(n6552) );
  XNOR U6734 ( .A(n6555), .B(n6556), .Z(n6551) );
  XOR U6735 ( .A(n6557), .B(n6558), .Z(n6556) );
  ANDN U6736 ( .B(n6559), .A(n6560), .Z(n6558) );
  XOR U6737 ( .A(n6561), .B(n6562), .Z(n2696) );
  XNOR U6738 ( .A(n6563), .B(n6564), .Z(n6562) );
  XNOR U6739 ( .A(n6565), .B(n6566), .Z(n6561) );
  XOR U6740 ( .A(n6567), .B(n6568), .Z(n6566) );
  ANDN U6741 ( .B(n6569), .A(n6570), .Z(n6568) );
  XNOR U6742 ( .A(key[405]), .B(n5076), .Z(n6549) );
  XNOR U6743 ( .A(n3633), .B(n3620), .Z(n5076) );
  XOR U6744 ( .A(n6571), .B(n6572), .Z(n3620) );
  XOR U6745 ( .A(n6546), .B(n6529), .Z(n3633) );
  XNOR U6746 ( .A(n6573), .B(n6574), .Z(n6529) );
  XNOR U6747 ( .A(n6575), .B(n6576), .Z(n6574) );
  NOR U6748 ( .A(n6577), .B(n6578), .Z(n6575) );
  XOR U6749 ( .A(n6579), .B(n6580), .Z(n6450) );
  XNOR U6750 ( .A(n6535), .B(n6533), .Z(n6580) );
  XNOR U6751 ( .A(n6581), .B(n6582), .Z(n6533) );
  XOR U6752 ( .A(n6538), .B(n3614), .Z(n6582) );
  XNOR U6753 ( .A(n5077), .B(n3634), .Z(n3614) );
  XNOR U6754 ( .A(n6583), .B(n6584), .Z(n3634) );
  XOR U6755 ( .A(n6585), .B(n6554), .Z(n6584) );
  XNOR U6756 ( .A(n6586), .B(n6587), .Z(n6554) );
  XNOR U6757 ( .A(n6588), .B(n6589), .Z(n6587) );
  NANDN U6758 ( .A(n6590), .B(n6591), .Z(n6589) );
  XNOR U6759 ( .A(n6592), .B(n6541), .Z(n6583) );
  XOR U6760 ( .A(n6593), .B(n6594), .Z(n5077) );
  XOR U6761 ( .A(n6539), .B(n6564), .Z(n6594) );
  XNOR U6762 ( .A(n6595), .B(n6596), .Z(n6564) );
  XNOR U6763 ( .A(n6597), .B(n6598), .Z(n6596) );
  OR U6764 ( .A(n6599), .B(n6600), .Z(n6598) );
  XOR U6765 ( .A(n6601), .B(n6602), .Z(n6593) );
  XNOR U6766 ( .A(n2728), .B(n5068), .Z(n6538) );
  XNOR U6767 ( .A(n6603), .B(n6604), .Z(n5068) );
  XOR U6768 ( .A(n6605), .B(n6606), .Z(n6604) );
  XOR U6769 ( .A(n6607), .B(n6571), .Z(n6603) );
  XOR U6770 ( .A(key[407]), .B(n5067), .Z(n6581) );
  XNOR U6771 ( .A(n6608), .B(n6609), .Z(n6535) );
  XOR U6772 ( .A(n5055), .B(n3601), .Z(n6609) );
  XNOR U6773 ( .A(n6610), .B(n6611), .Z(n3601) );
  XNOR U6774 ( .A(n3647), .B(n5072), .Z(n6611) );
  XNOR U6775 ( .A(n6612), .B(n6613), .Z(n5072) );
  XNOR U6776 ( .A(n6614), .B(n6606), .Z(n6613) );
  XNOR U6777 ( .A(n6615), .B(n6616), .Z(n6606) );
  XNOR U6778 ( .A(n6617), .B(n6618), .Z(n6616) );
  NANDN U6779 ( .A(n6619), .B(n6620), .Z(n6618) );
  XNOR U6780 ( .A(n6621), .B(n6622), .Z(n6612) );
  XOR U6781 ( .A(n6623), .B(n6624), .Z(n6622) );
  ANDN U6782 ( .B(n6625), .A(n6626), .Z(n6624) );
  XOR U6783 ( .A(n6555), .B(n3641), .Z(n3647) );
  XOR U6784 ( .A(n6627), .B(n6628), .Z(n3641) );
  XNOR U6785 ( .A(n2728), .B(n2710), .Z(n6610) );
  XOR U6786 ( .A(n6563), .B(n2681), .Z(n2710) );
  XNOR U6787 ( .A(n6601), .B(n6629), .Z(n2681) );
  IV U6788 ( .A(n6630), .Z(n6601) );
  XNOR U6789 ( .A(key[404]), .B(n5056), .Z(n6608) );
  XNOR U6790 ( .A(n5067), .B(n3618), .Z(n5056) );
  XNOR U6791 ( .A(n6631), .B(n6632), .Z(n3618) );
  XNOR U6792 ( .A(n6633), .B(n6547), .Z(n6632) );
  XNOR U6793 ( .A(n6634), .B(n6635), .Z(n6547) );
  XNOR U6794 ( .A(n6636), .B(n6637), .Z(n6635) );
  NANDN U6795 ( .A(n6638), .B(n6639), .Z(n6637) );
  XNOR U6796 ( .A(n6640), .B(n6641), .Z(n6631) );
  XOR U6797 ( .A(n6576), .B(n6642), .Z(n6641) );
  ANDN U6798 ( .B(n6643), .A(n6644), .Z(n6642) );
  ANDN U6799 ( .B(n6645), .A(n6646), .Z(n6576) );
  XOR U6800 ( .A(n6500), .B(n6514), .Z(n6579) );
  XOR U6801 ( .A(n6647), .B(n6648), .Z(n6514) );
  XNOR U6802 ( .A(n6519), .B(n6649), .Z(n6648) );
  XOR U6803 ( .A(n2680), .B(n3637), .Z(n6649) );
  XOR U6804 ( .A(n2728), .B(n5055), .Z(n3637) );
  XOR U6805 ( .A(n6621), .B(n3642), .Z(n5055) );
  XOR U6806 ( .A(n3651), .B(n2715), .Z(n2680) );
  XNOR U6807 ( .A(n6650), .B(n6651), .Z(n2715) );
  XOR U6808 ( .A(n6652), .B(n6540), .Z(n6651) );
  XNOR U6809 ( .A(n6653), .B(n6654), .Z(n6540) );
  XNOR U6810 ( .A(n6655), .B(n6567), .Z(n6654) );
  ANDN U6811 ( .B(n6656), .A(n6657), .Z(n6567) );
  NOR U6812 ( .A(n6658), .B(n6659), .Z(n6655) );
  XNOR U6813 ( .A(n6630), .B(n6602), .Z(n6650) );
  XNOR U6814 ( .A(n6660), .B(n6661), .Z(n3651) );
  XNOR U6815 ( .A(n6628), .B(n6542), .Z(n6661) );
  XNOR U6816 ( .A(n6662), .B(n6663), .Z(n6542) );
  XNOR U6817 ( .A(n6664), .B(n6557), .Z(n6663) );
  ANDN U6818 ( .B(n6665), .A(n6666), .Z(n6557) );
  NOR U6819 ( .A(n6667), .B(n6668), .Z(n6664) );
  XNOR U6820 ( .A(n6592), .B(n6669), .Z(n6660) );
  XOR U6821 ( .A(n6670), .B(n6671), .Z(n6519) );
  XOR U6822 ( .A(n2679), .B(n2727), .Z(n6671) );
  XNOR U6823 ( .A(n2720), .B(n3629), .Z(n2727) );
  XOR U6824 ( .A(n6628), .B(n6672), .Z(n3629) );
  XOR U6825 ( .A(n6592), .B(n6541), .Z(n6672) );
  XOR U6826 ( .A(n6627), .B(n6669), .Z(n6541) );
  XNOR U6827 ( .A(n6553), .B(n6673), .Z(n6669) );
  XNOR U6828 ( .A(n6674), .B(n6675), .Z(n6673) );
  NANDN U6829 ( .A(n6676), .B(n6677), .Z(n6675) );
  IV U6830 ( .A(n6678), .Z(n6627) );
  XNOR U6831 ( .A(n6674), .B(n6680), .Z(n6679) );
  NANDN U6832 ( .A(n6681), .B(n6591), .Z(n6680) );
  OR U6833 ( .A(n6682), .B(n6683), .Z(n6674) );
  XNOR U6834 ( .A(n6553), .B(n6684), .Z(n6662) );
  XNOR U6835 ( .A(n6685), .B(n6686), .Z(n6684) );
  NAND U6836 ( .A(n6687), .B(n6688), .Z(n6686) );
  XOR U6837 ( .A(n6689), .B(n6685), .Z(n6553) );
  NANDN U6838 ( .A(n6690), .B(n6691), .Z(n6685) );
  ANDN U6839 ( .B(n6692), .A(n6693), .Z(n6689) );
  IV U6840 ( .A(n6585), .Z(n6628) );
  XOR U6841 ( .A(n6694), .B(n6695), .Z(n6585) );
  XNOR U6842 ( .A(n6696), .B(n6697), .Z(n6695) );
  NANDN U6843 ( .A(n6698), .B(n6559), .Z(n6697) );
  XOR U6844 ( .A(n6539), .B(n6699), .Z(n2720) );
  XOR U6845 ( .A(n6630), .B(n6602), .Z(n6699) );
  XNOR U6846 ( .A(n6701), .B(n6702), .Z(n6700) );
  OR U6847 ( .A(n6599), .B(n6703), .Z(n6702) );
  XNOR U6848 ( .A(n6565), .B(n6704), .Z(n6653) );
  XNOR U6849 ( .A(n6705), .B(n6706), .Z(n6704) );
  NAND U6850 ( .A(n6707), .B(n6708), .Z(n6706) );
  XNOR U6851 ( .A(n6709), .B(n6710), .Z(n6630) );
  XNOR U6852 ( .A(n6711), .B(n6712), .Z(n6710) );
  NAND U6853 ( .A(n6713), .B(n6569), .Z(n6712) );
  XOR U6854 ( .A(n6714), .B(n6652), .Z(n6539) );
  XOR U6855 ( .A(n6565), .B(n6715), .Z(n6652) );
  XNOR U6856 ( .A(n6701), .B(n6716), .Z(n6715) );
  NANDN U6857 ( .A(n6717), .B(n6718), .Z(n6716) );
  OR U6858 ( .A(n6719), .B(n6720), .Z(n6701) );
  XOR U6859 ( .A(n6721), .B(n6705), .Z(n6565) );
  NANDN U6860 ( .A(n6722), .B(n6723), .Z(n6705) );
  AND U6861 ( .A(n6724), .B(n6725), .Z(n6721) );
  XOR U6862 ( .A(n3653), .B(n3642), .Z(n2679) );
  XNOR U6863 ( .A(n6726), .B(n6605), .Z(n3642) );
  XOR U6864 ( .A(key[401]), .B(n6727), .Z(n6670) );
  XNOR U6865 ( .A(n3650), .B(n6728), .Z(n6647) );
  XNOR U6866 ( .A(key[403]), .B(n5089), .Z(n6728) );
  XOR U6867 ( .A(n5067), .B(n3604), .Z(n5089) );
  XNOR U6868 ( .A(n6640), .B(n3653), .Z(n3604) );
  XOR U6869 ( .A(n6729), .B(n6530), .Z(n3653) );
  XOR U6870 ( .A(n6640), .B(n6730), .Z(n5067) );
  XNOR U6871 ( .A(n6634), .B(n6731), .Z(n6640) );
  XOR U6872 ( .A(n6732), .B(n6733), .Z(n6731) );
  NOR U6873 ( .A(n6734), .B(n6578), .Z(n6732) );
  XNOR U6874 ( .A(n6735), .B(n6736), .Z(n6634) );
  XNOR U6875 ( .A(n6737), .B(n6738), .Z(n6736) );
  NAND U6876 ( .A(n6739), .B(n6740), .Z(n6738) );
  XOR U6877 ( .A(n6741), .B(n6742), .Z(n3650) );
  XNOR U6878 ( .A(n6743), .B(n6744), .Z(n6572) );
  XNOR U6879 ( .A(n6745), .B(n6623), .Z(n6744) );
  ANDN U6880 ( .B(n6746), .A(n6747), .Z(n6623) );
  NOR U6881 ( .A(n6748), .B(n6749), .Z(n6745) );
  XOR U6882 ( .A(n6607), .B(n6750), .Z(n6741) );
  XOR U6883 ( .A(n6751), .B(n6752), .Z(n6500) );
  XNOR U6884 ( .A(n5091), .B(n2718), .Z(n6752) );
  XNOR U6885 ( .A(n3644), .B(n6727), .Z(n2718) );
  IV U6886 ( .A(n3630), .Z(n6727) );
  XOR U6887 ( .A(n6605), .B(n6753), .Z(n3630) );
  XOR U6888 ( .A(n6614), .B(n6754), .Z(n6750) );
  XNOR U6889 ( .A(n6755), .B(n6756), .Z(n6754) );
  NANDN U6890 ( .A(n6757), .B(n6758), .Z(n6756) );
  XNOR U6891 ( .A(n6755), .B(n6760), .Z(n6759) );
  NANDN U6892 ( .A(n6761), .B(n6620), .Z(n6760) );
  OR U6893 ( .A(n6762), .B(n6763), .Z(n6755) );
  XNOR U6894 ( .A(n6614), .B(n6764), .Z(n6743) );
  XNOR U6895 ( .A(n6765), .B(n6766), .Z(n6764) );
  NAND U6896 ( .A(n6767), .B(n6768), .Z(n6766) );
  XOR U6897 ( .A(n6769), .B(n6765), .Z(n6614) );
  NANDN U6898 ( .A(n6770), .B(n6771), .Z(n6765) );
  ANDN U6899 ( .B(n6772), .A(n6773), .Z(n6769) );
  XOR U6900 ( .A(n6774), .B(n6775), .Z(n6605) );
  XNOR U6901 ( .A(n6776), .B(n6777), .Z(n6775) );
  NANDN U6902 ( .A(n6778), .B(n6625), .Z(n6777) );
  XNOR U6903 ( .A(n6546), .B(n6779), .Z(n3644) );
  XOR U6904 ( .A(n6530), .B(n6531), .Z(n6779) );
  XNOR U6905 ( .A(n6781), .B(n6782), .Z(n6780) );
  NANDN U6906 ( .A(n6783), .B(n6639), .Z(n6782) );
  XNOR U6907 ( .A(n6633), .B(n6784), .Z(n6573) );
  XNOR U6908 ( .A(n6785), .B(n6786), .Z(n6784) );
  NAND U6909 ( .A(n6787), .B(n6739), .Z(n6786) );
  IV U6910 ( .A(n6548), .Z(n6530) );
  XOR U6911 ( .A(n6735), .B(n6788), .Z(n6548) );
  XNOR U6912 ( .A(n6733), .B(n6789), .Z(n6788) );
  NANDN U6913 ( .A(n6790), .B(n6643), .Z(n6789) );
  XNOR U6914 ( .A(n6578), .B(n6643), .Z(n6645) );
  XOR U6915 ( .A(n6729), .B(n6528), .Z(n6546) );
  XOR U6916 ( .A(n6633), .B(n6792), .Z(n6528) );
  XNOR U6917 ( .A(n6781), .B(n6793), .Z(n6792) );
  NANDN U6918 ( .A(n6794), .B(n6795), .Z(n6793) );
  OR U6919 ( .A(n6796), .B(n6797), .Z(n6781) );
  XOR U6920 ( .A(n6798), .B(n6785), .Z(n6633) );
  NANDN U6921 ( .A(n6799), .B(n6800), .Z(n6785) );
  ANDN U6922 ( .B(n6801), .A(n6802), .Z(n6798) );
  IV U6923 ( .A(n6730), .Z(n6729) );
  XNOR U6924 ( .A(n6735), .B(n6803), .Z(n6730) );
  XOR U6925 ( .A(n6804), .B(n6636), .Z(n6803) );
  OR U6926 ( .A(n6805), .B(n6796), .Z(n6636) );
  XNOR U6927 ( .A(n6639), .B(n6795), .Z(n6796) );
  ANDN U6928 ( .B(n6795), .A(n6806), .Z(n6804) );
  XOR U6929 ( .A(n6807), .B(n6737), .Z(n6735) );
  OR U6930 ( .A(n6799), .B(n6808), .Z(n6737) );
  XNOR U6931 ( .A(n6809), .B(n6739), .Z(n6799) );
  XOR U6932 ( .A(n6795), .B(n6643), .Z(n6739) );
  XOR U6933 ( .A(n6810), .B(n6811), .Z(n6643) );
  NANDN U6934 ( .A(n6812), .B(n6813), .Z(n6811) );
  XOR U6935 ( .A(n6814), .B(n6815), .Z(n6795) );
  NANDN U6936 ( .A(n6812), .B(n6816), .Z(n6815) );
  ANDN U6937 ( .B(n6809), .A(n6817), .Z(n6807) );
  IV U6938 ( .A(n6802), .Z(n6809) );
  XOR U6939 ( .A(n6578), .B(n6639), .Z(n6802) );
  XNOR U6940 ( .A(n6818), .B(n6814), .Z(n6639) );
  NANDN U6941 ( .A(n6819), .B(n6820), .Z(n6814) );
  XOR U6942 ( .A(n6816), .B(n6821), .Z(n6820) );
  ANDN U6943 ( .B(n6821), .A(n6822), .Z(n6818) );
  XOR U6944 ( .A(n6823), .B(n6810), .Z(n6578) );
  NANDN U6945 ( .A(n6819), .B(n6824), .Z(n6810) );
  XOR U6946 ( .A(n6825), .B(n6813), .Z(n6824) );
  XNOR U6947 ( .A(n6826), .B(n6827), .Z(n6812) );
  XOR U6948 ( .A(n6828), .B(n6829), .Z(n6827) );
  XNOR U6949 ( .A(n6830), .B(n6831), .Z(n6826) );
  XNOR U6950 ( .A(n6832), .B(n6833), .Z(n6831) );
  ANDN U6951 ( .B(n6825), .A(n6829), .Z(n6832) );
  ANDN U6952 ( .B(n6825), .A(n6822), .Z(n6823) );
  XNOR U6953 ( .A(n6828), .B(n6834), .Z(n6822) );
  XOR U6954 ( .A(n6835), .B(n6833), .Z(n6834) );
  NAND U6955 ( .A(n6836), .B(n6837), .Z(n6833) );
  XNOR U6956 ( .A(n6830), .B(n6813), .Z(n6837) );
  IV U6957 ( .A(n6825), .Z(n6830) );
  XNOR U6958 ( .A(n6816), .B(n6829), .Z(n6836) );
  IV U6959 ( .A(n6821), .Z(n6829) );
  XOR U6960 ( .A(n6838), .B(n6839), .Z(n6821) );
  XNOR U6961 ( .A(n6840), .B(n6841), .Z(n6839) );
  XNOR U6962 ( .A(n6842), .B(n6843), .Z(n6838) );
  NOR U6963 ( .A(n6577), .B(n6734), .Z(n6842) );
  AND U6964 ( .A(n6813), .B(n6816), .Z(n6835) );
  XNOR U6965 ( .A(n6813), .B(n6816), .Z(n6828) );
  XNOR U6966 ( .A(n6844), .B(n6845), .Z(n6816) );
  XNOR U6967 ( .A(n6846), .B(n6841), .Z(n6845) );
  XOR U6968 ( .A(n6847), .B(n6848), .Z(n6844) );
  XNOR U6969 ( .A(n6849), .B(n6843), .Z(n6848) );
  OR U6970 ( .A(n6646), .B(n6791), .Z(n6843) );
  XNOR U6971 ( .A(n6734), .B(n6790), .Z(n6791) );
  XNOR U6972 ( .A(n6577), .B(n6644), .Z(n6646) );
  ANDN U6973 ( .B(n6850), .A(n6790), .Z(n6849) );
  XNOR U6974 ( .A(n6851), .B(n6852), .Z(n6813) );
  XNOR U6975 ( .A(n6841), .B(n6853), .Z(n6852) );
  XOR U6976 ( .A(n6783), .B(n6847), .Z(n6853) );
  XNOR U6977 ( .A(n6734), .B(n6854), .Z(n6841) );
  XOR U6978 ( .A(n6638), .B(n6855), .Z(n6851) );
  XNOR U6979 ( .A(n6856), .B(n6857), .Z(n6855) );
  ANDN U6980 ( .B(n6858), .A(n6806), .Z(n6856) );
  XNOR U6981 ( .A(n6859), .B(n6860), .Z(n6825) );
  XNOR U6982 ( .A(n6846), .B(n6861), .Z(n6860) );
  XNOR U6983 ( .A(n6794), .B(n6840), .Z(n6861) );
  XOR U6984 ( .A(n6847), .B(n6862), .Z(n6840) );
  XNOR U6985 ( .A(n6863), .B(n6864), .Z(n6862) );
  NAND U6986 ( .A(n6740), .B(n6787), .Z(n6864) );
  XNOR U6987 ( .A(n6865), .B(n6863), .Z(n6847) );
  NANDN U6988 ( .A(n6808), .B(n6800), .Z(n6863) );
  XOR U6989 ( .A(n6801), .B(n6787), .Z(n6800) );
  XNOR U6990 ( .A(n6858), .B(n6644), .Z(n6787) );
  XOR U6991 ( .A(n6817), .B(n6740), .Z(n6808) );
  XNOR U6992 ( .A(n6806), .B(n6866), .Z(n6740) );
  ANDN U6993 ( .B(n6801), .A(n6817), .Z(n6865) );
  XNOR U6994 ( .A(n6638), .B(n6734), .Z(n6817) );
  XOR U6995 ( .A(n6867), .B(n6868), .Z(n6734) );
  XNOR U6996 ( .A(n6869), .B(n6870), .Z(n6868) );
  XOR U6997 ( .A(n6866), .B(n6850), .Z(n6846) );
  IV U6998 ( .A(n6644), .Z(n6850) );
  XOR U6999 ( .A(n6871), .B(n6872), .Z(n6644) );
  XNOR U7000 ( .A(n6873), .B(n6870), .Z(n6872) );
  IV U7001 ( .A(n6790), .Z(n6866) );
  XOR U7002 ( .A(n6870), .B(n6874), .Z(n6790) );
  XNOR U7003 ( .A(n6875), .B(n6876), .Z(n6859) );
  XNOR U7004 ( .A(n6877), .B(n6857), .Z(n6876) );
  OR U7005 ( .A(n6797), .B(n6805), .Z(n6857) );
  XNOR U7006 ( .A(n6638), .B(n6806), .Z(n6805) );
  IV U7007 ( .A(n6875), .Z(n6806) );
  XOR U7008 ( .A(n6783), .B(n6858), .Z(n6797) );
  IV U7009 ( .A(n6794), .Z(n6858) );
  XOR U7010 ( .A(n6854), .B(n6878), .Z(n6794) );
  XNOR U7011 ( .A(n6873), .B(n6867), .Z(n6878) );
  XOR U7012 ( .A(n6879), .B(n6880), .Z(n6867) );
  XNOR U7013 ( .A(n6881), .B(n6882), .Z(n6880) );
  XNOR U7014 ( .A(key[370]), .B(n6883), .Z(n6879) );
  IV U7015 ( .A(n6577), .Z(n6854) );
  XOR U7016 ( .A(n6871), .B(n6884), .Z(n6577) );
  XOR U7017 ( .A(n6870), .B(n6885), .Z(n6884) );
  NOR U7018 ( .A(n6783), .B(n6638), .Z(n6877) );
  XOR U7019 ( .A(n6871), .B(n6886), .Z(n6783) );
  XOR U7020 ( .A(n6870), .B(n6887), .Z(n6886) );
  XOR U7021 ( .A(n6888), .B(n6889), .Z(n6870) );
  XNOR U7022 ( .A(n6890), .B(n6073), .Z(n6889) );
  XOR U7023 ( .A(n6113), .B(n6891), .Z(n6073) );
  XNOR U7024 ( .A(n6892), .B(n6893), .Z(n6888) );
  XOR U7025 ( .A(key[374]), .B(n6638), .Z(n6893) );
  IV U7026 ( .A(n6874), .Z(n6871) );
  XOR U7027 ( .A(n6894), .B(n6895), .Z(n6874) );
  XNOR U7028 ( .A(n6896), .B(n6897), .Z(n6895) );
  XNOR U7029 ( .A(key[373]), .B(n6898), .Z(n6894) );
  XOR U7030 ( .A(n6899), .B(n6900), .Z(n6875) );
  XNOR U7031 ( .A(n6887), .B(n6885), .Z(n6900) );
  XNOR U7032 ( .A(n6901), .B(n6902), .Z(n6885) );
  XNOR U7033 ( .A(n6903), .B(n6904), .Z(n6902) );
  XNOR U7034 ( .A(key[375]), .B(n6113), .Z(n6901) );
  XNOR U7035 ( .A(n6905), .B(n6906), .Z(n6887) );
  XOR U7036 ( .A(n6907), .B(n6092), .Z(n6906) );
  XNOR U7037 ( .A(n6113), .B(n6908), .Z(n6092) );
  XNOR U7038 ( .A(n6909), .B(n6910), .Z(n6905) );
  XNOR U7039 ( .A(key[372]), .B(n6911), .Z(n6910) );
  XNOR U7040 ( .A(n6638), .B(n6869), .Z(n6899) );
  XOR U7041 ( .A(n6912), .B(n6913), .Z(n6869) );
  XNOR U7042 ( .A(n6914), .B(n6915), .Z(n6913) );
  XOR U7043 ( .A(n6873), .B(n6109), .Z(n6915) );
  XNOR U7044 ( .A(n6113), .B(n6916), .Z(n6109) );
  XOR U7045 ( .A(n6917), .B(n6918), .Z(n6873) );
  XOR U7046 ( .A(n6919), .B(n6065), .Z(n6918) );
  IV U7047 ( .A(n6920), .Z(n6065) );
  XNOR U7048 ( .A(key[369]), .B(n6921), .Z(n6917) );
  XNOR U7049 ( .A(n6922), .B(n6923), .Z(n6912) );
  XNOR U7050 ( .A(key[371]), .B(n6924), .Z(n6923) );
  XNOR U7051 ( .A(n6925), .B(n6926), .Z(n6638) );
  XOR U7052 ( .A(n6106), .B(n6114), .Z(n6926) );
  IV U7053 ( .A(n6927), .Z(n6114) );
  XNOR U7054 ( .A(key[368]), .B(n6928), .Z(n6925) );
  XOR U7055 ( .A(n6714), .B(n6563), .Z(n5091) );
  XNOR U7056 ( .A(n6595), .B(n6929), .Z(n6563) );
  XOR U7057 ( .A(n6930), .B(n6711), .Z(n6929) );
  XNOR U7058 ( .A(n6659), .B(n6569), .Z(n6656) );
  NOR U7059 ( .A(n6932), .B(n6659), .Z(n6930) );
  XNOR U7060 ( .A(n6709), .B(n6933), .Z(n6595) );
  XNOR U7061 ( .A(n6934), .B(n6935), .Z(n6933) );
  NAND U7062 ( .A(n6708), .B(n6936), .Z(n6935) );
  IV U7063 ( .A(n6629), .Z(n6714) );
  XNOR U7064 ( .A(n6709), .B(n6937), .Z(n6629) );
  XOR U7065 ( .A(n6938), .B(n6597), .Z(n6937) );
  OR U7066 ( .A(n6719), .B(n6939), .Z(n6597) );
  XNOR U7067 ( .A(n6599), .B(n6717), .Z(n6719) );
  NOR U7068 ( .A(n6940), .B(n6717), .Z(n6938) );
  XOR U7069 ( .A(n6941), .B(n6934), .Z(n6709) );
  OR U7070 ( .A(n6722), .B(n6942), .Z(n6934) );
  XNOR U7071 ( .A(n6724), .B(n6708), .Z(n6722) );
  XNOR U7072 ( .A(n6717), .B(n6569), .Z(n6708) );
  XOR U7073 ( .A(n6943), .B(n6944), .Z(n6569) );
  NANDN U7074 ( .A(n6945), .B(n6946), .Z(n6944) );
  XNOR U7075 ( .A(n6947), .B(n6948), .Z(n6717) );
  OR U7076 ( .A(n6945), .B(n6949), .Z(n6948) );
  ANDN U7077 ( .B(n6724), .A(n6950), .Z(n6941) );
  XOR U7078 ( .A(n6599), .B(n6659), .Z(n6724) );
  XOR U7079 ( .A(n6951), .B(n6943), .Z(n6659) );
  NANDN U7080 ( .A(n6952), .B(n6953), .Z(n6943) );
  ANDN U7081 ( .B(n6954), .A(n6955), .Z(n6951) );
  NANDN U7082 ( .A(n6952), .B(n6957), .Z(n6947) );
  XOR U7083 ( .A(n6958), .B(n6945), .Z(n6952) );
  XNOR U7084 ( .A(n6959), .B(n6960), .Z(n6945) );
  XOR U7085 ( .A(n6961), .B(n6954), .Z(n6960) );
  XNOR U7086 ( .A(n6962), .B(n6963), .Z(n6959) );
  XNOR U7087 ( .A(n6964), .B(n6965), .Z(n6963) );
  ANDN U7088 ( .B(n6954), .A(n6966), .Z(n6964) );
  IV U7089 ( .A(n6967), .Z(n6954) );
  ANDN U7090 ( .B(n6958), .A(n6966), .Z(n6956) );
  IV U7091 ( .A(n6962), .Z(n6966) );
  IV U7092 ( .A(n6955), .Z(n6958) );
  XNOR U7093 ( .A(n6961), .B(n6968), .Z(n6955) );
  XOR U7094 ( .A(n6969), .B(n6965), .Z(n6968) );
  NAND U7095 ( .A(n6957), .B(n6953), .Z(n6965) );
  XNOR U7096 ( .A(n6946), .B(n6967), .Z(n6953) );
  XOR U7097 ( .A(n6970), .B(n6971), .Z(n6967) );
  XOR U7098 ( .A(n6972), .B(n6973), .Z(n6971) );
  XNOR U7099 ( .A(n6718), .B(n6974), .Z(n6973) );
  XNOR U7100 ( .A(n6975), .B(n6976), .Z(n6970) );
  XNOR U7101 ( .A(n6977), .B(n6978), .Z(n6976) );
  ANDN U7102 ( .B(n6979), .A(n6600), .Z(n6977) );
  XNOR U7103 ( .A(n6962), .B(n6949), .Z(n6957) );
  XOR U7104 ( .A(n6980), .B(n6981), .Z(n6962) );
  XNOR U7105 ( .A(n6982), .B(n6974), .Z(n6981) );
  XOR U7106 ( .A(n6983), .B(n6984), .Z(n6974) );
  XNOR U7107 ( .A(n6985), .B(n6986), .Z(n6984) );
  NAND U7108 ( .A(n6936), .B(n6707), .Z(n6986) );
  XNOR U7109 ( .A(n6987), .B(n6988), .Z(n6980) );
  ANDN U7110 ( .B(n6989), .A(n6932), .Z(n6987) );
  ANDN U7111 ( .B(n6946), .A(n6949), .Z(n6969) );
  XOR U7112 ( .A(n6949), .B(n6946), .Z(n6961) );
  XNOR U7113 ( .A(n6990), .B(n6991), .Z(n6946) );
  XNOR U7114 ( .A(n6983), .B(n6992), .Z(n6991) );
  XOR U7115 ( .A(n6982), .B(n6703), .Z(n6992) );
  XOR U7116 ( .A(n6600), .B(n6993), .Z(n6990) );
  XNOR U7117 ( .A(n6994), .B(n6978), .Z(n6993) );
  OR U7118 ( .A(n6720), .B(n6939), .Z(n6978) );
  XNOR U7119 ( .A(n6600), .B(n6940), .Z(n6939) );
  XOR U7120 ( .A(n6703), .B(n6718), .Z(n6720) );
  ANDN U7121 ( .B(n6718), .A(n6940), .Z(n6994) );
  XOR U7122 ( .A(n6995), .B(n6996), .Z(n6949) );
  XOR U7123 ( .A(n6983), .B(n6972), .Z(n6996) );
  XOR U7124 ( .A(n6713), .B(n6570), .Z(n6972) );
  XOR U7125 ( .A(n6997), .B(n6985), .Z(n6983) );
  NANDN U7126 ( .A(n6942), .B(n6723), .Z(n6985) );
  XOR U7127 ( .A(n6725), .B(n6707), .Z(n6723) );
  XNOR U7128 ( .A(n6989), .B(n6998), .Z(n6718) );
  XNOR U7129 ( .A(n6999), .B(n7000), .Z(n6998) );
  XOR U7130 ( .A(n6950), .B(n6936), .Z(n6942) );
  XNOR U7131 ( .A(n6940), .B(n6713), .Z(n6936) );
  IV U7132 ( .A(n6975), .Z(n6940) );
  XOR U7133 ( .A(n7001), .B(n7002), .Z(n6975) );
  XOR U7134 ( .A(n7003), .B(n7004), .Z(n7002) );
  XNOR U7135 ( .A(n6600), .B(n7005), .Z(n7001) );
  ANDN U7136 ( .B(n6725), .A(n6950), .Z(n6997) );
  XNOR U7137 ( .A(n6600), .B(n6932), .Z(n6950) );
  XOR U7138 ( .A(n6989), .B(n6979), .Z(n6725) );
  IV U7139 ( .A(n6703), .Z(n6979) );
  XOR U7140 ( .A(n7006), .B(n7007), .Z(n6703) );
  XOR U7141 ( .A(n7008), .B(n7004), .Z(n7007) );
  XNOR U7142 ( .A(n7009), .B(n7010), .Z(n7004) );
  XNOR U7143 ( .A(n7011), .B(n6415), .Z(n7010) );
  XOR U7144 ( .A(n7012), .B(n7013), .Z(n6415) );
  XNOR U7145 ( .A(n7014), .B(n7015), .Z(n7009) );
  XNOR U7146 ( .A(key[284]), .B(n6417), .Z(n7015) );
  XOR U7147 ( .A(n7016), .B(n6405), .Z(n6417) );
  IV U7148 ( .A(n6658), .Z(n6989) );
  XOR U7149 ( .A(n6982), .B(n7017), .Z(n6995) );
  XNOR U7150 ( .A(n7018), .B(n6988), .Z(n7017) );
  OR U7151 ( .A(n6657), .B(n6931), .Z(n6988) );
  XNOR U7152 ( .A(n7019), .B(n6713), .Z(n6931) );
  XNOR U7153 ( .A(n6658), .B(n6570), .Z(n6657) );
  ANDN U7154 ( .B(n6713), .A(n6570), .Z(n7018) );
  XOR U7155 ( .A(n7006), .B(n7020), .Z(n6570) );
  XOR U7156 ( .A(n6999), .B(n7021), .Z(n7020) );
  XOR U7157 ( .A(n7008), .B(n7006), .Z(n6713) );
  XNOR U7158 ( .A(n6932), .B(n6658), .Z(n6982) );
  XOR U7159 ( .A(n7006), .B(n7022), .Z(n6658) );
  XNOR U7160 ( .A(n7008), .B(n7003), .Z(n7022) );
  XOR U7161 ( .A(n7023), .B(n7024), .Z(n7003) );
  XNOR U7162 ( .A(n6435), .B(n7025), .Z(n7024) );
  XNOR U7163 ( .A(key[287]), .B(n6411), .Z(n7023) );
  XOR U7164 ( .A(n7026), .B(n7027), .Z(n6411) );
  XNOR U7165 ( .A(n7028), .B(n7029), .Z(n7006) );
  XNOR U7166 ( .A(n6398), .B(n7030), .Z(n7029) );
  XNOR U7167 ( .A(n6403), .B(n7031), .Z(n7028) );
  XNOR U7168 ( .A(key[285]), .B(n7032), .Z(n7031) );
  XNOR U7169 ( .A(n7033), .B(n7034), .Z(n6403) );
  IV U7170 ( .A(n7019), .Z(n6932) );
  XNOR U7171 ( .A(n7000), .B(n7035), .Z(n7019) );
  XOR U7172 ( .A(n7005), .B(n7021), .Z(n7035) );
  IV U7173 ( .A(n7008), .Z(n7021) );
  XOR U7174 ( .A(n7036), .B(n7037), .Z(n7008) );
  XNOR U7175 ( .A(n7038), .B(n6410), .Z(n6400) );
  XOR U7176 ( .A(n7016), .B(n7039), .Z(n6410) );
  XNOR U7177 ( .A(n7041), .B(n7042), .Z(n7036) );
  XOR U7178 ( .A(key[286]), .B(n6600), .Z(n7042) );
  XNOR U7179 ( .A(n7043), .B(n7044), .Z(n6600) );
  XOR U7180 ( .A(n7045), .B(n6429), .Z(n7044) );
  XNOR U7181 ( .A(n7046), .B(n7047), .Z(n7043) );
  XOR U7182 ( .A(n7049), .B(n7050), .Z(n7005) );
  XOR U7183 ( .A(n6430), .B(n7051), .Z(n7050) );
  XOR U7184 ( .A(n7053), .B(n7054), .Z(n6999) );
  XOR U7185 ( .A(n6427), .B(n7055), .Z(n7054) );
  XNOR U7186 ( .A(n7056), .B(n7057), .Z(n7053) );
  XNOR U7187 ( .A(n7058), .B(n7059), .Z(n7049) );
  XNOR U7188 ( .A(key[283]), .B(n6432), .Z(n7059) );
  XOR U7189 ( .A(n7016), .B(n6419), .Z(n6432) );
  XOR U7190 ( .A(n7060), .B(n7061), .Z(n7000) );
  XOR U7191 ( .A(n6423), .B(n7062), .Z(n7061) );
  XNOR U7192 ( .A(n6388), .B(n7063), .Z(n7060) );
  XNOR U7193 ( .A(key[282]), .B(n7064), .Z(n7063) );
  XNOR U7194 ( .A(key[400]), .B(n3615), .Z(n6751) );
  XNOR U7195 ( .A(n2728), .B(n3602), .Z(n3615) );
  XOR U7196 ( .A(n6555), .B(n6678), .Z(n3602) );
  XNOR U7197 ( .A(n6694), .B(n7065), .Z(n6678) );
  XOR U7198 ( .A(n7066), .B(n6588), .Z(n7065) );
  OR U7199 ( .A(n7067), .B(n6682), .Z(n6588) );
  XNOR U7200 ( .A(n6591), .B(n6677), .Z(n6682) );
  ANDN U7201 ( .B(n6677), .A(n7068), .Z(n7066) );
  XNOR U7202 ( .A(n6586), .B(n7069), .Z(n6555) );
  XOR U7203 ( .A(n7070), .B(n6696), .Z(n7069) );
  XNOR U7204 ( .A(n6668), .B(n6559), .Z(n6665) );
  NOR U7205 ( .A(n7072), .B(n6668), .Z(n7070) );
  XNOR U7206 ( .A(n6694), .B(n7073), .Z(n6586) );
  XNOR U7207 ( .A(n7074), .B(n7075), .Z(n7073) );
  NAND U7208 ( .A(n6688), .B(n7076), .Z(n7075) );
  XOR U7209 ( .A(n7077), .B(n7074), .Z(n6694) );
  OR U7210 ( .A(n6690), .B(n7078), .Z(n7074) );
  XNOR U7211 ( .A(n7079), .B(n6688), .Z(n6690) );
  XOR U7212 ( .A(n6677), .B(n6559), .Z(n6688) );
  XOR U7213 ( .A(n7080), .B(n7081), .Z(n6559) );
  NANDN U7214 ( .A(n7082), .B(n7083), .Z(n7081) );
  XOR U7215 ( .A(n7084), .B(n7085), .Z(n6677) );
  NANDN U7216 ( .A(n7082), .B(n7086), .Z(n7085) );
  ANDN U7217 ( .B(n7079), .A(n7087), .Z(n7077) );
  IV U7218 ( .A(n6693), .Z(n7079) );
  XOR U7219 ( .A(n6668), .B(n6591), .Z(n6693) );
  XNOR U7220 ( .A(n7088), .B(n7084), .Z(n6591) );
  NANDN U7221 ( .A(n7089), .B(n7090), .Z(n7084) );
  XOR U7222 ( .A(n7086), .B(n7091), .Z(n7090) );
  ANDN U7223 ( .B(n7091), .A(n7092), .Z(n7088) );
  XOR U7224 ( .A(n7093), .B(n7080), .Z(n6668) );
  NANDN U7225 ( .A(n7089), .B(n7094), .Z(n7080) );
  XOR U7226 ( .A(n7095), .B(n7083), .Z(n7094) );
  XNOR U7227 ( .A(n7096), .B(n7097), .Z(n7082) );
  XOR U7228 ( .A(n7098), .B(n7099), .Z(n7097) );
  XNOR U7229 ( .A(n7100), .B(n7101), .Z(n7096) );
  XNOR U7230 ( .A(n7102), .B(n7103), .Z(n7101) );
  ANDN U7231 ( .B(n7095), .A(n7099), .Z(n7102) );
  ANDN U7232 ( .B(n7095), .A(n7092), .Z(n7093) );
  XNOR U7233 ( .A(n7098), .B(n7104), .Z(n7092) );
  XOR U7234 ( .A(n7105), .B(n7103), .Z(n7104) );
  NAND U7235 ( .A(n7106), .B(n7107), .Z(n7103) );
  XNOR U7236 ( .A(n7100), .B(n7083), .Z(n7107) );
  IV U7237 ( .A(n7095), .Z(n7100) );
  XNOR U7238 ( .A(n7086), .B(n7099), .Z(n7106) );
  IV U7239 ( .A(n7091), .Z(n7099) );
  XOR U7240 ( .A(n7108), .B(n7109), .Z(n7091) );
  XNOR U7241 ( .A(n7110), .B(n7111), .Z(n7109) );
  XNOR U7242 ( .A(n7112), .B(n7113), .Z(n7108) );
  NOR U7243 ( .A(n6667), .B(n7072), .Z(n7112) );
  AND U7244 ( .A(n7083), .B(n7086), .Z(n7105) );
  XNOR U7245 ( .A(n7083), .B(n7086), .Z(n7098) );
  XNOR U7246 ( .A(n7114), .B(n7115), .Z(n7086) );
  XNOR U7247 ( .A(n7116), .B(n7111), .Z(n7115) );
  XOR U7248 ( .A(n7117), .B(n7118), .Z(n7114) );
  XNOR U7249 ( .A(n7119), .B(n7113), .Z(n7118) );
  OR U7250 ( .A(n6666), .B(n7071), .Z(n7113) );
  XNOR U7251 ( .A(n7072), .B(n6698), .Z(n7071) );
  XNOR U7252 ( .A(n6667), .B(n6560), .Z(n6666) );
  ANDN U7253 ( .B(n7120), .A(n6698), .Z(n7119) );
  XNOR U7254 ( .A(n7121), .B(n7122), .Z(n7083) );
  XNOR U7255 ( .A(n7111), .B(n7123), .Z(n7122) );
  XOR U7256 ( .A(n6681), .B(n7117), .Z(n7123) );
  XNOR U7257 ( .A(n7072), .B(n7124), .Z(n7111) );
  XOR U7258 ( .A(n6590), .B(n7125), .Z(n7121) );
  XNOR U7259 ( .A(n7126), .B(n7127), .Z(n7125) );
  ANDN U7260 ( .B(n7128), .A(n7068), .Z(n7126) );
  XNOR U7261 ( .A(n7129), .B(n7130), .Z(n7095) );
  XNOR U7262 ( .A(n7116), .B(n7131), .Z(n7130) );
  XNOR U7263 ( .A(n6676), .B(n7110), .Z(n7131) );
  XOR U7264 ( .A(n7117), .B(n7132), .Z(n7110) );
  XNOR U7265 ( .A(n7133), .B(n7134), .Z(n7132) );
  NAND U7266 ( .A(n7076), .B(n6687), .Z(n7134) );
  XNOR U7267 ( .A(n7135), .B(n7133), .Z(n7117) );
  NANDN U7268 ( .A(n7078), .B(n6691), .Z(n7133) );
  XOR U7269 ( .A(n6692), .B(n6687), .Z(n6691) );
  XNOR U7270 ( .A(n7128), .B(n6560), .Z(n6687) );
  XOR U7271 ( .A(n7087), .B(n7076), .Z(n7078) );
  XNOR U7272 ( .A(n7068), .B(n7136), .Z(n7076) );
  ANDN U7273 ( .B(n6692), .A(n7087), .Z(n7135) );
  XNOR U7274 ( .A(n6590), .B(n7072), .Z(n7087) );
  XOR U7275 ( .A(n7137), .B(n7138), .Z(n7072) );
  XNOR U7276 ( .A(n7139), .B(n7140), .Z(n7138) );
  XOR U7277 ( .A(n7136), .B(n7120), .Z(n7116) );
  IV U7278 ( .A(n6560), .Z(n7120) );
  XOR U7279 ( .A(n7141), .B(n7142), .Z(n6560) );
  XNOR U7280 ( .A(n7143), .B(n7140), .Z(n7142) );
  IV U7281 ( .A(n6698), .Z(n7136) );
  XOR U7282 ( .A(n7140), .B(n7144), .Z(n6698) );
  XNOR U7283 ( .A(n7145), .B(n7146), .Z(n7129) );
  XNOR U7284 ( .A(n7147), .B(n7127), .Z(n7146) );
  OR U7285 ( .A(n6683), .B(n7067), .Z(n7127) );
  XNOR U7286 ( .A(n6590), .B(n7068), .Z(n7067) );
  IV U7287 ( .A(n7145), .Z(n7068) );
  XOR U7288 ( .A(n6681), .B(n7128), .Z(n6683) );
  IV U7289 ( .A(n6676), .Z(n7128) );
  XOR U7290 ( .A(n7124), .B(n7148), .Z(n6676) );
  XNOR U7291 ( .A(n7143), .B(n7137), .Z(n7148) );
  XOR U7292 ( .A(n7149), .B(n7150), .Z(n7137) );
  XNOR U7293 ( .A(n6281), .B(n7151), .Z(n7150) );
  XNOR U7294 ( .A(key[290]), .B(n7152), .Z(n7149) );
  IV U7295 ( .A(n6667), .Z(n7124) );
  XOR U7296 ( .A(n7141), .B(n7153), .Z(n6667) );
  XOR U7297 ( .A(n7140), .B(n7154), .Z(n7153) );
  NOR U7298 ( .A(n6681), .B(n6590), .Z(n7147) );
  XOR U7299 ( .A(n7141), .B(n7155), .Z(n6681) );
  XOR U7300 ( .A(n7140), .B(n7156), .Z(n7155) );
  XOR U7301 ( .A(n7157), .B(n7158), .Z(n7140) );
  XOR U7302 ( .A(n7159), .B(n7160), .Z(n7158) );
  XNOR U7303 ( .A(n6277), .B(n7161), .Z(n7157) );
  XOR U7304 ( .A(key[294]), .B(n6590), .Z(n7161) );
  XOR U7305 ( .A(n7162), .B(n7163), .Z(n6277) );
  IV U7306 ( .A(n7144), .Z(n7141) );
  XOR U7307 ( .A(n7164), .B(n7165), .Z(n7144) );
  XNOR U7308 ( .A(n7166), .B(n7167), .Z(n7165) );
  XNOR U7309 ( .A(key[293]), .B(n7168), .Z(n7164) );
  XOR U7310 ( .A(n7169), .B(n7170), .Z(n7145) );
  XNOR U7311 ( .A(n7156), .B(n7154), .Z(n7170) );
  XNOR U7312 ( .A(n7171), .B(n7172), .Z(n7154) );
  XNOR U7313 ( .A(n7173), .B(n7174), .Z(n7172) );
  XNOR U7314 ( .A(key[295]), .B(n6270), .Z(n7171) );
  XNOR U7315 ( .A(n7175), .B(n7176), .Z(n7156) );
  XOR U7316 ( .A(n7177), .B(n7178), .Z(n7176) );
  XNOR U7317 ( .A(n6246), .B(n7179), .Z(n7175) );
  XOR U7318 ( .A(key[292]), .B(n7180), .Z(n7179) );
  XOR U7319 ( .A(n7162), .B(n7181), .Z(n6246) );
  XNOR U7320 ( .A(n6590), .B(n7139), .Z(n7169) );
  XOR U7321 ( .A(n7182), .B(n7183), .Z(n7139) );
  XNOR U7322 ( .A(n7184), .B(n7185), .Z(n7183) );
  XOR U7323 ( .A(n7143), .B(n7186), .Z(n7185) );
  XOR U7324 ( .A(n7187), .B(n7188), .Z(n7143) );
  XNOR U7325 ( .A(n6299), .B(n7189), .Z(n7188) );
  XNOR U7326 ( .A(key[289]), .B(n7190), .Z(n7187) );
  XNOR U7327 ( .A(n7191), .B(n7192), .Z(n7182) );
  XNOR U7328 ( .A(key[291]), .B(n6292), .Z(n7192) );
  XOR U7329 ( .A(n7162), .B(n7193), .Z(n6292) );
  XNOR U7330 ( .A(n7194), .B(n7195), .Z(n6590) );
  XOR U7331 ( .A(n7196), .B(n6272), .Z(n7195) );
  IV U7332 ( .A(n7197), .Z(n6272) );
  XNOR U7333 ( .A(key[288]), .B(n6289), .Z(n7194) );
  XOR U7334 ( .A(n6621), .B(n6726), .Z(n2728) );
  XNOR U7335 ( .A(n6774), .B(n7198), .Z(n6726) );
  XOR U7336 ( .A(n7199), .B(n6617), .Z(n7198) );
  OR U7337 ( .A(n7200), .B(n6762), .Z(n6617) );
  XNOR U7338 ( .A(n6620), .B(n6758), .Z(n6762) );
  ANDN U7339 ( .B(n6758), .A(n7201), .Z(n7199) );
  XNOR U7340 ( .A(n6615), .B(n7202), .Z(n6621) );
  XOR U7341 ( .A(n7203), .B(n6776), .Z(n7202) );
  XNOR U7342 ( .A(n6749), .B(n6625), .Z(n6746) );
  NOR U7343 ( .A(n7205), .B(n6749), .Z(n7203) );
  XNOR U7344 ( .A(n6774), .B(n7206), .Z(n6615) );
  XNOR U7345 ( .A(n7207), .B(n7208), .Z(n7206) );
  NAND U7346 ( .A(n6768), .B(n7209), .Z(n7208) );
  XOR U7347 ( .A(n7210), .B(n7207), .Z(n6774) );
  OR U7348 ( .A(n6770), .B(n7211), .Z(n7207) );
  XNOR U7349 ( .A(n7212), .B(n6768), .Z(n6770) );
  XOR U7350 ( .A(n6758), .B(n6625), .Z(n6768) );
  XOR U7351 ( .A(n7213), .B(n7214), .Z(n6625) );
  NANDN U7352 ( .A(n7215), .B(n7216), .Z(n7214) );
  XOR U7353 ( .A(n7217), .B(n7218), .Z(n6758) );
  NANDN U7354 ( .A(n7215), .B(n7219), .Z(n7218) );
  ANDN U7355 ( .B(n7212), .A(n7220), .Z(n7210) );
  IV U7356 ( .A(n6773), .Z(n7212) );
  XOR U7357 ( .A(n6749), .B(n6620), .Z(n6773) );
  XNOR U7358 ( .A(n7221), .B(n7217), .Z(n6620) );
  NANDN U7359 ( .A(n7222), .B(n7223), .Z(n7217) );
  XOR U7360 ( .A(n7219), .B(n7224), .Z(n7223) );
  ANDN U7361 ( .B(n7224), .A(n7225), .Z(n7221) );
  XOR U7362 ( .A(n7226), .B(n7213), .Z(n6749) );
  NANDN U7363 ( .A(n7222), .B(n7227), .Z(n7213) );
  XOR U7364 ( .A(n7228), .B(n7216), .Z(n7227) );
  XNOR U7365 ( .A(n7229), .B(n7230), .Z(n7215) );
  XOR U7366 ( .A(n7231), .B(n7232), .Z(n7230) );
  XNOR U7367 ( .A(n7233), .B(n7234), .Z(n7229) );
  XNOR U7368 ( .A(n7235), .B(n7236), .Z(n7234) );
  ANDN U7369 ( .B(n7228), .A(n7232), .Z(n7235) );
  ANDN U7370 ( .B(n7228), .A(n7225), .Z(n7226) );
  XNOR U7371 ( .A(n7231), .B(n7237), .Z(n7225) );
  XOR U7372 ( .A(n7238), .B(n7236), .Z(n7237) );
  NAND U7373 ( .A(n7239), .B(n7240), .Z(n7236) );
  XNOR U7374 ( .A(n7233), .B(n7216), .Z(n7240) );
  IV U7375 ( .A(n7228), .Z(n7233) );
  XNOR U7376 ( .A(n7219), .B(n7232), .Z(n7239) );
  IV U7377 ( .A(n7224), .Z(n7232) );
  XOR U7378 ( .A(n7241), .B(n7242), .Z(n7224) );
  XNOR U7379 ( .A(n7243), .B(n7244), .Z(n7242) );
  XNOR U7380 ( .A(n7245), .B(n7246), .Z(n7241) );
  NOR U7381 ( .A(n6748), .B(n7205), .Z(n7245) );
  AND U7382 ( .A(n7216), .B(n7219), .Z(n7238) );
  XNOR U7383 ( .A(n7216), .B(n7219), .Z(n7231) );
  XNOR U7384 ( .A(n7247), .B(n7248), .Z(n7219) );
  XNOR U7385 ( .A(n7249), .B(n7244), .Z(n7248) );
  XOR U7386 ( .A(n7250), .B(n7251), .Z(n7247) );
  XNOR U7387 ( .A(n7252), .B(n7246), .Z(n7251) );
  OR U7388 ( .A(n6747), .B(n7204), .Z(n7246) );
  XNOR U7389 ( .A(n7205), .B(n6778), .Z(n7204) );
  XNOR U7390 ( .A(n6748), .B(n6626), .Z(n6747) );
  ANDN U7391 ( .B(n7253), .A(n6778), .Z(n7252) );
  XNOR U7392 ( .A(n7254), .B(n7255), .Z(n7216) );
  XNOR U7393 ( .A(n7244), .B(n7256), .Z(n7255) );
  XOR U7394 ( .A(n6761), .B(n7250), .Z(n7256) );
  XNOR U7395 ( .A(n7205), .B(n7257), .Z(n7244) );
  XOR U7396 ( .A(n6619), .B(n7258), .Z(n7254) );
  XNOR U7397 ( .A(n7259), .B(n7260), .Z(n7258) );
  ANDN U7398 ( .B(n7261), .A(n7201), .Z(n7259) );
  XNOR U7399 ( .A(n7262), .B(n7263), .Z(n7228) );
  XNOR U7400 ( .A(n7249), .B(n7264), .Z(n7263) );
  XNOR U7401 ( .A(n6757), .B(n7243), .Z(n7264) );
  XOR U7402 ( .A(n7250), .B(n7265), .Z(n7243) );
  XNOR U7403 ( .A(n7266), .B(n7267), .Z(n7265) );
  NAND U7404 ( .A(n7209), .B(n6767), .Z(n7267) );
  XNOR U7405 ( .A(n7268), .B(n7266), .Z(n7250) );
  NANDN U7406 ( .A(n7211), .B(n6771), .Z(n7266) );
  XOR U7407 ( .A(n6772), .B(n6767), .Z(n6771) );
  XNOR U7408 ( .A(n7261), .B(n6626), .Z(n6767) );
  XOR U7409 ( .A(n7220), .B(n7209), .Z(n7211) );
  XNOR U7410 ( .A(n7201), .B(n7269), .Z(n7209) );
  ANDN U7411 ( .B(n6772), .A(n7220), .Z(n7268) );
  XNOR U7412 ( .A(n6619), .B(n7205), .Z(n7220) );
  XOR U7413 ( .A(n7270), .B(n7271), .Z(n7205) );
  XNOR U7414 ( .A(n7272), .B(n7273), .Z(n7271) );
  XOR U7415 ( .A(n7269), .B(n7253), .Z(n7249) );
  IV U7416 ( .A(n6626), .Z(n7253) );
  XOR U7417 ( .A(n7274), .B(n7275), .Z(n6626) );
  XNOR U7418 ( .A(n7276), .B(n7273), .Z(n7275) );
  IV U7419 ( .A(n6778), .Z(n7269) );
  XOR U7420 ( .A(n7273), .B(n7277), .Z(n6778) );
  XNOR U7421 ( .A(n7278), .B(n7279), .Z(n7262) );
  XNOR U7422 ( .A(n7280), .B(n7260), .Z(n7279) );
  OR U7423 ( .A(n6763), .B(n7200), .Z(n7260) );
  XNOR U7424 ( .A(n6619), .B(n7201), .Z(n7200) );
  IV U7425 ( .A(n7278), .Z(n7201) );
  XOR U7426 ( .A(n6761), .B(n7261), .Z(n6763) );
  IV U7427 ( .A(n6757), .Z(n7261) );
  XOR U7428 ( .A(n7257), .B(n7281), .Z(n6757) );
  XNOR U7429 ( .A(n7276), .B(n7270), .Z(n7281) );
  XOR U7430 ( .A(n7282), .B(n7283), .Z(n7270) );
  XOR U7431 ( .A(n5958), .B(n7284), .Z(n7283) );
  XNOR U7432 ( .A(n5970), .B(n7285), .Z(n7282) );
  XNOR U7433 ( .A(key[330]), .B(n7286), .Z(n7285) );
  IV U7434 ( .A(n6748), .Z(n7257) );
  XOR U7435 ( .A(n7274), .B(n7287), .Z(n6748) );
  XOR U7436 ( .A(n7273), .B(n7288), .Z(n7287) );
  NOR U7437 ( .A(n6761), .B(n6619), .Z(n7280) );
  XOR U7438 ( .A(n7274), .B(n7289), .Z(n6761) );
  XOR U7439 ( .A(n7273), .B(n7290), .Z(n7289) );
  XOR U7440 ( .A(n7291), .B(n7292), .Z(n7273) );
  XOR U7441 ( .A(n7293), .B(n5954), .Z(n7292) );
  XNOR U7442 ( .A(n7294), .B(n5935), .Z(n5954) );
  XOR U7443 ( .A(n7295), .B(n7296), .Z(n5935) );
  XNOR U7444 ( .A(n7297), .B(n7298), .Z(n7291) );
  XOR U7445 ( .A(key[334]), .B(n6619), .Z(n7298) );
  IV U7446 ( .A(n7277), .Z(n7274) );
  XOR U7447 ( .A(n7299), .B(n7300), .Z(n7277) );
  XNOR U7448 ( .A(n5952), .B(n7301), .Z(n7300) );
  XNOR U7449 ( .A(n5940), .B(n7302), .Z(n7299) );
  XNOR U7450 ( .A(key[333]), .B(n7303), .Z(n7302) );
  XOR U7451 ( .A(n7304), .B(n7305), .Z(n5940) );
  XOR U7452 ( .A(n7306), .B(n7307), .Z(n7278) );
  XNOR U7453 ( .A(n7290), .B(n7288), .Z(n7307) );
  XNOR U7454 ( .A(n7308), .B(n7309), .Z(n7288) );
  XNOR U7455 ( .A(n5949), .B(n7310), .Z(n7309) );
  XNOR U7456 ( .A(key[335]), .B(n5936), .Z(n7308) );
  XNOR U7457 ( .A(n7311), .B(n7312), .Z(n5936) );
  XNOR U7458 ( .A(n7313), .B(n7314), .Z(n7290) );
  XOR U7459 ( .A(n7315), .B(n5923), .Z(n7314) );
  XNOR U7460 ( .A(n7316), .B(n7317), .Z(n5923) );
  XNOR U7461 ( .A(n7318), .B(n7319), .Z(n7313) );
  XNOR U7462 ( .A(key[332]), .B(n5925), .Z(n7319) );
  XOR U7463 ( .A(n7295), .B(n5942), .Z(n5925) );
  XNOR U7464 ( .A(n6619), .B(n7272), .Z(n7306) );
  XOR U7465 ( .A(n7320), .B(n7321), .Z(n7272) );
  XNOR U7466 ( .A(n7322), .B(n7323), .Z(n7321) );
  XNOR U7467 ( .A(n7276), .B(n7324), .Z(n7323) );
  XOR U7468 ( .A(n7325), .B(n7326), .Z(n7276) );
  XOR U7469 ( .A(n5962), .B(n7327), .Z(n7326) );
  XNOR U7470 ( .A(n7328), .B(n7329), .Z(n7325) );
  XNOR U7471 ( .A(n7330), .B(n7331), .Z(n7320) );
  XNOR U7472 ( .A(key[331]), .B(n5967), .Z(n7331) );
  XOR U7473 ( .A(n7295), .B(n5927), .Z(n5967) );
  XNOR U7474 ( .A(n7332), .B(n7333), .Z(n6619) );
  XOR U7475 ( .A(n7334), .B(n5964), .Z(n7333) );
  XNOR U7476 ( .A(n7335), .B(n7336), .Z(n7332) );
  XNOR U7477 ( .A(key[328]), .B(n7337), .Z(n7336) );
  XNOR U7478 ( .A(n5410), .B(n7338), .Z(n5416) );
  XNOR U7479 ( .A(n7339), .B(n7340), .Z(n7338) );
  ANDN U7480 ( .B(n7341), .A(n5444), .Z(n7339) );
  IV U7481 ( .A(n7342), .Z(n5444) );
  XNOR U7482 ( .A(n7343), .B(n7344), .Z(n5410) );
  XNOR U7483 ( .A(n7345), .B(n7346), .Z(n7344) );
  NANDN U7484 ( .A(n7347), .B(n7348), .Z(n7346) );
  XNOR U7485 ( .A(n1034), .B(n1039), .Z(n413) );
  XOR U7486 ( .A(n5363), .B(n7349), .Z(n1039) );
  XNOR U7487 ( .A(n5365), .B(n5350), .Z(n7349) );
  XOR U7488 ( .A(n5520), .B(n5445), .Z(n5350) );
  XNOR U7489 ( .A(n5409), .B(n7350), .Z(n5445) );
  XNOR U7490 ( .A(n7351), .B(n7352), .Z(n7350) );
  NANDN U7491 ( .A(n7353), .B(n7354), .Z(n7352) );
  XNOR U7492 ( .A(n7343), .B(n7355), .Z(n5520) );
  XOR U7493 ( .A(n7356), .B(n5412), .Z(n7355) );
  OR U7494 ( .A(n7357), .B(n7358), .Z(n5412) );
  ANDN U7495 ( .B(n7359), .A(n7360), .Z(n7356) );
  XOR U7496 ( .A(n7343), .B(n7361), .Z(n5365) );
  XOR U7497 ( .A(n7340), .B(n7362), .Z(n7361) );
  NANDN U7498 ( .A(n7363), .B(n5420), .Z(n7362) );
  XOR U7499 ( .A(n7342), .B(n5420), .Z(n5441) );
  XOR U7500 ( .A(n7365), .B(n7345), .Z(n7343) );
  OR U7501 ( .A(n7366), .B(n7367), .Z(n7345) );
  NOR U7502 ( .A(n7368), .B(n7369), .Z(n7365) );
  XOR U7503 ( .A(n5438), .B(n7370), .Z(n5363) );
  XNOR U7504 ( .A(n7351), .B(n7371), .Z(n7370) );
  NANDN U7505 ( .A(n7372), .B(n5415), .Z(n7371) );
  OR U7506 ( .A(n7358), .B(n7373), .Z(n7351) );
  XNOR U7507 ( .A(n5415), .B(n7354), .Z(n7358) );
  XNOR U7508 ( .A(n5409), .B(n7374), .Z(n5438) );
  XNOR U7509 ( .A(n7375), .B(n7376), .Z(n7374) );
  NANDN U7510 ( .A(n7347), .B(n7377), .Z(n7376) );
  XOR U7511 ( .A(n7378), .B(n7375), .Z(n5409) );
  NANDN U7512 ( .A(n7366), .B(n7379), .Z(n7375) );
  XNOR U7513 ( .A(n7368), .B(n7347), .Z(n7366) );
  XNOR U7514 ( .A(n7354), .B(n5420), .Z(n7347) );
  XOR U7515 ( .A(n7380), .B(n7381), .Z(n5420) );
  NANDN U7516 ( .A(n7382), .B(n7383), .Z(n7381) );
  IV U7517 ( .A(n7360), .Z(n7354) );
  XNOR U7518 ( .A(n7384), .B(n7385), .Z(n7360) );
  NANDN U7519 ( .A(n7382), .B(n7386), .Z(n7385) );
  ANDN U7520 ( .B(n7387), .A(n7368), .Z(n7378) );
  XNOR U7521 ( .A(n7342), .B(n5415), .Z(n7368) );
  XNOR U7522 ( .A(n7388), .B(n7384), .Z(n5415) );
  NANDN U7523 ( .A(n7389), .B(n7390), .Z(n7384) );
  XOR U7524 ( .A(n7386), .B(n7391), .Z(n7390) );
  ANDN U7525 ( .B(n7391), .A(n7392), .Z(n7388) );
  XNOR U7526 ( .A(n7393), .B(n7380), .Z(n7342) );
  NANDN U7527 ( .A(n7389), .B(n7394), .Z(n7380) );
  XOR U7528 ( .A(n7395), .B(n7383), .Z(n7394) );
  XNOR U7529 ( .A(n7396), .B(n7397), .Z(n7382) );
  XOR U7530 ( .A(n7398), .B(n7399), .Z(n7397) );
  XNOR U7531 ( .A(n7400), .B(n7401), .Z(n7396) );
  XNOR U7532 ( .A(n7402), .B(n7403), .Z(n7401) );
  ANDN U7533 ( .B(n7395), .A(n7399), .Z(n7402) );
  ANDN U7534 ( .B(n7395), .A(n7392), .Z(n7393) );
  XNOR U7535 ( .A(n7398), .B(n7404), .Z(n7392) );
  XOR U7536 ( .A(n7405), .B(n7403), .Z(n7404) );
  NAND U7537 ( .A(n7406), .B(n7407), .Z(n7403) );
  XNOR U7538 ( .A(n7400), .B(n7383), .Z(n7407) );
  IV U7539 ( .A(n7395), .Z(n7400) );
  XNOR U7540 ( .A(n7386), .B(n7399), .Z(n7406) );
  IV U7541 ( .A(n7391), .Z(n7399) );
  XOR U7542 ( .A(n7408), .B(n7409), .Z(n7391) );
  XNOR U7543 ( .A(n7410), .B(n7411), .Z(n7409) );
  XNOR U7544 ( .A(n7412), .B(n7413), .Z(n7408) );
  ANDN U7545 ( .B(n7341), .A(n7414), .Z(n7412) );
  AND U7546 ( .A(n7383), .B(n7386), .Z(n7405) );
  XNOR U7547 ( .A(n7383), .B(n7386), .Z(n7398) );
  XNOR U7548 ( .A(n7415), .B(n7416), .Z(n7386) );
  XNOR U7549 ( .A(n7417), .B(n7411), .Z(n7416) );
  XOR U7550 ( .A(n7418), .B(n7419), .Z(n7415) );
  XNOR U7551 ( .A(n7420), .B(n7413), .Z(n7419) );
  OR U7552 ( .A(n5442), .B(n7364), .Z(n7413) );
  XNOR U7553 ( .A(n7341), .B(n7421), .Z(n7364) );
  XNOR U7554 ( .A(n7414), .B(n5421), .Z(n5442) );
  ANDN U7555 ( .B(n7422), .A(n7363), .Z(n7420) );
  XNOR U7556 ( .A(n7423), .B(n7424), .Z(n7383) );
  XNOR U7557 ( .A(n7411), .B(n7425), .Z(n7424) );
  XOR U7558 ( .A(n7372), .B(n7418), .Z(n7425) );
  XNOR U7559 ( .A(n7341), .B(n7414), .Z(n7411) );
  XNOR U7560 ( .A(n7426), .B(n7427), .Z(n7423) );
  XNOR U7561 ( .A(n7428), .B(n7429), .Z(n7427) );
  ANDN U7562 ( .B(n7359), .A(n7353), .Z(n7428) );
  XNOR U7563 ( .A(n7430), .B(n7431), .Z(n7395) );
  XNOR U7564 ( .A(n7417), .B(n7432), .Z(n7431) );
  XNOR U7565 ( .A(n7353), .B(n7410), .Z(n7432) );
  XOR U7566 ( .A(n7418), .B(n7433), .Z(n7410) );
  XNOR U7567 ( .A(n7434), .B(n7435), .Z(n7433) );
  NAND U7568 ( .A(n7348), .B(n7377), .Z(n7435) );
  XNOR U7569 ( .A(n7436), .B(n7434), .Z(n7418) );
  NANDN U7570 ( .A(n7367), .B(n7379), .Z(n7434) );
  XOR U7571 ( .A(n7387), .B(n7377), .Z(n7379) );
  XNOR U7572 ( .A(n7437), .B(n5421), .Z(n7377) );
  XOR U7573 ( .A(n7369), .B(n7348), .Z(n7367) );
  XOR U7574 ( .A(n7359), .B(n7421), .Z(n7348) );
  ANDN U7575 ( .B(n7387), .A(n7369), .Z(n7436) );
  XNOR U7576 ( .A(n7426), .B(n7341), .Z(n7369) );
  XNOR U7577 ( .A(n7438), .B(n7439), .Z(n7341) );
  XNOR U7578 ( .A(n7440), .B(n7441), .Z(n7439) );
  XOR U7579 ( .A(n7421), .B(n7422), .Z(n7417) );
  IV U7580 ( .A(n5421), .Z(n7422) );
  XOR U7581 ( .A(n7442), .B(n7443), .Z(n5421) );
  XNOR U7582 ( .A(n7444), .B(n7441), .Z(n7443) );
  IV U7583 ( .A(n7363), .Z(n7421) );
  XOR U7584 ( .A(n7441), .B(n7445), .Z(n7363) );
  XNOR U7585 ( .A(n7359), .B(n7446), .Z(n7430) );
  XNOR U7586 ( .A(n7447), .B(n7429), .Z(n7446) );
  OR U7587 ( .A(n7373), .B(n7357), .Z(n7429) );
  XNOR U7588 ( .A(n7426), .B(n7359), .Z(n7357) );
  XOR U7589 ( .A(n7372), .B(n7437), .Z(n7373) );
  IV U7590 ( .A(n7353), .Z(n7437) );
  XOR U7591 ( .A(n5443), .B(n7448), .Z(n7353) );
  XNOR U7592 ( .A(n7444), .B(n7438), .Z(n7448) );
  XOR U7593 ( .A(n7449), .B(n7450), .Z(n7438) );
  XNOR U7594 ( .A(n2582), .B(n3813), .Z(n7450) );
  XNOR U7595 ( .A(n2560), .B(n7451), .Z(n3813) );
  XNOR U7596 ( .A(n4929), .B(n7452), .Z(n7449) );
  XOR U7597 ( .A(key[442]), .B(n2581), .Z(n7452) );
  XOR U7598 ( .A(n7453), .B(n7454), .Z(n4929) );
  XNOR U7599 ( .A(n7455), .B(n7456), .Z(n7454) );
  ANDN U7600 ( .B(n7457), .A(n5414), .Z(n7447) );
  XOR U7601 ( .A(n7458), .B(n7459), .Z(n7359) );
  XNOR U7602 ( .A(n7460), .B(n7461), .Z(n7459) );
  XOR U7603 ( .A(n7426), .B(n7440), .Z(n7458) );
  XOR U7604 ( .A(n7462), .B(n7463), .Z(n7440) );
  XNOR U7605 ( .A(n7444), .B(n7464), .Z(n7463) );
  XNOR U7606 ( .A(n2559), .B(n3809), .Z(n7464) );
  XNOR U7607 ( .A(n3798), .B(n2538), .Z(n3809) );
  XOR U7608 ( .A(n7465), .B(n7466), .Z(n2559) );
  XOR U7609 ( .A(n7467), .B(n7468), .Z(n7466) );
  XOR U7610 ( .A(n7469), .B(n7470), .Z(n7444) );
  XOR U7611 ( .A(n3819), .B(n2560), .Z(n7470) );
  XOR U7612 ( .A(n7471), .B(n2588), .Z(n3819) );
  XOR U7613 ( .A(n7472), .B(n7473), .Z(n2588) );
  XOR U7614 ( .A(n4926), .B(n7476), .Z(n7469) );
  XNOR U7615 ( .A(key[441]), .B(n2591), .Z(n7476) );
  XOR U7616 ( .A(n7477), .B(n7478), .Z(n2591) );
  XNOR U7617 ( .A(n7479), .B(n7480), .Z(n7478) );
  XOR U7618 ( .A(n4928), .B(n7481), .Z(n7462) );
  XOR U7619 ( .A(key[443]), .B(n4923), .Z(n7481) );
  XOR U7620 ( .A(n3820), .B(n3803), .Z(n4923) );
  XNOR U7621 ( .A(n7482), .B(n4926), .Z(n3803) );
  XNOR U7622 ( .A(n7483), .B(n7484), .Z(n4926) );
  XOR U7623 ( .A(n2582), .B(n2561), .Z(n4928) );
  XOR U7624 ( .A(n7485), .B(n7486), .Z(n2561) );
  XNOR U7625 ( .A(n7472), .B(n7487), .Z(n7486) );
  IV U7626 ( .A(n7488), .Z(n7472) );
  XOR U7627 ( .A(n7474), .B(n7489), .Z(n7485) );
  XOR U7628 ( .A(n7490), .B(n7491), .Z(n2582) );
  XNOR U7629 ( .A(n7492), .B(n7493), .Z(n7491) );
  XOR U7630 ( .A(n7494), .B(n7495), .Z(n7490) );
  XOR U7631 ( .A(n7457), .B(n5443), .Z(n7387) );
  IV U7632 ( .A(n7414), .Z(n5443) );
  XOR U7633 ( .A(n7442), .B(n7496), .Z(n7414) );
  XOR U7634 ( .A(n7441), .B(n7461), .Z(n7496) );
  XNOR U7635 ( .A(n7497), .B(n7498), .Z(n7461) );
  XNOR U7636 ( .A(n3796), .B(n4944), .Z(n7498) );
  XNOR U7637 ( .A(n7499), .B(n3795), .Z(n4944) );
  XNOR U7638 ( .A(n7500), .B(n7501), .Z(n3795) );
  XOR U7639 ( .A(n7488), .B(n7502), .Z(n7501) );
  XOR U7640 ( .A(n7474), .B(n7475), .Z(n7500) );
  XNOR U7641 ( .A(n7504), .B(n7505), .Z(n7503) );
  NANDN U7642 ( .A(n7506), .B(n7507), .Z(n7505) );
  XOR U7643 ( .A(n7465), .B(n7509), .Z(n3796) );
  XOR U7644 ( .A(n7477), .B(n7510), .Z(n7509) );
  XNOR U7645 ( .A(n7511), .B(n7480), .Z(n7465) );
  XNOR U7646 ( .A(n7513), .B(n7514), .Z(n7512) );
  OR U7647 ( .A(n7515), .B(n7516), .Z(n7514) );
  XOR U7648 ( .A(key[447]), .B(n2589), .Z(n7497) );
  XOR U7649 ( .A(n7518), .B(n3820), .Z(n2589) );
  IV U7650 ( .A(n7372), .Z(n7457) );
  XOR U7651 ( .A(n7442), .B(n7519), .Z(n7372) );
  XOR U7652 ( .A(n7441), .B(n7460), .Z(n7519) );
  XNOR U7653 ( .A(n7520), .B(n7521), .Z(n7460) );
  XOR U7654 ( .A(n4938), .B(n3801), .Z(n7521) );
  XOR U7655 ( .A(n7518), .B(n2548), .Z(n3801) );
  XNOR U7656 ( .A(n7522), .B(n2578), .Z(n3805) );
  IV U7657 ( .A(n7451), .Z(n2578) );
  XNOR U7658 ( .A(n7523), .B(n7488), .Z(n7451) );
  XOR U7659 ( .A(n7524), .B(n7525), .Z(n7488) );
  XNOR U7660 ( .A(n7526), .B(n7527), .Z(n7525) );
  NANDN U7661 ( .A(n7528), .B(n7529), .Z(n7527) );
  XNOR U7662 ( .A(n7530), .B(n2560), .Z(n2538) );
  XOR U7663 ( .A(n7531), .B(n7492), .Z(n2560) );
  IV U7664 ( .A(n7532), .Z(n7492) );
  XNOR U7665 ( .A(n4937), .B(n7533), .Z(n7520) );
  XNOR U7666 ( .A(key[444]), .B(n3802), .Z(n7533) );
  XOR U7667 ( .A(n7534), .B(n2581), .Z(n3802) );
  XNOR U7668 ( .A(n7479), .B(n7535), .Z(n2581) );
  IV U7669 ( .A(n7511), .Z(n7479) );
  XNOR U7670 ( .A(n7536), .B(n7537), .Z(n7511) );
  XNOR U7671 ( .A(n7538), .B(n7539), .Z(n7537) );
  NAND U7672 ( .A(n7540), .B(n7541), .Z(n7539) );
  XOR U7673 ( .A(n7542), .B(n7543), .Z(n3788) );
  XNOR U7674 ( .A(n7482), .B(n7544), .Z(n7543) );
  XNOR U7675 ( .A(n7545), .B(n7546), .Z(n7542) );
  XOR U7676 ( .A(n7547), .B(n7548), .Z(n7546) );
  ANDN U7677 ( .B(n7549), .A(n7550), .Z(n7548) );
  XOR U7678 ( .A(n7551), .B(n7552), .Z(n7441) );
  XOR U7679 ( .A(n3780), .B(n5414), .Z(n7552) );
  IV U7680 ( .A(n7426), .Z(n5414) );
  XOR U7681 ( .A(n7553), .B(n7554), .Z(n7426) );
  XNOR U7682 ( .A(n7471), .B(n2554), .Z(n7554) );
  XNOR U7683 ( .A(n3806), .B(n2587), .Z(n2554) );
  XOR U7684 ( .A(n7555), .B(n7534), .Z(n2587) );
  XOR U7685 ( .A(n7522), .B(n7556), .Z(n3806) );
  IV U7686 ( .A(n2577), .Z(n7471) );
  XOR U7687 ( .A(n7532), .B(n7557), .Z(n2577) );
  XOR U7688 ( .A(n7518), .B(n7559), .Z(n7553) );
  XNOR U7689 ( .A(key[440]), .B(n4927), .Z(n7559) );
  XNOR U7690 ( .A(n7560), .B(n7561), .Z(n4927) );
  XOR U7691 ( .A(n7483), .B(n7562), .Z(n7561) );
  XOR U7692 ( .A(n3798), .B(n7499), .Z(n3780) );
  IV U7693 ( .A(n2555), .Z(n7499) );
  XOR U7694 ( .A(n7563), .B(n7564), .Z(n2555) );
  XOR U7695 ( .A(n7532), .B(n7565), .Z(n7564) );
  XOR U7696 ( .A(n7566), .B(n7567), .Z(n7532) );
  XNOR U7697 ( .A(n7568), .B(n7569), .Z(n7567) );
  NANDN U7698 ( .A(n7570), .B(n7571), .Z(n7569) );
  XOR U7699 ( .A(n7494), .B(n7558), .Z(n7563) );
  XNOR U7700 ( .A(n7573), .B(n7574), .Z(n7572) );
  NANDN U7701 ( .A(n7575), .B(n7576), .Z(n7574) );
  IV U7702 ( .A(n7518), .Z(n3798) );
  XOR U7703 ( .A(n7530), .B(n7578), .Z(n7518) );
  XOR U7704 ( .A(n4955), .B(n7579), .Z(n7551) );
  XNOR U7705 ( .A(key[446]), .B(n4947), .Z(n7579) );
  XNOR U7706 ( .A(n3789), .B(n4943), .Z(n4947) );
  XNOR U7707 ( .A(n3820), .B(n3797), .Z(n4943) );
  XNOR U7708 ( .A(n7453), .B(n7580), .Z(n3797) );
  XNOR U7709 ( .A(n7560), .B(n7544), .Z(n7580) );
  XNOR U7710 ( .A(n7581), .B(n7582), .Z(n7544) );
  XNOR U7711 ( .A(n7583), .B(n7584), .Z(n7582) );
  OR U7712 ( .A(n7585), .B(n7586), .Z(n7584) );
  XNOR U7713 ( .A(n7483), .B(n7562), .Z(n7453) );
  XNOR U7714 ( .A(n7588), .B(n7589), .Z(n7587) );
  OR U7715 ( .A(n7585), .B(n7590), .Z(n7589) );
  XNOR U7716 ( .A(n7592), .B(n7593), .Z(n7483) );
  XNOR U7717 ( .A(n7594), .B(n7595), .Z(n7593) );
  NAND U7718 ( .A(n7596), .B(n7549), .Z(n7595) );
  XNOR U7719 ( .A(n7484), .B(n7482), .Z(n3820) );
  XNOR U7720 ( .A(n7581), .B(n7597), .Z(n7482) );
  XOR U7721 ( .A(n7598), .B(n7594), .Z(n7597) );
  NOR U7722 ( .A(n7601), .B(n7602), .Z(n7598) );
  XNOR U7723 ( .A(n7592), .B(n7603), .Z(n7581) );
  XNOR U7724 ( .A(n7604), .B(n7605), .Z(n7603) );
  NAND U7725 ( .A(n7606), .B(n7607), .Z(n7605) );
  XNOR U7726 ( .A(n2567), .B(n2550), .Z(n3789) );
  XOR U7727 ( .A(n7475), .B(n7487), .Z(n2550) );
  XNOR U7728 ( .A(n7508), .B(n7608), .Z(n7487) );
  XNOR U7729 ( .A(n7609), .B(n7610), .Z(n7608) );
  NOR U7730 ( .A(n7611), .B(n7612), .Z(n7609) );
  XNOR U7731 ( .A(n7613), .B(n7614), .Z(n7508) );
  XNOR U7732 ( .A(n7615), .B(n7616), .Z(n7614) );
  NAND U7733 ( .A(n7617), .B(n7618), .Z(n7616) );
  XOR U7734 ( .A(n7523), .B(n7489), .Z(n7475) );
  XOR U7735 ( .A(n7613), .B(n7619), .Z(n7489) );
  XNOR U7736 ( .A(n7504), .B(n7620), .Z(n7619) );
  NANDN U7737 ( .A(n7621), .B(n7622), .Z(n7620) );
  OR U7738 ( .A(n7623), .B(n7624), .Z(n7504) );
  IV U7739 ( .A(n7556), .Z(n7523) );
  XNOR U7740 ( .A(n7524), .B(n7625), .Z(n7556) );
  XOR U7741 ( .A(n7626), .B(n7627), .Z(n7625) );
  ANDN U7742 ( .B(n7622), .A(n7628), .Z(n7626) );
  IV U7743 ( .A(n2546), .Z(n4955) );
  XOR U7744 ( .A(n7477), .B(n7468), .Z(n2546) );
  XNOR U7745 ( .A(n7517), .B(n7629), .Z(n7468) );
  XNOR U7746 ( .A(n7630), .B(n7631), .Z(n7629) );
  NOR U7747 ( .A(n7632), .B(n7633), .Z(n7630) );
  XNOR U7748 ( .A(n7634), .B(n7635), .Z(n7517) );
  XNOR U7749 ( .A(n7636), .B(n7637), .Z(n7635) );
  NAND U7750 ( .A(n7638), .B(n7639), .Z(n7637) );
  XOR U7751 ( .A(n7555), .B(n7467), .Z(n7477) );
  XOR U7752 ( .A(n7634), .B(n7640), .Z(n7467) );
  XNOR U7753 ( .A(n7513), .B(n7641), .Z(n7640) );
  NANDN U7754 ( .A(n7642), .B(n7643), .Z(n7641) );
  OR U7755 ( .A(n7644), .B(n7645), .Z(n7513) );
  IV U7756 ( .A(n7535), .Z(n7555) );
  XNOR U7757 ( .A(n7536), .B(n7646), .Z(n7535) );
  XOR U7758 ( .A(n7647), .B(n7648), .Z(n7646) );
  NOR U7759 ( .A(n7649), .B(n7642), .Z(n7647) );
  IV U7760 ( .A(n7445), .Z(n7442) );
  XOR U7761 ( .A(n7650), .B(n7651), .Z(n7445) );
  XNOR U7762 ( .A(n3787), .B(n4954), .Z(n7651) );
  XNOR U7763 ( .A(n2548), .B(n3786), .Z(n4954) );
  XNOR U7764 ( .A(n7652), .B(n7653), .Z(n3786) );
  XNOR U7765 ( .A(n7613), .B(n7502), .Z(n7653) );
  XNOR U7766 ( .A(n7654), .B(n7655), .Z(n7502) );
  XNOR U7767 ( .A(n7627), .B(n7656), .Z(n7655) );
  NANDN U7768 ( .A(n7657), .B(n7507), .Z(n7656) );
  OR U7769 ( .A(n7658), .B(n7623), .Z(n7627) );
  XNOR U7770 ( .A(n7507), .B(n7622), .Z(n7623) );
  XOR U7771 ( .A(n7659), .B(n7615), .Z(n7613) );
  NANDN U7772 ( .A(n7660), .B(n7661), .Z(n7615) );
  ANDN U7773 ( .B(n7662), .A(n7663), .Z(n7659) );
  XNOR U7774 ( .A(n7522), .B(n7664), .Z(n7652) );
  XOR U7775 ( .A(n7610), .B(n7665), .Z(n7664) );
  ANDN U7776 ( .B(n7529), .A(n7666), .Z(n7665) );
  ANDN U7777 ( .B(n7667), .A(n7668), .Z(n7610) );
  XNOR U7778 ( .A(n7654), .B(n7669), .Z(n7522) );
  XOR U7779 ( .A(n7670), .B(n7526), .Z(n7669) );
  XNOR U7780 ( .A(n7612), .B(n7529), .Z(n7667) );
  NOR U7781 ( .A(n7672), .B(n7612), .Z(n7670) );
  XNOR U7782 ( .A(n7524), .B(n7673), .Z(n7654) );
  XNOR U7783 ( .A(n7674), .B(n7675), .Z(n7673) );
  NAND U7784 ( .A(n7618), .B(n7676), .Z(n7675) );
  XOR U7785 ( .A(n7677), .B(n7674), .Z(n7524) );
  OR U7786 ( .A(n7660), .B(n7678), .Z(n7674) );
  XNOR U7787 ( .A(n7679), .B(n7618), .Z(n7660) );
  XOR U7788 ( .A(n7622), .B(n7529), .Z(n7618) );
  XOR U7789 ( .A(n7680), .B(n7681), .Z(n7529) );
  NANDN U7790 ( .A(n7682), .B(n7683), .Z(n7681) );
  XOR U7791 ( .A(n7684), .B(n7685), .Z(n7622) );
  NANDN U7792 ( .A(n7682), .B(n7686), .Z(n7685) );
  ANDN U7793 ( .B(n7679), .A(n7687), .Z(n7677) );
  IV U7794 ( .A(n7663), .Z(n7679) );
  XOR U7795 ( .A(n7612), .B(n7507), .Z(n7663) );
  XNOR U7796 ( .A(n7688), .B(n7684), .Z(n7507) );
  NANDN U7797 ( .A(n7689), .B(n7690), .Z(n7684) );
  XOR U7798 ( .A(n7686), .B(n7691), .Z(n7690) );
  ANDN U7799 ( .B(n7691), .A(n7692), .Z(n7688) );
  XOR U7800 ( .A(n7693), .B(n7680), .Z(n7612) );
  NANDN U7801 ( .A(n7689), .B(n7694), .Z(n7680) );
  XOR U7802 ( .A(n7695), .B(n7683), .Z(n7694) );
  XNOR U7803 ( .A(n7696), .B(n7697), .Z(n7682) );
  XOR U7804 ( .A(n7698), .B(n7699), .Z(n7697) );
  XNOR U7805 ( .A(n7700), .B(n7701), .Z(n7696) );
  XNOR U7806 ( .A(n7702), .B(n7703), .Z(n7701) );
  ANDN U7807 ( .B(n7695), .A(n7699), .Z(n7702) );
  ANDN U7808 ( .B(n7695), .A(n7692), .Z(n7693) );
  XNOR U7809 ( .A(n7698), .B(n7704), .Z(n7692) );
  XOR U7810 ( .A(n7705), .B(n7703), .Z(n7704) );
  NAND U7811 ( .A(n7706), .B(n7707), .Z(n7703) );
  XNOR U7812 ( .A(n7700), .B(n7683), .Z(n7707) );
  IV U7813 ( .A(n7695), .Z(n7700) );
  XNOR U7814 ( .A(n7686), .B(n7699), .Z(n7706) );
  IV U7815 ( .A(n7691), .Z(n7699) );
  XOR U7816 ( .A(n7708), .B(n7709), .Z(n7691) );
  XNOR U7817 ( .A(n7710), .B(n7711), .Z(n7709) );
  XNOR U7818 ( .A(n7712), .B(n7713), .Z(n7708) );
  NOR U7819 ( .A(n7611), .B(n7672), .Z(n7712) );
  AND U7820 ( .A(n7683), .B(n7686), .Z(n7705) );
  XNOR U7821 ( .A(n7683), .B(n7686), .Z(n7698) );
  XNOR U7822 ( .A(n7714), .B(n7715), .Z(n7686) );
  XNOR U7823 ( .A(n7716), .B(n7711), .Z(n7715) );
  XOR U7824 ( .A(n7717), .B(n7718), .Z(n7714) );
  XNOR U7825 ( .A(n7719), .B(n7713), .Z(n7718) );
  OR U7826 ( .A(n7668), .B(n7671), .Z(n7713) );
  XNOR U7827 ( .A(n7672), .B(n7528), .Z(n7671) );
  XNOR U7828 ( .A(n7611), .B(n7666), .Z(n7668) );
  ANDN U7829 ( .B(n7720), .A(n7528), .Z(n7719) );
  XNOR U7830 ( .A(n7721), .B(n7722), .Z(n7683) );
  XNOR U7831 ( .A(n7711), .B(n7723), .Z(n7722) );
  XOR U7832 ( .A(n7506), .B(n7717), .Z(n7723) );
  XNOR U7833 ( .A(n7672), .B(n7724), .Z(n7711) );
  XOR U7834 ( .A(n7657), .B(n7725), .Z(n7721) );
  XNOR U7835 ( .A(n7726), .B(n7727), .Z(n7725) );
  ANDN U7836 ( .B(n7728), .A(n7628), .Z(n7726) );
  XNOR U7837 ( .A(n7729), .B(n7730), .Z(n7695) );
  XNOR U7838 ( .A(n7716), .B(n7731), .Z(n7730) );
  XNOR U7839 ( .A(n7621), .B(n7710), .Z(n7731) );
  XOR U7840 ( .A(n7717), .B(n7732), .Z(n7710) );
  XNOR U7841 ( .A(n7733), .B(n7734), .Z(n7732) );
  NAND U7842 ( .A(n7676), .B(n7617), .Z(n7734) );
  XNOR U7843 ( .A(n7735), .B(n7733), .Z(n7717) );
  NANDN U7844 ( .A(n7678), .B(n7661), .Z(n7733) );
  XOR U7845 ( .A(n7662), .B(n7617), .Z(n7661) );
  XNOR U7846 ( .A(n7728), .B(n7666), .Z(n7617) );
  XOR U7847 ( .A(n7687), .B(n7676), .Z(n7678) );
  XNOR U7848 ( .A(n7628), .B(n7736), .Z(n7676) );
  ANDN U7849 ( .B(n7662), .A(n7687), .Z(n7735) );
  XNOR U7850 ( .A(n7657), .B(n7672), .Z(n7687) );
  XOR U7851 ( .A(n7737), .B(n7738), .Z(n7672) );
  XNOR U7852 ( .A(n7739), .B(n7740), .Z(n7738) );
  XOR U7853 ( .A(n7736), .B(n7720), .Z(n7716) );
  IV U7854 ( .A(n7666), .Z(n7720) );
  XOR U7855 ( .A(n7741), .B(n7742), .Z(n7666) );
  XOR U7856 ( .A(n7743), .B(n7740), .Z(n7742) );
  IV U7857 ( .A(n7528), .Z(n7736) );
  XOR U7858 ( .A(n7740), .B(n7744), .Z(n7528) );
  XNOR U7859 ( .A(n7745), .B(n7746), .Z(n7729) );
  XNOR U7860 ( .A(n7747), .B(n7727), .Z(n7746) );
  OR U7861 ( .A(n7624), .B(n7658), .Z(n7727) );
  XNOR U7862 ( .A(n7657), .B(n7628), .Z(n7658) );
  IV U7863 ( .A(n7745), .Z(n7628) );
  XOR U7864 ( .A(n7506), .B(n7728), .Z(n7624) );
  IV U7865 ( .A(n7621), .Z(n7728) );
  XOR U7866 ( .A(n7724), .B(n7748), .Z(n7621) );
  XNOR U7867 ( .A(n7749), .B(n7737), .Z(n7748) );
  XOR U7868 ( .A(n7750), .B(n7751), .Z(n7737) );
  XNOR U7869 ( .A(n6107), .B(n6881), .Z(n7751) );
  XNOR U7870 ( .A(n7752), .B(n7753), .Z(n7750) );
  XNOR U7871 ( .A(key[362]), .B(n6922), .Z(n7753) );
  IV U7872 ( .A(n7611), .Z(n7724) );
  XOR U7873 ( .A(n7741), .B(n7754), .Z(n7611) );
  XOR U7874 ( .A(n7740), .B(n7755), .Z(n7754) );
  NOR U7875 ( .A(n7506), .B(n7657), .Z(n7747) );
  XOR U7876 ( .A(n7741), .B(n7756), .Z(n7506) );
  XOR U7877 ( .A(n7740), .B(n7757), .Z(n7756) );
  XOR U7878 ( .A(n7758), .B(n7759), .Z(n7740) );
  XNOR U7879 ( .A(n7657), .B(n7760), .Z(n7759) );
  XNOR U7880 ( .A(n7761), .B(n7762), .Z(n7758) );
  XNOR U7881 ( .A(key[366]), .B(n6892), .Z(n7762) );
  XNOR U7882 ( .A(n7763), .B(n6903), .Z(n6892) );
  XNOR U7883 ( .A(n7764), .B(n7765), .Z(n6903) );
  IV U7884 ( .A(n7744), .Z(n7741) );
  XOR U7885 ( .A(n7766), .B(n7767), .Z(n7744) );
  XOR U7886 ( .A(n6908), .B(n6896), .Z(n7767) );
  XNOR U7887 ( .A(n7768), .B(n6080), .Z(n6896) );
  XNOR U7888 ( .A(n6890), .B(n7769), .Z(n7766) );
  XNOR U7889 ( .A(key[365]), .B(n7770), .Z(n7769) );
  XOR U7890 ( .A(n7771), .B(n7772), .Z(n7745) );
  XNOR U7891 ( .A(n7757), .B(n7755), .Z(n7772) );
  XNOR U7892 ( .A(n7773), .B(n7774), .Z(n7755) );
  XOR U7893 ( .A(n6891), .B(n6904), .Z(n7774) );
  XNOR U7894 ( .A(n7775), .B(n7776), .Z(n6904) );
  XNOR U7895 ( .A(key[367]), .B(n6927), .Z(n7773) );
  XOR U7896 ( .A(n7764), .B(n7777), .Z(n6927) );
  XNOR U7897 ( .A(n7778), .B(n7779), .Z(n7757) );
  XNOR U7898 ( .A(n6907), .B(n7780), .Z(n7779) );
  XNOR U7899 ( .A(n6094), .B(n7781), .Z(n6907) );
  XNOR U7900 ( .A(n6909), .B(n7782), .Z(n7778) );
  XOR U7901 ( .A(key[364]), .B(n6916), .Z(n7782) );
  XNOR U7902 ( .A(n7764), .B(n6898), .Z(n6909) );
  XNOR U7903 ( .A(n7657), .B(n7739), .Z(n7771) );
  XOR U7904 ( .A(n7783), .B(n7784), .Z(n7739) );
  XNOR U7905 ( .A(n7785), .B(n7786), .Z(n7784) );
  XOR U7906 ( .A(n6062), .B(n7749), .Z(n7786) );
  IV U7907 ( .A(n7743), .Z(n7749) );
  XNOR U7908 ( .A(n7787), .B(n7788), .Z(n7743) );
  XNOR U7909 ( .A(n6919), .B(n6061), .Z(n7788) );
  XNOR U7910 ( .A(n6883), .B(n7789), .Z(n7787) );
  XOR U7911 ( .A(key[361]), .B(n6116), .Z(n7789) );
  XNOR U7912 ( .A(n6914), .B(n7790), .Z(n7783) );
  XNOR U7913 ( .A(key[363]), .B(n6924), .Z(n7790) );
  XNOR U7914 ( .A(n7764), .B(n6911), .Z(n6924) );
  IV U7915 ( .A(n7791), .Z(n6914) );
  XNOR U7916 ( .A(n7792), .B(n7793), .Z(n7657) );
  XOR U7917 ( .A(n7794), .B(n6087), .Z(n7793) );
  XNOR U7918 ( .A(n7795), .B(n7796), .Z(n7792) );
  XOR U7919 ( .A(key[360]), .B(n7797), .Z(n7796) );
  XNOR U7920 ( .A(n7798), .B(n7799), .Z(n2548) );
  XNOR U7921 ( .A(n7800), .B(n7565), .Z(n7799) );
  XNOR U7922 ( .A(n7801), .B(n7802), .Z(n7565) );
  XNOR U7923 ( .A(n7803), .B(n7804), .Z(n7802) );
  NANDN U7924 ( .A(n7805), .B(n7576), .Z(n7804) );
  XNOR U7925 ( .A(n7530), .B(n7806), .Z(n7798) );
  XOR U7926 ( .A(n7807), .B(n7808), .Z(n7806) );
  ANDN U7927 ( .B(n7571), .A(n7809), .Z(n7808) );
  XNOR U7928 ( .A(n7801), .B(n7810), .Z(n7530) );
  XOR U7929 ( .A(n7811), .B(n7568), .Z(n7810) );
  NOR U7930 ( .A(n7814), .B(n7815), .Z(n7811) );
  XNOR U7931 ( .A(n7566), .B(n7816), .Z(n7801) );
  XNOR U7932 ( .A(n7817), .B(n7818), .Z(n7816) );
  NAND U7933 ( .A(n7819), .B(n7820), .Z(n7818) );
  XOR U7934 ( .A(n7821), .B(n7822), .Z(n3787) );
  XNOR U7935 ( .A(n7534), .B(n7510), .Z(n7822) );
  XNOR U7936 ( .A(n7823), .B(n7824), .Z(n7510) );
  XNOR U7937 ( .A(n7648), .B(n7825), .Z(n7824) );
  OR U7938 ( .A(n7515), .B(n7826), .Z(n7825) );
  OR U7939 ( .A(n7644), .B(n7827), .Z(n7648) );
  XNOR U7940 ( .A(n7515), .B(n7642), .Z(n7644) );
  XNOR U7941 ( .A(n7823), .B(n7828), .Z(n7534) );
  XOR U7942 ( .A(n7829), .B(n7538), .Z(n7828) );
  NOR U7943 ( .A(n7832), .B(n7633), .Z(n7829) );
  XNOR U7944 ( .A(n7536), .B(n7833), .Z(n7823) );
  XNOR U7945 ( .A(n7834), .B(n7835), .Z(n7833) );
  NAND U7946 ( .A(n7639), .B(n7836), .Z(n7835) );
  XOR U7947 ( .A(n7837), .B(n7834), .Z(n7536) );
  OR U7948 ( .A(n7838), .B(n7839), .Z(n7834) );
  ANDN U7949 ( .B(n7840), .A(n7841), .Z(n7837) );
  XNOR U7950 ( .A(n7634), .B(n7842), .Z(n7821) );
  XOR U7951 ( .A(n7631), .B(n7843), .Z(n7842) );
  ANDN U7952 ( .B(n7541), .A(n7844), .Z(n7843) );
  ANDN U7953 ( .B(n7831), .A(n7845), .Z(n7631) );
  XNOR U7954 ( .A(n7633), .B(n7541), .Z(n7831) );
  XOR U7955 ( .A(n7846), .B(n7636), .Z(n7634) );
  NANDN U7956 ( .A(n7838), .B(n7847), .Z(n7636) );
  XNOR U7957 ( .A(n7840), .B(n7639), .Z(n7838) );
  XNOR U7958 ( .A(n7642), .B(n7541), .Z(n7639) );
  XOR U7959 ( .A(n7848), .B(n7849), .Z(n7541) );
  NANDN U7960 ( .A(n7850), .B(n7851), .Z(n7849) );
  XNOR U7961 ( .A(n7852), .B(n7853), .Z(n7642) );
  OR U7962 ( .A(n7850), .B(n7854), .Z(n7853) );
  AND U7963 ( .A(n7840), .B(n7855), .Z(n7846) );
  XOR U7964 ( .A(n7515), .B(n7633), .Z(n7840) );
  XOR U7965 ( .A(n7856), .B(n7848), .Z(n7633) );
  NANDN U7966 ( .A(n7857), .B(n7858), .Z(n7848) );
  ANDN U7967 ( .B(n7859), .A(n7860), .Z(n7856) );
  NANDN U7968 ( .A(n7857), .B(n7862), .Z(n7852) );
  XOR U7969 ( .A(n7863), .B(n7850), .Z(n7857) );
  XNOR U7970 ( .A(n7864), .B(n7865), .Z(n7850) );
  XOR U7971 ( .A(n7866), .B(n7859), .Z(n7865) );
  XNOR U7972 ( .A(n7867), .B(n7868), .Z(n7864) );
  XNOR U7973 ( .A(n7869), .B(n7870), .Z(n7868) );
  ANDN U7974 ( .B(n7859), .A(n7871), .Z(n7869) );
  IV U7975 ( .A(n7872), .Z(n7859) );
  ANDN U7976 ( .B(n7863), .A(n7871), .Z(n7861) );
  IV U7977 ( .A(n7867), .Z(n7871) );
  IV U7978 ( .A(n7860), .Z(n7863) );
  XNOR U7979 ( .A(n7866), .B(n7873), .Z(n7860) );
  XOR U7980 ( .A(n7874), .B(n7870), .Z(n7873) );
  NAND U7981 ( .A(n7862), .B(n7858), .Z(n7870) );
  XNOR U7982 ( .A(n7851), .B(n7872), .Z(n7858) );
  XOR U7983 ( .A(n7875), .B(n7876), .Z(n7872) );
  XOR U7984 ( .A(n7877), .B(n7878), .Z(n7876) );
  XNOR U7985 ( .A(n7643), .B(n7879), .Z(n7878) );
  XNOR U7986 ( .A(n7880), .B(n7881), .Z(n7875) );
  XNOR U7987 ( .A(n7882), .B(n7883), .Z(n7881) );
  ANDN U7988 ( .B(n7884), .A(n7826), .Z(n7882) );
  XNOR U7989 ( .A(n7867), .B(n7854), .Z(n7862) );
  XOR U7990 ( .A(n7885), .B(n7886), .Z(n7867) );
  XNOR U7991 ( .A(n7887), .B(n7879), .Z(n7886) );
  XOR U7992 ( .A(n7888), .B(n7889), .Z(n7879) );
  XNOR U7993 ( .A(n7890), .B(n7891), .Z(n7889) );
  NAND U7994 ( .A(n7836), .B(n7638), .Z(n7891) );
  XNOR U7995 ( .A(n7892), .B(n7893), .Z(n7885) );
  ANDN U7996 ( .B(n7894), .A(n7832), .Z(n7892) );
  ANDN U7997 ( .B(n7851), .A(n7854), .Z(n7874) );
  XOR U7998 ( .A(n7854), .B(n7851), .Z(n7866) );
  XNOR U7999 ( .A(n7895), .B(n7896), .Z(n7851) );
  XNOR U8000 ( .A(n7888), .B(n7897), .Z(n7896) );
  XOR U8001 ( .A(n7887), .B(n7516), .Z(n7897) );
  XOR U8002 ( .A(n7826), .B(n7898), .Z(n7895) );
  XNOR U8003 ( .A(n7899), .B(n7883), .Z(n7898) );
  OR U8004 ( .A(n7645), .B(n7827), .Z(n7883) );
  XNOR U8005 ( .A(n7826), .B(n7649), .Z(n7827) );
  XOR U8006 ( .A(n7516), .B(n7643), .Z(n7645) );
  ANDN U8007 ( .B(n7643), .A(n7649), .Z(n7899) );
  XOR U8008 ( .A(n7900), .B(n7901), .Z(n7854) );
  XOR U8009 ( .A(n7888), .B(n7877), .Z(n7901) );
  XOR U8010 ( .A(n7540), .B(n7844), .Z(n7877) );
  XOR U8011 ( .A(n7902), .B(n7890), .Z(n7888) );
  NANDN U8012 ( .A(n7839), .B(n7847), .Z(n7890) );
  XOR U8013 ( .A(n7855), .B(n7638), .Z(n7847) );
  XNOR U8014 ( .A(n7894), .B(n7903), .Z(n7643) );
  XNOR U8015 ( .A(n7904), .B(n7905), .Z(n7903) );
  XOR U8016 ( .A(n7841), .B(n7836), .Z(n7839) );
  XNOR U8017 ( .A(n7649), .B(n7540), .Z(n7836) );
  IV U8018 ( .A(n7880), .Z(n7649) );
  XOR U8019 ( .A(n7906), .B(n7907), .Z(n7880) );
  XOR U8020 ( .A(n7908), .B(n7909), .Z(n7907) );
  XNOR U8021 ( .A(n7826), .B(n7910), .Z(n7906) );
  ANDN U8022 ( .B(n7855), .A(n7841), .Z(n7902) );
  XNOR U8023 ( .A(n7826), .B(n7832), .Z(n7841) );
  XOR U8024 ( .A(n7894), .B(n7884), .Z(n7855) );
  IV U8025 ( .A(n7516), .Z(n7884) );
  XOR U8026 ( .A(n7911), .B(n7912), .Z(n7516) );
  XOR U8027 ( .A(n7913), .B(n7909), .Z(n7912) );
  XNOR U8028 ( .A(n7914), .B(n7915), .Z(n7909) );
  XOR U8029 ( .A(n7916), .B(n7917), .Z(n7915) );
  XOR U8030 ( .A(n7317), .B(n7918), .Z(n7914) );
  XNOR U8031 ( .A(key[324]), .B(n7318), .Z(n7918) );
  XOR U8032 ( .A(n7919), .B(n7304), .Z(n7318) );
  IV U8033 ( .A(n7632), .Z(n7894) );
  XOR U8034 ( .A(n7887), .B(n7920), .Z(n7900) );
  XNOR U8035 ( .A(n7921), .B(n7893), .Z(n7920) );
  OR U8036 ( .A(n7845), .B(n7830), .Z(n7893) );
  XNOR U8037 ( .A(n7922), .B(n7540), .Z(n7830) );
  XNOR U8038 ( .A(n7632), .B(n7844), .Z(n7845) );
  ANDN U8039 ( .B(n7540), .A(n7844), .Z(n7921) );
  XOR U8040 ( .A(n7911), .B(n7923), .Z(n7844) );
  XOR U8041 ( .A(n7904), .B(n7924), .Z(n7923) );
  XOR U8042 ( .A(n7913), .B(n7911), .Z(n7540) );
  XNOR U8043 ( .A(n7832), .B(n7632), .Z(n7887) );
  XOR U8044 ( .A(n7911), .B(n7925), .Z(n7632) );
  XNOR U8045 ( .A(n7913), .B(n7908), .Z(n7925) );
  XOR U8046 ( .A(n7926), .B(n7927), .Z(n7908) );
  XOR U8047 ( .A(n7928), .B(n7929), .Z(n7927) );
  XOR U8048 ( .A(key[327]), .B(n7919), .Z(n7926) );
  XNOR U8049 ( .A(n7930), .B(n7931), .Z(n7911) );
  XNOR U8050 ( .A(n7932), .B(n7933), .Z(n7931) );
  XNOR U8051 ( .A(key[325]), .B(n7294), .Z(n7930) );
  XNOR U8052 ( .A(n7303), .B(n7934), .Z(n7294) );
  IV U8053 ( .A(n7922), .Z(n7832) );
  XNOR U8054 ( .A(n7905), .B(n7935), .Z(n7922) );
  XOR U8055 ( .A(n7910), .B(n7924), .Z(n7935) );
  IV U8056 ( .A(n7913), .Z(n7924) );
  XOR U8057 ( .A(n7936), .B(n7937), .Z(n7913) );
  XNOR U8058 ( .A(n7826), .B(n7938), .Z(n7937) );
  XNOR U8059 ( .A(n7939), .B(n7940), .Z(n7826) );
  XNOR U8060 ( .A(n7941), .B(n5962), .Z(n7940) );
  XOR U8061 ( .A(n7334), .B(n7942), .Z(n5962) );
  XNOR U8062 ( .A(key[320]), .B(n7335), .Z(n7939) );
  XNOR U8063 ( .A(n7934), .B(n7943), .Z(n7936) );
  XNOR U8064 ( .A(key[326]), .B(n7297), .Z(n7943) );
  XOR U8065 ( .A(n7337), .B(n7311), .Z(n7297) );
  IV U8066 ( .A(n7919), .Z(n7337) );
  XOR U8067 ( .A(n7944), .B(n7945), .Z(n7910) );
  XNOR U8068 ( .A(n5971), .B(n7946), .Z(n7945) );
  XNOR U8069 ( .A(n7904), .B(n7947), .Z(n7946) );
  XOR U8070 ( .A(n7948), .B(n7949), .Z(n7904) );
  XOR U8071 ( .A(n5970), .B(n5950), .Z(n7949) );
  XNOR U8072 ( .A(n7950), .B(n7951), .Z(n5970) );
  XNOR U8073 ( .A(key[321]), .B(n7952), .Z(n7948) );
  XNOR U8074 ( .A(n7953), .B(n7954), .Z(n7944) );
  XNOR U8075 ( .A(key[323]), .B(n7330), .Z(n7954) );
  XOR U8076 ( .A(n7919), .B(n7316), .Z(n7330) );
  XOR U8077 ( .A(n7955), .B(n7956), .Z(n7905) );
  XOR U8078 ( .A(n7951), .B(n5963), .Z(n7956) );
  XNOR U8079 ( .A(key[322]), .B(n7324), .Z(n7955) );
  IV U8080 ( .A(n5965), .Z(n7324) );
  XOR U8081 ( .A(n7286), .B(n7953), .Z(n5965) );
  XNOR U8082 ( .A(n4948), .B(n7957), .Z(n7650) );
  XNOR U8083 ( .A(key[445]), .B(n2567), .Z(n7957) );
  XOR U8084 ( .A(n7558), .B(n7493), .Z(n2567) );
  XNOR U8085 ( .A(n7577), .B(n7958), .Z(n7493) );
  XNOR U8086 ( .A(n7959), .B(n7807), .Z(n7958) );
  ANDN U8087 ( .B(n7813), .A(n7960), .Z(n7807) );
  XNOR U8088 ( .A(n7815), .B(n7571), .Z(n7813) );
  NOR U8089 ( .A(n7961), .B(n7815), .Z(n7959) );
  XNOR U8090 ( .A(n7800), .B(n7962), .Z(n7577) );
  XNOR U8091 ( .A(n7963), .B(n7964), .Z(n7962) );
  NAND U8092 ( .A(n7965), .B(n7819), .Z(n7964) );
  XOR U8093 ( .A(n7531), .B(n7495), .Z(n7558) );
  XOR U8094 ( .A(n7800), .B(n7966), .Z(n7495) );
  XNOR U8095 ( .A(n7573), .B(n7967), .Z(n7966) );
  NANDN U8096 ( .A(n7968), .B(n7969), .Z(n7967) );
  OR U8097 ( .A(n7970), .B(n7971), .Z(n7573) );
  XOR U8098 ( .A(n7972), .B(n7963), .Z(n7800) );
  NANDN U8099 ( .A(n7973), .B(n7974), .Z(n7963) );
  ANDN U8100 ( .B(n7975), .A(n7976), .Z(n7972) );
  IV U8101 ( .A(n7578), .Z(n7531) );
  XNOR U8102 ( .A(n7566), .B(n7977), .Z(n7578) );
  XOR U8103 ( .A(n7978), .B(n7803), .Z(n7977) );
  OR U8104 ( .A(n7979), .B(n7970), .Z(n7803) );
  XNOR U8105 ( .A(n7576), .B(n7969), .Z(n7970) );
  ANDN U8106 ( .B(n7969), .A(n7980), .Z(n7978) );
  XOR U8107 ( .A(n7981), .B(n7817), .Z(n7566) );
  OR U8108 ( .A(n7973), .B(n7982), .Z(n7817) );
  XNOR U8109 ( .A(n7983), .B(n7819), .Z(n7973) );
  XOR U8110 ( .A(n7969), .B(n7571), .Z(n7819) );
  XOR U8111 ( .A(n7984), .B(n7985), .Z(n7571) );
  NANDN U8112 ( .A(n7986), .B(n7987), .Z(n7985) );
  XOR U8113 ( .A(n7988), .B(n7989), .Z(n7969) );
  NANDN U8114 ( .A(n7986), .B(n7990), .Z(n7989) );
  ANDN U8115 ( .B(n7983), .A(n7991), .Z(n7981) );
  IV U8116 ( .A(n7976), .Z(n7983) );
  XOR U8117 ( .A(n7815), .B(n7576), .Z(n7976) );
  XNOR U8118 ( .A(n7992), .B(n7988), .Z(n7576) );
  NANDN U8119 ( .A(n7993), .B(n7994), .Z(n7988) );
  XOR U8120 ( .A(n7990), .B(n7995), .Z(n7994) );
  ANDN U8121 ( .B(n7995), .A(n7996), .Z(n7992) );
  XOR U8122 ( .A(n7997), .B(n7984), .Z(n7815) );
  NANDN U8123 ( .A(n7993), .B(n7998), .Z(n7984) );
  XOR U8124 ( .A(n7999), .B(n7987), .Z(n7998) );
  XNOR U8125 ( .A(n8000), .B(n8001), .Z(n7986) );
  XOR U8126 ( .A(n8002), .B(n8003), .Z(n8001) );
  XNOR U8127 ( .A(n8004), .B(n8005), .Z(n8000) );
  XNOR U8128 ( .A(n8006), .B(n8007), .Z(n8005) );
  ANDN U8129 ( .B(n7999), .A(n8003), .Z(n8006) );
  ANDN U8130 ( .B(n7999), .A(n7996), .Z(n7997) );
  XNOR U8131 ( .A(n8002), .B(n8008), .Z(n7996) );
  XOR U8132 ( .A(n8009), .B(n8007), .Z(n8008) );
  NAND U8133 ( .A(n8010), .B(n8011), .Z(n8007) );
  XNOR U8134 ( .A(n8004), .B(n7987), .Z(n8011) );
  IV U8135 ( .A(n7999), .Z(n8004) );
  XNOR U8136 ( .A(n7990), .B(n8003), .Z(n8010) );
  IV U8137 ( .A(n7995), .Z(n8003) );
  XOR U8138 ( .A(n8012), .B(n8013), .Z(n7995) );
  XNOR U8139 ( .A(n8014), .B(n8015), .Z(n8013) );
  XNOR U8140 ( .A(n8016), .B(n8017), .Z(n8012) );
  NOR U8141 ( .A(n7961), .B(n7814), .Z(n8016) );
  AND U8142 ( .A(n7987), .B(n7990), .Z(n8009) );
  XNOR U8143 ( .A(n7987), .B(n7990), .Z(n8002) );
  XNOR U8144 ( .A(n8018), .B(n8019), .Z(n7990) );
  XNOR U8145 ( .A(n8020), .B(n8015), .Z(n8019) );
  XOR U8146 ( .A(n8021), .B(n8022), .Z(n8018) );
  XNOR U8147 ( .A(n8023), .B(n8017), .Z(n8022) );
  OR U8148 ( .A(n7960), .B(n7812), .Z(n8017) );
  XNOR U8149 ( .A(n7814), .B(n7570), .Z(n7812) );
  XNOR U8150 ( .A(n7961), .B(n7809), .Z(n7960) );
  ANDN U8151 ( .B(n8024), .A(n7570), .Z(n8023) );
  XNOR U8152 ( .A(n8025), .B(n8026), .Z(n7987) );
  XNOR U8153 ( .A(n8015), .B(n8027), .Z(n8026) );
  XOR U8154 ( .A(n7575), .B(n8021), .Z(n8027) );
  XNOR U8155 ( .A(n7814), .B(n8028), .Z(n8015) );
  XOR U8156 ( .A(n7805), .B(n8029), .Z(n8025) );
  XNOR U8157 ( .A(n8030), .B(n8031), .Z(n8029) );
  ANDN U8158 ( .B(n8032), .A(n7980), .Z(n8030) );
  XNOR U8159 ( .A(n8033), .B(n8034), .Z(n7999) );
  XNOR U8160 ( .A(n8020), .B(n8035), .Z(n8034) );
  XNOR U8161 ( .A(n7968), .B(n8014), .Z(n8035) );
  XOR U8162 ( .A(n8021), .B(n8036), .Z(n8014) );
  XNOR U8163 ( .A(n8037), .B(n8038), .Z(n8036) );
  NAND U8164 ( .A(n7820), .B(n7965), .Z(n8038) );
  XNOR U8165 ( .A(n8039), .B(n8037), .Z(n8021) );
  NANDN U8166 ( .A(n7982), .B(n7974), .Z(n8037) );
  XOR U8167 ( .A(n7975), .B(n7965), .Z(n7974) );
  XNOR U8168 ( .A(n8032), .B(n7809), .Z(n7965) );
  XOR U8169 ( .A(n7991), .B(n7820), .Z(n7982) );
  XNOR U8170 ( .A(n7980), .B(n8040), .Z(n7820) );
  ANDN U8171 ( .B(n7975), .A(n7991), .Z(n8039) );
  XNOR U8172 ( .A(n7805), .B(n7814), .Z(n7991) );
  XOR U8173 ( .A(n8041), .B(n8042), .Z(n7814) );
  XNOR U8174 ( .A(n8043), .B(n8044), .Z(n8042) );
  XOR U8175 ( .A(n8040), .B(n8024), .Z(n8020) );
  IV U8176 ( .A(n7809), .Z(n8024) );
  XOR U8177 ( .A(n8045), .B(n8046), .Z(n7809) );
  XNOR U8178 ( .A(n8047), .B(n8044), .Z(n8046) );
  IV U8179 ( .A(n7570), .Z(n8040) );
  XOR U8180 ( .A(n8044), .B(n8048), .Z(n7570) );
  XNOR U8181 ( .A(n8049), .B(n8050), .Z(n8033) );
  XNOR U8182 ( .A(n8051), .B(n8031), .Z(n8050) );
  OR U8183 ( .A(n7971), .B(n7979), .Z(n8031) );
  XNOR U8184 ( .A(n7805), .B(n7980), .Z(n7979) );
  IV U8185 ( .A(n8049), .Z(n7980) );
  XOR U8186 ( .A(n7575), .B(n8032), .Z(n7971) );
  IV U8187 ( .A(n7968), .Z(n8032) );
  XOR U8188 ( .A(n8028), .B(n8052), .Z(n7968) );
  XNOR U8189 ( .A(n8047), .B(n8041), .Z(n8052) );
  XOR U8190 ( .A(n8053), .B(n8054), .Z(n8041) );
  XNOR U8191 ( .A(n8055), .B(n6428), .Z(n8054) );
  IV U8192 ( .A(n8056), .Z(n6428) );
  XOR U8193 ( .A(key[274]), .B(n6430), .Z(n8053) );
  XOR U8194 ( .A(n7064), .B(n8057), .Z(n6430) );
  IV U8195 ( .A(n7961), .Z(n8028) );
  XOR U8196 ( .A(n8045), .B(n8058), .Z(n7961) );
  XOR U8197 ( .A(n8044), .B(n8059), .Z(n8058) );
  NOR U8198 ( .A(n7575), .B(n7805), .Z(n8051) );
  XOR U8199 ( .A(n8045), .B(n8060), .Z(n7575) );
  XOR U8200 ( .A(n8044), .B(n8061), .Z(n8060) );
  XOR U8201 ( .A(n8062), .B(n8063), .Z(n8044) );
  XOR U8202 ( .A(n7805), .B(n8064), .Z(n8063) );
  XNOR U8203 ( .A(n8065), .B(n8066), .Z(n8062) );
  XNOR U8204 ( .A(key[278]), .B(n7041), .Z(n8066) );
  XOR U8205 ( .A(n7048), .B(n7026), .Z(n7041) );
  IV U8206 ( .A(n8048), .Z(n8045) );
  XOR U8207 ( .A(n8067), .B(n8068), .Z(n8048) );
  XOR U8208 ( .A(n7034), .B(n8069), .Z(n8068) );
  XNOR U8209 ( .A(key[277]), .B(n7038), .Z(n8067) );
  XNOR U8210 ( .A(n7032), .B(n8065), .Z(n7038) );
  XOR U8211 ( .A(n8070), .B(n8071), .Z(n8049) );
  XNOR U8212 ( .A(n8061), .B(n8059), .Z(n8071) );
  XNOR U8213 ( .A(n8072), .B(n8073), .Z(n8059) );
  XNOR U8214 ( .A(n8074), .B(n8075), .Z(n8073) );
  XOR U8215 ( .A(key[279]), .B(n7048), .Z(n8072) );
  XNOR U8216 ( .A(n8076), .B(n8077), .Z(n8061) );
  XNOR U8217 ( .A(n7013), .B(n8078), .Z(n8077) );
  XNOR U8218 ( .A(key[276]), .B(n7014), .Z(n8076) );
  XNOR U8219 ( .A(n7048), .B(n7033), .Z(n7014) );
  XNOR U8220 ( .A(n7805), .B(n8043), .Z(n8070) );
  XOR U8221 ( .A(n8079), .B(n8080), .Z(n8043) );
  XNOR U8222 ( .A(n8047), .B(n8082), .Z(n8081) );
  XOR U8223 ( .A(n8083), .B(n8084), .Z(n8047) );
  XOR U8224 ( .A(n6388), .B(n6436), .Z(n8084) );
  XOR U8225 ( .A(n7056), .B(n8055), .Z(n6388) );
  XNOR U8226 ( .A(key[273]), .B(n8085), .Z(n8083) );
  XNOR U8227 ( .A(n8057), .B(n8086), .Z(n8079) );
  XNOR U8228 ( .A(key[275]), .B(n7058), .Z(n8086) );
  XOR U8229 ( .A(n7048), .B(n7012), .Z(n7058) );
  XNOR U8230 ( .A(n8087), .B(n8088), .Z(n7805) );
  XNOR U8231 ( .A(n8089), .B(n6427), .Z(n8088) );
  XNOR U8232 ( .A(n7045), .B(n8090), .Z(n6427) );
  XNOR U8233 ( .A(key[272]), .B(n7046), .Z(n8087) );
  XNOR U8234 ( .A(n7560), .B(n7456), .Z(n4948) );
  XNOR U8235 ( .A(n7591), .B(n8091), .Z(n7456) );
  XNOR U8236 ( .A(n8092), .B(n7547), .Z(n8091) );
  ANDN U8237 ( .B(n7600), .A(n8093), .Z(n7547) );
  XNOR U8238 ( .A(n7602), .B(n7549), .Z(n7600) );
  NOR U8239 ( .A(n8094), .B(n7602), .Z(n8092) );
  XNOR U8240 ( .A(n7545), .B(n8095), .Z(n7591) );
  XNOR U8241 ( .A(n8096), .B(n8097), .Z(n8095) );
  NAND U8242 ( .A(n8098), .B(n7606), .Z(n8097) );
  XOR U8243 ( .A(n7455), .B(n7484), .Z(n7560) );
  XOR U8244 ( .A(n7592), .B(n8099), .Z(n7484) );
  XOR U8245 ( .A(n8100), .B(n7583), .Z(n8099) );
  OR U8246 ( .A(n8101), .B(n8102), .Z(n7583) );
  NOR U8247 ( .A(n8103), .B(n8104), .Z(n8100) );
  XOR U8248 ( .A(n8105), .B(n7604), .Z(n7592) );
  OR U8249 ( .A(n8106), .B(n8107), .Z(n7604) );
  ANDN U8250 ( .B(n8108), .A(n8109), .Z(n8105) );
  XNOR U8251 ( .A(n7545), .B(n8110), .Z(n7455) );
  XNOR U8252 ( .A(n7588), .B(n8111), .Z(n8110) );
  NANDN U8253 ( .A(n8104), .B(n8112), .Z(n8111) );
  OR U8254 ( .A(n8102), .B(n8113), .Z(n7588) );
  XNOR U8255 ( .A(n7585), .B(n8104), .Z(n8102) );
  XOR U8256 ( .A(n8114), .B(n8096), .Z(n7545) );
  NANDN U8257 ( .A(n8106), .B(n8115), .Z(n8096) );
  XNOR U8258 ( .A(n8108), .B(n7606), .Z(n8106) );
  XNOR U8259 ( .A(n8104), .B(n7549), .Z(n7606) );
  XOR U8260 ( .A(n8116), .B(n8117), .Z(n7549) );
  NANDN U8261 ( .A(n8118), .B(n8119), .Z(n8117) );
  XNOR U8262 ( .A(n8120), .B(n8121), .Z(n8104) );
  OR U8263 ( .A(n8118), .B(n8122), .Z(n8121) );
  AND U8264 ( .A(n8108), .B(n8123), .Z(n8114) );
  XOR U8265 ( .A(n7585), .B(n7602), .Z(n8108) );
  XOR U8266 ( .A(n8124), .B(n8116), .Z(n7602) );
  NANDN U8267 ( .A(n8125), .B(n8126), .Z(n8116) );
  ANDN U8268 ( .B(n8127), .A(n8128), .Z(n8124) );
  NANDN U8269 ( .A(n8125), .B(n8130), .Z(n8120) );
  XOR U8270 ( .A(n8131), .B(n8118), .Z(n8125) );
  XNOR U8271 ( .A(n8132), .B(n8133), .Z(n8118) );
  XOR U8272 ( .A(n8134), .B(n8127), .Z(n8133) );
  XNOR U8273 ( .A(n8135), .B(n8136), .Z(n8132) );
  XNOR U8274 ( .A(n8137), .B(n8138), .Z(n8136) );
  ANDN U8275 ( .B(n8127), .A(n8139), .Z(n8137) );
  IV U8276 ( .A(n8140), .Z(n8127) );
  ANDN U8277 ( .B(n8131), .A(n8139), .Z(n8129) );
  IV U8278 ( .A(n8135), .Z(n8139) );
  IV U8279 ( .A(n8128), .Z(n8131) );
  XNOR U8280 ( .A(n8134), .B(n8141), .Z(n8128) );
  XOR U8281 ( .A(n8142), .B(n8138), .Z(n8141) );
  NAND U8282 ( .A(n8130), .B(n8126), .Z(n8138) );
  XNOR U8283 ( .A(n8119), .B(n8140), .Z(n8126) );
  XOR U8284 ( .A(n8143), .B(n8144), .Z(n8140) );
  XOR U8285 ( .A(n8145), .B(n8146), .Z(n8144) );
  XNOR U8286 ( .A(n8112), .B(n8147), .Z(n8146) );
  XNOR U8287 ( .A(n8148), .B(n8149), .Z(n8143) );
  XNOR U8288 ( .A(n8150), .B(n8151), .Z(n8149) );
  ANDN U8289 ( .B(n8152), .A(n7586), .Z(n8150) );
  XNOR U8290 ( .A(n8135), .B(n8122), .Z(n8130) );
  XOR U8291 ( .A(n8153), .B(n8154), .Z(n8135) );
  XNOR U8292 ( .A(n8155), .B(n8147), .Z(n8154) );
  XOR U8293 ( .A(n8156), .B(n8157), .Z(n8147) );
  XNOR U8294 ( .A(n8158), .B(n8159), .Z(n8157) );
  NAND U8295 ( .A(n7607), .B(n8098), .Z(n8159) );
  XNOR U8296 ( .A(n8160), .B(n8161), .Z(n8153) );
  ANDN U8297 ( .B(n8162), .A(n7601), .Z(n8160) );
  ANDN U8298 ( .B(n8119), .A(n8122), .Z(n8142) );
  XOR U8299 ( .A(n8122), .B(n8119), .Z(n8134) );
  XNOR U8300 ( .A(n8163), .B(n8164), .Z(n8119) );
  XNOR U8301 ( .A(n8156), .B(n8165), .Z(n8164) );
  XOR U8302 ( .A(n8155), .B(n7590), .Z(n8165) );
  XOR U8303 ( .A(n7586), .B(n8166), .Z(n8163) );
  XNOR U8304 ( .A(n8167), .B(n8151), .Z(n8166) );
  OR U8305 ( .A(n8113), .B(n8101), .Z(n8151) );
  XNOR U8306 ( .A(n7586), .B(n8103), .Z(n8101) );
  XOR U8307 ( .A(n7590), .B(n8112), .Z(n8113) );
  ANDN U8308 ( .B(n8112), .A(n8103), .Z(n8167) );
  XOR U8309 ( .A(n8168), .B(n8169), .Z(n8122) );
  XOR U8310 ( .A(n8156), .B(n8145), .Z(n8169) );
  XOR U8311 ( .A(n7596), .B(n7550), .Z(n8145) );
  XOR U8312 ( .A(n8170), .B(n8158), .Z(n8156) );
  NANDN U8313 ( .A(n8107), .B(n8115), .Z(n8158) );
  XOR U8314 ( .A(n8123), .B(n8098), .Z(n8115) );
  XNOR U8315 ( .A(n8162), .B(n8171), .Z(n8112) );
  XOR U8316 ( .A(n8172), .B(n8173), .Z(n8171) );
  XOR U8317 ( .A(n8109), .B(n7607), .Z(n8107) );
  XNOR U8318 ( .A(n8103), .B(n7596), .Z(n7607) );
  IV U8319 ( .A(n8148), .Z(n8103) );
  XOR U8320 ( .A(n8174), .B(n8175), .Z(n8148) );
  XOR U8321 ( .A(n8176), .B(n8177), .Z(n8175) );
  XNOR U8322 ( .A(n7586), .B(n8178), .Z(n8174) );
  ANDN U8323 ( .B(n8123), .A(n8109), .Z(n8170) );
  XNOR U8324 ( .A(n7586), .B(n7601), .Z(n8109) );
  XOR U8325 ( .A(n8162), .B(n8152), .Z(n8123) );
  IV U8326 ( .A(n7590), .Z(n8152) );
  XOR U8327 ( .A(n8179), .B(n8180), .Z(n7590) );
  XOR U8328 ( .A(n8181), .B(n8177), .Z(n8180) );
  XNOR U8329 ( .A(n8182), .B(n8183), .Z(n8177) );
  XNOR U8330 ( .A(n7178), .B(n8184), .Z(n8183) );
  XOR U8331 ( .A(n6244), .B(n8185), .Z(n7178) );
  XNOR U8332 ( .A(n7177), .B(n8186), .Z(n8182) );
  XNOR U8333 ( .A(key[316]), .B(n7193), .Z(n8186) );
  XNOR U8334 ( .A(n8187), .B(n7168), .Z(n7177) );
  IV U8335 ( .A(n8094), .Z(n8162) );
  XOR U8336 ( .A(n8155), .B(n8188), .Z(n8168) );
  XNOR U8337 ( .A(n8189), .B(n8161), .Z(n8188) );
  OR U8338 ( .A(n8093), .B(n7599), .Z(n8161) );
  XNOR U8339 ( .A(n8190), .B(n7596), .Z(n7599) );
  XNOR U8340 ( .A(n8094), .B(n7550), .Z(n8093) );
  ANDN U8341 ( .B(n7596), .A(n7550), .Z(n8189) );
  XOR U8342 ( .A(n8179), .B(n8191), .Z(n7550) );
  XNOR U8343 ( .A(n8192), .B(n8181), .Z(n8191) );
  XOR U8344 ( .A(n8181), .B(n8179), .Z(n7596) );
  XNOR U8345 ( .A(n7601), .B(n8094), .Z(n8155) );
  XOR U8346 ( .A(n8179), .B(n8193), .Z(n8094) );
  XNOR U8347 ( .A(n8181), .B(n8176), .Z(n8193) );
  XOR U8348 ( .A(n8194), .B(n8195), .Z(n8176) );
  XNOR U8349 ( .A(n7163), .B(n7174), .Z(n8195) );
  XNOR U8350 ( .A(n8196), .B(n8197), .Z(n7174) );
  XNOR U8351 ( .A(key[319]), .B(n7197), .Z(n8194) );
  XNOR U8352 ( .A(n8198), .B(n8199), .Z(n7197) );
  XNOR U8353 ( .A(n8200), .B(n8201), .Z(n8179) );
  XNOR U8354 ( .A(n7181), .B(n7166), .Z(n8201) );
  XNOR U8355 ( .A(n6261), .B(n8202), .Z(n7166) );
  XNOR U8356 ( .A(n8203), .B(n8204), .Z(n8200) );
  XNOR U8357 ( .A(key[317]), .B(n8205), .Z(n8204) );
  IV U8358 ( .A(n8190), .Z(n7601) );
  XNOR U8359 ( .A(n8173), .B(n8206), .Z(n8190) );
  XOR U8360 ( .A(n8207), .B(n8208), .Z(n8181) );
  XNOR U8361 ( .A(n7586), .B(n8209), .Z(n8208) );
  XNOR U8362 ( .A(n8210), .B(n8211), .Z(n7586) );
  XOR U8363 ( .A(n8212), .B(n6254), .Z(n8211) );
  XOR U8364 ( .A(key[312]), .B(n8214), .Z(n8213) );
  XNOR U8365 ( .A(n6259), .B(n8215), .Z(n8207) );
  XNOR U8366 ( .A(key[318]), .B(n7159), .Z(n8215) );
  XNOR U8367 ( .A(n8216), .B(n7173), .Z(n7159) );
  XOR U8368 ( .A(n8187), .B(n8217), .Z(n7173) );
  XOR U8369 ( .A(n8218), .B(n8219), .Z(n8178) );
  XNOR U8370 ( .A(n8220), .B(n8221), .Z(n8219) );
  XNOR U8371 ( .A(n6295), .B(n8192), .Z(n8221) );
  IV U8372 ( .A(n8172), .Z(n8192) );
  XNOR U8373 ( .A(n8222), .B(n8223), .Z(n8172) );
  XNOR U8374 ( .A(n7189), .B(n6296), .Z(n8223) );
  XNOR U8375 ( .A(n7152), .B(n8224), .Z(n8222) );
  XOR U8376 ( .A(key[313]), .B(n6274), .Z(n8224) );
  XNOR U8377 ( .A(n7184), .B(n8225), .Z(n8218) );
  XOR U8378 ( .A(key[315]), .B(n7186), .Z(n8225) );
  XOR U8379 ( .A(n8199), .B(n7180), .Z(n7186) );
  IV U8380 ( .A(n8226), .Z(n7184) );
  XOR U8381 ( .A(n8227), .B(n8228), .Z(n8173) );
  XOR U8382 ( .A(n6290), .B(n7151), .Z(n8228) );
  XNOR U8383 ( .A(n7191), .B(n8229), .Z(n8227) );
  XOR U8384 ( .A(n5309), .B(n8230), .Z(n1034) );
  XNOR U8385 ( .A(n5311), .B(n5327), .Z(n8230) );
  XOR U8386 ( .A(n5430), .B(n8231), .Z(n5425) );
  XOR U8387 ( .A(n8232), .B(n5400), .Z(n8231) );
  OR U8388 ( .A(n8233), .B(n8234), .Z(n5400) );
  ANDN U8389 ( .B(n8235), .A(n8236), .Z(n8232) );
  XNOR U8390 ( .A(n5391), .B(n8237), .Z(n5312) );
  XNOR U8391 ( .A(n8238), .B(n8239), .Z(n8237) );
  NANDN U8392 ( .A(n8240), .B(n8241), .Z(n8239) );
  XOR U8393 ( .A(n5430), .B(n8242), .Z(n5311) );
  XNOR U8394 ( .A(n5428), .B(n8243), .Z(n8242) );
  NANDN U8395 ( .A(n8244), .B(n5395), .Z(n8243) );
  XNOR U8396 ( .A(n5357), .B(n5395), .Z(n5397) );
  XOR U8397 ( .A(n8246), .B(n5432), .Z(n5430) );
  OR U8398 ( .A(n8247), .B(n8248), .Z(n5432) );
  ANDN U8399 ( .B(n8249), .A(n8250), .Z(n8246) );
  XOR U8400 ( .A(n5352), .B(n8251), .Z(n5309) );
  XNOR U8401 ( .A(n8238), .B(n8252), .Z(n8251) );
  NANDN U8402 ( .A(n8253), .B(n5403), .Z(n8252) );
  OR U8403 ( .A(n8234), .B(n8254), .Z(n8238) );
  XNOR U8404 ( .A(n5403), .B(n8241), .Z(n8234) );
  XNOR U8405 ( .A(n5391), .B(n8255), .Z(n5352) );
  XNOR U8406 ( .A(n8256), .B(n8257), .Z(n8255) );
  NANDN U8407 ( .A(n5434), .B(n8258), .Z(n8257) );
  XOR U8408 ( .A(n8259), .B(n8256), .Z(n5391) );
  NANDN U8409 ( .A(n8247), .B(n8260), .Z(n8256) );
  XOR U8410 ( .A(n8249), .B(n5434), .Z(n8247) );
  XNOR U8411 ( .A(n8241), .B(n5395), .Z(n5434) );
  XOR U8412 ( .A(n8261), .B(n8262), .Z(n5395) );
  NANDN U8413 ( .A(n8263), .B(n8264), .Z(n8262) );
  IV U8414 ( .A(n8236), .Z(n8241) );
  XNOR U8415 ( .A(n8265), .B(n8266), .Z(n8236) );
  NANDN U8416 ( .A(n8263), .B(n8267), .Z(n8266) );
  IV U8417 ( .A(n8268), .Z(n8249) );
  ANDN U8418 ( .B(n8269), .A(n8268), .Z(n8259) );
  XOR U8419 ( .A(n5357), .B(n5403), .Z(n8268) );
  XNOR U8420 ( .A(n8270), .B(n8265), .Z(n5403) );
  NANDN U8421 ( .A(n8271), .B(n8272), .Z(n8265) );
  XOR U8422 ( .A(n8267), .B(n8273), .Z(n8272) );
  ANDN U8423 ( .B(n8273), .A(n8274), .Z(n8270) );
  XOR U8424 ( .A(n8275), .B(n8261), .Z(n5357) );
  NANDN U8425 ( .A(n8271), .B(n8276), .Z(n8261) );
  XOR U8426 ( .A(n8277), .B(n8264), .Z(n8276) );
  XNOR U8427 ( .A(n8278), .B(n8279), .Z(n8263) );
  XOR U8428 ( .A(n8280), .B(n8281), .Z(n8279) );
  XNOR U8429 ( .A(n8282), .B(n8283), .Z(n8278) );
  XNOR U8430 ( .A(n8284), .B(n8285), .Z(n8283) );
  ANDN U8431 ( .B(n8277), .A(n8281), .Z(n8284) );
  ANDN U8432 ( .B(n8277), .A(n8274), .Z(n8275) );
  XNOR U8433 ( .A(n8280), .B(n8286), .Z(n8274) );
  XOR U8434 ( .A(n8287), .B(n8285), .Z(n8286) );
  NAND U8435 ( .A(n8288), .B(n8289), .Z(n8285) );
  XNOR U8436 ( .A(n8282), .B(n8264), .Z(n8289) );
  IV U8437 ( .A(n8277), .Z(n8282) );
  XNOR U8438 ( .A(n8267), .B(n8281), .Z(n8288) );
  IV U8439 ( .A(n8273), .Z(n8281) );
  XOR U8440 ( .A(n8290), .B(n8291), .Z(n8273) );
  XNOR U8441 ( .A(n8292), .B(n8293), .Z(n8291) );
  XNOR U8442 ( .A(n8294), .B(n8295), .Z(n8290) );
  NOR U8443 ( .A(n5356), .B(n5429), .Z(n8294) );
  AND U8444 ( .A(n8264), .B(n8267), .Z(n8287) );
  XNOR U8445 ( .A(n8264), .B(n8267), .Z(n8280) );
  XNOR U8446 ( .A(n8296), .B(n8297), .Z(n8267) );
  XNOR U8447 ( .A(n8298), .B(n8293), .Z(n8297) );
  XOR U8448 ( .A(n8299), .B(n8300), .Z(n8296) );
  XNOR U8449 ( .A(n8301), .B(n8295), .Z(n8300) );
  OR U8450 ( .A(n5398), .B(n8245), .Z(n8295) );
  XNOR U8451 ( .A(n5429), .B(n8244), .Z(n8245) );
  XNOR U8452 ( .A(n5356), .B(n5396), .Z(n5398) );
  ANDN U8453 ( .B(n8302), .A(n8244), .Z(n8301) );
  XNOR U8454 ( .A(n8303), .B(n8304), .Z(n8264) );
  XNOR U8455 ( .A(n8293), .B(n8305), .Z(n8304) );
  XOR U8456 ( .A(n8253), .B(n8299), .Z(n8305) );
  XNOR U8457 ( .A(n5429), .B(n8306), .Z(n8293) );
  XNOR U8458 ( .A(n8307), .B(n8308), .Z(n8303) );
  XNOR U8459 ( .A(n8309), .B(n8310), .Z(n8308) );
  ANDN U8460 ( .B(n8235), .A(n8240), .Z(n8309) );
  XNOR U8461 ( .A(n8311), .B(n8312), .Z(n8277) );
  XNOR U8462 ( .A(n8298), .B(n8313), .Z(n8312) );
  XNOR U8463 ( .A(n8240), .B(n8292), .Z(n8313) );
  XOR U8464 ( .A(n8299), .B(n8314), .Z(n8292) );
  XNOR U8465 ( .A(n8315), .B(n8316), .Z(n8314) );
  NAND U8466 ( .A(n5435), .B(n8258), .Z(n8316) );
  XNOR U8467 ( .A(n8317), .B(n8315), .Z(n8299) );
  NANDN U8468 ( .A(n8248), .B(n8260), .Z(n8315) );
  XOR U8469 ( .A(n8269), .B(n8258), .Z(n8260) );
  XNOR U8470 ( .A(n8318), .B(n5396), .Z(n8258) );
  XOR U8471 ( .A(n8250), .B(n5435), .Z(n8248) );
  XOR U8472 ( .A(n8235), .B(n8319), .Z(n5435) );
  ANDN U8473 ( .B(n8269), .A(n8250), .Z(n8317) );
  XOR U8474 ( .A(n8307), .B(n5429), .Z(n8250) );
  XOR U8475 ( .A(n8320), .B(n8321), .Z(n5429) );
  XNOR U8476 ( .A(n8322), .B(n8323), .Z(n8321) );
  XOR U8477 ( .A(n8319), .B(n8302), .Z(n8298) );
  IV U8478 ( .A(n5396), .Z(n8302) );
  XOR U8479 ( .A(n8324), .B(n8325), .Z(n5396) );
  XNOR U8480 ( .A(n8326), .B(n8323), .Z(n8325) );
  IV U8481 ( .A(n8244), .Z(n8319) );
  XOR U8482 ( .A(n8323), .B(n8327), .Z(n8244) );
  XNOR U8483 ( .A(n8235), .B(n8328), .Z(n8311) );
  XNOR U8484 ( .A(n8329), .B(n8310), .Z(n8328) );
  OR U8485 ( .A(n8254), .B(n8233), .Z(n8310) );
  XNOR U8486 ( .A(n8307), .B(n8235), .Z(n8233) );
  XOR U8487 ( .A(n8253), .B(n8318), .Z(n8254) );
  IV U8488 ( .A(n8240), .Z(n8318) );
  XOR U8489 ( .A(n8306), .B(n8330), .Z(n8240) );
  XNOR U8490 ( .A(n8326), .B(n8320), .Z(n8330) );
  XOR U8491 ( .A(n8331), .B(n8332), .Z(n8320) );
  XNOR U8492 ( .A(n5211), .B(n3019), .Z(n8332) );
  XOR U8493 ( .A(n3976), .B(n3045), .Z(n3019) );
  XOR U8494 ( .A(n3981), .B(n3935), .Z(n5211) );
  XOR U8495 ( .A(n8333), .B(n8334), .Z(n3981) );
  XNOR U8496 ( .A(n8335), .B(n8336), .Z(n8334) );
  XOR U8497 ( .A(n8337), .B(n8338), .Z(n8333) );
  XOR U8498 ( .A(key[450]), .B(n3975), .Z(n8331) );
  ANDN U8499 ( .B(n8339), .A(n5402), .Z(n8329) );
  XOR U8500 ( .A(n8340), .B(n8341), .Z(n8235) );
  XNOR U8501 ( .A(n8342), .B(n8343), .Z(n8341) );
  XOR U8502 ( .A(n8307), .B(n8322), .Z(n8340) );
  XOR U8503 ( .A(n8344), .B(n8345), .Z(n8322) );
  XNOR U8504 ( .A(n8326), .B(n8346), .Z(n8345) );
  XOR U8505 ( .A(n3982), .B(n3971), .Z(n8346) );
  XOR U8506 ( .A(n8347), .B(n5204), .Z(n3971) );
  XOR U8507 ( .A(n3005), .B(n3936), .Z(n3982) );
  XNOR U8508 ( .A(n8348), .B(n8349), .Z(n3936) );
  XOR U8509 ( .A(n8350), .B(n8351), .Z(n8349) );
  XNOR U8510 ( .A(n8352), .B(n8353), .Z(n8348) );
  XNOR U8511 ( .A(n8354), .B(n8355), .Z(n3005) );
  XOR U8512 ( .A(n8356), .B(n8357), .Z(n8355) );
  XOR U8513 ( .A(n8358), .B(n8359), .Z(n8354) );
  XOR U8514 ( .A(n8360), .B(n8361), .Z(n8326) );
  XNOR U8515 ( .A(n8362), .B(n3038), .Z(n8361) );
  XNOR U8516 ( .A(n3020), .B(n3985), .Z(n3038) );
  XNOR U8517 ( .A(n8351), .B(n8363), .Z(n3985) );
  XNOR U8518 ( .A(n8352), .B(n8364), .Z(n8363) );
  XOR U8519 ( .A(n8356), .B(n8365), .Z(n3020) );
  XOR U8520 ( .A(n8366), .B(n8359), .Z(n8365) );
  IV U8521 ( .A(n8367), .Z(n8356) );
  XOR U8522 ( .A(key[449]), .B(n5180), .Z(n8360) );
  XOR U8523 ( .A(n5217), .B(n3975), .Z(n5180) );
  XNOR U8524 ( .A(n3935), .B(n8368), .Z(n8344) );
  XNOR U8525 ( .A(key[451]), .B(n5213), .Z(n8368) );
  XOR U8526 ( .A(n5200), .B(n3967), .Z(n5213) );
  XOR U8527 ( .A(n8369), .B(n5217), .Z(n3967) );
  XOR U8528 ( .A(n8370), .B(n8335), .Z(n5217) );
  XOR U8529 ( .A(n8371), .B(n8372), .Z(n3935) );
  XOR U8530 ( .A(n8373), .B(n8374), .Z(n8372) );
  XOR U8531 ( .A(n8375), .B(n8376), .Z(n8371) );
  XOR U8532 ( .A(n8339), .B(n8306), .Z(n8269) );
  IV U8533 ( .A(n5356), .Z(n8306) );
  XOR U8534 ( .A(n8324), .B(n8377), .Z(n5356) );
  XOR U8535 ( .A(n8323), .B(n8343), .Z(n8377) );
  XNOR U8536 ( .A(n8378), .B(n8379), .Z(n8343) );
  XOR U8537 ( .A(n8380), .B(n3962), .Z(n8379) );
  XNOR U8538 ( .A(n5193), .B(n3949), .Z(n3962) );
  XNOR U8539 ( .A(n8381), .B(n8382), .Z(n3949) );
  XOR U8540 ( .A(n8351), .B(n8383), .Z(n8382) );
  XOR U8541 ( .A(n8384), .B(n8385), .Z(n8351) );
  XNOR U8542 ( .A(n8386), .B(n8387), .Z(n8385) );
  OR U8543 ( .A(n8388), .B(n8389), .Z(n8387) );
  XOR U8544 ( .A(n8352), .B(n8364), .Z(n8381) );
  XOR U8545 ( .A(n8390), .B(n8391), .Z(n5193) );
  XNOR U8546 ( .A(n8367), .B(n8392), .Z(n8391) );
  XNOR U8547 ( .A(n8393), .B(n8394), .Z(n8367) );
  XNOR U8548 ( .A(n8395), .B(n8396), .Z(n8394) );
  ANDN U8549 ( .B(n8397), .A(n8398), .Z(n8395) );
  XNOR U8550 ( .A(n8366), .B(n8359), .Z(n8390) );
  XOR U8551 ( .A(key[455]), .B(n5200), .Z(n8378) );
  IV U8552 ( .A(n8253), .Z(n8339) );
  XOR U8553 ( .A(n8324), .B(n8399), .Z(n8253) );
  XOR U8554 ( .A(n8323), .B(n8342), .Z(n8399) );
  XNOR U8555 ( .A(n8400), .B(n3965), .Z(n8342) );
  XNOR U8556 ( .A(n8401), .B(n8402), .Z(n3965) );
  XNOR U8557 ( .A(n3014), .B(n3979), .Z(n8402) );
  XOR U8558 ( .A(n8403), .B(n3976), .Z(n3979) );
  IV U8559 ( .A(n5181), .Z(n3976) );
  XOR U8560 ( .A(n8404), .B(n8352), .Z(n5181) );
  XOR U8561 ( .A(n8405), .B(n8406), .Z(n8352) );
  XOR U8562 ( .A(n8407), .B(n8408), .Z(n8406) );
  NAND U8563 ( .A(n8409), .B(n8410), .Z(n8408) );
  XOR U8564 ( .A(n8411), .B(n3045), .Z(n3014) );
  XNOR U8565 ( .A(n8412), .B(n8359), .Z(n3045) );
  XOR U8566 ( .A(n8413), .B(n8414), .Z(n8359) );
  XNOR U8567 ( .A(n8415), .B(n8416), .Z(n8414) );
  NANDN U8568 ( .A(n8417), .B(n8418), .Z(n8416) );
  XNOR U8569 ( .A(n3039), .B(n5188), .Z(n8401) );
  IV U8570 ( .A(n8347), .Z(n3039) );
  XNOR U8571 ( .A(n5204), .B(n8419), .Z(n8400) );
  XNOR U8572 ( .A(key[452]), .B(n5205), .Z(n8419) );
  XOR U8573 ( .A(n8420), .B(n3952), .Z(n5205) );
  XNOR U8574 ( .A(n8421), .B(n8422), .Z(n3952) );
  XNOR U8575 ( .A(n8369), .B(n8423), .Z(n8422) );
  XNOR U8576 ( .A(n8424), .B(n8425), .Z(n8421) );
  XNOR U8577 ( .A(n8426), .B(n8427), .Z(n8425) );
  ANDN U8578 ( .B(n8428), .A(n8429), .Z(n8426) );
  XOR U8579 ( .A(n8430), .B(n3975), .Z(n5204) );
  XNOR U8580 ( .A(n8431), .B(n8432), .Z(n3975) );
  XOR U8581 ( .A(n8433), .B(n8434), .Z(n8323) );
  XNOR U8582 ( .A(n3945), .B(n5402), .Z(n8434) );
  IV U8583 ( .A(n8307), .Z(n5402) );
  XOR U8584 ( .A(n8435), .B(n8436), .Z(n8307) );
  XNOR U8585 ( .A(n5207), .B(n3018), .Z(n8436) );
  XOR U8586 ( .A(n3978), .B(n8362), .Z(n3018) );
  IV U8587 ( .A(n3986), .Z(n8362) );
  XOR U8588 ( .A(n8374), .B(n8437), .Z(n3986) );
  XOR U8589 ( .A(n8375), .B(n8438), .Z(n8437) );
  IV U8590 ( .A(n8439), .Z(n8374) );
  XNOR U8591 ( .A(n8337), .B(n8441), .Z(n8440) );
  IV U8592 ( .A(n5192), .Z(n5207) );
  XOR U8593 ( .A(n8412), .B(n8411), .Z(n5192) );
  XNOR U8594 ( .A(key[448]), .B(n3963), .Z(n8435) );
  XNOR U8595 ( .A(n8347), .B(n3948), .Z(n3963) );
  IV U8596 ( .A(n3031), .Z(n3948) );
  XOR U8597 ( .A(n3025), .B(n8380), .Z(n3945) );
  XNOR U8598 ( .A(n8347), .B(n5201), .Z(n8380) );
  XNOR U8599 ( .A(n8442), .B(n8443), .Z(n5201) );
  XNOR U8600 ( .A(n8439), .B(n8444), .Z(n8443) );
  XNOR U8601 ( .A(n8445), .B(n8446), .Z(n8439) );
  XNOR U8602 ( .A(n8447), .B(n8448), .Z(n8446) );
  OR U8603 ( .A(n8449), .B(n8450), .Z(n8448) );
  XNOR U8604 ( .A(n8375), .B(n8438), .Z(n8442) );
  IV U8605 ( .A(n8432), .Z(n8375) );
  XOR U8606 ( .A(n8451), .B(n8452), .Z(n8432) );
  XOR U8607 ( .A(n8453), .B(n8454), .Z(n8452) );
  NAND U8608 ( .A(n8455), .B(n8456), .Z(n8454) );
  XOR U8609 ( .A(n8431), .B(n8430), .Z(n8347) );
  XOR U8610 ( .A(n3956), .B(n3040), .Z(n3025) );
  XOR U8611 ( .A(n8357), .B(n8366), .Z(n3040) );
  XOR U8612 ( .A(n8412), .B(n8358), .Z(n8366) );
  XOR U8613 ( .A(n8457), .B(n8458), .Z(n8358) );
  XOR U8614 ( .A(n8396), .B(n8459), .Z(n8458) );
  OR U8615 ( .A(n8460), .B(n8461), .Z(n8459) );
  NOR U8616 ( .A(n8462), .B(n8463), .Z(n8396) );
  XNOR U8617 ( .A(n8413), .B(n8464), .Z(n8412) );
  XNOR U8618 ( .A(n8465), .B(n8466), .Z(n8464) );
  NOR U8619 ( .A(n8467), .B(n8460), .Z(n8465) );
  XNOR U8620 ( .A(n8393), .B(n8468), .Z(n8357) );
  XOR U8621 ( .A(n8469), .B(n8470), .Z(n8468) );
  NOR U8622 ( .A(n8471), .B(n8472), .Z(n8469) );
  XNOR U8623 ( .A(n8457), .B(n8473), .Z(n8393) );
  XNOR U8624 ( .A(n8474), .B(n8475), .Z(n8473) );
  NANDN U8625 ( .A(n8476), .B(n8477), .Z(n8475) );
  XOR U8626 ( .A(n8364), .B(n8350), .Z(n3956) );
  XNOR U8627 ( .A(n8384), .B(n8478), .Z(n8350) );
  XNOR U8628 ( .A(n8479), .B(n8480), .Z(n8478) );
  ANDN U8629 ( .B(n8481), .A(n8482), .Z(n8479) );
  XNOR U8630 ( .A(n8483), .B(n8484), .Z(n8384) );
  XNOR U8631 ( .A(n8485), .B(n8486), .Z(n8484) );
  NANDN U8632 ( .A(n8487), .B(n8488), .Z(n8486) );
  XOR U8633 ( .A(n8404), .B(n8353), .Z(n8364) );
  XNOR U8634 ( .A(n8483), .B(n8489), .Z(n8353) );
  XNOR U8635 ( .A(n8386), .B(n8490), .Z(n8489) );
  NANDN U8636 ( .A(n8491), .B(n8492), .Z(n8490) );
  OR U8637 ( .A(n8493), .B(n8494), .Z(n8386) );
  XNOR U8638 ( .A(n8405), .B(n8495), .Z(n8404) );
  XOR U8639 ( .A(n8496), .B(n8497), .Z(n8495) );
  NOR U8640 ( .A(n8498), .B(n8491), .Z(n8496) );
  XNOR U8641 ( .A(n3954), .B(n8499), .Z(n8433) );
  XNOR U8642 ( .A(key[454]), .B(n5194), .Z(n8499) );
  XOR U8643 ( .A(n8420), .B(n3961), .Z(n5194) );
  XNOR U8644 ( .A(n8500), .B(n8501), .Z(n3961) );
  XNOR U8645 ( .A(n8335), .B(n8423), .Z(n8501) );
  XNOR U8646 ( .A(n8502), .B(n8503), .Z(n8423) );
  XNOR U8647 ( .A(n8504), .B(n8505), .Z(n8503) );
  NANDN U8648 ( .A(n8506), .B(n8507), .Z(n8505) );
  XNOR U8649 ( .A(n8508), .B(n8509), .Z(n8335) );
  XNOR U8650 ( .A(n8510), .B(n8511), .Z(n8509) );
  NANDN U8651 ( .A(n8512), .B(n8428), .Z(n8511) );
  XOR U8652 ( .A(n8337), .B(n8441), .Z(n8500) );
  XNOR U8653 ( .A(n8370), .B(n8338), .Z(n8441) );
  XNOR U8654 ( .A(n8514), .B(n8515), .Z(n8513) );
  NANDN U8655 ( .A(n8506), .B(n8516), .Z(n8515) );
  IV U8656 ( .A(n5200), .Z(n8420) );
  XOR U8657 ( .A(n8370), .B(n8369), .Z(n5200) );
  XNOR U8658 ( .A(n8502), .B(n8518), .Z(n8369) );
  XOR U8659 ( .A(n8519), .B(n8510), .Z(n8518) );
  NANDN U8660 ( .A(n8520), .B(n8521), .Z(n8510) );
  ANDN U8661 ( .B(n8522), .A(n8523), .Z(n8519) );
  XNOR U8662 ( .A(n8508), .B(n8524), .Z(n8502) );
  XNOR U8663 ( .A(n8525), .B(n8526), .Z(n8524) );
  NAND U8664 ( .A(n8527), .B(n8528), .Z(n8526) );
  IV U8665 ( .A(n8327), .Z(n8324) );
  XOR U8666 ( .A(n8529), .B(n8530), .Z(n8327) );
  XOR U8667 ( .A(n5188), .B(n3953), .Z(n8530) );
  XNOR U8668 ( .A(n3968), .B(n3024), .Z(n3953) );
  XOR U8669 ( .A(n8531), .B(n8532), .Z(n3024) );
  XNOR U8670 ( .A(n8411), .B(n8392), .Z(n8532) );
  XNOR U8671 ( .A(n8533), .B(n8534), .Z(n8392) );
  XOR U8672 ( .A(n8466), .B(n8535), .Z(n8534) );
  NANDN U8673 ( .A(n8536), .B(n8397), .Z(n8535) );
  NOR U8674 ( .A(n8462), .B(n8537), .Z(n8466) );
  XOR U8675 ( .A(n8397), .B(n8460), .Z(n8462) );
  XNOR U8676 ( .A(n8533), .B(n8538), .Z(n8411) );
  XNOR U8677 ( .A(n8415), .B(n8539), .Z(n8538) );
  NANDN U8678 ( .A(n8472), .B(n8540), .Z(n8539) );
  OR U8679 ( .A(n8541), .B(n8542), .Z(n8415) );
  XNOR U8680 ( .A(n8413), .B(n8543), .Z(n8533) );
  XNOR U8681 ( .A(n8544), .B(n8545), .Z(n8543) );
  NANDN U8682 ( .A(n8476), .B(n8546), .Z(n8545) );
  XOR U8683 ( .A(n8547), .B(n8544), .Z(n8413) );
  OR U8684 ( .A(n8548), .B(n8549), .Z(n8544) );
  ANDN U8685 ( .B(n8550), .A(n8551), .Z(n8547) );
  XNOR U8686 ( .A(n8457), .B(n8552), .Z(n8531) );
  XNOR U8687 ( .A(n8470), .B(n8553), .Z(n8552) );
  ANDN U8688 ( .B(n8418), .A(n8554), .Z(n8553) );
  OR U8689 ( .A(n8541), .B(n8555), .Z(n8470) );
  XOR U8690 ( .A(n8472), .B(n8418), .Z(n8541) );
  XOR U8691 ( .A(n8556), .B(n8474), .Z(n8457) );
  NANDN U8692 ( .A(n8548), .B(n8557), .Z(n8474) );
  XOR U8693 ( .A(n8550), .B(n8476), .Z(n8548) );
  XOR U8694 ( .A(n8418), .B(n8460), .Z(n8476) );
  XOR U8695 ( .A(n8558), .B(n8559), .Z(n8460) );
  OR U8696 ( .A(n8560), .B(n8561), .Z(n8559) );
  XOR U8697 ( .A(n8562), .B(n8563), .Z(n8418) );
  NANDN U8698 ( .A(n8560), .B(n8564), .Z(n8563) );
  AND U8699 ( .A(n8565), .B(n8550), .Z(n8556) );
  XNOR U8700 ( .A(n8472), .B(n8397), .Z(n8550) );
  XOR U8701 ( .A(n8566), .B(n8558), .Z(n8397) );
  ANDN U8702 ( .B(n8567), .A(n8568), .Z(n8558) );
  NOR U8703 ( .A(n8569), .B(n8570), .Z(n8566) );
  XNOR U8704 ( .A(n8562), .B(n8571), .Z(n8472) );
  NANDN U8705 ( .A(n8569), .B(n8572), .Z(n8571) );
  NANDN U8706 ( .A(n8568), .B(n8573), .Z(n8562) );
  XNOR U8707 ( .A(n8574), .B(n8575), .Z(n8560) );
  XOR U8708 ( .A(n8576), .B(n8570), .Z(n8575) );
  XOR U8709 ( .A(n8572), .B(n8577), .Z(n8574) );
  XNOR U8710 ( .A(n8578), .B(n8579), .Z(n8577) );
  ANDN U8711 ( .B(n8572), .A(n8570), .Z(n8578) );
  XNOR U8712 ( .A(n8576), .B(n8580), .Z(n8569) );
  XNOR U8713 ( .A(n8579), .B(n8581), .Z(n8580) );
  NANDN U8714 ( .A(n8561), .B(n8564), .Z(n8581) );
  XOR U8715 ( .A(n8572), .B(n8564), .Z(n8573) );
  XNOR U8716 ( .A(n8582), .B(n8583), .Z(n8572) );
  XNOR U8717 ( .A(n8584), .B(n8585), .Z(n8583) );
  XNOR U8718 ( .A(n8461), .B(n8586), .Z(n8585) );
  XNOR U8719 ( .A(n8587), .B(n8588), .Z(n8582) );
  XNOR U8720 ( .A(n8589), .B(n8590), .Z(n8588) );
  NOR U8721 ( .A(n8398), .B(n8536), .Z(n8589) );
  XOR U8722 ( .A(n8561), .B(n8570), .Z(n8567) );
  XNOR U8723 ( .A(n8591), .B(n8592), .Z(n8570) );
  XNOR U8724 ( .A(n8586), .B(n8593), .Z(n8592) );
  XOR U8725 ( .A(n8594), .B(n8595), .Z(n8586) );
  XNOR U8726 ( .A(n8596), .B(n8597), .Z(n8595) );
  NAND U8727 ( .A(n8546), .B(n8477), .Z(n8597) );
  XNOR U8728 ( .A(n8598), .B(n8599), .Z(n8591) );
  ANDN U8729 ( .B(n8540), .A(n8471), .Z(n8598) );
  XOR U8730 ( .A(n8564), .B(n8561), .Z(n8576) );
  XOR U8731 ( .A(n8600), .B(n8601), .Z(n8561) );
  XNOR U8732 ( .A(n8584), .B(n8593), .Z(n8601) );
  XOR U8733 ( .A(n8602), .B(n8603), .Z(n8584) );
  XOR U8734 ( .A(n8594), .B(n8604), .Z(n8600) );
  XNOR U8735 ( .A(n8605), .B(n8599), .Z(n8604) );
  OR U8736 ( .A(n8555), .B(n8542), .Z(n8599) );
  XNOR U8737 ( .A(n8540), .B(n8602), .Z(n8542) );
  XNOR U8738 ( .A(n8471), .B(n8554), .Z(n8555) );
  ANDN U8739 ( .B(n8603), .A(n8417), .Z(n8605) );
  IV U8740 ( .A(n8554), .Z(n8603) );
  XNOR U8741 ( .A(n8606), .B(n8607), .Z(n8564) );
  XNOR U8742 ( .A(n8593), .B(n8608), .Z(n8607) );
  XOR U8743 ( .A(n8398), .B(n8594), .Z(n8608) );
  XNOR U8744 ( .A(n8609), .B(n8596), .Z(n8594) );
  NANDN U8745 ( .A(n8549), .B(n8557), .Z(n8596) );
  XOR U8746 ( .A(n8565), .B(n8477), .Z(n8557) );
  XNOR U8747 ( .A(n8610), .B(n8554), .Z(n8477) );
  XOR U8748 ( .A(n8611), .B(n8612), .Z(n8554) );
  XOR U8749 ( .A(n8613), .B(n8614), .Z(n8612) );
  XOR U8750 ( .A(n8551), .B(n8546), .Z(n8549) );
  XNOR U8751 ( .A(n8467), .B(n8602), .Z(n8546) );
  IV U8752 ( .A(n8417), .Z(n8602) );
  XOR U8753 ( .A(n8614), .B(n8615), .Z(n8417) );
  ANDN U8754 ( .B(n8565), .A(n8551), .Z(n8609) );
  XOR U8755 ( .A(n8536), .B(n8540), .Z(n8551) );
  XNOR U8756 ( .A(n8540), .B(n8471), .Z(n8593) );
  XNOR U8757 ( .A(n8614), .B(n8616), .Z(n8540) );
  XOR U8758 ( .A(n8617), .B(n8618), .Z(n8616) );
  XOR U8759 ( .A(n8536), .B(n8619), .Z(n8606) );
  XNOR U8760 ( .A(n8620), .B(n8590), .Z(n8619) );
  OR U8761 ( .A(n8463), .B(n8537), .Z(n8590) );
  XNOR U8762 ( .A(n8536), .B(n8467), .Z(n8537) );
  XOR U8763 ( .A(n8398), .B(n8610), .Z(n8463) );
  ANDN U8764 ( .B(n8610), .A(n8467), .Z(n8620) );
  IV U8765 ( .A(n8587), .Z(n8467) );
  XOR U8766 ( .A(n8621), .B(n8622), .Z(n8587) );
  XNOR U8767 ( .A(n8623), .B(n8624), .Z(n8622) );
  XOR U8768 ( .A(n8536), .B(n8618), .Z(n8621) );
  XNOR U8769 ( .A(n8625), .B(n8626), .Z(n8618) );
  XNOR U8770 ( .A(n6424), .B(n8627), .Z(n8626) );
  XNOR U8771 ( .A(n6389), .B(n8613), .Z(n8627) );
  XOR U8772 ( .A(n7052), .B(n6423), .Z(n6389) );
  XNOR U8773 ( .A(n8628), .B(n8629), .Z(n6423) );
  XOR U8774 ( .A(n8630), .B(n8631), .Z(n8629) );
  XNOR U8775 ( .A(n8632), .B(n8633), .Z(n8628) );
  XOR U8776 ( .A(n8634), .B(n7011), .Z(n6424) );
  XNOR U8777 ( .A(n8082), .B(n8635), .Z(n8625) );
  XNOR U8778 ( .A(key[267]), .B(n7064), .Z(n8635) );
  XOR U8779 ( .A(n8636), .B(n8637), .Z(n7064) );
  XOR U8780 ( .A(n8638), .B(n8639), .Z(n8637) );
  XNOR U8781 ( .A(n8640), .B(n8641), .Z(n8636) );
  XOR U8782 ( .A(n6437), .B(n7013), .Z(n8082) );
  XOR U8783 ( .A(n8642), .B(n8055), .Z(n7013) );
  IV U8784 ( .A(n8461), .Z(n8610) );
  XOR U8785 ( .A(n8643), .B(n8644), .Z(n8461) );
  XOR U8786 ( .A(n8617), .B(n8613), .Z(n8644) );
  XNOR U8787 ( .A(n8645), .B(n8646), .Z(n8613) );
  XOR U8788 ( .A(n7062), .B(n6436), .Z(n8646) );
  XNOR U8789 ( .A(n6429), .B(n7055), .Z(n6436) );
  XOR U8790 ( .A(n8647), .B(n8648), .Z(n6429) );
  XOR U8791 ( .A(n8632), .B(n8633), .Z(n8648) );
  XOR U8792 ( .A(n8055), .B(n8649), .Z(n8645) );
  XOR U8793 ( .A(key[265]), .B(n7045), .Z(n8649) );
  XNOR U8794 ( .A(n8650), .B(n8651), .Z(n7045) );
  XOR U8795 ( .A(n8640), .B(n8641), .Z(n8651) );
  XNOR U8796 ( .A(n8652), .B(n8653), .Z(n8055) );
  XOR U8797 ( .A(n8654), .B(n8655), .Z(n8617) );
  XNOR U8798 ( .A(n8057), .B(n8056), .Z(n8655) );
  XOR U8799 ( .A(n6390), .B(n7062), .Z(n8056) );
  XOR U8800 ( .A(n8656), .B(n8657), .Z(n8057) );
  XOR U8801 ( .A(n8659), .B(n8660), .Z(n8656) );
  XOR U8802 ( .A(n7052), .B(n8661), .Z(n8654) );
  XNOR U8803 ( .A(key[266]), .B(n7056), .Z(n8661) );
  XNOR U8804 ( .A(n8662), .B(n8663), .Z(n7052) );
  XNOR U8805 ( .A(n8664), .B(n8665), .Z(n8663) );
  XNOR U8806 ( .A(n8666), .B(n8667), .Z(n8662) );
  IV U8807 ( .A(n8471), .Z(n8643) );
  XOR U8808 ( .A(n8611), .B(n8668), .Z(n8471) );
  XOR U8809 ( .A(n8614), .B(n8623), .Z(n8668) );
  XNOR U8810 ( .A(n8669), .B(n8670), .Z(n8623) );
  XOR U8811 ( .A(n7026), .B(n8075), .Z(n8670) );
  XNOR U8812 ( .A(n7039), .B(n7025), .Z(n8075) );
  XOR U8813 ( .A(n8671), .B(n8672), .Z(n7039) );
  XOR U8814 ( .A(n8647), .B(n8673), .Z(n8672) );
  XOR U8815 ( .A(n8674), .B(n8633), .Z(n8671) );
  XNOR U8816 ( .A(n8676), .B(n8677), .Z(n8675) );
  NANDN U8817 ( .A(n8678), .B(n8679), .Z(n8677) );
  XOR U8818 ( .A(n8681), .B(n8682), .Z(n7026) );
  XOR U8819 ( .A(n8650), .B(n8683), .Z(n8682) );
  XOR U8820 ( .A(n8684), .B(n8641), .Z(n8681) );
  XNOR U8821 ( .A(n8686), .B(n8687), .Z(n8685) );
  NANDN U8822 ( .A(n8688), .B(n8689), .Z(n8687) );
  XNOR U8823 ( .A(key[271]), .B(n7046), .Z(n8669) );
  XNOR U8824 ( .A(n6437), .B(n6412), .Z(n7046) );
  XOR U8825 ( .A(n8611), .B(n8691), .Z(n8398) );
  XOR U8826 ( .A(n8614), .B(n8624), .Z(n8691) );
  XNOR U8827 ( .A(n8692), .B(n8693), .Z(n8624) );
  XOR U8828 ( .A(n8078), .B(n6416), .Z(n8693) );
  XNOR U8829 ( .A(n8634), .B(n7030), .Z(n6416) );
  XOR U8830 ( .A(n8694), .B(n8695), .Z(n8078) );
  XNOR U8831 ( .A(n7011), .B(n7034), .Z(n8695) );
  XNOR U8832 ( .A(n8696), .B(n8697), .Z(n7034) );
  XNOR U8833 ( .A(n8698), .B(n8699), .Z(n8697) );
  XNOR U8834 ( .A(n8642), .B(n8700), .Z(n8696) );
  XOR U8835 ( .A(n8701), .B(n8702), .Z(n8700) );
  ANDN U8836 ( .B(n8703), .A(n8704), .Z(n8702) );
  XOR U8837 ( .A(n8705), .B(n7062), .Z(n7011) );
  XOR U8838 ( .A(n8706), .B(n8664), .Z(n7062) );
  XOR U8839 ( .A(n8707), .B(n6419), .Z(n8694) );
  XOR U8840 ( .A(n8708), .B(n6390), .Z(n6419) );
  XNOR U8841 ( .A(n8674), .B(n8709), .Z(n6390) );
  IV U8842 ( .A(n8632), .Z(n8674) );
  XNOR U8843 ( .A(n8710), .B(n8711), .Z(n8632) );
  XNOR U8844 ( .A(n8712), .B(n8713), .Z(n8711) );
  NAND U8845 ( .A(n8714), .B(n8715), .Z(n8713) );
  XNOR U8846 ( .A(key[268]), .B(n7012), .Z(n8692) );
  XNOR U8847 ( .A(n8716), .B(n7056), .Z(n7012) );
  XOR U8848 ( .A(n8717), .B(n8640), .Z(n7056) );
  IV U8849 ( .A(n8684), .Z(n8640) );
  XOR U8850 ( .A(n8718), .B(n8719), .Z(n8684) );
  XNOR U8851 ( .A(n8720), .B(n8721), .Z(n8719) );
  NANDN U8852 ( .A(n8722), .B(n8723), .Z(n8721) );
  XOR U8853 ( .A(n8724), .B(n8725), .Z(n8614) );
  XOR U8854 ( .A(n8536), .B(n6397), .Z(n8725) );
  XNOR U8855 ( .A(n6412), .B(n7025), .Z(n6397) );
  XNOR U8856 ( .A(n8726), .B(n8727), .Z(n7025) );
  XOR U8857 ( .A(n8728), .B(n8729), .Z(n8727) );
  XNOR U8858 ( .A(n8666), .B(n8730), .Z(n8726) );
  XNOR U8859 ( .A(n8731), .B(n8732), .Z(n8536) );
  XNOR U8860 ( .A(n7055), .B(n6435), .Z(n8732) );
  XOR U8861 ( .A(n7048), .B(n7016), .Z(n6435) );
  IV U8862 ( .A(n8089), .Z(n7016) );
  XOR U8863 ( .A(n8733), .B(n8708), .Z(n8089) );
  XOR U8864 ( .A(n8716), .B(n8734), .Z(n7048) );
  XOR U8865 ( .A(n8664), .B(n8735), .Z(n7055) );
  XOR U8866 ( .A(n8666), .B(n8730), .Z(n8735) );
  XNOR U8867 ( .A(n8737), .B(n8738), .Z(n8736) );
  NANDN U8868 ( .A(n8739), .B(n8740), .Z(n8738) );
  IV U8869 ( .A(n8728), .Z(n8664) );
  XOR U8870 ( .A(n8742), .B(n8743), .Z(n8728) );
  XNOR U8871 ( .A(n8744), .B(n8745), .Z(n8743) );
  NANDN U8872 ( .A(n8746), .B(n8747), .Z(n8745) );
  XOR U8873 ( .A(n8090), .B(n8748), .Z(n8731) );
  XNOR U8874 ( .A(key[264]), .B(n8634), .Z(n8748) );
  IV U8875 ( .A(n6412), .Z(n8634) );
  XOR U8876 ( .A(n8705), .B(n8749), .Z(n6412) );
  IV U8877 ( .A(n8085), .Z(n8090) );
  XOR U8878 ( .A(n8653), .B(n8750), .Z(n8085) );
  XNOR U8879 ( .A(n8064), .B(n8752), .Z(n8724) );
  XNOR U8880 ( .A(key[270]), .B(n7032), .Z(n8752) );
  XOR U8881 ( .A(n8650), .B(n8639), .Z(n7032) );
  XNOR U8882 ( .A(n8690), .B(n8753), .Z(n8639) );
  XNOR U8883 ( .A(n8754), .B(n8755), .Z(n8753) );
  NOR U8884 ( .A(n8756), .B(n8757), .Z(n8754) );
  XNOR U8885 ( .A(n8758), .B(n8759), .Z(n8690) );
  XNOR U8886 ( .A(n8760), .B(n8761), .Z(n8759) );
  NAND U8887 ( .A(n8762), .B(n8763), .Z(n8761) );
  XOR U8888 ( .A(n8717), .B(n8638), .Z(n8650) );
  XOR U8889 ( .A(n8758), .B(n8764), .Z(n8638) );
  XNOR U8890 ( .A(n8686), .B(n8765), .Z(n8764) );
  NANDN U8891 ( .A(n8766), .B(n8767), .Z(n8765) );
  OR U8892 ( .A(n8768), .B(n8769), .Z(n8686) );
  IV U8893 ( .A(n8734), .Z(n8717) );
  XNOR U8894 ( .A(n8718), .B(n8770), .Z(n8734) );
  XOR U8895 ( .A(n8771), .B(n8772), .Z(n8770) );
  ANDN U8896 ( .B(n8773), .A(n8774), .Z(n8771) );
  XNOR U8897 ( .A(n8074), .B(n6404), .Z(n8064) );
  XOR U8898 ( .A(n7040), .B(n6398), .Z(n6404) );
  XNOR U8899 ( .A(n8647), .B(n8631), .Z(n6398) );
  XNOR U8900 ( .A(n8680), .B(n8775), .Z(n8631) );
  XNOR U8901 ( .A(n8776), .B(n8777), .Z(n8775) );
  NOR U8902 ( .A(n8778), .B(n8779), .Z(n8776) );
  XNOR U8903 ( .A(n8780), .B(n8781), .Z(n8680) );
  XNOR U8904 ( .A(n8782), .B(n8783), .Z(n8781) );
  NAND U8905 ( .A(n8784), .B(n8785), .Z(n8783) );
  XOR U8906 ( .A(n8733), .B(n8630), .Z(n8647) );
  XOR U8907 ( .A(n8780), .B(n8786), .Z(n8630) );
  XNOR U8908 ( .A(n8676), .B(n8787), .Z(n8786) );
  NANDN U8909 ( .A(n8788), .B(n8789), .Z(n8787) );
  OR U8910 ( .A(n8790), .B(n8791), .Z(n8676) );
  IV U8911 ( .A(n8709), .Z(n8733) );
  XNOR U8912 ( .A(n8710), .B(n8792), .Z(n8709) );
  XOR U8913 ( .A(n8793), .B(n8794), .Z(n8792) );
  NOR U8914 ( .A(n8795), .B(n8788), .Z(n8793) );
  XNOR U8915 ( .A(n8707), .B(n7027), .Z(n8074) );
  XNOR U8916 ( .A(n8796), .B(n8797), .Z(n7027) );
  XOR U8917 ( .A(n8653), .B(n8699), .Z(n8797) );
  XNOR U8918 ( .A(n8798), .B(n8799), .Z(n8699) );
  XNOR U8919 ( .A(n8800), .B(n8801), .Z(n8799) );
  NANDN U8920 ( .A(n8802), .B(n8803), .Z(n8801) );
  XOR U8921 ( .A(n8804), .B(n8805), .Z(n8653) );
  XNOR U8922 ( .A(n8806), .B(n8807), .Z(n8805) );
  NANDN U8923 ( .A(n8808), .B(n8703), .Z(n8807) );
  XOR U8924 ( .A(n8659), .B(n8751), .Z(n8796) );
  XNOR U8925 ( .A(n8810), .B(n8811), .Z(n8809) );
  NANDN U8926 ( .A(n8812), .B(n8803), .Z(n8811) );
  IV U8927 ( .A(n6437), .Z(n8707) );
  XOR U8928 ( .A(n8642), .B(n8652), .Z(n6437) );
  XNOR U8929 ( .A(n8798), .B(n8814), .Z(n8642) );
  XOR U8930 ( .A(n8815), .B(n8806), .Z(n8814) );
  NOR U8931 ( .A(n8818), .B(n8819), .Z(n8815) );
  XNOR U8932 ( .A(n8804), .B(n8820), .Z(n8798) );
  XNOR U8933 ( .A(n8821), .B(n8822), .Z(n8820) );
  NAND U8934 ( .A(n8823), .B(n8824), .Z(n8822) );
  IV U8935 ( .A(n8615), .Z(n8611) );
  XOR U8936 ( .A(n8825), .B(n8826), .Z(n8615) );
  XOR U8937 ( .A(n7033), .B(n8069), .Z(n8826) );
  XOR U8938 ( .A(n6405), .B(n7030), .Z(n8069) );
  XNOR U8939 ( .A(n8827), .B(n8828), .Z(n7030) );
  XNOR U8940 ( .A(n8829), .B(n8729), .Z(n8828) );
  XNOR U8941 ( .A(n8830), .B(n8831), .Z(n8729) );
  XNOR U8942 ( .A(n8832), .B(n8833), .Z(n8831) );
  NANDN U8943 ( .A(n8834), .B(n8740), .Z(n8833) );
  XNOR U8944 ( .A(n8705), .B(n8835), .Z(n8827) );
  XOR U8945 ( .A(n8836), .B(n8837), .Z(n8835) );
  ANDN U8946 ( .B(n8747), .A(n8838), .Z(n8837) );
  XNOR U8947 ( .A(n8830), .B(n8839), .Z(n8705) );
  XOR U8948 ( .A(n8840), .B(n8744), .Z(n8839) );
  NOR U8949 ( .A(n8843), .B(n8844), .Z(n8840) );
  XNOR U8950 ( .A(n8742), .B(n8845), .Z(n8830) );
  XNOR U8951 ( .A(n8846), .B(n8847), .Z(n8845) );
  NAND U8952 ( .A(n8848), .B(n8849), .Z(n8847) );
  XOR U8953 ( .A(n8850), .B(n8851), .Z(n6405) );
  XNOR U8954 ( .A(n8708), .B(n8673), .Z(n8851) );
  XNOR U8955 ( .A(n8852), .B(n8853), .Z(n8673) );
  XNOR U8956 ( .A(n8794), .B(n8854), .Z(n8853) );
  OR U8957 ( .A(n8678), .B(n8855), .Z(n8854) );
  OR U8958 ( .A(n8790), .B(n8856), .Z(n8794) );
  XNOR U8959 ( .A(n8678), .B(n8788), .Z(n8790) );
  XNOR U8960 ( .A(n8852), .B(n8857), .Z(n8708) );
  XOR U8961 ( .A(n8858), .B(n8712), .Z(n8857) );
  NOR U8962 ( .A(n8861), .B(n8779), .Z(n8858) );
  XNOR U8963 ( .A(n8710), .B(n8862), .Z(n8852) );
  XNOR U8964 ( .A(n8863), .B(n8864), .Z(n8862) );
  NAND U8965 ( .A(n8785), .B(n8865), .Z(n8864) );
  XOR U8966 ( .A(n8866), .B(n8863), .Z(n8710) );
  OR U8967 ( .A(n8867), .B(n8868), .Z(n8863) );
  ANDN U8968 ( .B(n8869), .A(n8870), .Z(n8866) );
  XNOR U8969 ( .A(n8780), .B(n8871), .Z(n8850) );
  XOR U8970 ( .A(n8777), .B(n8872), .Z(n8871) );
  ANDN U8971 ( .B(n8715), .A(n8873), .Z(n8872) );
  ANDN U8972 ( .B(n8860), .A(n8874), .Z(n8777) );
  XNOR U8973 ( .A(n8779), .B(n8715), .Z(n8860) );
  XOR U8974 ( .A(n8875), .B(n8782), .Z(n8780) );
  NANDN U8975 ( .A(n8867), .B(n8876), .Z(n8782) );
  XNOR U8976 ( .A(n8869), .B(n8785), .Z(n8867) );
  XNOR U8977 ( .A(n8788), .B(n8715), .Z(n8785) );
  XOR U8978 ( .A(n8877), .B(n8878), .Z(n8715) );
  NANDN U8979 ( .A(n8879), .B(n8880), .Z(n8878) );
  XNOR U8980 ( .A(n8881), .B(n8882), .Z(n8788) );
  OR U8981 ( .A(n8879), .B(n8883), .Z(n8882) );
  AND U8982 ( .A(n8869), .B(n8884), .Z(n8875) );
  XOR U8983 ( .A(n8678), .B(n8779), .Z(n8869) );
  XOR U8984 ( .A(n8885), .B(n8877), .Z(n8779) );
  NANDN U8985 ( .A(n8886), .B(n8887), .Z(n8877) );
  ANDN U8986 ( .B(n8888), .A(n8889), .Z(n8885) );
  NANDN U8987 ( .A(n8886), .B(n8891), .Z(n8881) );
  XOR U8988 ( .A(n8892), .B(n8879), .Z(n8886) );
  XNOR U8989 ( .A(n8893), .B(n8894), .Z(n8879) );
  XOR U8990 ( .A(n8895), .B(n8888), .Z(n8894) );
  XNOR U8991 ( .A(n8896), .B(n8897), .Z(n8893) );
  XNOR U8992 ( .A(n8898), .B(n8899), .Z(n8897) );
  ANDN U8993 ( .B(n8888), .A(n8900), .Z(n8898) );
  IV U8994 ( .A(n8901), .Z(n8888) );
  ANDN U8995 ( .B(n8892), .A(n8900), .Z(n8890) );
  IV U8996 ( .A(n8896), .Z(n8900) );
  IV U8997 ( .A(n8889), .Z(n8892) );
  XNOR U8998 ( .A(n8895), .B(n8902), .Z(n8889) );
  XOR U8999 ( .A(n8903), .B(n8899), .Z(n8902) );
  NAND U9000 ( .A(n8891), .B(n8887), .Z(n8899) );
  XNOR U9001 ( .A(n8880), .B(n8901), .Z(n8887) );
  XOR U9002 ( .A(n8904), .B(n8905), .Z(n8901) );
  XOR U9003 ( .A(n8906), .B(n8907), .Z(n8905) );
  XNOR U9004 ( .A(n8789), .B(n8908), .Z(n8907) );
  XNOR U9005 ( .A(n8909), .B(n8910), .Z(n8904) );
  XNOR U9006 ( .A(n8911), .B(n8912), .Z(n8910) );
  ANDN U9007 ( .B(n8679), .A(n8855), .Z(n8911) );
  XNOR U9008 ( .A(n8896), .B(n8883), .Z(n8891) );
  XOR U9009 ( .A(n8913), .B(n8914), .Z(n8896) );
  XNOR U9010 ( .A(n8915), .B(n8908), .Z(n8914) );
  XOR U9011 ( .A(n8916), .B(n8917), .Z(n8908) );
  XNOR U9012 ( .A(n8918), .B(n8919), .Z(n8917) );
  NAND U9013 ( .A(n8865), .B(n8784), .Z(n8919) );
  XNOR U9014 ( .A(n8920), .B(n8921), .Z(n8913) );
  ANDN U9015 ( .B(n8922), .A(n8861), .Z(n8920) );
  ANDN U9016 ( .B(n8880), .A(n8883), .Z(n8903) );
  XOR U9017 ( .A(n8883), .B(n8880), .Z(n8895) );
  XNOR U9018 ( .A(n8923), .B(n8924), .Z(n8880) );
  XNOR U9019 ( .A(n8916), .B(n8925), .Z(n8924) );
  XNOR U9020 ( .A(n8915), .B(n8679), .Z(n8925) );
  XNOR U9021 ( .A(n8926), .B(n8927), .Z(n8923) );
  XNOR U9022 ( .A(n8928), .B(n8912), .Z(n8927) );
  OR U9023 ( .A(n8791), .B(n8856), .Z(n8912) );
  XNOR U9024 ( .A(n8926), .B(n8909), .Z(n8856) );
  XNOR U9025 ( .A(n8679), .B(n8789), .Z(n8791) );
  ANDN U9026 ( .B(n8789), .A(n8795), .Z(n8928) );
  XOR U9027 ( .A(n8929), .B(n8930), .Z(n8883) );
  XOR U9028 ( .A(n8916), .B(n8906), .Z(n8930) );
  XOR U9029 ( .A(n8714), .B(n8873), .Z(n8906) );
  XOR U9030 ( .A(n8931), .B(n8918), .Z(n8916) );
  NANDN U9031 ( .A(n8868), .B(n8876), .Z(n8918) );
  XOR U9032 ( .A(n8884), .B(n8784), .Z(n8876) );
  XNOR U9033 ( .A(n8922), .B(n8932), .Z(n8789) );
  XNOR U9034 ( .A(n8933), .B(n8934), .Z(n8932) );
  XOR U9035 ( .A(n8870), .B(n8865), .Z(n8868) );
  XNOR U9036 ( .A(n8795), .B(n8714), .Z(n8865) );
  IV U9037 ( .A(n8909), .Z(n8795) );
  XOR U9038 ( .A(n8935), .B(n8936), .Z(n8909) );
  XOR U9039 ( .A(n8937), .B(n8938), .Z(n8936) );
  XOR U9040 ( .A(n8926), .B(n8939), .Z(n8935) );
  ANDN U9041 ( .B(n8884), .A(n8870), .Z(n8931) );
  XNOR U9042 ( .A(n8926), .B(n8940), .Z(n8870) );
  XOR U9043 ( .A(n8922), .B(n8679), .Z(n8884) );
  XNOR U9044 ( .A(n8941), .B(n8942), .Z(n8679) );
  XOR U9045 ( .A(n8943), .B(n8938), .Z(n8942) );
  XNOR U9046 ( .A(n8944), .B(n8945), .Z(n8938) );
  XNOR U9047 ( .A(n8946), .B(n8947), .Z(n8945) );
  XNOR U9048 ( .A(n8948), .B(n8949), .Z(n8944) );
  XNOR U9049 ( .A(key[156]), .B(n8950), .Z(n8949) );
  IV U9050 ( .A(n8778), .Z(n8922) );
  XOR U9051 ( .A(n8915), .B(n8951), .Z(n8929) );
  XNOR U9052 ( .A(n8952), .B(n8921), .Z(n8951) );
  OR U9053 ( .A(n8874), .B(n8859), .Z(n8921) );
  XNOR U9054 ( .A(n8940), .B(n8714), .Z(n8859) );
  XNOR U9055 ( .A(n8778), .B(n8873), .Z(n8874) );
  ANDN U9056 ( .B(n8714), .A(n8873), .Z(n8952) );
  XOR U9057 ( .A(n8941), .B(n8953), .Z(n8873) );
  XOR U9058 ( .A(n8933), .B(n8954), .Z(n8953) );
  XOR U9059 ( .A(n8943), .B(n8941), .Z(n8714) );
  XNOR U9060 ( .A(n8861), .B(n8778), .Z(n8915) );
  XOR U9061 ( .A(n8941), .B(n8955), .Z(n8778) );
  XNOR U9062 ( .A(n8943), .B(n8937), .Z(n8955) );
  XOR U9063 ( .A(n8956), .B(n8957), .Z(n8937) );
  XNOR U9064 ( .A(n8958), .B(n8959), .Z(n8957) );
  XNOR U9065 ( .A(key[159]), .B(n8960), .Z(n8956) );
  XNOR U9066 ( .A(n8961), .B(n8962), .Z(n8941) );
  XOR U9067 ( .A(n8963), .B(n8964), .Z(n8962) );
  XNOR U9068 ( .A(n8965), .B(n8966), .Z(n8961) );
  XNOR U9069 ( .A(key[157]), .B(n8967), .Z(n8966) );
  IV U9070 ( .A(n8940), .Z(n8861) );
  XNOR U9071 ( .A(n8934), .B(n8968), .Z(n8940) );
  XOR U9072 ( .A(n8939), .B(n8954), .Z(n8968) );
  IV U9073 ( .A(n8943), .Z(n8954) );
  XOR U9074 ( .A(n8969), .B(n8970), .Z(n8943) );
  XOR U9075 ( .A(n8971), .B(n8855), .Z(n8970) );
  IV U9076 ( .A(n8926), .Z(n8855) );
  XOR U9077 ( .A(n8972), .B(n8973), .Z(n8926) );
  XOR U9078 ( .A(n8974), .B(n8975), .Z(n8973) );
  XOR U9079 ( .A(n8976), .B(n8977), .Z(n8972) );
  XNOR U9080 ( .A(key[152]), .B(n8978), .Z(n8977) );
  XOR U9081 ( .A(n8979), .B(n8980), .Z(n8969) );
  XOR U9082 ( .A(key[158]), .B(n8981), .Z(n8980) );
  XOR U9083 ( .A(n8982), .B(n8983), .Z(n8939) );
  XNOR U9084 ( .A(n8933), .B(n8984), .Z(n8983) );
  XOR U9085 ( .A(n8985), .B(n8986), .Z(n8984) );
  XOR U9086 ( .A(n8987), .B(n8988), .Z(n8933) );
  XNOR U9087 ( .A(n8989), .B(n8990), .Z(n8988) );
  XOR U9088 ( .A(n8991), .B(n8992), .Z(n8987) );
  XOR U9089 ( .A(key[153]), .B(n8993), .Z(n8992) );
  XNOR U9090 ( .A(n8994), .B(n8995), .Z(n8982) );
  XNOR U9091 ( .A(key[155]), .B(n8996), .Z(n8995) );
  XOR U9092 ( .A(n8997), .B(n8998), .Z(n8934) );
  XOR U9093 ( .A(n8999), .B(n9000), .Z(n8998) );
  XNOR U9094 ( .A(n9001), .B(n9002), .Z(n8997) );
  XOR U9095 ( .A(key[154]), .B(n9003), .Z(n9002) );
  XNOR U9096 ( .A(n9004), .B(n9005), .Z(n7033) );
  XNOR U9097 ( .A(n8758), .B(n8683), .Z(n9005) );
  XNOR U9098 ( .A(n9006), .B(n9007), .Z(n8683) );
  XNOR U9099 ( .A(n8772), .B(n9008), .Z(n9007) );
  NANDN U9100 ( .A(n9009), .B(n8689), .Z(n9008) );
  OR U9101 ( .A(n9010), .B(n8768), .Z(n8772) );
  XNOR U9102 ( .A(n8689), .B(n8767), .Z(n8768) );
  XOR U9103 ( .A(n9011), .B(n8760), .Z(n8758) );
  NANDN U9104 ( .A(n9012), .B(n9013), .Z(n8760) );
  ANDN U9105 ( .B(n9014), .A(n9015), .Z(n9011) );
  XNOR U9106 ( .A(n8716), .B(n9016), .Z(n9004) );
  XOR U9107 ( .A(n8755), .B(n9017), .Z(n9016) );
  ANDN U9108 ( .B(n8723), .A(n9018), .Z(n9017) );
  ANDN U9109 ( .B(n9019), .A(n9020), .Z(n8755) );
  XNOR U9110 ( .A(n9006), .B(n9021), .Z(n8716) );
  XOR U9111 ( .A(n9022), .B(n8720), .Z(n9021) );
  XNOR U9112 ( .A(n8757), .B(n8723), .Z(n9019) );
  NOR U9113 ( .A(n9024), .B(n8757), .Z(n9022) );
  XNOR U9114 ( .A(n8718), .B(n9025), .Z(n9006) );
  XNOR U9115 ( .A(n9026), .B(n9027), .Z(n9025) );
  NAND U9116 ( .A(n8763), .B(n9028), .Z(n9027) );
  XOR U9117 ( .A(n9029), .B(n9026), .Z(n8718) );
  OR U9118 ( .A(n9012), .B(n9030), .Z(n9026) );
  XNOR U9119 ( .A(n9031), .B(n8763), .Z(n9012) );
  XOR U9120 ( .A(n8767), .B(n8723), .Z(n8763) );
  XOR U9121 ( .A(n9032), .B(n9033), .Z(n8723) );
  NANDN U9122 ( .A(n9034), .B(n9035), .Z(n9033) );
  IV U9123 ( .A(n8774), .Z(n8767) );
  XNOR U9124 ( .A(n9036), .B(n9037), .Z(n8774) );
  NANDN U9125 ( .A(n9034), .B(n9038), .Z(n9037) );
  ANDN U9126 ( .B(n9031), .A(n9039), .Z(n9029) );
  IV U9127 ( .A(n9015), .Z(n9031) );
  XOR U9128 ( .A(n8757), .B(n8689), .Z(n9015) );
  XNOR U9129 ( .A(n9040), .B(n9036), .Z(n8689) );
  NANDN U9130 ( .A(n9041), .B(n9042), .Z(n9036) );
  XOR U9131 ( .A(n9038), .B(n9043), .Z(n9042) );
  ANDN U9132 ( .B(n9043), .A(n9044), .Z(n9040) );
  XOR U9133 ( .A(n9045), .B(n9032), .Z(n8757) );
  NANDN U9134 ( .A(n9041), .B(n9046), .Z(n9032) );
  XOR U9135 ( .A(n9047), .B(n9035), .Z(n9046) );
  XNOR U9136 ( .A(n9048), .B(n9049), .Z(n9034) );
  XOR U9137 ( .A(n9050), .B(n9051), .Z(n9049) );
  XNOR U9138 ( .A(n9052), .B(n9053), .Z(n9048) );
  XNOR U9139 ( .A(n9054), .B(n9055), .Z(n9053) );
  ANDN U9140 ( .B(n9047), .A(n9051), .Z(n9054) );
  ANDN U9141 ( .B(n9047), .A(n9044), .Z(n9045) );
  XNOR U9142 ( .A(n9050), .B(n9056), .Z(n9044) );
  XOR U9143 ( .A(n9057), .B(n9055), .Z(n9056) );
  NAND U9144 ( .A(n9058), .B(n9059), .Z(n9055) );
  XNOR U9145 ( .A(n9052), .B(n9035), .Z(n9059) );
  IV U9146 ( .A(n9047), .Z(n9052) );
  XNOR U9147 ( .A(n9038), .B(n9051), .Z(n9058) );
  IV U9148 ( .A(n9043), .Z(n9051) );
  XOR U9149 ( .A(n9060), .B(n9061), .Z(n9043) );
  XNOR U9150 ( .A(n9062), .B(n9063), .Z(n9061) );
  XNOR U9151 ( .A(n9064), .B(n9065), .Z(n9060) );
  NOR U9152 ( .A(n8756), .B(n9024), .Z(n9064) );
  AND U9153 ( .A(n9035), .B(n9038), .Z(n9057) );
  XNOR U9154 ( .A(n9035), .B(n9038), .Z(n9050) );
  XNOR U9155 ( .A(n9066), .B(n9067), .Z(n9038) );
  XNOR U9156 ( .A(n9068), .B(n9063), .Z(n9067) );
  XOR U9157 ( .A(n9069), .B(n9070), .Z(n9066) );
  XNOR U9158 ( .A(n9071), .B(n9065), .Z(n9070) );
  OR U9159 ( .A(n9020), .B(n9023), .Z(n9065) );
  XNOR U9160 ( .A(n9024), .B(n8722), .Z(n9023) );
  XNOR U9161 ( .A(n8756), .B(n9018), .Z(n9020) );
  ANDN U9162 ( .B(n9072), .A(n8722), .Z(n9071) );
  XNOR U9163 ( .A(n9073), .B(n9074), .Z(n9035) );
  XNOR U9164 ( .A(n9063), .B(n9075), .Z(n9074) );
  XOR U9165 ( .A(n8688), .B(n9069), .Z(n9075) );
  XNOR U9166 ( .A(n9024), .B(n9076), .Z(n9063) );
  XNOR U9167 ( .A(n9077), .B(n9078), .Z(n9073) );
  XNOR U9168 ( .A(n9079), .B(n9080), .Z(n9078) );
  ANDN U9169 ( .B(n8773), .A(n8766), .Z(n9079) );
  XNOR U9170 ( .A(n9081), .B(n9082), .Z(n9047) );
  XNOR U9171 ( .A(n9068), .B(n9083), .Z(n9082) );
  XNOR U9172 ( .A(n8766), .B(n9062), .Z(n9083) );
  XOR U9173 ( .A(n9069), .B(n9084), .Z(n9062) );
  XNOR U9174 ( .A(n9085), .B(n9086), .Z(n9084) );
  NAND U9175 ( .A(n9028), .B(n8762), .Z(n9086) );
  XNOR U9176 ( .A(n9087), .B(n9085), .Z(n9069) );
  NANDN U9177 ( .A(n9030), .B(n9013), .Z(n9085) );
  XOR U9178 ( .A(n9014), .B(n8762), .Z(n9013) );
  XNOR U9179 ( .A(n9088), .B(n9018), .Z(n8762) );
  XOR U9180 ( .A(n9039), .B(n9028), .Z(n9030) );
  XOR U9181 ( .A(n8773), .B(n9089), .Z(n9028) );
  ANDN U9182 ( .B(n9014), .A(n9039), .Z(n9087) );
  XOR U9183 ( .A(n9077), .B(n9024), .Z(n9039) );
  XOR U9184 ( .A(n9090), .B(n9091), .Z(n9024) );
  XNOR U9185 ( .A(n9092), .B(n9093), .Z(n9091) );
  XOR U9186 ( .A(n9094), .B(n9076), .Z(n9014) );
  XOR U9187 ( .A(n9089), .B(n9072), .Z(n9068) );
  IV U9188 ( .A(n9018), .Z(n9072) );
  XOR U9189 ( .A(n9095), .B(n9096), .Z(n9018) );
  XNOR U9190 ( .A(n9097), .B(n9093), .Z(n9096) );
  IV U9191 ( .A(n8722), .Z(n9089) );
  XOR U9192 ( .A(n9093), .B(n9098), .Z(n8722) );
  XNOR U9193 ( .A(n8773), .B(n9099), .Z(n9081) );
  XNOR U9194 ( .A(n9100), .B(n9080), .Z(n9099) );
  OR U9195 ( .A(n8769), .B(n9010), .Z(n9080) );
  XNOR U9196 ( .A(n9077), .B(n8773), .Z(n9010) );
  XOR U9197 ( .A(n8688), .B(n9088), .Z(n8769) );
  IV U9198 ( .A(n8766), .Z(n9088) );
  XOR U9199 ( .A(n9076), .B(n9101), .Z(n8766) );
  XNOR U9200 ( .A(n9097), .B(n9090), .Z(n9101) );
  XOR U9201 ( .A(n9102), .B(n9103), .Z(n9090) );
  XOR U9202 ( .A(n9104), .B(n9105), .Z(n9103) );
  XOR U9203 ( .A(key[242]), .B(n9106), .Z(n9102) );
  IV U9204 ( .A(n8756), .Z(n9076) );
  XOR U9205 ( .A(n9095), .B(n9107), .Z(n8756) );
  XOR U9206 ( .A(n9093), .B(n9108), .Z(n9107) );
  ANDN U9207 ( .B(n9094), .A(n9009), .Z(n9100) );
  IV U9208 ( .A(n8688), .Z(n9094) );
  XOR U9209 ( .A(n9095), .B(n9109), .Z(n8688) );
  XOR U9210 ( .A(n9093), .B(n9110), .Z(n9109) );
  XOR U9211 ( .A(n9111), .B(n9112), .Z(n9093) );
  XOR U9212 ( .A(n9113), .B(n9009), .Z(n9112) );
  IV U9213 ( .A(n9077), .Z(n9009) );
  XOR U9214 ( .A(n9114), .B(n9115), .Z(n9111) );
  XNOR U9215 ( .A(key[246]), .B(n9116), .Z(n9115) );
  IV U9216 ( .A(n9098), .Z(n9095) );
  XOR U9217 ( .A(n9117), .B(n9118), .Z(n9098) );
  XOR U9218 ( .A(n9119), .B(n9120), .Z(n9118) );
  XNOR U9219 ( .A(key[245]), .B(n9121), .Z(n9117) );
  XOR U9220 ( .A(n9122), .B(n9123), .Z(n8773) );
  XNOR U9221 ( .A(n9110), .B(n9108), .Z(n9123) );
  XNOR U9222 ( .A(n9124), .B(n9125), .Z(n9108) );
  XNOR U9223 ( .A(n9126), .B(n9127), .Z(n9125) );
  XNOR U9224 ( .A(key[247]), .B(n9128), .Z(n9124) );
  XNOR U9225 ( .A(n9129), .B(n9130), .Z(n9110) );
  XNOR U9226 ( .A(n9131), .B(n9132), .Z(n9129) );
  XNOR U9227 ( .A(key[244]), .B(n9133), .Z(n9132) );
  XOR U9228 ( .A(n9077), .B(n9092), .Z(n9122) );
  XOR U9229 ( .A(n9134), .B(n9135), .Z(n9092) );
  XNOR U9230 ( .A(n9097), .B(n9136), .Z(n9135) );
  XOR U9231 ( .A(n9137), .B(n9138), .Z(n9136) );
  XOR U9232 ( .A(n9139), .B(n9140), .Z(n9097) );
  XOR U9233 ( .A(n9141), .B(n9142), .Z(n9140) );
  XNOR U9234 ( .A(key[241]), .B(n9143), .Z(n9139) );
  XNOR U9235 ( .A(n9144), .B(n9145), .Z(n9134) );
  XNOR U9236 ( .A(key[243]), .B(n9146), .Z(n9145) );
  XOR U9237 ( .A(n9147), .B(n9148), .Z(n9077) );
  XNOR U9238 ( .A(n9149), .B(n9150), .Z(n9148) );
  XNOR U9239 ( .A(key[240]), .B(n9151), .Z(n9147) );
  XNOR U9240 ( .A(n8065), .B(n9152), .Z(n8825) );
  XOR U9241 ( .A(key[269]), .B(n7040), .Z(n9152) );
  XOR U9242 ( .A(n8730), .B(n8665), .Z(n7040) );
  XNOR U9243 ( .A(n8741), .B(n9153), .Z(n8665) );
  XNOR U9244 ( .A(n9154), .B(n8836), .Z(n9153) );
  ANDN U9245 ( .B(n8842), .A(n9155), .Z(n8836) );
  XNOR U9246 ( .A(n8844), .B(n8747), .Z(n8842) );
  NOR U9247 ( .A(n9156), .B(n8844), .Z(n9154) );
  XNOR U9248 ( .A(n8829), .B(n9157), .Z(n8741) );
  XNOR U9249 ( .A(n9158), .B(n9159), .Z(n9157) );
  NAND U9250 ( .A(n9160), .B(n8848), .Z(n9159) );
  XOR U9251 ( .A(n8706), .B(n8667), .Z(n8730) );
  XNOR U9252 ( .A(n8829), .B(n9161), .Z(n8667) );
  XNOR U9253 ( .A(n8737), .B(n9162), .Z(n9161) );
  NANDN U9254 ( .A(n9163), .B(n9164), .Z(n9162) );
  OR U9255 ( .A(n9165), .B(n9166), .Z(n8737) );
  XOR U9256 ( .A(n9167), .B(n9158), .Z(n8829) );
  NANDN U9257 ( .A(n9168), .B(n9169), .Z(n9158) );
  ANDN U9258 ( .B(n9170), .A(n9171), .Z(n9167) );
  IV U9259 ( .A(n8749), .Z(n8706) );
  XNOR U9260 ( .A(n8742), .B(n9172), .Z(n8749) );
  XOR U9261 ( .A(n9173), .B(n8832), .Z(n9172) );
  OR U9262 ( .A(n9174), .B(n9165), .Z(n8832) );
  XNOR U9263 ( .A(n8740), .B(n9164), .Z(n9165) );
  ANDN U9264 ( .B(n9175), .A(n9176), .Z(n9173) );
  XOR U9265 ( .A(n9177), .B(n8846), .Z(n8742) );
  OR U9266 ( .A(n9168), .B(n9178), .Z(n8846) );
  XNOR U9267 ( .A(n9179), .B(n8848), .Z(n9168) );
  XOR U9268 ( .A(n9164), .B(n8747), .Z(n8848) );
  XOR U9269 ( .A(n9180), .B(n9181), .Z(n8747) );
  NANDN U9270 ( .A(n9182), .B(n9183), .Z(n9181) );
  IV U9271 ( .A(n9176), .Z(n9164) );
  XNOR U9272 ( .A(n9184), .B(n9185), .Z(n9176) );
  NANDN U9273 ( .A(n9182), .B(n9186), .Z(n9185) );
  ANDN U9274 ( .B(n9179), .A(n9187), .Z(n9177) );
  IV U9275 ( .A(n9171), .Z(n9179) );
  XOR U9276 ( .A(n8844), .B(n8740), .Z(n9171) );
  XNOR U9277 ( .A(n9188), .B(n9184), .Z(n8740) );
  NANDN U9278 ( .A(n9189), .B(n9190), .Z(n9184) );
  XOR U9279 ( .A(n9186), .B(n9191), .Z(n9190) );
  ANDN U9280 ( .B(n9191), .A(n9192), .Z(n9188) );
  XOR U9281 ( .A(n9193), .B(n9180), .Z(n8844) );
  NANDN U9282 ( .A(n9189), .B(n9194), .Z(n9180) );
  XOR U9283 ( .A(n9195), .B(n9183), .Z(n9194) );
  XNOR U9284 ( .A(n9196), .B(n9197), .Z(n9182) );
  XOR U9285 ( .A(n9198), .B(n9199), .Z(n9197) );
  XNOR U9286 ( .A(n9200), .B(n9201), .Z(n9196) );
  XNOR U9287 ( .A(n9202), .B(n9203), .Z(n9201) );
  ANDN U9288 ( .B(n9195), .A(n9199), .Z(n9202) );
  ANDN U9289 ( .B(n9195), .A(n9192), .Z(n9193) );
  XNOR U9290 ( .A(n9198), .B(n9204), .Z(n9192) );
  XOR U9291 ( .A(n9205), .B(n9203), .Z(n9204) );
  NAND U9292 ( .A(n9206), .B(n9207), .Z(n9203) );
  XNOR U9293 ( .A(n9200), .B(n9183), .Z(n9207) );
  IV U9294 ( .A(n9195), .Z(n9200) );
  XNOR U9295 ( .A(n9186), .B(n9199), .Z(n9206) );
  IV U9296 ( .A(n9191), .Z(n9199) );
  XOR U9297 ( .A(n9208), .B(n9209), .Z(n9191) );
  XNOR U9298 ( .A(n9210), .B(n9211), .Z(n9209) );
  XNOR U9299 ( .A(n9212), .B(n9213), .Z(n9208) );
  NOR U9300 ( .A(n9156), .B(n8843), .Z(n9212) );
  AND U9301 ( .A(n9183), .B(n9186), .Z(n9205) );
  XNOR U9302 ( .A(n9183), .B(n9186), .Z(n9198) );
  XNOR U9303 ( .A(n9214), .B(n9215), .Z(n9186) );
  XNOR U9304 ( .A(n9216), .B(n9211), .Z(n9215) );
  XOR U9305 ( .A(n9217), .B(n9218), .Z(n9214) );
  XNOR U9306 ( .A(n9219), .B(n9213), .Z(n9218) );
  OR U9307 ( .A(n9155), .B(n8841), .Z(n9213) );
  XNOR U9308 ( .A(n8843), .B(n8746), .Z(n8841) );
  XNOR U9309 ( .A(n9156), .B(n8838), .Z(n9155) );
  ANDN U9310 ( .B(n9220), .A(n8746), .Z(n9219) );
  XNOR U9311 ( .A(n9221), .B(n9222), .Z(n9183) );
  XNOR U9312 ( .A(n9211), .B(n9223), .Z(n9222) );
  XOR U9313 ( .A(n8739), .B(n9217), .Z(n9223) );
  XNOR U9314 ( .A(n8843), .B(n9224), .Z(n9211) );
  XNOR U9315 ( .A(n9225), .B(n9226), .Z(n9221) );
  XNOR U9316 ( .A(n9227), .B(n9228), .Z(n9226) );
  ANDN U9317 ( .B(n9175), .A(n9163), .Z(n9227) );
  XNOR U9318 ( .A(n9229), .B(n9230), .Z(n9195) );
  XNOR U9319 ( .A(n9216), .B(n9231), .Z(n9230) );
  XNOR U9320 ( .A(n9163), .B(n9210), .Z(n9231) );
  XOR U9321 ( .A(n9217), .B(n9232), .Z(n9210) );
  XNOR U9322 ( .A(n9233), .B(n9234), .Z(n9232) );
  NAND U9323 ( .A(n8849), .B(n9160), .Z(n9234) );
  XNOR U9324 ( .A(n9235), .B(n9233), .Z(n9217) );
  NANDN U9325 ( .A(n9178), .B(n9169), .Z(n9233) );
  XOR U9326 ( .A(n9170), .B(n9160), .Z(n9169) );
  XNOR U9327 ( .A(n9236), .B(n8838), .Z(n9160) );
  XOR U9328 ( .A(n9187), .B(n8849), .Z(n9178) );
  XOR U9329 ( .A(n9175), .B(n9237), .Z(n8849) );
  ANDN U9330 ( .B(n9170), .A(n9187), .Z(n9235) );
  XOR U9331 ( .A(n9225), .B(n8843), .Z(n9187) );
  XOR U9332 ( .A(n9238), .B(n9239), .Z(n8843) );
  XNOR U9333 ( .A(n9240), .B(n9241), .Z(n9239) );
  XOR U9334 ( .A(n9242), .B(n9224), .Z(n9170) );
  XOR U9335 ( .A(n9237), .B(n9220), .Z(n9216) );
  IV U9336 ( .A(n8838), .Z(n9220) );
  XOR U9337 ( .A(n9243), .B(n9244), .Z(n8838) );
  XNOR U9338 ( .A(n9245), .B(n9241), .Z(n9244) );
  IV U9339 ( .A(n8746), .Z(n9237) );
  XOR U9340 ( .A(n9241), .B(n9246), .Z(n8746) );
  XNOR U9341 ( .A(n9175), .B(n9247), .Z(n9229) );
  XNOR U9342 ( .A(n9248), .B(n9228), .Z(n9247) );
  OR U9343 ( .A(n9166), .B(n9174), .Z(n9228) );
  XNOR U9344 ( .A(n9225), .B(n9175), .Z(n9174) );
  XOR U9345 ( .A(n8739), .B(n9236), .Z(n9166) );
  IV U9346 ( .A(n9163), .Z(n9236) );
  XOR U9347 ( .A(n9224), .B(n9249), .Z(n9163) );
  XNOR U9348 ( .A(n9245), .B(n9238), .Z(n9249) );
  XOR U9349 ( .A(n9250), .B(n9251), .Z(n9238) );
  XOR U9350 ( .A(n9252), .B(n9253), .Z(n9251) );
  XOR U9351 ( .A(key[162]), .B(n9254), .Z(n9250) );
  IV U9352 ( .A(n9156), .Z(n9224) );
  XOR U9353 ( .A(n9243), .B(n9255), .Z(n9156) );
  XOR U9354 ( .A(n9241), .B(n9256), .Z(n9255) );
  ANDN U9355 ( .B(n9242), .A(n8834), .Z(n9248) );
  IV U9356 ( .A(n8739), .Z(n9242) );
  XOR U9357 ( .A(n9243), .B(n9257), .Z(n8739) );
  XOR U9358 ( .A(n9241), .B(n9258), .Z(n9257) );
  XOR U9359 ( .A(n9259), .B(n9260), .Z(n9241) );
  XOR U9360 ( .A(n9261), .B(n8834), .Z(n9260) );
  IV U9361 ( .A(n9225), .Z(n8834) );
  XNOR U9362 ( .A(n9262), .B(n9263), .Z(n9259) );
  XNOR U9363 ( .A(key[166]), .B(n9264), .Z(n9263) );
  IV U9364 ( .A(n9246), .Z(n9243) );
  XOR U9365 ( .A(n9265), .B(n9266), .Z(n9246) );
  XOR U9366 ( .A(n9267), .B(n9268), .Z(n9266) );
  XNOR U9367 ( .A(key[165]), .B(n9269), .Z(n9265) );
  XOR U9368 ( .A(n9270), .B(n9271), .Z(n9175) );
  XNOR U9369 ( .A(n9258), .B(n9256), .Z(n9271) );
  XNOR U9370 ( .A(n9272), .B(n9273), .Z(n9256) );
  XNOR U9371 ( .A(n9274), .B(n9275), .Z(n9273) );
  XOR U9372 ( .A(key[167]), .B(n9276), .Z(n9272) );
  XNOR U9373 ( .A(n9277), .B(n9278), .Z(n9258) );
  XNOR U9374 ( .A(n9279), .B(n9280), .Z(n9277) );
  XNOR U9375 ( .A(key[164]), .B(n9281), .Z(n9280) );
  XOR U9376 ( .A(n9225), .B(n9240), .Z(n9270) );
  XOR U9377 ( .A(n9282), .B(n9283), .Z(n9240) );
  XNOR U9378 ( .A(n9245), .B(n9284), .Z(n9283) );
  XNOR U9379 ( .A(n9285), .B(n9286), .Z(n9284) );
  XOR U9380 ( .A(n9287), .B(n9288), .Z(n9245) );
  XNOR U9381 ( .A(key[161]), .B(n9291), .Z(n9287) );
  XNOR U9382 ( .A(n9292), .B(n9293), .Z(n9282) );
  XNOR U9383 ( .A(key[163]), .B(n9294), .Z(n9293) );
  XOR U9384 ( .A(n9295), .B(n9296), .Z(n9225) );
  XOR U9385 ( .A(n9297), .B(n9298), .Z(n9296) );
  XNOR U9386 ( .A(key[160]), .B(n9299), .Z(n9295) );
  XOR U9387 ( .A(n8751), .B(n8658), .Z(n8065) );
  XNOR U9388 ( .A(n8813), .B(n9300), .Z(n8658) );
  XNOR U9389 ( .A(n9301), .B(n8701), .Z(n9300) );
  ANDN U9390 ( .B(n8817), .A(n9302), .Z(n8701) );
  XNOR U9391 ( .A(n8819), .B(n8703), .Z(n8817) );
  NOR U9392 ( .A(n9303), .B(n8819), .Z(n9301) );
  XNOR U9393 ( .A(n8698), .B(n9304), .Z(n8813) );
  XNOR U9394 ( .A(n9305), .B(n9306), .Z(n9304) );
  NAND U9395 ( .A(n9307), .B(n8823), .Z(n9306) );
  XOR U9396 ( .A(n8698), .B(n9308), .Z(n8660) );
  XNOR U9397 ( .A(n8810), .B(n9309), .Z(n9308) );
  NANDN U9398 ( .A(n9310), .B(n9311), .Z(n9309) );
  OR U9399 ( .A(n9312), .B(n9313), .Z(n8810) );
  XOR U9400 ( .A(n9314), .B(n9305), .Z(n8698) );
  NANDN U9401 ( .A(n9315), .B(n9316), .Z(n9305) );
  ANDN U9402 ( .B(n9317), .A(n9318), .Z(n9314) );
  XNOR U9403 ( .A(n8804), .B(n9319), .Z(n8652) );
  XOR U9404 ( .A(n9320), .B(n8800), .Z(n9319) );
  OR U9405 ( .A(n9321), .B(n9312), .Z(n8800) );
  XNOR U9406 ( .A(n8803), .B(n9311), .Z(n9312) );
  ANDN U9407 ( .B(n9322), .A(n9323), .Z(n9320) );
  XOR U9408 ( .A(n9324), .B(n8821), .Z(n8804) );
  OR U9409 ( .A(n9315), .B(n9325), .Z(n8821) );
  XNOR U9410 ( .A(n9326), .B(n8823), .Z(n9315) );
  XOR U9411 ( .A(n9311), .B(n8703), .Z(n8823) );
  XOR U9412 ( .A(n9327), .B(n9328), .Z(n8703) );
  NANDN U9413 ( .A(n9329), .B(n9330), .Z(n9328) );
  IV U9414 ( .A(n9323), .Z(n9311) );
  XNOR U9415 ( .A(n9331), .B(n9332), .Z(n9323) );
  NANDN U9416 ( .A(n9329), .B(n9333), .Z(n9332) );
  ANDN U9417 ( .B(n9326), .A(n9334), .Z(n9324) );
  IV U9418 ( .A(n9318), .Z(n9326) );
  XOR U9419 ( .A(n8819), .B(n8803), .Z(n9318) );
  XNOR U9420 ( .A(n9335), .B(n9331), .Z(n8803) );
  NANDN U9421 ( .A(n9336), .B(n9337), .Z(n9331) );
  XOR U9422 ( .A(n9333), .B(n9338), .Z(n9337) );
  ANDN U9423 ( .B(n9338), .A(n9339), .Z(n9335) );
  XOR U9424 ( .A(n9340), .B(n9327), .Z(n8819) );
  NANDN U9425 ( .A(n9336), .B(n9341), .Z(n9327) );
  XOR U9426 ( .A(n9342), .B(n9330), .Z(n9341) );
  XNOR U9427 ( .A(n9343), .B(n9344), .Z(n9329) );
  XOR U9428 ( .A(n9345), .B(n9346), .Z(n9344) );
  XNOR U9429 ( .A(n9347), .B(n9348), .Z(n9343) );
  XNOR U9430 ( .A(n9349), .B(n9350), .Z(n9348) );
  ANDN U9431 ( .B(n9342), .A(n9346), .Z(n9349) );
  ANDN U9432 ( .B(n9342), .A(n9339), .Z(n9340) );
  XNOR U9433 ( .A(n9345), .B(n9351), .Z(n9339) );
  XOR U9434 ( .A(n9352), .B(n9350), .Z(n9351) );
  NAND U9435 ( .A(n9353), .B(n9354), .Z(n9350) );
  XNOR U9436 ( .A(n9347), .B(n9330), .Z(n9354) );
  IV U9437 ( .A(n9342), .Z(n9347) );
  XNOR U9438 ( .A(n9333), .B(n9346), .Z(n9353) );
  IV U9439 ( .A(n9338), .Z(n9346) );
  XOR U9440 ( .A(n9355), .B(n9356), .Z(n9338) );
  XNOR U9441 ( .A(n9357), .B(n9358), .Z(n9356) );
  XNOR U9442 ( .A(n9359), .B(n9360), .Z(n9355) );
  NOR U9443 ( .A(n9303), .B(n8818), .Z(n9359) );
  AND U9444 ( .A(n9330), .B(n9333), .Z(n9352) );
  XNOR U9445 ( .A(n9330), .B(n9333), .Z(n9345) );
  XNOR U9446 ( .A(n9361), .B(n9362), .Z(n9333) );
  XNOR U9447 ( .A(n9363), .B(n9358), .Z(n9362) );
  XOR U9448 ( .A(n9364), .B(n9365), .Z(n9361) );
  XNOR U9449 ( .A(n9366), .B(n9360), .Z(n9365) );
  OR U9450 ( .A(n9302), .B(n8816), .Z(n9360) );
  XNOR U9451 ( .A(n8818), .B(n8808), .Z(n8816) );
  XNOR U9452 ( .A(n9303), .B(n8704), .Z(n9302) );
  ANDN U9453 ( .B(n9367), .A(n8808), .Z(n9366) );
  XNOR U9454 ( .A(n9368), .B(n9369), .Z(n9330) );
  XNOR U9455 ( .A(n9358), .B(n9370), .Z(n9369) );
  XOR U9456 ( .A(n8812), .B(n9364), .Z(n9370) );
  XNOR U9457 ( .A(n8818), .B(n9371), .Z(n9358) );
  XNOR U9458 ( .A(n9372), .B(n9373), .Z(n9368) );
  XNOR U9459 ( .A(n9374), .B(n9375), .Z(n9373) );
  ANDN U9460 ( .B(n9322), .A(n9310), .Z(n9374) );
  XNOR U9461 ( .A(n9376), .B(n9377), .Z(n9342) );
  XNOR U9462 ( .A(n9363), .B(n9378), .Z(n9377) );
  XNOR U9463 ( .A(n9310), .B(n9357), .Z(n9378) );
  XOR U9464 ( .A(n9364), .B(n9379), .Z(n9357) );
  XNOR U9465 ( .A(n9380), .B(n9381), .Z(n9379) );
  NAND U9466 ( .A(n8824), .B(n9307), .Z(n9381) );
  XNOR U9467 ( .A(n9382), .B(n9380), .Z(n9364) );
  NANDN U9468 ( .A(n9325), .B(n9316), .Z(n9380) );
  XOR U9469 ( .A(n9317), .B(n9307), .Z(n9316) );
  XNOR U9470 ( .A(n9383), .B(n8704), .Z(n9307) );
  XOR U9471 ( .A(n9334), .B(n8824), .Z(n9325) );
  XOR U9472 ( .A(n9322), .B(n9384), .Z(n8824) );
  ANDN U9473 ( .B(n9317), .A(n9334), .Z(n9382) );
  XOR U9474 ( .A(n9372), .B(n8818), .Z(n9334) );
  XOR U9475 ( .A(n9385), .B(n9386), .Z(n8818) );
  XNOR U9476 ( .A(n9387), .B(n9388), .Z(n9386) );
  XOR U9477 ( .A(n9389), .B(n9371), .Z(n9317) );
  XOR U9478 ( .A(n9384), .B(n9367), .Z(n9363) );
  IV U9479 ( .A(n8704), .Z(n9367) );
  XOR U9480 ( .A(n9390), .B(n9391), .Z(n8704) );
  XNOR U9481 ( .A(n9392), .B(n9388), .Z(n9391) );
  IV U9482 ( .A(n8808), .Z(n9384) );
  XOR U9483 ( .A(n9388), .B(n9393), .Z(n8808) );
  XNOR U9484 ( .A(n9322), .B(n9394), .Z(n9376) );
  XNOR U9485 ( .A(n9395), .B(n9375), .Z(n9394) );
  OR U9486 ( .A(n9313), .B(n9321), .Z(n9375) );
  XNOR U9487 ( .A(n9372), .B(n9322), .Z(n9321) );
  XOR U9488 ( .A(n8812), .B(n9383), .Z(n9313) );
  IV U9489 ( .A(n9310), .Z(n9383) );
  XOR U9490 ( .A(n9371), .B(n9396), .Z(n9310) );
  XNOR U9491 ( .A(n9392), .B(n9385), .Z(n9396) );
  XOR U9492 ( .A(n9397), .B(n9398), .Z(n9385) );
  XNOR U9493 ( .A(n9399), .B(n9400), .Z(n9398) );
  XOR U9494 ( .A(n9401), .B(n9402), .Z(n9397) );
  XNOR U9495 ( .A(key[202]), .B(n9403), .Z(n9402) );
  IV U9496 ( .A(n9303), .Z(n9371) );
  XOR U9497 ( .A(n9390), .B(n9404), .Z(n9303) );
  XOR U9498 ( .A(n9388), .B(n9405), .Z(n9404) );
  ANDN U9499 ( .B(n9389), .A(n8802), .Z(n9395) );
  IV U9500 ( .A(n8812), .Z(n9389) );
  XOR U9501 ( .A(n9390), .B(n9406), .Z(n8812) );
  XOR U9502 ( .A(n9388), .B(n9407), .Z(n9406) );
  XOR U9503 ( .A(n9408), .B(n9409), .Z(n9388) );
  XOR U9504 ( .A(n9410), .B(n8802), .Z(n9409) );
  IV U9505 ( .A(n9372), .Z(n8802) );
  XOR U9506 ( .A(n9411), .B(n9412), .Z(n9408) );
  XNOR U9507 ( .A(key[206]), .B(n9413), .Z(n9412) );
  IV U9508 ( .A(n9393), .Z(n9390) );
  XOR U9509 ( .A(n9414), .B(n9415), .Z(n9393) );
  XOR U9510 ( .A(n9416), .B(n9417), .Z(n9415) );
  XNOR U9511 ( .A(n9418), .B(n9419), .Z(n9414) );
  XNOR U9512 ( .A(key[205]), .B(n9420), .Z(n9419) );
  XOR U9513 ( .A(n9421), .B(n9422), .Z(n9322) );
  XNOR U9514 ( .A(n9407), .B(n9405), .Z(n9422) );
  XNOR U9515 ( .A(n9423), .B(n9424), .Z(n9405) );
  XOR U9516 ( .A(n9425), .B(n9426), .Z(n9424) );
  XOR U9517 ( .A(key[207]), .B(n9427), .Z(n9423) );
  XNOR U9518 ( .A(n9428), .B(n9429), .Z(n9407) );
  XNOR U9519 ( .A(n9430), .B(n9431), .Z(n9429) );
  XNOR U9520 ( .A(n9432), .B(n9433), .Z(n9428) );
  XNOR U9521 ( .A(key[204]), .B(n9434), .Z(n9433) );
  XOR U9522 ( .A(n9372), .B(n9387), .Z(n9421) );
  XOR U9523 ( .A(n9435), .B(n9436), .Z(n9387) );
  XNOR U9524 ( .A(n9392), .B(n9437), .Z(n9436) );
  XOR U9525 ( .A(n9438), .B(n9439), .Z(n9437) );
  XOR U9526 ( .A(n9440), .B(n9441), .Z(n9392) );
  XNOR U9527 ( .A(n9442), .B(n9443), .Z(n9441) );
  XOR U9528 ( .A(n9444), .B(n9445), .Z(n9440) );
  XOR U9529 ( .A(key[201]), .B(n9446), .Z(n9445) );
  XNOR U9530 ( .A(n9447), .B(n9448), .Z(n9435) );
  XNOR U9531 ( .A(key[203]), .B(n9449), .Z(n9448) );
  XOR U9532 ( .A(n9450), .B(n9451), .Z(n9372) );
  XOR U9533 ( .A(n9452), .B(n9453), .Z(n9451) );
  XOR U9534 ( .A(n9454), .B(n9455), .Z(n9450) );
  XNOR U9535 ( .A(key[200]), .B(n9456), .Z(n9455) );
  XNOR U9536 ( .A(n9457), .B(n9458), .Z(n3968) );
  XNOR U9537 ( .A(n8483), .B(n8383), .Z(n9458) );
  XNOR U9538 ( .A(n9459), .B(n9460), .Z(n8383) );
  XNOR U9539 ( .A(n8497), .B(n9461), .Z(n9460) );
  OR U9540 ( .A(n8388), .B(n9462), .Z(n9461) );
  OR U9541 ( .A(n9463), .B(n8493), .Z(n8497) );
  XNOR U9542 ( .A(n8388), .B(n8491), .Z(n8493) );
  XOR U9543 ( .A(n9464), .B(n8485), .Z(n8483) );
  NANDN U9544 ( .A(n9465), .B(n9466), .Z(n8485) );
  ANDN U9545 ( .B(n9467), .A(n9468), .Z(n9464) );
  XNOR U9546 ( .A(n8403), .B(n9469), .Z(n9457) );
  XOR U9547 ( .A(n8480), .B(n9470), .Z(n9469) );
  ANDN U9548 ( .B(n8410), .A(n9471), .Z(n9470) );
  ANDN U9549 ( .B(n9472), .A(n9473), .Z(n8480) );
  XNOR U9550 ( .A(n9459), .B(n9474), .Z(n8403) );
  XNOR U9551 ( .A(n9475), .B(n8407), .Z(n9474) );
  XOR U9552 ( .A(n8481), .B(n8410), .Z(n9472) );
  ANDN U9553 ( .B(n8481), .A(n9477), .Z(n9475) );
  XNOR U9554 ( .A(n8405), .B(n9478), .Z(n9459) );
  XNOR U9555 ( .A(n9479), .B(n9480), .Z(n9478) );
  NANDN U9556 ( .A(n8487), .B(n9481), .Z(n9480) );
  XOR U9557 ( .A(n9482), .B(n9479), .Z(n8405) );
  OR U9558 ( .A(n9465), .B(n9483), .Z(n9479) );
  XOR U9559 ( .A(n9484), .B(n8487), .Z(n9465) );
  XOR U9560 ( .A(n8491), .B(n8410), .Z(n8487) );
  XOR U9561 ( .A(n9485), .B(n9486), .Z(n8410) );
  NANDN U9562 ( .A(n9487), .B(n9488), .Z(n9486) );
  XNOR U9563 ( .A(n9489), .B(n9490), .Z(n8491) );
  OR U9564 ( .A(n9487), .B(n9491), .Z(n9490) );
  ANDN U9565 ( .B(n9484), .A(n9492), .Z(n9482) );
  IV U9566 ( .A(n9468), .Z(n9484) );
  XOR U9567 ( .A(n8388), .B(n8481), .Z(n9468) );
  XNOR U9568 ( .A(n9493), .B(n9485), .Z(n8481) );
  NANDN U9569 ( .A(n9494), .B(n9495), .Z(n9485) );
  ANDN U9570 ( .B(n9496), .A(n9497), .Z(n9493) );
  NANDN U9571 ( .A(n9494), .B(n9499), .Z(n9489) );
  XOR U9572 ( .A(n9500), .B(n9487), .Z(n9494) );
  XNOR U9573 ( .A(n9501), .B(n9502), .Z(n9487) );
  XOR U9574 ( .A(n9503), .B(n9496), .Z(n9502) );
  XNOR U9575 ( .A(n9504), .B(n9505), .Z(n9501) );
  XNOR U9576 ( .A(n9506), .B(n9507), .Z(n9505) );
  ANDN U9577 ( .B(n9496), .A(n9508), .Z(n9506) );
  IV U9578 ( .A(n9509), .Z(n9496) );
  ANDN U9579 ( .B(n9500), .A(n9508), .Z(n9498) );
  IV U9580 ( .A(n9504), .Z(n9508) );
  IV U9581 ( .A(n9497), .Z(n9500) );
  XNOR U9582 ( .A(n9503), .B(n9510), .Z(n9497) );
  XOR U9583 ( .A(n9511), .B(n9507), .Z(n9510) );
  NAND U9584 ( .A(n9499), .B(n9495), .Z(n9507) );
  XNOR U9585 ( .A(n9488), .B(n9509), .Z(n9495) );
  XOR U9586 ( .A(n9512), .B(n9513), .Z(n9509) );
  XOR U9587 ( .A(n9514), .B(n9515), .Z(n9513) );
  XNOR U9588 ( .A(n8492), .B(n9516), .Z(n9515) );
  XNOR U9589 ( .A(n9517), .B(n9518), .Z(n9512) );
  XNOR U9590 ( .A(n9519), .B(n9520), .Z(n9518) );
  ANDN U9591 ( .B(n9521), .A(n9462), .Z(n9519) );
  XNOR U9592 ( .A(n9504), .B(n9491), .Z(n9499) );
  XOR U9593 ( .A(n9522), .B(n9523), .Z(n9504) );
  XNOR U9594 ( .A(n9524), .B(n9516), .Z(n9523) );
  XOR U9595 ( .A(n9525), .B(n9526), .Z(n9516) );
  XNOR U9596 ( .A(n9527), .B(n9528), .Z(n9526) );
  NAND U9597 ( .A(n9481), .B(n8488), .Z(n9528) );
  XNOR U9598 ( .A(n9529), .B(n9530), .Z(n9522) );
  ANDN U9599 ( .B(n9531), .A(n9477), .Z(n9529) );
  ANDN U9600 ( .B(n9488), .A(n9491), .Z(n9511) );
  XOR U9601 ( .A(n9491), .B(n9488), .Z(n9503) );
  XNOR U9602 ( .A(n9532), .B(n9533), .Z(n9488) );
  XNOR U9603 ( .A(n9525), .B(n9534), .Z(n9533) );
  XOR U9604 ( .A(n9524), .B(n8389), .Z(n9534) );
  XOR U9605 ( .A(n9462), .B(n9535), .Z(n9532) );
  XNOR U9606 ( .A(n9536), .B(n9520), .Z(n9535) );
  OR U9607 ( .A(n8494), .B(n9463), .Z(n9520) );
  XNOR U9608 ( .A(n9462), .B(n8498), .Z(n9463) );
  XOR U9609 ( .A(n8389), .B(n8492), .Z(n8494) );
  ANDN U9610 ( .B(n8492), .A(n8498), .Z(n9536) );
  XOR U9611 ( .A(n9537), .B(n9538), .Z(n9491) );
  XOR U9612 ( .A(n9525), .B(n9514), .Z(n9538) );
  XOR U9613 ( .A(n8409), .B(n9471), .Z(n9514) );
  XOR U9614 ( .A(n9539), .B(n9527), .Z(n9525) );
  NANDN U9615 ( .A(n9483), .B(n9466), .Z(n9527) );
  XOR U9616 ( .A(n9467), .B(n8488), .Z(n9466) );
  XNOR U9617 ( .A(n9531), .B(n9540), .Z(n8492) );
  XOR U9618 ( .A(n9541), .B(n9542), .Z(n9540) );
  XOR U9619 ( .A(n9492), .B(n9481), .Z(n9483) );
  XNOR U9620 ( .A(n8498), .B(n8409), .Z(n9481) );
  IV U9621 ( .A(n9517), .Z(n8498) );
  XOR U9622 ( .A(n9543), .B(n9544), .Z(n9517) );
  XOR U9623 ( .A(n9545), .B(n9546), .Z(n9544) );
  XNOR U9624 ( .A(n9462), .B(n9547), .Z(n9543) );
  ANDN U9625 ( .B(n9467), .A(n9492), .Z(n9539) );
  XNOR U9626 ( .A(n9462), .B(n9477), .Z(n9492) );
  XOR U9627 ( .A(n9531), .B(n9521), .Z(n9467) );
  IV U9628 ( .A(n8389), .Z(n9521) );
  XOR U9629 ( .A(n9548), .B(n9549), .Z(n8389) );
  XOR U9630 ( .A(n9550), .B(n9546), .Z(n9549) );
  XNOR U9631 ( .A(n9551), .B(n6243), .Z(n9546) );
  XNOR U9632 ( .A(n9552), .B(n9553), .Z(n6243) );
  XOR U9633 ( .A(n7193), .B(n7180), .Z(n9553) );
  XOR U9634 ( .A(n9554), .B(n7152), .Z(n7180) );
  XOR U9635 ( .A(n9555), .B(n6287), .Z(n7193) );
  XOR U9636 ( .A(n7196), .B(n8202), .Z(n9552) );
  IV U9637 ( .A(n9556), .Z(n8202) );
  IV U9638 ( .A(n9557), .Z(n7196) );
  XOR U9639 ( .A(n8184), .B(n9558), .Z(n9551) );
  XOR U9640 ( .A(key[308]), .B(n8185), .Z(n9558) );
  XOR U9641 ( .A(n8198), .B(n6261), .Z(n8184) );
  XNOR U9642 ( .A(n9559), .B(n9560), .Z(n6261) );
  XNOR U9643 ( .A(n9561), .B(n9562), .Z(n9560) );
  XNOR U9644 ( .A(n9563), .B(n9564), .Z(n9559) );
  XOR U9645 ( .A(n9565), .B(n9566), .Z(n9564) );
  ANDN U9646 ( .B(n9567), .A(n9568), .Z(n9566) );
  IV U9647 ( .A(n8482), .Z(n9531) );
  XOR U9648 ( .A(n9524), .B(n9569), .Z(n9537) );
  XNOR U9649 ( .A(n9570), .B(n9530), .Z(n9569) );
  OR U9650 ( .A(n9473), .B(n9476), .Z(n9530) );
  XNOR U9651 ( .A(n9571), .B(n8409), .Z(n9476) );
  XNOR U9652 ( .A(n8482), .B(n9471), .Z(n9473) );
  ANDN U9653 ( .B(n8409), .A(n9471), .Z(n9570) );
  XOR U9654 ( .A(n9548), .B(n9572), .Z(n9471) );
  XNOR U9655 ( .A(n9573), .B(n9550), .Z(n9572) );
  XOR U9656 ( .A(n9550), .B(n9548), .Z(n8409) );
  XNOR U9657 ( .A(n9477), .B(n8482), .Z(n9524) );
  XOR U9658 ( .A(n9548), .B(n9574), .Z(n8482) );
  XNOR U9659 ( .A(n9550), .B(n9545), .Z(n9574) );
  XOR U9660 ( .A(n9575), .B(n9576), .Z(n9545) );
  XOR U9661 ( .A(n9577), .B(n6255), .Z(n9576) );
  XNOR U9662 ( .A(n7163), .B(n8217), .Z(n6255) );
  XNOR U9663 ( .A(n9578), .B(n9579), .Z(n8217) );
  XOR U9664 ( .A(n9580), .B(n9581), .Z(n9579) );
  XOR U9665 ( .A(n9582), .B(n9583), .Z(n7163) );
  XNOR U9666 ( .A(n9584), .B(n9585), .Z(n9583) );
  XOR U9667 ( .A(n9586), .B(n9587), .Z(n9582) );
  XOR U9668 ( .A(key[311]), .B(n8198), .Z(n9575) );
  XNOR U9669 ( .A(n9588), .B(n9589), .Z(n9548) );
  XNOR U9670 ( .A(n9556), .B(n6260), .Z(n9589) );
  XNOR U9671 ( .A(n7181), .B(n7168), .Z(n6260) );
  XOR U9672 ( .A(n9590), .B(n9591), .Z(n7168) );
  XNOR U9673 ( .A(n9554), .B(n9581), .Z(n9591) );
  XNOR U9674 ( .A(n9592), .B(n9593), .Z(n9581) );
  XNOR U9675 ( .A(n9594), .B(n9595), .Z(n9593) );
  OR U9676 ( .A(n9596), .B(n9597), .Z(n9595) );
  XNOR U9677 ( .A(n9598), .B(n9599), .Z(n9590) );
  XOR U9678 ( .A(n9600), .B(n9601), .Z(n9599) );
  ANDN U9679 ( .B(n9602), .A(n9603), .Z(n9601) );
  XOR U9680 ( .A(n9604), .B(n9605), .Z(n7181) );
  XNOR U9681 ( .A(n9555), .B(n9585), .Z(n9605) );
  XNOR U9682 ( .A(n9606), .B(n9607), .Z(n9585) );
  XNOR U9683 ( .A(n9608), .B(n9609), .Z(n9607) );
  OR U9684 ( .A(n9610), .B(n9611), .Z(n9609) );
  XNOR U9685 ( .A(n9612), .B(n9613), .Z(n9604) );
  XNOR U9686 ( .A(n9614), .B(n9615), .Z(n9613) );
  ANDN U9687 ( .B(n9616), .A(n9617), .Z(n9615) );
  XOR U9688 ( .A(n9618), .B(n9619), .Z(n9556) );
  XNOR U9689 ( .A(n9620), .B(n9621), .Z(n9619) );
  XNOR U9690 ( .A(n9622), .B(n9623), .Z(n9618) );
  XOR U9691 ( .A(n9624), .B(n9625), .Z(n9623) );
  ANDN U9692 ( .B(n9626), .A(n9627), .Z(n9625) );
  XNOR U9693 ( .A(key[309]), .B(n8216), .Z(n9588) );
  XOR U9694 ( .A(n6275), .B(n6263), .Z(n8216) );
  IV U9695 ( .A(n8205), .Z(n6275) );
  XOR U9696 ( .A(n9628), .B(n9629), .Z(n8205) );
  IV U9697 ( .A(n9571), .Z(n9477) );
  XNOR U9698 ( .A(n9542), .B(n9630), .Z(n9571) );
  XOR U9699 ( .A(n9631), .B(n9632), .Z(n9550) );
  XNOR U9700 ( .A(n9462), .B(n6267), .Z(n9632) );
  XOR U9701 ( .A(n7167), .B(n9577), .Z(n6267) );
  XNOR U9702 ( .A(n9557), .B(n8197), .Z(n9577) );
  XNOR U9703 ( .A(n9633), .B(n9634), .Z(n8197) );
  XNOR U9704 ( .A(n9635), .B(n9621), .Z(n9634) );
  XNOR U9705 ( .A(n9636), .B(n9637), .Z(n9621) );
  XNOR U9706 ( .A(n9638), .B(n9639), .Z(n9637) );
  NANDN U9707 ( .A(n9640), .B(n9641), .Z(n9639) );
  XOR U9708 ( .A(n9642), .B(n9643), .Z(n9633) );
  XOR U9709 ( .A(n7160), .B(n6259), .Z(n7167) );
  XOR U9710 ( .A(n9584), .B(n9644), .Z(n6259) );
  IV U9711 ( .A(n8203), .Z(n7160) );
  XOR U9712 ( .A(n9580), .B(n9645), .Z(n8203) );
  XNOR U9713 ( .A(n9646), .B(n9647), .Z(n9462) );
  XNOR U9714 ( .A(n7189), .B(n6254), .Z(n9647) );
  XOR U9715 ( .A(n9557), .B(n7162), .Z(n6254) );
  IV U9716 ( .A(n6270), .Z(n7162) );
  XOR U9717 ( .A(n9648), .B(n9555), .Z(n6270) );
  XNOR U9718 ( .A(n9606), .B(n9649), .Z(n9555) );
  XOR U9719 ( .A(n9650), .B(n9651), .Z(n9649) );
  ANDN U9720 ( .B(n9652), .A(n9653), .Z(n9650) );
  XNOR U9721 ( .A(n9654), .B(n9655), .Z(n9606) );
  XNOR U9722 ( .A(n9656), .B(n9657), .Z(n9655) );
  NAND U9723 ( .A(n9658), .B(n9659), .Z(n9657) );
  XOR U9724 ( .A(n6285), .B(n6271), .Z(n7189) );
  IV U9725 ( .A(n8212), .Z(n6285) );
  XOR U9726 ( .A(n9660), .B(n9661), .Z(n8212) );
  XNOR U9727 ( .A(n9662), .B(n9628), .Z(n9661) );
  XOR U9728 ( .A(key[304]), .B(n8199), .Z(n9646) );
  IV U9729 ( .A(n8187), .Z(n8199) );
  XNOR U9730 ( .A(n9592), .B(n9663), .Z(n9554) );
  XOR U9731 ( .A(n9664), .B(n9665), .Z(n9663) );
  ANDN U9732 ( .B(n9666), .A(n9667), .Z(n9664) );
  XNOR U9733 ( .A(n9668), .B(n9669), .Z(n9592) );
  XNOR U9734 ( .A(n9670), .B(n9671), .Z(n9669) );
  NAND U9735 ( .A(n9672), .B(n9673), .Z(n9671) );
  XOR U9736 ( .A(n8209), .B(n9675), .Z(n9631) );
  XNOR U9737 ( .A(key[310]), .B(n6263), .Z(n9675) );
  XOR U9738 ( .A(n9643), .B(n9676), .Z(n6263) );
  XOR U9739 ( .A(n8198), .B(n8196), .Z(n8209) );
  IV U9740 ( .A(n6256), .Z(n8196) );
  XOR U9741 ( .A(n9677), .B(n9678), .Z(n6256) );
  XNOR U9742 ( .A(n9679), .B(n9562), .Z(n9678) );
  XNOR U9743 ( .A(n9680), .B(n9681), .Z(n9562) );
  XNOR U9744 ( .A(n9682), .B(n9683), .Z(n9681) );
  NANDN U9745 ( .A(n9684), .B(n9685), .Z(n9683) );
  XOR U9746 ( .A(n9662), .B(n9628), .Z(n9677) );
  XNOR U9747 ( .A(n9686), .B(n9687), .Z(n9628) );
  XOR U9748 ( .A(n9688), .B(n9689), .Z(n9547) );
  XNOR U9749 ( .A(n6282), .B(n9690), .Z(n9689) );
  XNOR U9750 ( .A(n8220), .B(n9573), .Z(n9690) );
  IV U9751 ( .A(n9541), .Z(n9573) );
  XNOR U9752 ( .A(n9691), .B(n9692), .Z(n9541) );
  XNOR U9753 ( .A(n6271), .B(n7151), .Z(n9692) );
  XNOR U9754 ( .A(n6296), .B(n9693), .Z(n7151) );
  XNOR U9755 ( .A(n9694), .B(n9695), .Z(n6271) );
  XNOR U9756 ( .A(n9642), .B(n9643), .Z(n9695) );
  XNOR U9757 ( .A(n9696), .B(n9697), .Z(n9643) );
  XNOR U9758 ( .A(key[305]), .B(n6289), .Z(n9691) );
  XNOR U9759 ( .A(n8214), .B(n6274), .Z(n6289) );
  XOR U9760 ( .A(n9584), .B(n9698), .Z(n6274) );
  XOR U9761 ( .A(n9699), .B(n9587), .Z(n9698) );
  XOR U9762 ( .A(n9648), .B(n9700), .Z(n9584) );
  IV U9763 ( .A(n9701), .Z(n9648) );
  IV U9764 ( .A(n7190), .Z(n8214) );
  XOR U9765 ( .A(n9580), .B(n9702), .Z(n7190) );
  XOR U9766 ( .A(n9703), .B(n9704), .Z(n9702) );
  XOR U9767 ( .A(n9705), .B(n9674), .Z(n9580) );
  XNOR U9768 ( .A(n8198), .B(n6244), .Z(n8220) );
  XOR U9769 ( .A(n9686), .B(n9679), .Z(n6296) );
  XOR U9770 ( .A(n9563), .B(n9686), .Z(n8198) );
  XNOR U9771 ( .A(n9706), .B(n9707), .Z(n9686) );
  XOR U9772 ( .A(n9708), .B(n9682), .Z(n9707) );
  OR U9773 ( .A(n9709), .B(n9710), .Z(n9682) );
  ANDN U9774 ( .B(n9711), .A(n9712), .Z(n9708) );
  XNOR U9775 ( .A(n9680), .B(n9713), .Z(n9563) );
  XNOR U9776 ( .A(n9714), .B(n9715), .Z(n9713) );
  ANDN U9777 ( .B(n9716), .A(n9717), .Z(n9714) );
  XNOR U9778 ( .A(n9706), .B(n9718), .Z(n9680) );
  XNOR U9779 ( .A(n9719), .B(n9720), .Z(n9718) );
  NANDN U9780 ( .A(n9721), .B(n9722), .Z(n9720) );
  XNOR U9781 ( .A(n9557), .B(n8185), .Z(n6282) );
  XOR U9782 ( .A(n9622), .B(n9693), .Z(n8185) );
  XOR U9783 ( .A(n9622), .B(n9696), .Z(n9557) );
  XNOR U9784 ( .A(n9636), .B(n9723), .Z(n9622) );
  XNOR U9785 ( .A(n9724), .B(n9725), .Z(n9723) );
  ANDN U9786 ( .B(n9726), .A(n9727), .Z(n9724) );
  XNOR U9787 ( .A(n9728), .B(n9729), .Z(n9636) );
  XNOR U9788 ( .A(n9730), .B(n9731), .Z(n9729) );
  NANDN U9789 ( .A(n9732), .B(n9733), .Z(n9731) );
  XOR U9790 ( .A(n6281), .B(n9734), .Z(n9688) );
  XNOR U9791 ( .A(key[307]), .B(n6297), .Z(n9734) );
  XOR U9792 ( .A(n7191), .B(n6295), .Z(n6281) );
  XOR U9793 ( .A(n9735), .B(n9736), .Z(n6295) );
  XOR U9794 ( .A(n9700), .B(n9644), .Z(n9736) );
  XOR U9795 ( .A(n9737), .B(n9738), .Z(n9644) );
  XOR U9796 ( .A(n9739), .B(n9614), .Z(n9738) );
  NANDN U9797 ( .A(n9740), .B(n9741), .Z(n9614) );
  ANDN U9798 ( .B(n9652), .A(n9742), .Z(n9739) );
  XNOR U9799 ( .A(n9612), .B(n9743), .Z(n9700) );
  XNOR U9800 ( .A(n9744), .B(n9745), .Z(n9743) );
  NANDN U9801 ( .A(n9746), .B(n9747), .Z(n9745) );
  XNOR U9802 ( .A(n9699), .B(n9587), .Z(n9735) );
  XOR U9803 ( .A(n9737), .B(n9748), .Z(n9587) );
  XNOR U9804 ( .A(n9744), .B(n9749), .Z(n9748) );
  OR U9805 ( .A(n9610), .B(n9750), .Z(n9749) );
  OR U9806 ( .A(n9751), .B(n9752), .Z(n9744) );
  XNOR U9807 ( .A(n9612), .B(n9753), .Z(n9737) );
  XNOR U9808 ( .A(n9754), .B(n9755), .Z(n9753) );
  NAND U9809 ( .A(n9756), .B(n9658), .Z(n9755) );
  XOR U9810 ( .A(n9757), .B(n9754), .Z(n9612) );
  NANDN U9811 ( .A(n9758), .B(n9759), .Z(n9754) );
  ANDN U9812 ( .B(n9760), .A(n9761), .Z(n9757) );
  IV U9813 ( .A(n9586), .Z(n9699) );
  XOR U9814 ( .A(n9578), .B(n9762), .Z(n7191) );
  XNOR U9815 ( .A(n9705), .B(n9645), .Z(n9762) );
  XNOR U9816 ( .A(n9763), .B(n9764), .Z(n9645) );
  XNOR U9817 ( .A(n9765), .B(n9600), .Z(n9764) );
  ANDN U9818 ( .B(n9766), .A(n9767), .Z(n9600) );
  ANDN U9819 ( .B(n9666), .A(n9768), .Z(n9765) );
  XNOR U9820 ( .A(n9598), .B(n9769), .Z(n9705) );
  XNOR U9821 ( .A(n9770), .B(n9771), .Z(n9769) );
  NANDN U9822 ( .A(n9772), .B(n9773), .Z(n9771) );
  XNOR U9823 ( .A(n9703), .B(n9704), .Z(n9578) );
  XOR U9824 ( .A(n9763), .B(n9774), .Z(n9704) );
  XNOR U9825 ( .A(n9770), .B(n9775), .Z(n9774) );
  NANDN U9826 ( .A(n9596), .B(n9776), .Z(n9775) );
  OR U9827 ( .A(n9777), .B(n9778), .Z(n9770) );
  XNOR U9828 ( .A(n9598), .B(n9779), .Z(n9763) );
  XNOR U9829 ( .A(n9780), .B(n9781), .Z(n9779) );
  NAND U9830 ( .A(n9782), .B(n9672), .Z(n9781) );
  XOR U9831 ( .A(n9783), .B(n9780), .Z(n9598) );
  NANDN U9832 ( .A(n9784), .B(n9785), .Z(n9780) );
  ANDN U9833 ( .B(n9786), .A(n9787), .Z(n9783) );
  XOR U9834 ( .A(n9788), .B(n9789), .Z(n9542) );
  XOR U9835 ( .A(n8226), .B(n9693), .Z(n9789) );
  IV U9836 ( .A(n6286), .Z(n9693) );
  XOR U9837 ( .A(n9696), .B(n9635), .Z(n6286) );
  XNOR U9838 ( .A(n9728), .B(n9790), .Z(n9696) );
  XOR U9839 ( .A(n9791), .B(n9638), .Z(n9790) );
  OR U9840 ( .A(n9792), .B(n9793), .Z(n9638) );
  ANDN U9841 ( .B(n9794), .A(n9795), .Z(n9791) );
  XOR U9842 ( .A(n6290), .B(n6297), .Z(n8226) );
  XOR U9843 ( .A(n9796), .B(n9797), .Z(n6297) );
  XNOR U9844 ( .A(n9635), .B(n9676), .Z(n9797) );
  XNOR U9845 ( .A(n9798), .B(n9799), .Z(n9676) );
  XNOR U9846 ( .A(n9800), .B(n9624), .Z(n9799) );
  ANDN U9847 ( .B(n9801), .A(n9802), .Z(n9624) );
  ANDN U9848 ( .B(n9803), .A(n9727), .Z(n9800) );
  IV U9849 ( .A(n9804), .Z(n9727) );
  IV U9850 ( .A(n9694), .Z(n9635) );
  XOR U9851 ( .A(n9728), .B(n9805), .Z(n9694) );
  XOR U9852 ( .A(n9725), .B(n9806), .Z(n9805) );
  NANDN U9853 ( .A(n9807), .B(n9626), .Z(n9806) );
  XOR U9854 ( .A(n9804), .B(n9626), .Z(n9801) );
  XOR U9855 ( .A(n9809), .B(n9730), .Z(n9728) );
  OR U9856 ( .A(n9810), .B(n9811), .Z(n9730) );
  NOR U9857 ( .A(n9812), .B(n9813), .Z(n9809) );
  XOR U9858 ( .A(n9642), .B(n9697), .Z(n9796) );
  XOR U9859 ( .A(n9620), .B(n9814), .Z(n9697) );
  XNOR U9860 ( .A(n9815), .B(n9816), .Z(n9814) );
  NANDN U9861 ( .A(n9817), .B(n9794), .Z(n9816) );
  XNOR U9862 ( .A(n9815), .B(n9819), .Z(n9818) );
  NANDN U9863 ( .A(n9820), .B(n9641), .Z(n9819) );
  OR U9864 ( .A(n9793), .B(n9821), .Z(n9815) );
  XNOR U9865 ( .A(n9641), .B(n9794), .Z(n9793) );
  XNOR U9866 ( .A(n9620), .B(n9822), .Z(n9798) );
  XNOR U9867 ( .A(n9823), .B(n9824), .Z(n9822) );
  NANDN U9868 ( .A(n9732), .B(n9825), .Z(n9824) );
  XOR U9869 ( .A(n9826), .B(n9823), .Z(n9620) );
  NANDN U9870 ( .A(n9810), .B(n9827), .Z(n9823) );
  XNOR U9871 ( .A(n9812), .B(n9732), .Z(n9810) );
  XNOR U9872 ( .A(n9794), .B(n9626), .Z(n9732) );
  XOR U9873 ( .A(n9828), .B(n9829), .Z(n9626) );
  NANDN U9874 ( .A(n9830), .B(n9831), .Z(n9829) );
  XOR U9875 ( .A(n9832), .B(n9833), .Z(n9794) );
  NANDN U9876 ( .A(n9830), .B(n9834), .Z(n9833) );
  ANDN U9877 ( .B(n9835), .A(n9812), .Z(n9826) );
  XNOR U9878 ( .A(n9804), .B(n9641), .Z(n9812) );
  XNOR U9879 ( .A(n9836), .B(n9832), .Z(n9641) );
  NANDN U9880 ( .A(n9837), .B(n9838), .Z(n9832) );
  XOR U9881 ( .A(n9834), .B(n9839), .Z(n9838) );
  ANDN U9882 ( .B(n9839), .A(n9840), .Z(n9836) );
  XNOR U9883 ( .A(n9841), .B(n9828), .Z(n9804) );
  NANDN U9884 ( .A(n9837), .B(n9842), .Z(n9828) );
  XOR U9885 ( .A(n9843), .B(n9831), .Z(n9842) );
  XNOR U9886 ( .A(n9844), .B(n9845), .Z(n9830) );
  XOR U9887 ( .A(n9846), .B(n9847), .Z(n9845) );
  XNOR U9888 ( .A(n9848), .B(n9849), .Z(n9844) );
  XNOR U9889 ( .A(n9850), .B(n9851), .Z(n9849) );
  ANDN U9890 ( .B(n9843), .A(n9847), .Z(n9850) );
  ANDN U9891 ( .B(n9843), .A(n9840), .Z(n9841) );
  XNOR U9892 ( .A(n9846), .B(n9852), .Z(n9840) );
  XOR U9893 ( .A(n9853), .B(n9851), .Z(n9852) );
  NAND U9894 ( .A(n9854), .B(n9855), .Z(n9851) );
  XNOR U9895 ( .A(n9848), .B(n9831), .Z(n9855) );
  IV U9896 ( .A(n9843), .Z(n9848) );
  XNOR U9897 ( .A(n9834), .B(n9847), .Z(n9854) );
  IV U9898 ( .A(n9839), .Z(n9847) );
  XOR U9899 ( .A(n9856), .B(n9857), .Z(n9839) );
  XNOR U9900 ( .A(n9858), .B(n9859), .Z(n9857) );
  XNOR U9901 ( .A(n9860), .B(n9861), .Z(n9856) );
  ANDN U9902 ( .B(n9726), .A(n9862), .Z(n9860) );
  AND U9903 ( .A(n9831), .B(n9834), .Z(n9853) );
  XNOR U9904 ( .A(n9831), .B(n9834), .Z(n9846) );
  XNOR U9905 ( .A(n9863), .B(n9864), .Z(n9834) );
  XNOR U9906 ( .A(n9865), .B(n9859), .Z(n9864) );
  XOR U9907 ( .A(n9866), .B(n9867), .Z(n9863) );
  XNOR U9908 ( .A(n9868), .B(n9861), .Z(n9867) );
  OR U9909 ( .A(n9802), .B(n9808), .Z(n9861) );
  XNOR U9910 ( .A(n9726), .B(n9869), .Z(n9808) );
  XNOR U9911 ( .A(n9862), .B(n9627), .Z(n9802) );
  ANDN U9912 ( .B(n9870), .A(n9807), .Z(n9868) );
  XNOR U9913 ( .A(n9871), .B(n9872), .Z(n9831) );
  XNOR U9914 ( .A(n9859), .B(n9873), .Z(n9872) );
  XOR U9915 ( .A(n9820), .B(n9866), .Z(n9873) );
  XNOR U9916 ( .A(n9726), .B(n9862), .Z(n9859) );
  XOR U9917 ( .A(n9640), .B(n9874), .Z(n9871) );
  XNOR U9918 ( .A(n9875), .B(n9876), .Z(n9874) );
  ANDN U9919 ( .B(n9877), .A(n9795), .Z(n9875) );
  XNOR U9920 ( .A(n9878), .B(n9879), .Z(n9843) );
  XNOR U9921 ( .A(n9865), .B(n9880), .Z(n9879) );
  XNOR U9922 ( .A(n9817), .B(n9858), .Z(n9880) );
  XOR U9923 ( .A(n9866), .B(n9881), .Z(n9858) );
  XNOR U9924 ( .A(n9882), .B(n9883), .Z(n9881) );
  NAND U9925 ( .A(n9733), .B(n9825), .Z(n9883) );
  XNOR U9926 ( .A(n9884), .B(n9882), .Z(n9866) );
  NANDN U9927 ( .A(n9811), .B(n9827), .Z(n9882) );
  XOR U9928 ( .A(n9835), .B(n9825), .Z(n9827) );
  XNOR U9929 ( .A(n9877), .B(n9627), .Z(n9825) );
  XOR U9930 ( .A(n9813), .B(n9733), .Z(n9811) );
  XNOR U9931 ( .A(n9795), .B(n9869), .Z(n9733) );
  ANDN U9932 ( .B(n9835), .A(n9813), .Z(n9884) );
  XOR U9933 ( .A(n9640), .B(n9726), .Z(n9813) );
  XNOR U9934 ( .A(n9885), .B(n9886), .Z(n9726) );
  XNOR U9935 ( .A(n9887), .B(n9888), .Z(n9886) );
  XOR U9936 ( .A(n9869), .B(n9870), .Z(n9865) );
  IV U9937 ( .A(n9627), .Z(n9870) );
  XOR U9938 ( .A(n9889), .B(n9890), .Z(n9627) );
  XOR U9939 ( .A(n9891), .B(n9888), .Z(n9890) );
  IV U9940 ( .A(n9807), .Z(n9869) );
  XOR U9941 ( .A(n9888), .B(n9892), .Z(n9807) );
  XNOR U9942 ( .A(n9893), .B(n9894), .Z(n9878) );
  XNOR U9943 ( .A(n9895), .B(n9876), .Z(n9894) );
  OR U9944 ( .A(n9821), .B(n9792), .Z(n9876) );
  XNOR U9945 ( .A(n9640), .B(n9795), .Z(n9792) );
  IV U9946 ( .A(n9893), .Z(n9795) );
  XOR U9947 ( .A(n9820), .B(n9877), .Z(n9821) );
  IV U9948 ( .A(n9817), .Z(n9877) );
  XOR U9949 ( .A(n9803), .B(n9896), .Z(n9817) );
  XNOR U9950 ( .A(n9897), .B(n9885), .Z(n9896) );
  XOR U9951 ( .A(n9898), .B(n9899), .Z(n9885) );
  XOR U9952 ( .A(n9900), .B(n9105), .Z(n9899) );
  XOR U9953 ( .A(n9901), .B(n9902), .Z(n9898) );
  XNOR U9954 ( .A(key[234]), .B(n9146), .Z(n9902) );
  NOR U9955 ( .A(n9820), .B(n9640), .Z(n9895) );
  XOR U9956 ( .A(n9903), .B(n9904), .Z(n9893) );
  XNOR U9957 ( .A(n9905), .B(n9906), .Z(n9904) );
  XNOR U9958 ( .A(n9640), .B(n9887), .Z(n9903) );
  XOR U9959 ( .A(n9907), .B(n9908), .Z(n9887) );
  XNOR U9960 ( .A(n9138), .B(n9909), .Z(n9908) );
  XOR U9961 ( .A(n9910), .B(n9897), .Z(n9909) );
  IV U9962 ( .A(n9891), .Z(n9897) );
  XNOR U9963 ( .A(n9911), .B(n9912), .Z(n9891) );
  XOR U9964 ( .A(n9104), .B(n9142), .Z(n9912) );
  XOR U9965 ( .A(n9913), .B(n9914), .Z(n9911) );
  XNOR U9966 ( .A(key[233]), .B(n9915), .Z(n9914) );
  XOR U9967 ( .A(n9916), .B(n9133), .Z(n9138) );
  XOR U9968 ( .A(n9137), .B(n9917), .Z(n9907) );
  XNOR U9969 ( .A(key[235]), .B(n9918), .Z(n9917) );
  IV U9970 ( .A(n9862), .Z(n9803) );
  XOR U9971 ( .A(n9889), .B(n9919), .Z(n9862) );
  XOR U9972 ( .A(n9888), .B(n9906), .Z(n9919) );
  XNOR U9973 ( .A(n9920), .B(n9921), .Z(n9906) );
  XNOR U9974 ( .A(n9922), .B(n9127), .Z(n9921) );
  XNOR U9975 ( .A(n9923), .B(n9924), .Z(n9127) );
  XOR U9976 ( .A(key[239]), .B(n9925), .Z(n9920) );
  XOR U9977 ( .A(n9889), .B(n9926), .Z(n9820) );
  XOR U9978 ( .A(n9888), .B(n9905), .Z(n9926) );
  XNOR U9979 ( .A(n9927), .B(n9130), .Z(n9905) );
  XNOR U9980 ( .A(n9928), .B(n9929), .Z(n9130) );
  XNOR U9981 ( .A(n9930), .B(n9931), .Z(n9929) );
  XNOR U9982 ( .A(n9916), .B(n9119), .Z(n9928) );
  XOR U9983 ( .A(n9932), .B(n9933), .Z(n9927) );
  XNOR U9984 ( .A(key[236]), .B(n9934), .Z(n9933) );
  XOR U9985 ( .A(n9935), .B(n9936), .Z(n9888) );
  XOR U9986 ( .A(n9640), .B(n9113), .Z(n9936) );
  XOR U9987 ( .A(n9937), .B(n9126), .Z(n9113) );
  XNOR U9988 ( .A(n9938), .B(n9939), .Z(n9126) );
  XNOR U9989 ( .A(n9940), .B(n9941), .Z(n9640) );
  XOR U9990 ( .A(n9942), .B(n9943), .Z(n9941) );
  XOR U9991 ( .A(n9944), .B(n9945), .Z(n9940) );
  XOR U9992 ( .A(key[232]), .B(n9946), .Z(n9945) );
  XNOR U9993 ( .A(n9947), .B(n9948), .Z(n9935) );
  XOR U9994 ( .A(key[238]), .B(n9949), .Z(n9948) );
  IV U9995 ( .A(n9892), .Z(n9889) );
  XOR U9996 ( .A(n9950), .B(n9951), .Z(n9892) );
  XNOR U9997 ( .A(n9952), .B(n9120), .Z(n9951) );
  XOR U9998 ( .A(n9953), .B(n9954), .Z(n9120) );
  XNOR U9999 ( .A(n9116), .B(n9955), .Z(n9950) );
  XOR U10000 ( .A(key[237]), .B(n9956), .Z(n9955) );
  XOR U10001 ( .A(n9957), .B(n9958), .Z(n6290) );
  XNOR U10002 ( .A(n9679), .B(n9629), .Z(n9958) );
  XNOR U10003 ( .A(n9959), .B(n9960), .Z(n9629) );
  XNOR U10004 ( .A(n9961), .B(n9565), .Z(n9960) );
  ANDN U10005 ( .B(n9962), .A(n9963), .Z(n9565) );
  ANDN U10006 ( .B(n9964), .A(n9717), .Z(n9961) );
  IV U10007 ( .A(n9965), .Z(n9717) );
  IV U10008 ( .A(n9660), .Z(n9679) );
  XOR U10009 ( .A(n9706), .B(n9966), .Z(n9660) );
  XOR U10010 ( .A(n9715), .B(n9967), .Z(n9966) );
  NANDN U10011 ( .A(n9968), .B(n9567), .Z(n9967) );
  XOR U10012 ( .A(n9965), .B(n9567), .Z(n9962) );
  XOR U10013 ( .A(n9970), .B(n9719), .Z(n9706) );
  OR U10014 ( .A(n9971), .B(n9972), .Z(n9719) );
  NOR U10015 ( .A(n9973), .B(n9974), .Z(n9970) );
  XOR U10016 ( .A(n9662), .B(n9687), .Z(n9957) );
  XOR U10017 ( .A(n9561), .B(n9975), .Z(n9687) );
  XNOR U10018 ( .A(n9976), .B(n9977), .Z(n9975) );
  NANDN U10019 ( .A(n9978), .B(n9711), .Z(n9977) );
  XNOR U10020 ( .A(n9976), .B(n9980), .Z(n9979) );
  NANDN U10021 ( .A(n9981), .B(n9685), .Z(n9980) );
  OR U10022 ( .A(n9710), .B(n9982), .Z(n9976) );
  XNOR U10023 ( .A(n9685), .B(n9711), .Z(n9710) );
  XNOR U10024 ( .A(n9561), .B(n9983), .Z(n9959) );
  XNOR U10025 ( .A(n9984), .B(n9985), .Z(n9983) );
  NANDN U10026 ( .A(n9721), .B(n9986), .Z(n9985) );
  XOR U10027 ( .A(n9987), .B(n9984), .Z(n9561) );
  NANDN U10028 ( .A(n9971), .B(n9988), .Z(n9984) );
  XNOR U10029 ( .A(n9973), .B(n9721), .Z(n9971) );
  XNOR U10030 ( .A(n9711), .B(n9567), .Z(n9721) );
  XOR U10031 ( .A(n9989), .B(n9990), .Z(n9567) );
  NANDN U10032 ( .A(n9991), .B(n9992), .Z(n9990) );
  XOR U10033 ( .A(n9993), .B(n9994), .Z(n9711) );
  NANDN U10034 ( .A(n9991), .B(n9995), .Z(n9994) );
  ANDN U10035 ( .B(n9996), .A(n9973), .Z(n9987) );
  XNOR U10036 ( .A(n9965), .B(n9685), .Z(n9973) );
  XNOR U10037 ( .A(n9997), .B(n9993), .Z(n9685) );
  NANDN U10038 ( .A(n9998), .B(n9999), .Z(n9993) );
  XOR U10039 ( .A(n9995), .B(n10000), .Z(n9999) );
  ANDN U10040 ( .B(n10000), .A(n10001), .Z(n9997) );
  XNOR U10041 ( .A(n10002), .B(n9989), .Z(n9965) );
  NANDN U10042 ( .A(n9998), .B(n10003), .Z(n9989) );
  XOR U10043 ( .A(n10004), .B(n9992), .Z(n10003) );
  XNOR U10044 ( .A(n10005), .B(n10006), .Z(n9991) );
  XOR U10045 ( .A(n10007), .B(n10008), .Z(n10006) );
  XNOR U10046 ( .A(n10009), .B(n10010), .Z(n10005) );
  XNOR U10047 ( .A(n10011), .B(n10012), .Z(n10010) );
  ANDN U10048 ( .B(n10004), .A(n10008), .Z(n10011) );
  ANDN U10049 ( .B(n10004), .A(n10001), .Z(n10002) );
  XNOR U10050 ( .A(n10007), .B(n10013), .Z(n10001) );
  XOR U10051 ( .A(n10014), .B(n10012), .Z(n10013) );
  NAND U10052 ( .A(n10015), .B(n10016), .Z(n10012) );
  XNOR U10053 ( .A(n10009), .B(n9992), .Z(n10016) );
  IV U10054 ( .A(n10004), .Z(n10009) );
  XNOR U10055 ( .A(n9995), .B(n10008), .Z(n10015) );
  IV U10056 ( .A(n10000), .Z(n10008) );
  XOR U10057 ( .A(n10017), .B(n10018), .Z(n10000) );
  XNOR U10058 ( .A(n10019), .B(n10020), .Z(n10018) );
  XNOR U10059 ( .A(n10021), .B(n10022), .Z(n10017) );
  ANDN U10060 ( .B(n9716), .A(n10023), .Z(n10021) );
  AND U10061 ( .A(n9992), .B(n9995), .Z(n10014) );
  XNOR U10062 ( .A(n9992), .B(n9995), .Z(n10007) );
  XNOR U10063 ( .A(n10024), .B(n10025), .Z(n9995) );
  XNOR U10064 ( .A(n10026), .B(n10020), .Z(n10025) );
  XOR U10065 ( .A(n10027), .B(n10028), .Z(n10024) );
  XNOR U10066 ( .A(n10029), .B(n10022), .Z(n10028) );
  OR U10067 ( .A(n9963), .B(n9969), .Z(n10022) );
  XNOR U10068 ( .A(n9716), .B(n10030), .Z(n9969) );
  XNOR U10069 ( .A(n10023), .B(n9568), .Z(n9963) );
  ANDN U10070 ( .B(n10031), .A(n9968), .Z(n10029) );
  XNOR U10071 ( .A(n10032), .B(n10033), .Z(n9992) );
  XNOR U10072 ( .A(n10020), .B(n10034), .Z(n10033) );
  XOR U10073 ( .A(n9981), .B(n10027), .Z(n10034) );
  XNOR U10074 ( .A(n9716), .B(n10023), .Z(n10020) );
  XOR U10075 ( .A(n9684), .B(n10035), .Z(n10032) );
  XNOR U10076 ( .A(n10036), .B(n10037), .Z(n10035) );
  ANDN U10077 ( .B(n10038), .A(n9712), .Z(n10036) );
  XNOR U10078 ( .A(n10039), .B(n10040), .Z(n10004) );
  XNOR U10079 ( .A(n10026), .B(n10041), .Z(n10040) );
  XNOR U10080 ( .A(n9978), .B(n10019), .Z(n10041) );
  XOR U10081 ( .A(n10027), .B(n10042), .Z(n10019) );
  XNOR U10082 ( .A(n10043), .B(n10044), .Z(n10042) );
  NAND U10083 ( .A(n9722), .B(n9986), .Z(n10044) );
  XNOR U10084 ( .A(n10045), .B(n10043), .Z(n10027) );
  NANDN U10085 ( .A(n9972), .B(n9988), .Z(n10043) );
  XOR U10086 ( .A(n9996), .B(n9986), .Z(n9988) );
  XNOR U10087 ( .A(n10038), .B(n9568), .Z(n9986) );
  XOR U10088 ( .A(n9974), .B(n9722), .Z(n9972) );
  XNOR U10089 ( .A(n9712), .B(n10030), .Z(n9722) );
  ANDN U10090 ( .B(n9996), .A(n9974), .Z(n10045) );
  XOR U10091 ( .A(n9684), .B(n9716), .Z(n9974) );
  XNOR U10092 ( .A(n10046), .B(n10047), .Z(n9716) );
  XNOR U10093 ( .A(n10048), .B(n10049), .Z(n10047) );
  XOR U10094 ( .A(n10030), .B(n10031), .Z(n10026) );
  IV U10095 ( .A(n9568), .Z(n10031) );
  XOR U10096 ( .A(n10050), .B(n10051), .Z(n9568) );
  XOR U10097 ( .A(n10052), .B(n10049), .Z(n10051) );
  IV U10098 ( .A(n9968), .Z(n10030) );
  XOR U10099 ( .A(n10049), .B(n10053), .Z(n9968) );
  XNOR U10100 ( .A(n10054), .B(n10055), .Z(n10039) );
  XNOR U10101 ( .A(n10056), .B(n10037), .Z(n10055) );
  OR U10102 ( .A(n9982), .B(n9709), .Z(n10037) );
  XNOR U10103 ( .A(n9684), .B(n9712), .Z(n9709) );
  IV U10104 ( .A(n10054), .Z(n9712) );
  XOR U10105 ( .A(n9981), .B(n10038), .Z(n9982) );
  IV U10106 ( .A(n9978), .Z(n10038) );
  XOR U10107 ( .A(n9964), .B(n10057), .Z(n9978) );
  XNOR U10108 ( .A(n10058), .B(n10046), .Z(n10057) );
  XOR U10109 ( .A(n10059), .B(n10060), .Z(n10046) );
  XNOR U10110 ( .A(n10061), .B(n10062), .Z(n10060) );
  XOR U10111 ( .A(key[146]), .B(n10063), .Z(n10059) );
  NOR U10112 ( .A(n9981), .B(n9684), .Z(n10056) );
  XOR U10113 ( .A(n10064), .B(n10065), .Z(n10054) );
  XNOR U10114 ( .A(n10066), .B(n10067), .Z(n10065) );
  XNOR U10115 ( .A(n9684), .B(n10048), .Z(n10064) );
  XOR U10116 ( .A(n10068), .B(n10069), .Z(n10048) );
  XOR U10117 ( .A(n8986), .B(n10070), .Z(n10069) );
  XNOR U10118 ( .A(n10071), .B(n10058), .Z(n10070) );
  IV U10119 ( .A(n10052), .Z(n10058) );
  XNOR U10120 ( .A(n10072), .B(n10073), .Z(n10052) );
  XOR U10121 ( .A(n10074), .B(n9000), .Z(n10073) );
  XOR U10122 ( .A(key[145]), .B(n10075), .Z(n10072) );
  XOR U10123 ( .A(n10076), .B(n10077), .Z(n8986) );
  XOR U10124 ( .A(n10078), .B(n10079), .Z(n10068) );
  XNOR U10125 ( .A(key[147]), .B(n10080), .Z(n10079) );
  IV U10126 ( .A(n10023), .Z(n9964) );
  XOR U10127 ( .A(n10050), .B(n10081), .Z(n10023) );
  XOR U10128 ( .A(n10049), .B(n10067), .Z(n10081) );
  XNOR U10129 ( .A(n10082), .B(n10083), .Z(n10067) );
  XNOR U10130 ( .A(n10084), .B(n10085), .Z(n10083) );
  XOR U10131 ( .A(key[151]), .B(n10076), .Z(n10082) );
  XOR U10132 ( .A(n10050), .B(n10086), .Z(n9981) );
  XOR U10133 ( .A(n10049), .B(n10066), .Z(n10086) );
  XNOR U10134 ( .A(n10087), .B(n10088), .Z(n10066) );
  XOR U10135 ( .A(n10089), .B(n8947), .Z(n10088) );
  XOR U10136 ( .A(n10076), .B(n10090), .Z(n8947) );
  XOR U10137 ( .A(key[148]), .B(n10091), .Z(n10087) );
  XOR U10138 ( .A(n10092), .B(n10093), .Z(n10049) );
  XOR U10139 ( .A(n9684), .B(n8971), .Z(n10093) );
  XNOR U10140 ( .A(n8978), .B(n10094), .Z(n8971) );
  XNOR U10141 ( .A(n10095), .B(n10096), .Z(n9684) );
  XNOR U10142 ( .A(n10097), .B(n8975), .Z(n10096) );
  XOR U10143 ( .A(key[144]), .B(n10098), .Z(n10095) );
  XOR U10144 ( .A(n10099), .B(n10100), .Z(n10092) );
  XOR U10145 ( .A(key[150]), .B(n10101), .Z(n10100) );
  IV U10146 ( .A(n10053), .Z(n10050) );
  XOR U10147 ( .A(n10102), .B(n10103), .Z(n10053) );
  XOR U10148 ( .A(n10104), .B(n10105), .Z(n10103) );
  XNOR U10149 ( .A(key[149]), .B(n10106), .Z(n10102) );
  XOR U10150 ( .A(key[306]), .B(n6299), .Z(n9788) );
  XNOR U10151 ( .A(n6287), .B(n7152), .Z(n6299) );
  XNOR U10152 ( .A(n9703), .B(n9674), .Z(n7152) );
  XNOR U10153 ( .A(n9668), .B(n10107), .Z(n9674) );
  XOR U10154 ( .A(n10108), .B(n9594), .Z(n10107) );
  OR U10155 ( .A(n9777), .B(n10109), .Z(n9594) );
  XNOR U10156 ( .A(n9596), .B(n9772), .Z(n9777) );
  NOR U10157 ( .A(n10110), .B(n9772), .Z(n10108) );
  XNOR U10158 ( .A(n9668), .B(n10111), .Z(n9703) );
  XNOR U10159 ( .A(n9665), .B(n10112), .Z(n10111) );
  NAND U10160 ( .A(n10113), .B(n9602), .Z(n10112) );
  XOR U10161 ( .A(n9666), .B(n9602), .Z(n9766) );
  XOR U10162 ( .A(n10115), .B(n9670), .Z(n9668) );
  OR U10163 ( .A(n9784), .B(n10116), .Z(n9670) );
  XOR U10164 ( .A(n9787), .B(n9672), .Z(n9784) );
  XNOR U10165 ( .A(n9772), .B(n9602), .Z(n9672) );
  XOR U10166 ( .A(n10117), .B(n10118), .Z(n9602) );
  NANDN U10167 ( .A(n10119), .B(n10120), .Z(n10118) );
  XNOR U10168 ( .A(n10121), .B(n10122), .Z(n9772) );
  OR U10169 ( .A(n10119), .B(n10123), .Z(n10122) );
  ANDN U10170 ( .B(n10124), .A(n9787), .Z(n10115) );
  XOR U10171 ( .A(n9596), .B(n9666), .Z(n9787) );
  XNOR U10172 ( .A(n10125), .B(n10117), .Z(n9666) );
  NANDN U10173 ( .A(n10126), .B(n10127), .Z(n10117) );
  ANDN U10174 ( .B(n10128), .A(n10129), .Z(n10125) );
  NANDN U10175 ( .A(n10126), .B(n10131), .Z(n10121) );
  XOR U10176 ( .A(n10132), .B(n10119), .Z(n10126) );
  XNOR U10177 ( .A(n10133), .B(n10134), .Z(n10119) );
  XOR U10178 ( .A(n10135), .B(n10128), .Z(n10134) );
  XNOR U10179 ( .A(n10136), .B(n10137), .Z(n10133) );
  XNOR U10180 ( .A(n10138), .B(n10139), .Z(n10137) );
  ANDN U10181 ( .B(n10128), .A(n10140), .Z(n10138) );
  IV U10182 ( .A(n10141), .Z(n10128) );
  ANDN U10183 ( .B(n10132), .A(n10140), .Z(n10130) );
  IV U10184 ( .A(n10136), .Z(n10140) );
  IV U10185 ( .A(n10129), .Z(n10132) );
  XNOR U10186 ( .A(n10135), .B(n10142), .Z(n10129) );
  XOR U10187 ( .A(n10143), .B(n10139), .Z(n10142) );
  NAND U10188 ( .A(n10131), .B(n10127), .Z(n10139) );
  XNOR U10189 ( .A(n10120), .B(n10141), .Z(n10127) );
  XOR U10190 ( .A(n10144), .B(n10145), .Z(n10141) );
  XOR U10191 ( .A(n10146), .B(n10147), .Z(n10145) );
  XNOR U10192 ( .A(n9773), .B(n10148), .Z(n10147) );
  XNOR U10193 ( .A(n10149), .B(n10150), .Z(n10144) );
  XNOR U10194 ( .A(n10151), .B(n10152), .Z(n10150) );
  ANDN U10195 ( .B(n9776), .A(n9597), .Z(n10151) );
  XNOR U10196 ( .A(n10136), .B(n10123), .Z(n10131) );
  XOR U10197 ( .A(n10153), .B(n10154), .Z(n10136) );
  XNOR U10198 ( .A(n10155), .B(n10148), .Z(n10154) );
  XOR U10199 ( .A(n10156), .B(n10157), .Z(n10148) );
  XNOR U10200 ( .A(n10158), .B(n10159), .Z(n10157) );
  NAND U10201 ( .A(n9673), .B(n9782), .Z(n10159) );
  XNOR U10202 ( .A(n10160), .B(n10161), .Z(n10153) );
  ANDN U10203 ( .B(n10162), .A(n9667), .Z(n10160) );
  ANDN U10204 ( .B(n10120), .A(n10123), .Z(n10143) );
  XOR U10205 ( .A(n10123), .B(n10120), .Z(n10135) );
  XNOR U10206 ( .A(n10163), .B(n10164), .Z(n10120) );
  XNOR U10207 ( .A(n10156), .B(n10165), .Z(n10164) );
  XNOR U10208 ( .A(n10155), .B(n9776), .Z(n10165) );
  XNOR U10209 ( .A(n10166), .B(n10167), .Z(n10163) );
  XNOR U10210 ( .A(n10168), .B(n10152), .Z(n10167) );
  OR U10211 ( .A(n9778), .B(n10109), .Z(n10152) );
  XNOR U10212 ( .A(n10166), .B(n10149), .Z(n10109) );
  XNOR U10213 ( .A(n9776), .B(n9773), .Z(n9778) );
  ANDN U10214 ( .B(n9773), .A(n10110), .Z(n10168) );
  XOR U10215 ( .A(n10169), .B(n10170), .Z(n10123) );
  XOR U10216 ( .A(n10156), .B(n10146), .Z(n10170) );
  XOR U10217 ( .A(n10113), .B(n9603), .Z(n10146) );
  XOR U10218 ( .A(n10171), .B(n10158), .Z(n10156) );
  NANDN U10219 ( .A(n10116), .B(n9785), .Z(n10158) );
  XOR U10220 ( .A(n9786), .B(n9782), .Z(n9785) );
  XNOR U10221 ( .A(n10162), .B(n10172), .Z(n9773) );
  XOR U10222 ( .A(n10173), .B(n10174), .Z(n10172) );
  XNOR U10223 ( .A(n10124), .B(n9673), .Z(n10116) );
  XNOR U10224 ( .A(n10110), .B(n10113), .Z(n9673) );
  IV U10225 ( .A(n10149), .Z(n10110) );
  XOR U10226 ( .A(n10175), .B(n10176), .Z(n10149) );
  XOR U10227 ( .A(n10177), .B(n10178), .Z(n10176) );
  XOR U10228 ( .A(n10166), .B(n10179), .Z(n10175) );
  AND U10229 ( .A(n9786), .B(n10124), .Z(n10171) );
  XOR U10230 ( .A(n10162), .B(n9776), .Z(n9786) );
  XNOR U10231 ( .A(n10180), .B(n10181), .Z(n9776) );
  XOR U10232 ( .A(n10182), .B(n10178), .Z(n10181) );
  XNOR U10233 ( .A(n10183), .B(n9278), .Z(n10178) );
  XOR U10234 ( .A(n10184), .B(n10185), .Z(n9278) );
  XNOR U10235 ( .A(n10186), .B(n10187), .Z(n10185) );
  XNOR U10236 ( .A(n10188), .B(n9267), .Z(n10184) );
  XOR U10237 ( .A(n10189), .B(n10190), .Z(n10183) );
  XNOR U10238 ( .A(key[188]), .B(n10191), .Z(n10190) );
  IV U10239 ( .A(n9768), .Z(n10162) );
  XOR U10240 ( .A(n10155), .B(n10192), .Z(n10169) );
  XNOR U10241 ( .A(n10193), .B(n10161), .Z(n10192) );
  OR U10242 ( .A(n9767), .B(n10114), .Z(n10161) );
  XNOR U10243 ( .A(n10194), .B(n10113), .Z(n10114) );
  XNOR U10244 ( .A(n9768), .B(n9603), .Z(n9767) );
  ANDN U10245 ( .B(n10113), .A(n9603), .Z(n10193) );
  XOR U10246 ( .A(n10180), .B(n10195), .Z(n9603) );
  XOR U10247 ( .A(n10182), .B(n10180), .Z(n10113) );
  XNOR U10248 ( .A(n9667), .B(n9768), .Z(n10155) );
  XOR U10249 ( .A(n10180), .B(n10196), .Z(n9768) );
  XNOR U10250 ( .A(n10182), .B(n10177), .Z(n10196) );
  XOR U10251 ( .A(n10197), .B(n10198), .Z(n10177) );
  XNOR U10252 ( .A(n10199), .B(n9275), .Z(n10198) );
  XOR U10253 ( .A(n10200), .B(n10201), .Z(n9275) );
  XOR U10254 ( .A(key[191]), .B(n10202), .Z(n10197) );
  XNOR U10255 ( .A(n10203), .B(n10204), .Z(n10180) );
  XNOR U10256 ( .A(n10205), .B(n9268), .Z(n10204) );
  XOR U10257 ( .A(n10206), .B(n10207), .Z(n9268) );
  XNOR U10258 ( .A(n9264), .B(n10208), .Z(n10203) );
  XNOR U10259 ( .A(key[189]), .B(n10209), .Z(n10208) );
  XOR U10260 ( .A(n9597), .B(n9667), .Z(n10124) );
  IV U10261 ( .A(n10194), .Z(n9667) );
  XNOR U10262 ( .A(n10174), .B(n10210), .Z(n10194) );
  XOR U10263 ( .A(n10211), .B(n10212), .Z(n10182) );
  XNOR U10264 ( .A(n10166), .B(n9261), .Z(n10212) );
  XNOR U10265 ( .A(n10213), .B(n9274), .Z(n9261) );
  XNOR U10266 ( .A(n10214), .B(n10215), .Z(n9274) );
  XOR U10267 ( .A(n10216), .B(n10217), .Z(n10211) );
  XNOR U10268 ( .A(key[190]), .B(n10218), .Z(n10217) );
  XOR U10269 ( .A(n10219), .B(n10220), .Z(n10179) );
  XNOR U10270 ( .A(n9286), .B(n10221), .Z(n10220) );
  XNOR U10271 ( .A(n10222), .B(n10173), .Z(n10221) );
  XNOR U10272 ( .A(n10223), .B(n10224), .Z(n10173) );
  XOR U10273 ( .A(n10225), .B(n9290), .Z(n10224) );
  XOR U10274 ( .A(n9252), .B(n10226), .Z(n10223) );
  XOR U10275 ( .A(key[185]), .B(n10227), .Z(n10226) );
  XOR U10276 ( .A(n10214), .B(n9281), .Z(n9286) );
  XNOR U10277 ( .A(n10228), .B(n10229), .Z(n10219) );
  XNOR U10278 ( .A(key[187]), .B(n10230), .Z(n10229) );
  XOR U10279 ( .A(n10231), .B(n10232), .Z(n10174) );
  XOR U10280 ( .A(n10233), .B(n9253), .Z(n10232) );
  XNOR U10281 ( .A(n10234), .B(n10235), .Z(n10231) );
  XNOR U10282 ( .A(key[186]), .B(n9294), .Z(n10235) );
  IV U10283 ( .A(n10166), .Z(n9597) );
  XOR U10284 ( .A(n10236), .B(n10237), .Z(n10166) );
  XOR U10285 ( .A(n10238), .B(n10239), .Z(n10237) );
  XOR U10286 ( .A(n10240), .B(n10241), .Z(n10236) );
  XOR U10287 ( .A(key[184]), .B(n10242), .Z(n10241) );
  XNOR U10288 ( .A(n9586), .B(n9701), .Z(n6287) );
  XNOR U10289 ( .A(n9654), .B(n10243), .Z(n9701) );
  XOR U10290 ( .A(n10244), .B(n9608), .Z(n10243) );
  OR U10291 ( .A(n10245), .B(n9751), .Z(n9608) );
  XNOR U10292 ( .A(n9610), .B(n9746), .Z(n9751) );
  NOR U10293 ( .A(n10246), .B(n9746), .Z(n10244) );
  XOR U10294 ( .A(n9654), .B(n10247), .Z(n9586) );
  XNOR U10295 ( .A(n9651), .B(n10248), .Z(n10247) );
  NAND U10296 ( .A(n10249), .B(n9616), .Z(n10248) );
  NANDN U10297 ( .A(n10250), .B(n9741), .Z(n9651) );
  XOR U10298 ( .A(n9652), .B(n9616), .Z(n9741) );
  XOR U10299 ( .A(n10251), .B(n9656), .Z(n9654) );
  OR U10300 ( .A(n9758), .B(n10252), .Z(n9656) );
  XNOR U10301 ( .A(n10253), .B(n9658), .Z(n9758) );
  XNOR U10302 ( .A(n9746), .B(n9616), .Z(n9658) );
  XOR U10303 ( .A(n10254), .B(n10255), .Z(n9616) );
  NANDN U10304 ( .A(n10256), .B(n10257), .Z(n10255) );
  XNOR U10305 ( .A(n10258), .B(n10259), .Z(n9746) );
  OR U10306 ( .A(n10256), .B(n10260), .Z(n10259) );
  ANDN U10307 ( .B(n10253), .A(n10261), .Z(n10251) );
  IV U10308 ( .A(n9761), .Z(n10253) );
  XOR U10309 ( .A(n9610), .B(n9652), .Z(n9761) );
  XNOR U10310 ( .A(n10262), .B(n10254), .Z(n9652) );
  NANDN U10311 ( .A(n10263), .B(n10264), .Z(n10254) );
  ANDN U10312 ( .B(n10265), .A(n10266), .Z(n10262) );
  NANDN U10313 ( .A(n10263), .B(n10268), .Z(n10258) );
  XOR U10314 ( .A(n10269), .B(n10256), .Z(n10263) );
  XNOR U10315 ( .A(n10270), .B(n10271), .Z(n10256) );
  XOR U10316 ( .A(n10272), .B(n10265), .Z(n10271) );
  XNOR U10317 ( .A(n10273), .B(n10274), .Z(n10270) );
  XNOR U10318 ( .A(n10275), .B(n10276), .Z(n10274) );
  ANDN U10319 ( .B(n10265), .A(n10277), .Z(n10275) );
  IV U10320 ( .A(n10278), .Z(n10265) );
  ANDN U10321 ( .B(n10269), .A(n10277), .Z(n10267) );
  IV U10322 ( .A(n10273), .Z(n10277) );
  IV U10323 ( .A(n10266), .Z(n10269) );
  XNOR U10324 ( .A(n10272), .B(n10279), .Z(n10266) );
  XOR U10325 ( .A(n10280), .B(n10276), .Z(n10279) );
  NAND U10326 ( .A(n10268), .B(n10264), .Z(n10276) );
  XNOR U10327 ( .A(n10257), .B(n10278), .Z(n10264) );
  XOR U10328 ( .A(n10281), .B(n10282), .Z(n10278) );
  XOR U10329 ( .A(n10283), .B(n10284), .Z(n10282) );
  XNOR U10330 ( .A(n9747), .B(n10285), .Z(n10284) );
  XNOR U10331 ( .A(n10286), .B(n10287), .Z(n10281) );
  XNOR U10332 ( .A(n10288), .B(n10289), .Z(n10287) );
  ANDN U10333 ( .B(n10290), .A(n9611), .Z(n10288) );
  XNOR U10334 ( .A(n10273), .B(n10260), .Z(n10268) );
  XOR U10335 ( .A(n10291), .B(n10292), .Z(n10273) );
  XNOR U10336 ( .A(n10293), .B(n10285), .Z(n10292) );
  XOR U10337 ( .A(n10294), .B(n10295), .Z(n10285) );
  XNOR U10338 ( .A(n10296), .B(n10297), .Z(n10295) );
  NAND U10339 ( .A(n9659), .B(n9756), .Z(n10297) );
  XNOR U10340 ( .A(n10298), .B(n10299), .Z(n10291) );
  ANDN U10341 ( .B(n10300), .A(n9653), .Z(n10298) );
  ANDN U10342 ( .B(n10257), .A(n10260), .Z(n10280) );
  XOR U10343 ( .A(n10260), .B(n10257), .Z(n10272) );
  XNOR U10344 ( .A(n10301), .B(n10302), .Z(n10257) );
  XNOR U10345 ( .A(n10294), .B(n10303), .Z(n10302) );
  XOR U10346 ( .A(n10293), .B(n9750), .Z(n10303) );
  XOR U10347 ( .A(n9611), .B(n10304), .Z(n10301) );
  XNOR U10348 ( .A(n10305), .B(n10289), .Z(n10304) );
  OR U10349 ( .A(n9752), .B(n10245), .Z(n10289) );
  XNOR U10350 ( .A(n9611), .B(n10246), .Z(n10245) );
  XOR U10351 ( .A(n9750), .B(n9747), .Z(n9752) );
  ANDN U10352 ( .B(n9747), .A(n10246), .Z(n10305) );
  XOR U10353 ( .A(n10306), .B(n10307), .Z(n10260) );
  XOR U10354 ( .A(n10294), .B(n10283), .Z(n10307) );
  XOR U10355 ( .A(n10249), .B(n9617), .Z(n10283) );
  XOR U10356 ( .A(n10308), .B(n10296), .Z(n10294) );
  NANDN U10357 ( .A(n10252), .B(n9759), .Z(n10296) );
  XOR U10358 ( .A(n9760), .B(n9756), .Z(n9759) );
  XNOR U10359 ( .A(n10300), .B(n10309), .Z(n9747) );
  XOR U10360 ( .A(n10310), .B(n10311), .Z(n10309) );
  XOR U10361 ( .A(n10261), .B(n9659), .Z(n10252) );
  XNOR U10362 ( .A(n10246), .B(n10249), .Z(n9659) );
  IV U10363 ( .A(n10286), .Z(n10246) );
  XOR U10364 ( .A(n10312), .B(n10313), .Z(n10286) );
  XOR U10365 ( .A(n10314), .B(n10315), .Z(n10313) );
  XNOR U10366 ( .A(n9611), .B(n10316), .Z(n10312) );
  ANDN U10367 ( .B(n9760), .A(n10261), .Z(n10308) );
  XNOR U10368 ( .A(n9611), .B(n9653), .Z(n10261) );
  XOR U10369 ( .A(n10300), .B(n10290), .Z(n9760) );
  IV U10370 ( .A(n9750), .Z(n10290) );
  XOR U10371 ( .A(n10317), .B(n10318), .Z(n9750) );
  XOR U10372 ( .A(n10319), .B(n10315), .Z(n10318) );
  XNOR U10373 ( .A(n10320), .B(n10321), .Z(n10315) );
  XNOR U10374 ( .A(n10322), .B(n9431), .Z(n10321) );
  XOR U10375 ( .A(n10323), .B(n10324), .Z(n9431) );
  XNOR U10376 ( .A(n10325), .B(n10326), .Z(n10320) );
  XOR U10377 ( .A(key[196]), .B(n10327), .Z(n10326) );
  IV U10378 ( .A(n9742), .Z(n10300) );
  XOR U10379 ( .A(n10293), .B(n10328), .Z(n10306) );
  XNOR U10380 ( .A(n10329), .B(n10299), .Z(n10328) );
  OR U10381 ( .A(n9740), .B(n10250), .Z(n10299) );
  XNOR U10382 ( .A(n10330), .B(n10249), .Z(n10250) );
  XNOR U10383 ( .A(n9742), .B(n9617), .Z(n9740) );
  ANDN U10384 ( .B(n10249), .A(n9617), .Z(n10329) );
  XOR U10385 ( .A(n10317), .B(n10331), .Z(n9617) );
  XNOR U10386 ( .A(n10332), .B(n10319), .Z(n10331) );
  XOR U10387 ( .A(n10319), .B(n10317), .Z(n10249) );
  XNOR U10388 ( .A(n9653), .B(n9742), .Z(n10293) );
  XOR U10389 ( .A(n10317), .B(n10333), .Z(n9742) );
  XNOR U10390 ( .A(n10319), .B(n10314), .Z(n10333) );
  XOR U10391 ( .A(n10334), .B(n10335), .Z(n10314) );
  XNOR U10392 ( .A(n10336), .B(n10337), .Z(n10335) );
  XOR U10393 ( .A(key[199]), .B(n10323), .Z(n10334) );
  XNOR U10394 ( .A(n10338), .B(n10339), .Z(n10317) );
  XOR U10395 ( .A(n10340), .B(n10341), .Z(n10339) );
  XNOR U10396 ( .A(key[197]), .B(n10342), .Z(n10338) );
  IV U10397 ( .A(n10330), .Z(n9653) );
  XNOR U10398 ( .A(n10311), .B(n10343), .Z(n10330) );
  XOR U10399 ( .A(n10344), .B(n10345), .Z(n10319) );
  XOR U10400 ( .A(n9611), .B(n9410), .Z(n10345) );
  XOR U10401 ( .A(n9456), .B(n10346), .Z(n9410) );
  IV U10402 ( .A(n10323), .Z(n9456) );
  XNOR U10403 ( .A(n10347), .B(n10348), .Z(n9611) );
  XOR U10404 ( .A(n10349), .B(n9453), .Z(n10348) );
  XNOR U10405 ( .A(key[192]), .B(n10350), .Z(n10347) );
  XOR U10406 ( .A(n10351), .B(n10352), .Z(n10344) );
  XNOR U10407 ( .A(key[198]), .B(n10353), .Z(n10352) );
  XOR U10408 ( .A(n10354), .B(n10355), .Z(n10316) );
  XOR U10409 ( .A(n9439), .B(n10356), .Z(n10355) );
  XOR U10410 ( .A(n10357), .B(n10332), .Z(n10356) );
  IV U10411 ( .A(n10310), .Z(n10332) );
  XNOR U10412 ( .A(n10358), .B(n10359), .Z(n10310) );
  XNOR U10413 ( .A(n10360), .B(n9400), .Z(n10359) );
  XOR U10414 ( .A(key[193]), .B(n10361), .Z(n10358) );
  XOR U10415 ( .A(n10323), .B(n10362), .Z(n9439) );
  XOR U10416 ( .A(n10363), .B(n10364), .Z(n10354) );
  XNOR U10417 ( .A(key[195]), .B(n10365), .Z(n10364) );
  XOR U10418 ( .A(n10366), .B(n10367), .Z(n10311) );
  XNOR U10419 ( .A(n10368), .B(n10369), .Z(n10367) );
  XOR U10420 ( .A(key[194]), .B(n10370), .Z(n10366) );
  XOR U10421 ( .A(n10371), .B(n10372), .Z(n5188) );
  XNOR U10422 ( .A(n10373), .B(n8444), .Z(n10372) );
  XNOR U10423 ( .A(n10374), .B(n10375), .Z(n8444) );
  XNOR U10424 ( .A(n10376), .B(n10377), .Z(n10375) );
  OR U10425 ( .A(n8449), .B(n10378), .Z(n10377) );
  XNOR U10426 ( .A(n8430), .B(n10379), .Z(n10371) );
  XOR U10427 ( .A(n10380), .B(n10381), .Z(n10379) );
  ANDN U10428 ( .B(n8456), .A(n10382), .Z(n10381) );
  XNOR U10429 ( .A(n10374), .B(n10383), .Z(n8430) );
  XNOR U10430 ( .A(n10384), .B(n8453), .Z(n10383) );
  ANDN U10431 ( .B(n10387), .A(n10388), .Z(n10384) );
  XNOR U10432 ( .A(n8451), .B(n10389), .Z(n10374) );
  XNOR U10433 ( .A(n10390), .B(n10391), .Z(n10389) );
  NANDN U10434 ( .A(n10392), .B(n10393), .Z(n10391) );
  XNOR U10435 ( .A(key[453]), .B(n5191), .Z(n8529) );
  XNOR U10436 ( .A(n3947), .B(n3954), .Z(n5191) );
  XOR U10437 ( .A(n8438), .B(n8373), .Z(n3954) );
  XNOR U10438 ( .A(n8445), .B(n10394), .Z(n8373) );
  XNOR U10439 ( .A(n10395), .B(n10380), .Z(n10394) );
  ANDN U10440 ( .B(n10386), .A(n10396), .Z(n10380) );
  XOR U10441 ( .A(n10387), .B(n8456), .Z(n10386) );
  ANDN U10442 ( .B(n10387), .A(n10397), .Z(n10395) );
  XNOR U10443 ( .A(n10373), .B(n10398), .Z(n8445) );
  XNOR U10444 ( .A(n10399), .B(n10400), .Z(n10398) );
  NANDN U10445 ( .A(n10392), .B(n10401), .Z(n10400) );
  XOR U10446 ( .A(n8431), .B(n8376), .Z(n8438) );
  XNOR U10447 ( .A(n10373), .B(n10402), .Z(n8376) );
  XNOR U10448 ( .A(n8447), .B(n10403), .Z(n10402) );
  NANDN U10449 ( .A(n10404), .B(n10405), .Z(n10403) );
  OR U10450 ( .A(n10406), .B(n10407), .Z(n8447) );
  XOR U10451 ( .A(n10408), .B(n10399), .Z(n10373) );
  NANDN U10452 ( .A(n10409), .B(n10410), .Z(n10399) );
  ANDN U10453 ( .B(n10411), .A(n10412), .Z(n10408) );
  XNOR U10454 ( .A(n8451), .B(n10413), .Z(n8431) );
  XOR U10455 ( .A(n10414), .B(n10376), .Z(n10413) );
  OR U10456 ( .A(n10415), .B(n10406), .Z(n10376) );
  XNOR U10457 ( .A(n8449), .B(n10404), .Z(n10406) );
  NOR U10458 ( .A(n10416), .B(n10404), .Z(n10414) );
  XOR U10459 ( .A(n10417), .B(n10390), .Z(n8451) );
  OR U10460 ( .A(n10409), .B(n10418), .Z(n10390) );
  XOR U10461 ( .A(n10419), .B(n10392), .Z(n10409) );
  XOR U10462 ( .A(n10404), .B(n8456), .Z(n10392) );
  XOR U10463 ( .A(n10420), .B(n10421), .Z(n8456) );
  NANDN U10464 ( .A(n10422), .B(n10423), .Z(n10421) );
  XNOR U10465 ( .A(n10424), .B(n10425), .Z(n10404) );
  OR U10466 ( .A(n10422), .B(n10426), .Z(n10425) );
  ANDN U10467 ( .B(n10419), .A(n10427), .Z(n10417) );
  IV U10468 ( .A(n10412), .Z(n10419) );
  XOR U10469 ( .A(n8449), .B(n10387), .Z(n10412) );
  XNOR U10470 ( .A(n10428), .B(n10420), .Z(n10387) );
  NANDN U10471 ( .A(n10429), .B(n10430), .Z(n10420) );
  ANDN U10472 ( .B(n10431), .A(n10432), .Z(n10428) );
  NANDN U10473 ( .A(n10429), .B(n10434), .Z(n10424) );
  XOR U10474 ( .A(n10435), .B(n10422), .Z(n10429) );
  XNOR U10475 ( .A(n10436), .B(n10437), .Z(n10422) );
  XOR U10476 ( .A(n10438), .B(n10431), .Z(n10437) );
  XNOR U10477 ( .A(n10439), .B(n10440), .Z(n10436) );
  XNOR U10478 ( .A(n10441), .B(n10442), .Z(n10440) );
  ANDN U10479 ( .B(n10431), .A(n10443), .Z(n10441) );
  IV U10480 ( .A(n10444), .Z(n10431) );
  ANDN U10481 ( .B(n10435), .A(n10443), .Z(n10433) );
  IV U10482 ( .A(n10439), .Z(n10443) );
  IV U10483 ( .A(n10432), .Z(n10435) );
  XNOR U10484 ( .A(n10438), .B(n10445), .Z(n10432) );
  XOR U10485 ( .A(n10446), .B(n10442), .Z(n10445) );
  NAND U10486 ( .A(n10434), .B(n10430), .Z(n10442) );
  XNOR U10487 ( .A(n10423), .B(n10444), .Z(n10430) );
  XOR U10488 ( .A(n10447), .B(n10448), .Z(n10444) );
  XOR U10489 ( .A(n10449), .B(n10450), .Z(n10448) );
  XNOR U10490 ( .A(n10405), .B(n10451), .Z(n10450) );
  XNOR U10491 ( .A(n10452), .B(n10453), .Z(n10447) );
  XNOR U10492 ( .A(n10454), .B(n10455), .Z(n10453) );
  ANDN U10493 ( .B(n10456), .A(n10378), .Z(n10454) );
  XNOR U10494 ( .A(n10439), .B(n10426), .Z(n10434) );
  XOR U10495 ( .A(n10457), .B(n10458), .Z(n10439) );
  XNOR U10496 ( .A(n10459), .B(n10451), .Z(n10458) );
  XOR U10497 ( .A(n10460), .B(n10461), .Z(n10451) );
  XNOR U10498 ( .A(n10462), .B(n10463), .Z(n10461) );
  NAND U10499 ( .A(n10393), .B(n10401), .Z(n10463) );
  XNOR U10500 ( .A(n10464), .B(n10465), .Z(n10457) );
  ANDN U10501 ( .B(n10466), .A(n10388), .Z(n10464) );
  ANDN U10502 ( .B(n10423), .A(n10426), .Z(n10446) );
  XOR U10503 ( .A(n10426), .B(n10423), .Z(n10438) );
  XNOR U10504 ( .A(n10467), .B(n10468), .Z(n10423) );
  XNOR U10505 ( .A(n10460), .B(n10469), .Z(n10468) );
  XOR U10506 ( .A(n10459), .B(n8450), .Z(n10469) );
  XOR U10507 ( .A(n10378), .B(n10470), .Z(n10467) );
  XNOR U10508 ( .A(n10471), .B(n10455), .Z(n10470) );
  OR U10509 ( .A(n10407), .B(n10415), .Z(n10455) );
  XNOR U10510 ( .A(n10378), .B(n10416), .Z(n10415) );
  XOR U10511 ( .A(n8450), .B(n10405), .Z(n10407) );
  ANDN U10512 ( .B(n10405), .A(n10416), .Z(n10471) );
  XOR U10513 ( .A(n10472), .B(n10473), .Z(n10426) );
  XOR U10514 ( .A(n10460), .B(n10449), .Z(n10473) );
  XOR U10515 ( .A(n8455), .B(n10382), .Z(n10449) );
  XOR U10516 ( .A(n10474), .B(n10462), .Z(n10460) );
  NANDN U10517 ( .A(n10418), .B(n10410), .Z(n10462) );
  XOR U10518 ( .A(n10411), .B(n10401), .Z(n10410) );
  XNOR U10519 ( .A(n10466), .B(n10475), .Z(n10405) );
  XOR U10520 ( .A(n10476), .B(n10477), .Z(n10475) );
  XOR U10521 ( .A(n10427), .B(n10393), .Z(n10418) );
  XNOR U10522 ( .A(n10416), .B(n8455), .Z(n10393) );
  IV U10523 ( .A(n10452), .Z(n10416) );
  XOR U10524 ( .A(n10478), .B(n10479), .Z(n10452) );
  XOR U10525 ( .A(n10480), .B(n10481), .Z(n10479) );
  XNOR U10526 ( .A(n10378), .B(n10482), .Z(n10478) );
  ANDN U10527 ( .B(n10411), .A(n10427), .Z(n10474) );
  XNOR U10528 ( .A(n10378), .B(n10388), .Z(n10427) );
  XOR U10529 ( .A(n10466), .B(n10456), .Z(n10411) );
  IV U10530 ( .A(n8450), .Z(n10456) );
  XOR U10531 ( .A(n10483), .B(n10484), .Z(n8450) );
  XOR U10532 ( .A(n10485), .B(n10481), .Z(n10484) );
  XNOR U10533 ( .A(n10486), .B(n10487), .Z(n10481) );
  XNOR U10534 ( .A(n7917), .B(n5924), .Z(n10487) );
  XNOR U10535 ( .A(n10488), .B(n7301), .Z(n5924) );
  XOR U10536 ( .A(n5927), .B(n7315), .Z(n7917) );
  XOR U10537 ( .A(n10489), .B(n5972), .Z(n5927) );
  XNOR U10538 ( .A(n7916), .B(n10490), .Z(n10486) );
  XNOR U10539 ( .A(key[348]), .B(n7316), .Z(n10490) );
  XOR U10540 ( .A(n10491), .B(n7950), .Z(n7316) );
  XOR U10541 ( .A(n5951), .B(n7305), .Z(n7916) );
  IV U10542 ( .A(n7932), .Z(n7305) );
  XOR U10543 ( .A(n10492), .B(n10493), .Z(n7932) );
  XNOR U10544 ( .A(n10494), .B(n10495), .Z(n10493) );
  XNOR U10545 ( .A(n10496), .B(n10497), .Z(n10492) );
  XOR U10546 ( .A(n10498), .B(n10499), .Z(n10497) );
  ANDN U10547 ( .B(n10500), .A(n10501), .Z(n10499) );
  IV U10548 ( .A(n10397), .Z(n10466) );
  XOR U10549 ( .A(n10459), .B(n10502), .Z(n10472) );
  XNOR U10550 ( .A(n10503), .B(n10465), .Z(n10502) );
  OR U10551 ( .A(n10396), .B(n10385), .Z(n10465) );
  XNOR U10552 ( .A(n10504), .B(n8455), .Z(n10385) );
  XNOR U10553 ( .A(n10397), .B(n10382), .Z(n10396) );
  ANDN U10554 ( .B(n8455), .A(n10382), .Z(n10503) );
  XOR U10555 ( .A(n10483), .B(n10505), .Z(n10382) );
  XNOR U10556 ( .A(n10506), .B(n10485), .Z(n10505) );
  XOR U10557 ( .A(n10485), .B(n10483), .Z(n8455) );
  XNOR U10558 ( .A(n10388), .B(n10397), .Z(n10459) );
  XOR U10559 ( .A(n10483), .B(n10507), .Z(n10397) );
  XNOR U10560 ( .A(n10485), .B(n10480), .Z(n10507) );
  XOR U10561 ( .A(n10508), .B(n10509), .Z(n10480) );
  XNOR U10562 ( .A(n7311), .B(n7929), .Z(n10509) );
  XNOR U10563 ( .A(n7296), .B(n7310), .Z(n7929) );
  XOR U10564 ( .A(n10510), .B(n10511), .Z(n7296) );
  XNOR U10565 ( .A(n10512), .B(n10513), .Z(n10511) );
  XOR U10566 ( .A(n10514), .B(n10515), .Z(n10510) );
  XNOR U10567 ( .A(n10516), .B(n10517), .Z(n7311) );
  XOR U10568 ( .A(n10518), .B(n10519), .Z(n10517) );
  XOR U10569 ( .A(n10520), .B(n10521), .Z(n10516) );
  XNOR U10570 ( .A(key[351]), .B(n7335), .Z(n10508) );
  XOR U10571 ( .A(n5951), .B(n5937), .Z(n7335) );
  XNOR U10572 ( .A(n10522), .B(n10523), .Z(n10483) );
  XNOR U10573 ( .A(n7304), .B(n7933), .Z(n10523) );
  XOR U10574 ( .A(n5942), .B(n7301), .Z(n7933) );
  XNOR U10575 ( .A(n10524), .B(n10525), .Z(n7301) );
  XNOR U10576 ( .A(n10526), .B(n10527), .Z(n10525) );
  XOR U10577 ( .A(n10528), .B(n10529), .Z(n10524) );
  XOR U10578 ( .A(n10530), .B(n10531), .Z(n10529) );
  ANDN U10579 ( .B(n10532), .A(n10533), .Z(n10531) );
  XOR U10580 ( .A(n10534), .B(n10535), .Z(n5942) );
  XNOR U10581 ( .A(n10489), .B(n10513), .Z(n10535) );
  XNOR U10582 ( .A(n10536), .B(n10537), .Z(n10513) );
  XNOR U10583 ( .A(n10538), .B(n10539), .Z(n10537) );
  OR U10584 ( .A(n10540), .B(n10541), .Z(n10539) );
  XNOR U10585 ( .A(n10542), .B(n10543), .Z(n10534) );
  XNOR U10586 ( .A(n10544), .B(n10545), .Z(n10543) );
  ANDN U10587 ( .B(n10546), .A(n10547), .Z(n10545) );
  XOR U10588 ( .A(n10548), .B(n10549), .Z(n7304) );
  XNOR U10589 ( .A(n10550), .B(n10519), .Z(n10549) );
  XNOR U10590 ( .A(n10551), .B(n10552), .Z(n10519) );
  XNOR U10591 ( .A(n10553), .B(n10554), .Z(n10552) );
  OR U10592 ( .A(n10555), .B(n10556), .Z(n10554) );
  XNOR U10593 ( .A(n10491), .B(n10557), .Z(n10548) );
  XNOR U10594 ( .A(n10558), .B(n10559), .Z(n10557) );
  ANDN U10595 ( .B(n10560), .A(n10561), .Z(n10558) );
  XNOR U10596 ( .A(n7934), .B(n10562), .Z(n10522) );
  XOR U10597 ( .A(key[349]), .B(n7293), .Z(n10562) );
  XOR U10598 ( .A(n10563), .B(n10564), .Z(n7934) );
  IV U10599 ( .A(n10504), .Z(n10388) );
  XNOR U10600 ( .A(n10477), .B(n10565), .Z(n10504) );
  XOR U10601 ( .A(n10566), .B(n10567), .Z(n10485) );
  XOR U10602 ( .A(n10378), .B(n5946), .Z(n10567) );
  XNOR U10603 ( .A(n5937), .B(n7310), .Z(n5946) );
  XNOR U10604 ( .A(n10568), .B(n10569), .Z(n7310) );
  XOR U10605 ( .A(n10570), .B(n10527), .Z(n10569) );
  XNOR U10606 ( .A(n10571), .B(n10572), .Z(n10527) );
  XNOR U10607 ( .A(n10573), .B(n10574), .Z(n10572) );
  NANDN U10608 ( .A(n10575), .B(n10576), .Z(n10574) );
  XOR U10609 ( .A(n10577), .B(n10578), .Z(n10568) );
  IV U10610 ( .A(n10488), .Z(n5937) );
  XNOR U10611 ( .A(n10579), .B(n10580), .Z(n10378) );
  XNOR U10612 ( .A(n7327), .B(n5949), .Z(n10580) );
  XOR U10613 ( .A(n7919), .B(n7295), .Z(n5949) );
  IV U10614 ( .A(n7941), .Z(n7295) );
  XNOR U10615 ( .A(n10536), .B(n10581), .Z(n10489) );
  XNOR U10616 ( .A(n10582), .B(n10583), .Z(n10581) );
  OR U10617 ( .A(n10584), .B(n10585), .Z(n10583) );
  XNOR U10618 ( .A(n10586), .B(n10587), .Z(n10536) );
  XNOR U10619 ( .A(n10588), .B(n10589), .Z(n10587) );
  NAND U10620 ( .A(n10590), .B(n10591), .Z(n10589) );
  XOR U10621 ( .A(n10593), .B(n10491), .Z(n7919) );
  XNOR U10622 ( .A(n10551), .B(n10594), .Z(n10491) );
  XNOR U10623 ( .A(n10595), .B(n10596), .Z(n10594) );
  ANDN U10624 ( .B(n10597), .A(n10598), .Z(n10595) );
  XNOR U10625 ( .A(n10599), .B(n10600), .Z(n10551) );
  XNOR U10626 ( .A(n10601), .B(n10602), .Z(n10600) );
  NANDN U10627 ( .A(n10603), .B(n10604), .Z(n10602) );
  XOR U10628 ( .A(n7942), .B(n10605), .Z(n10579) );
  XNOR U10629 ( .A(key[344]), .B(n10488), .Z(n10605) );
  IV U10630 ( .A(n7952), .Z(n7942) );
  XOR U10631 ( .A(n10606), .B(n10607), .Z(n7952) );
  XNOR U10632 ( .A(n10608), .B(n10563), .Z(n10607) );
  XOR U10633 ( .A(n7938), .B(n10609), .Z(n10566) );
  XNOR U10634 ( .A(key[350]), .B(n7303), .Z(n10609) );
  XNOR U10635 ( .A(n10610), .B(n10611), .Z(n7303) );
  XOR U10636 ( .A(n10593), .B(n10612), .Z(n10611) );
  XOR U10637 ( .A(n5941), .B(n7928), .Z(n7938) );
  XOR U10638 ( .A(n5951), .B(n7312), .Z(n7928) );
  XNOR U10639 ( .A(n10613), .B(n10614), .Z(n7312) );
  XOR U10640 ( .A(n10606), .B(n10495), .Z(n10614) );
  XNOR U10641 ( .A(n10615), .B(n10616), .Z(n10495) );
  XNOR U10642 ( .A(n10617), .B(n10618), .Z(n10616) );
  NANDN U10643 ( .A(n10619), .B(n10620), .Z(n10618) );
  XOR U10644 ( .A(n10608), .B(n10563), .Z(n10613) );
  XOR U10645 ( .A(n10621), .B(n10622), .Z(n10563) );
  XNOR U10646 ( .A(n7293), .B(n5952), .Z(n5941) );
  XOR U10647 ( .A(n10623), .B(n10512), .Z(n5952) );
  XNOR U10648 ( .A(n10578), .B(n10624), .Z(n7293) );
  XOR U10649 ( .A(n10625), .B(n10626), .Z(n10482) );
  XNOR U10650 ( .A(n5959), .B(n10627), .Z(n10626) );
  XNOR U10651 ( .A(n5971), .B(n10506), .Z(n10627) );
  IV U10652 ( .A(n10476), .Z(n10506) );
  XNOR U10653 ( .A(n10628), .B(n10629), .Z(n10476) );
  XOR U10654 ( .A(n7284), .B(n5950), .Z(n10629) );
  XOR U10655 ( .A(n5964), .B(n7327), .Z(n5950) );
  XNOR U10656 ( .A(n10570), .B(n10630), .Z(n7327) );
  XNOR U10657 ( .A(n10577), .B(n10578), .Z(n10630) );
  XNOR U10658 ( .A(n10631), .B(n10632), .Z(n10578) );
  XOR U10659 ( .A(n10512), .B(n10633), .Z(n5964) );
  XOR U10660 ( .A(n10634), .B(n10515), .Z(n10633) );
  XOR U10661 ( .A(n10592), .B(n10635), .Z(n10512) );
  XOR U10662 ( .A(n7951), .B(n10636), .Z(n10628) );
  XNOR U10663 ( .A(key[345]), .B(n7334), .Z(n10636) );
  XOR U10664 ( .A(n10518), .B(n10637), .Z(n7334) );
  XNOR U10665 ( .A(n10520), .B(n10521), .Z(n10637) );
  XNOR U10666 ( .A(n10593), .B(n10612), .Z(n10521) );
  XOR U10667 ( .A(n7322), .B(n5958), .Z(n5971) );
  XNOR U10668 ( .A(n10638), .B(n10639), .Z(n5958) );
  XOR U10669 ( .A(n10635), .B(n10623), .Z(n10639) );
  XNOR U10670 ( .A(n10640), .B(n10641), .Z(n10623) );
  XOR U10671 ( .A(n10642), .B(n10544), .Z(n10641) );
  NANDN U10672 ( .A(n10643), .B(n10644), .Z(n10544) );
  NOR U10673 ( .A(n10645), .B(n10584), .Z(n10642) );
  XOR U10674 ( .A(n10542), .B(n10646), .Z(n10635) );
  XNOR U10675 ( .A(n10647), .B(n10648), .Z(n10646) );
  NANDN U10676 ( .A(n10649), .B(n10650), .Z(n10648) );
  XNOR U10677 ( .A(n10634), .B(n10515), .Z(n10638) );
  XOR U10678 ( .A(n10640), .B(n10651), .Z(n10515) );
  XOR U10679 ( .A(n10652), .B(n10647), .Z(n10651) );
  OR U10680 ( .A(n10653), .B(n10654), .Z(n10647) );
  NOR U10681 ( .A(n10655), .B(n10540), .Z(n10652) );
  XNOR U10682 ( .A(n10542), .B(n10656), .Z(n10640) );
  XNOR U10683 ( .A(n10657), .B(n10658), .Z(n10656) );
  NAND U10684 ( .A(n10659), .B(n10590), .Z(n10658) );
  XOR U10685 ( .A(n10660), .B(n10657), .Z(n10542) );
  NANDN U10686 ( .A(n10661), .B(n10662), .Z(n10657) );
  AND U10687 ( .A(n10663), .B(n10664), .Z(n10660) );
  IV U10688 ( .A(n10514), .Z(n10634) );
  XNOR U10689 ( .A(n10488), .B(n7315), .Z(n5959) );
  XNOR U10690 ( .A(n10665), .B(n7284), .Z(n7315) );
  XOR U10691 ( .A(n10528), .B(n10631), .Z(n10488) );
  IV U10692 ( .A(n10665), .Z(n10528) );
  XNOR U10693 ( .A(n10667), .B(n10668), .Z(n10666) );
  ANDN U10694 ( .B(n10669), .A(n10670), .Z(n10667) );
  XNOR U10695 ( .A(n10671), .B(n10672), .Z(n10571) );
  XNOR U10696 ( .A(n10673), .B(n10674), .Z(n10672) );
  NANDN U10697 ( .A(n10675), .B(n10676), .Z(n10674) );
  XNOR U10698 ( .A(n7947), .B(n10677), .Z(n10625) );
  XNOR U10699 ( .A(key[347]), .B(n7286), .Z(n10677) );
  XOR U10700 ( .A(n10678), .B(n10679), .Z(n7286) );
  XOR U10701 ( .A(n10518), .B(n10610), .Z(n10679) );
  XNOR U10702 ( .A(n10680), .B(n10681), .Z(n10610) );
  XNOR U10703 ( .A(n10559), .B(n10682), .Z(n10681) );
  NANDN U10704 ( .A(n10683), .B(n10597), .Z(n10682) );
  NANDN U10705 ( .A(n10684), .B(n10685), .Z(n10559) );
  XOR U10706 ( .A(n10520), .B(n10612), .Z(n10678) );
  XOR U10707 ( .A(n10550), .B(n10686), .Z(n10612) );
  XOR U10708 ( .A(n10687), .B(n10688), .Z(n10686) );
  AND U10709 ( .A(n10689), .B(n10690), .Z(n10687) );
  XNOR U10710 ( .A(n10688), .B(n10692), .Z(n10691) );
  OR U10711 ( .A(n10555), .B(n10693), .Z(n10692) );
  OR U10712 ( .A(n10694), .B(n10695), .Z(n10688) );
  XNOR U10713 ( .A(n10550), .B(n10696), .Z(n10680) );
  XNOR U10714 ( .A(n10697), .B(n10698), .Z(n10696) );
  NANDN U10715 ( .A(n10603), .B(n10699), .Z(n10698) );
  XOR U10716 ( .A(n10700), .B(n10697), .Z(n10550) );
  NANDN U10717 ( .A(n10701), .B(n10702), .Z(n10697) );
  ANDN U10718 ( .B(n10703), .A(n10704), .Z(n10700) );
  XOR U10719 ( .A(n5951), .B(n7317), .Z(n7947) );
  XNOR U10720 ( .A(n10496), .B(n7951), .Z(n7317) );
  XNOR U10721 ( .A(n10621), .B(n10606), .Z(n7951) );
  XNOR U10722 ( .A(n10496), .B(n10621), .Z(n5951) );
  XNOR U10723 ( .A(n10705), .B(n10706), .Z(n10621) );
  XOR U10724 ( .A(n10707), .B(n10617), .Z(n10706) );
  OR U10725 ( .A(n10708), .B(n10709), .Z(n10617) );
  ANDN U10726 ( .B(n10710), .A(n10711), .Z(n10707) );
  XNOR U10727 ( .A(n10615), .B(n10712), .Z(n10496) );
  XNOR U10728 ( .A(n10713), .B(n10714), .Z(n10712) );
  ANDN U10729 ( .B(n10715), .A(n10716), .Z(n10713) );
  XNOR U10730 ( .A(n10705), .B(n10717), .Z(n10615) );
  XNOR U10731 ( .A(n10718), .B(n10719), .Z(n10717) );
  NANDN U10732 ( .A(n10720), .B(n10721), .Z(n10719) );
  XOR U10733 ( .A(n10722), .B(n10723), .Z(n10477) );
  XNOR U10734 ( .A(n7322), .B(n5963), .Z(n10723) );
  XOR U10735 ( .A(n5972), .B(n7284), .Z(n5963) );
  XOR U10736 ( .A(n10631), .B(n10570), .Z(n7284) );
  XNOR U10737 ( .A(n10671), .B(n10724), .Z(n10631) );
  XOR U10738 ( .A(n10725), .B(n10573), .Z(n10724) );
  OR U10739 ( .A(n10726), .B(n10727), .Z(n10573) );
  ANDN U10740 ( .B(n10728), .A(n10729), .Z(n10725) );
  XNOR U10741 ( .A(n10514), .B(n10592), .Z(n5972) );
  XNOR U10742 ( .A(n10586), .B(n10730), .Z(n10592) );
  XOR U10743 ( .A(n10731), .B(n10538), .Z(n10730) );
  OR U10744 ( .A(n10732), .B(n10653), .Z(n10538) );
  XNOR U10745 ( .A(n10540), .B(n10649), .Z(n10653) );
  NOR U10746 ( .A(n10733), .B(n10649), .Z(n10731) );
  XOR U10747 ( .A(n10586), .B(n10734), .Z(n10514) );
  XNOR U10748 ( .A(n10582), .B(n10735), .Z(n10734) );
  NANDN U10749 ( .A(n10547), .B(n10736), .Z(n10735) );
  NANDN U10750 ( .A(n10737), .B(n10644), .Z(n10582) );
  XOR U10751 ( .A(n10584), .B(n10547), .Z(n10644) );
  XOR U10752 ( .A(n10738), .B(n10588), .Z(n10586) );
  OR U10753 ( .A(n10661), .B(n10739), .Z(n10588) );
  XNOR U10754 ( .A(n10663), .B(n10590), .Z(n10661) );
  XOR U10755 ( .A(n10649), .B(n10547), .Z(n10590) );
  XNOR U10756 ( .A(n10740), .B(n10741), .Z(n10547) );
  NANDN U10757 ( .A(n10742), .B(n10743), .Z(n10741) );
  XNOR U10758 ( .A(n10744), .B(n10745), .Z(n10649) );
  OR U10759 ( .A(n10742), .B(n10746), .Z(n10745) );
  ANDN U10760 ( .B(n10663), .A(n10747), .Z(n10738) );
  XOR U10761 ( .A(n10540), .B(n10584), .Z(n10663) );
  XNOR U10762 ( .A(n10740), .B(n10748), .Z(n10584) );
  NANDN U10763 ( .A(n10749), .B(n10750), .Z(n10748) );
  NANDN U10764 ( .A(n10751), .B(n10752), .Z(n10740) );
  OR U10765 ( .A(n10754), .B(n10751), .Z(n10744) );
  XOR U10766 ( .A(n10755), .B(n10742), .Z(n10751) );
  XNOR U10767 ( .A(n10756), .B(n10757), .Z(n10742) );
  XOR U10768 ( .A(n10758), .B(n10750), .Z(n10757) );
  XNOR U10769 ( .A(n10759), .B(n10760), .Z(n10756) );
  XNOR U10770 ( .A(n10761), .B(n10762), .Z(n10760) );
  ANDN U10771 ( .B(n10750), .A(n10763), .Z(n10761) );
  IV U10772 ( .A(n10764), .Z(n10750) );
  ANDN U10773 ( .B(n10755), .A(n10763), .Z(n10753) );
  IV U10774 ( .A(n10749), .Z(n10755) );
  XNOR U10775 ( .A(n10758), .B(n10765), .Z(n10749) );
  XNOR U10776 ( .A(n10762), .B(n10766), .Z(n10765) );
  NANDN U10777 ( .A(n10746), .B(n10743), .Z(n10766) );
  NANDN U10778 ( .A(n10754), .B(n10752), .Z(n10762) );
  XNOR U10779 ( .A(n10743), .B(n10764), .Z(n10752) );
  XOR U10780 ( .A(n10767), .B(n10768), .Z(n10764) );
  XOR U10781 ( .A(n10769), .B(n10770), .Z(n10768) );
  XNOR U10782 ( .A(n10650), .B(n10771), .Z(n10770) );
  XNOR U10783 ( .A(n10772), .B(n10773), .Z(n10767) );
  XNOR U10784 ( .A(n10774), .B(n10775), .Z(n10773) );
  ANDN U10785 ( .B(n10776), .A(n10541), .Z(n10774) );
  XNOR U10786 ( .A(n10763), .B(n10746), .Z(n10754) );
  IV U10787 ( .A(n10759), .Z(n10763) );
  XOR U10788 ( .A(n10777), .B(n10778), .Z(n10759) );
  XNOR U10789 ( .A(n10779), .B(n10771), .Z(n10778) );
  XOR U10790 ( .A(n10780), .B(n10781), .Z(n10771) );
  XNOR U10791 ( .A(n10782), .B(n10783), .Z(n10781) );
  NAND U10792 ( .A(n10591), .B(n10659), .Z(n10783) );
  XNOR U10793 ( .A(n10784), .B(n10785), .Z(n10777) );
  ANDN U10794 ( .B(n10786), .A(n10585), .Z(n10784) );
  XOR U10795 ( .A(n10746), .B(n10743), .Z(n10758) );
  XNOR U10796 ( .A(n10787), .B(n10788), .Z(n10743) );
  XNOR U10797 ( .A(n10780), .B(n10789), .Z(n10788) );
  XOR U10798 ( .A(n10779), .B(n10655), .Z(n10789) );
  XOR U10799 ( .A(n10541), .B(n10790), .Z(n10787) );
  XNOR U10800 ( .A(n10791), .B(n10775), .Z(n10790) );
  OR U10801 ( .A(n10654), .B(n10732), .Z(n10775) );
  XNOR U10802 ( .A(n10541), .B(n10733), .Z(n10732) );
  XOR U10803 ( .A(n10655), .B(n10650), .Z(n10654) );
  ANDN U10804 ( .B(n10650), .A(n10733), .Z(n10791) );
  XOR U10805 ( .A(n10792), .B(n10793), .Z(n10746) );
  XOR U10806 ( .A(n10780), .B(n10769), .Z(n10793) );
  XOR U10807 ( .A(n10794), .B(n10546), .Z(n10769) );
  XOR U10808 ( .A(n10795), .B(n10782), .Z(n10780) );
  NANDN U10809 ( .A(n10739), .B(n10662), .Z(n10782) );
  XOR U10810 ( .A(n10664), .B(n10659), .Z(n10662) );
  XOR U10811 ( .A(n10546), .B(n10650), .Z(n10659) );
  XNOR U10812 ( .A(n10786), .B(n10796), .Z(n10650) );
  XOR U10813 ( .A(n10797), .B(n10798), .Z(n10796) );
  XOR U10814 ( .A(n10747), .B(n10591), .Z(n10739) );
  XNOR U10815 ( .A(n10733), .B(n10736), .Z(n10591) );
  IV U10816 ( .A(n10772), .Z(n10733) );
  XOR U10817 ( .A(n10799), .B(n10800), .Z(n10772) );
  XOR U10818 ( .A(n10801), .B(n10802), .Z(n10800) );
  XNOR U10819 ( .A(n10541), .B(n10803), .Z(n10799) );
  ANDN U10820 ( .B(n10664), .A(n10747), .Z(n10795) );
  XNOR U10821 ( .A(n10541), .B(n10585), .Z(n10747) );
  XOR U10822 ( .A(n10786), .B(n10776), .Z(n10664) );
  IV U10823 ( .A(n10655), .Z(n10776) );
  XOR U10824 ( .A(n10804), .B(n10805), .Z(n10655) );
  XOR U10825 ( .A(n10806), .B(n10802), .Z(n10805) );
  XNOR U10826 ( .A(n10807), .B(n10808), .Z(n10802) );
  XOR U10827 ( .A(n10077), .B(n10089), .Z(n10808) );
  XOR U10828 ( .A(n10809), .B(n10810), .Z(n10089) );
  XOR U10829 ( .A(n10811), .B(n10812), .Z(n10810) );
  XNOR U10830 ( .A(n10813), .B(n8950), .Z(n10809) );
  XNOR U10831 ( .A(key[140]), .B(n10814), .Z(n10807) );
  XOR U10832 ( .A(n10779), .B(n10815), .Z(n10792) );
  XNOR U10833 ( .A(n10816), .B(n10785), .Z(n10815) );
  OR U10834 ( .A(n10643), .B(n10737), .Z(n10785) );
  XNOR U10835 ( .A(n10817), .B(n10736), .Z(n10737) );
  IV U10836 ( .A(n10794), .Z(n10736) );
  XNOR U10837 ( .A(n10786), .B(n10546), .Z(n10643) );
  IV U10838 ( .A(n10645), .Z(n10786) );
  ANDN U10839 ( .B(n10546), .A(n10794), .Z(n10816) );
  XNOR U10840 ( .A(n10818), .B(n10819), .Z(n10794) );
  XNOR U10841 ( .A(n10804), .B(n10820), .Z(n10546) );
  XNOR U10842 ( .A(n10798), .B(n10818), .Z(n10820) );
  XNOR U10843 ( .A(n10585), .B(n10645), .Z(n10779) );
  XOR U10844 ( .A(n10804), .B(n10821), .Z(n10645) );
  XNOR U10845 ( .A(n10806), .B(n10801), .Z(n10821) );
  XOR U10846 ( .A(n10822), .B(n10823), .Z(n10801) );
  XOR U10847 ( .A(n10085), .B(n8975), .Z(n10823) );
  XNOR U10848 ( .A(n10813), .B(n10824), .Z(n8975) );
  XOR U10849 ( .A(n8958), .B(n10825), .Z(n10085) );
  XNOR U10850 ( .A(key[143]), .B(n10094), .Z(n10822) );
  IV U10851 ( .A(n10819), .Z(n10804) );
  XOR U10852 ( .A(n10826), .B(n10827), .Z(n10819) );
  XNOR U10853 ( .A(n10090), .B(n10105), .Z(n10827) );
  XOR U10854 ( .A(n8963), .B(n10828), .Z(n10105) );
  XNOR U10855 ( .A(n10829), .B(n10830), .Z(n10826) );
  XNOR U10856 ( .A(key[141]), .B(n10831), .Z(n10830) );
  IV U10857 ( .A(n10817), .Z(n10585) );
  XOR U10858 ( .A(n10818), .B(n10832), .Z(n10817) );
  XNOR U10859 ( .A(n10797), .B(n10803), .Z(n10832) );
  XOR U10860 ( .A(n10833), .B(n10834), .Z(n10803) );
  XOR U10861 ( .A(n10798), .B(n10835), .Z(n10834) );
  XOR U10862 ( .A(n10078), .B(n10071), .Z(n10835) );
  XNOR U10863 ( .A(n10813), .B(n10091), .Z(n10071) );
  XNOR U10864 ( .A(n10836), .B(n10837), .Z(n10798) );
  XNOR U10865 ( .A(n8974), .B(n10838), .Z(n10837) );
  XNOR U10866 ( .A(n10839), .B(n10840), .Z(n10836) );
  XNOR U10867 ( .A(key[137]), .B(n10841), .Z(n10840) );
  XNOR U10868 ( .A(n8999), .B(n10842), .Z(n10833) );
  XNOR U10869 ( .A(key[139]), .B(n10843), .Z(n10842) );
  XOR U10870 ( .A(n10844), .B(n10845), .Z(n10797) );
  XNOR U10871 ( .A(n8985), .B(n8990), .Z(n10845) );
  XNOR U10872 ( .A(n10080), .B(n10846), .Z(n10844) );
  XNOR U10873 ( .A(key[138]), .B(n10847), .Z(n10846) );
  IV U10874 ( .A(n10806), .Z(n10818) );
  XOR U10875 ( .A(n10848), .B(n10849), .Z(n10806) );
  XNOR U10876 ( .A(n10541), .B(n10099), .Z(n10849) );
  XOR U10877 ( .A(n10850), .B(n10084), .Z(n10099) );
  XNOR U10878 ( .A(n10813), .B(n10851), .Z(n10084) );
  XNOR U10879 ( .A(n10852), .B(n10853), .Z(n10541) );
  XNOR U10880 ( .A(n10824), .B(n10074), .Z(n10853) );
  XNOR U10881 ( .A(n10854), .B(n10855), .Z(n10852) );
  XNOR U10882 ( .A(key[136]), .B(n8960), .Z(n10855) );
  XNOR U10883 ( .A(n8965), .B(n10856), .Z(n10848) );
  XNOR U10884 ( .A(key[142]), .B(n10857), .Z(n10856) );
  XOR U10885 ( .A(n10858), .B(n10859), .Z(n7322) );
  XOR U10886 ( .A(n10570), .B(n10624), .Z(n10859) );
  XNOR U10887 ( .A(n10860), .B(n10861), .Z(n10624) );
  XNOR U10888 ( .A(n10862), .B(n10530), .Z(n10861) );
  ANDN U10889 ( .B(n10863), .A(n10864), .Z(n10530) );
  ANDN U10890 ( .B(n10865), .A(n10670), .Z(n10862) );
  IV U10891 ( .A(n10866), .Z(n10670) );
  XOR U10892 ( .A(n10671), .B(n10867), .Z(n10570) );
  XOR U10893 ( .A(n10668), .B(n10868), .Z(n10867) );
  NANDN U10894 ( .A(n10869), .B(n10532), .Z(n10868) );
  XOR U10895 ( .A(n10866), .B(n10532), .Z(n10863) );
  XOR U10896 ( .A(n10871), .B(n10673), .Z(n10671) );
  OR U10897 ( .A(n10872), .B(n10873), .Z(n10673) );
  NOR U10898 ( .A(n10874), .B(n10875), .Z(n10871) );
  XOR U10899 ( .A(n10577), .B(n10632), .Z(n10858) );
  XOR U10900 ( .A(n10526), .B(n10876), .Z(n10632) );
  XNOR U10901 ( .A(n10877), .B(n10878), .Z(n10876) );
  NANDN U10902 ( .A(n10879), .B(n10728), .Z(n10878) );
  XNOR U10903 ( .A(n10877), .B(n10881), .Z(n10880) );
  NANDN U10904 ( .A(n10882), .B(n10576), .Z(n10881) );
  OR U10905 ( .A(n10727), .B(n10883), .Z(n10877) );
  XNOR U10906 ( .A(n10576), .B(n10728), .Z(n10727) );
  XNOR U10907 ( .A(n10526), .B(n10884), .Z(n10860) );
  XNOR U10908 ( .A(n10885), .B(n10886), .Z(n10884) );
  NANDN U10909 ( .A(n10675), .B(n10887), .Z(n10886) );
  XOR U10910 ( .A(n10888), .B(n10885), .Z(n10526) );
  NANDN U10911 ( .A(n10872), .B(n10889), .Z(n10885) );
  XNOR U10912 ( .A(n10874), .B(n10675), .Z(n10872) );
  XNOR U10913 ( .A(n10728), .B(n10532), .Z(n10675) );
  XOR U10914 ( .A(n10890), .B(n10891), .Z(n10532) );
  NANDN U10915 ( .A(n10892), .B(n10893), .Z(n10891) );
  XOR U10916 ( .A(n10894), .B(n10895), .Z(n10728) );
  NANDN U10917 ( .A(n10892), .B(n10896), .Z(n10895) );
  ANDN U10918 ( .B(n10897), .A(n10874), .Z(n10888) );
  XNOR U10919 ( .A(n10866), .B(n10576), .Z(n10874) );
  XNOR U10920 ( .A(n10898), .B(n10894), .Z(n10576) );
  NANDN U10921 ( .A(n10899), .B(n10900), .Z(n10894) );
  XOR U10922 ( .A(n10896), .B(n10901), .Z(n10900) );
  ANDN U10923 ( .B(n10901), .A(n10902), .Z(n10898) );
  XNOR U10924 ( .A(n10903), .B(n10890), .Z(n10866) );
  NANDN U10925 ( .A(n10899), .B(n10904), .Z(n10890) );
  XOR U10926 ( .A(n10905), .B(n10893), .Z(n10904) );
  XNOR U10927 ( .A(n10906), .B(n10907), .Z(n10892) );
  XOR U10928 ( .A(n10908), .B(n10909), .Z(n10907) );
  XNOR U10929 ( .A(n10910), .B(n10911), .Z(n10906) );
  XNOR U10930 ( .A(n10912), .B(n10913), .Z(n10911) );
  ANDN U10931 ( .B(n10905), .A(n10909), .Z(n10912) );
  ANDN U10932 ( .B(n10905), .A(n10902), .Z(n10903) );
  XNOR U10933 ( .A(n10908), .B(n10914), .Z(n10902) );
  XOR U10934 ( .A(n10915), .B(n10913), .Z(n10914) );
  NAND U10935 ( .A(n10916), .B(n10917), .Z(n10913) );
  XNOR U10936 ( .A(n10910), .B(n10893), .Z(n10917) );
  IV U10937 ( .A(n10905), .Z(n10910) );
  XNOR U10938 ( .A(n10896), .B(n10909), .Z(n10916) );
  IV U10939 ( .A(n10901), .Z(n10909) );
  XOR U10940 ( .A(n10918), .B(n10919), .Z(n10901) );
  XNOR U10941 ( .A(n10920), .B(n10921), .Z(n10919) );
  XNOR U10942 ( .A(n10922), .B(n10923), .Z(n10918) );
  ANDN U10943 ( .B(n10669), .A(n10924), .Z(n10922) );
  AND U10944 ( .A(n10893), .B(n10896), .Z(n10915) );
  XNOR U10945 ( .A(n10893), .B(n10896), .Z(n10908) );
  XNOR U10946 ( .A(n10925), .B(n10926), .Z(n10896) );
  XNOR U10947 ( .A(n10927), .B(n10921), .Z(n10926) );
  XOR U10948 ( .A(n10928), .B(n10929), .Z(n10925) );
  XNOR U10949 ( .A(n10930), .B(n10923), .Z(n10929) );
  OR U10950 ( .A(n10864), .B(n10870), .Z(n10923) );
  XNOR U10951 ( .A(n10669), .B(n10931), .Z(n10870) );
  XNOR U10952 ( .A(n10924), .B(n10533), .Z(n10864) );
  ANDN U10953 ( .B(n10932), .A(n10869), .Z(n10930) );
  XNOR U10954 ( .A(n10933), .B(n10934), .Z(n10893) );
  XNOR U10955 ( .A(n10921), .B(n10935), .Z(n10934) );
  XOR U10956 ( .A(n10882), .B(n10928), .Z(n10935) );
  XNOR U10957 ( .A(n10669), .B(n10924), .Z(n10921) );
  XOR U10958 ( .A(n10575), .B(n10936), .Z(n10933) );
  XNOR U10959 ( .A(n10937), .B(n10938), .Z(n10936) );
  ANDN U10960 ( .B(n10939), .A(n10729), .Z(n10937) );
  XNOR U10961 ( .A(n10940), .B(n10941), .Z(n10905) );
  XNOR U10962 ( .A(n10927), .B(n10942), .Z(n10941) );
  XNOR U10963 ( .A(n10879), .B(n10920), .Z(n10942) );
  XOR U10964 ( .A(n10928), .B(n10943), .Z(n10920) );
  XNOR U10965 ( .A(n10944), .B(n10945), .Z(n10943) );
  NAND U10966 ( .A(n10676), .B(n10887), .Z(n10945) );
  XNOR U10967 ( .A(n10946), .B(n10944), .Z(n10928) );
  NANDN U10968 ( .A(n10873), .B(n10889), .Z(n10944) );
  XOR U10969 ( .A(n10897), .B(n10887), .Z(n10889) );
  XNOR U10970 ( .A(n10939), .B(n10533), .Z(n10887) );
  XOR U10971 ( .A(n10875), .B(n10676), .Z(n10873) );
  XNOR U10972 ( .A(n10729), .B(n10931), .Z(n10676) );
  ANDN U10973 ( .B(n10897), .A(n10875), .Z(n10946) );
  XOR U10974 ( .A(n10575), .B(n10669), .Z(n10875) );
  XNOR U10975 ( .A(n10947), .B(n10948), .Z(n10669) );
  XNOR U10976 ( .A(n10949), .B(n10950), .Z(n10948) );
  XOR U10977 ( .A(n10931), .B(n10932), .Z(n10927) );
  IV U10978 ( .A(n10533), .Z(n10932) );
  XOR U10979 ( .A(n10951), .B(n10952), .Z(n10533) );
  XOR U10980 ( .A(n10953), .B(n10950), .Z(n10952) );
  IV U10981 ( .A(n10869), .Z(n10931) );
  XOR U10982 ( .A(n10950), .B(n10954), .Z(n10869) );
  XNOR U10983 ( .A(n10955), .B(n10956), .Z(n10940) );
  XNOR U10984 ( .A(n10957), .B(n10938), .Z(n10956) );
  OR U10985 ( .A(n10883), .B(n10726), .Z(n10938) );
  XNOR U10986 ( .A(n10575), .B(n10729), .Z(n10726) );
  IV U10987 ( .A(n10955), .Z(n10729) );
  XOR U10988 ( .A(n10882), .B(n10939), .Z(n10883) );
  IV U10989 ( .A(n10879), .Z(n10939) );
  XOR U10990 ( .A(n10865), .B(n10958), .Z(n10879) );
  XNOR U10991 ( .A(n10959), .B(n10947), .Z(n10958) );
  XOR U10992 ( .A(n10960), .B(n10961), .Z(n10947) );
  XNOR U10993 ( .A(n9289), .B(n9285), .Z(n10961) );
  IV U10994 ( .A(n10222), .Z(n9285) );
  XNOR U10995 ( .A(n10234), .B(n10962), .Z(n10222) );
  XNOR U10996 ( .A(key[178]), .B(n10963), .Z(n10960) );
  NOR U10997 ( .A(n10882), .B(n10575), .Z(n10957) );
  XOR U10998 ( .A(n10964), .B(n10965), .Z(n10955) );
  XNOR U10999 ( .A(n10966), .B(n10967), .Z(n10965) );
  XNOR U11000 ( .A(n10575), .B(n10949), .Z(n10964) );
  XOR U11001 ( .A(n10968), .B(n10969), .Z(n10949) );
  XNOR U11002 ( .A(n10228), .B(n10970), .Z(n10969) );
  XOR U11003 ( .A(n10962), .B(n10959), .Z(n10970) );
  IV U11004 ( .A(n10953), .Z(n10959) );
  XNOR U11005 ( .A(n10971), .B(n10972), .Z(n10953) );
  XNOR U11006 ( .A(n10973), .B(n9253), .Z(n10972) );
  XOR U11007 ( .A(n10963), .B(n10225), .Z(n9253) );
  XNOR U11008 ( .A(key[177]), .B(n10974), .Z(n10971) );
  XNOR U11009 ( .A(n10975), .B(n10187), .Z(n10228) );
  XNOR U11010 ( .A(n10976), .B(n10977), .Z(n10968) );
  XOR U11011 ( .A(key[179]), .B(n9254), .Z(n10977) );
  IV U11012 ( .A(n10924), .Z(n10865) );
  XOR U11013 ( .A(n10951), .B(n10978), .Z(n10924) );
  XOR U11014 ( .A(n10950), .B(n10967), .Z(n10978) );
  XNOR U11015 ( .A(n10979), .B(n10980), .Z(n10967) );
  XNOR U11016 ( .A(n10981), .B(n10982), .Z(n10980) );
  XNOR U11017 ( .A(key[183]), .B(n10975), .Z(n10979) );
  IV U11018 ( .A(n10242), .Z(n10975) );
  XOR U11019 ( .A(n10951), .B(n10983), .Z(n10882) );
  XOR U11020 ( .A(n10950), .B(n10966), .Z(n10983) );
  XNOR U11021 ( .A(n10984), .B(n10985), .Z(n10966) );
  XOR U11022 ( .A(n10986), .B(n10189), .Z(n10985) );
  XOR U11023 ( .A(n10242), .B(n10207), .Z(n10189) );
  XNOR U11024 ( .A(n10987), .B(n10988), .Z(n10984) );
  XNOR U11025 ( .A(key[180]), .B(n10186), .Z(n10988) );
  XOR U11026 ( .A(n10989), .B(n10990), .Z(n10950) );
  XNOR U11027 ( .A(n10575), .B(n10216), .Z(n10990) );
  XOR U11028 ( .A(n10242), .B(n10201), .Z(n10216) );
  XNOR U11029 ( .A(n10991), .B(n10992), .Z(n10575) );
  XOR U11030 ( .A(n10993), .B(n9290), .Z(n10992) );
  XOR U11031 ( .A(n10974), .B(n10240), .Z(n9290) );
  XNOR U11032 ( .A(key[176]), .B(n10188), .Z(n10991) );
  IV U11033 ( .A(n10214), .Z(n10188) );
  XOR U11034 ( .A(n10994), .B(n10995), .Z(n10989) );
  XNOR U11035 ( .A(key[182]), .B(n10996), .Z(n10995) );
  IV U11036 ( .A(n10954), .Z(n10951) );
  XOR U11037 ( .A(n10997), .B(n10998), .Z(n10954) );
  XNOR U11038 ( .A(n10999), .B(n10213), .Z(n10998) );
  XOR U11039 ( .A(n10209), .B(n10994), .Z(n10213) );
  XNOR U11040 ( .A(key[181]), .B(n10206), .Z(n10997) );
  XNOR U11041 ( .A(n7953), .B(n11000), .Z(n10722) );
  XOR U11042 ( .A(key[346]), .B(n7950), .Z(n11000) );
  IV U11043 ( .A(n7328), .Z(n7950) );
  XOR U11044 ( .A(n10593), .B(n10518), .Z(n7328) );
  XOR U11045 ( .A(n10599), .B(n11001), .Z(n10518) );
  XOR U11046 ( .A(n10596), .B(n11002), .Z(n11001) );
  NAND U11047 ( .A(n11003), .B(n10560), .Z(n11002) );
  ANDN U11048 ( .B(n10685), .A(n11004), .Z(n10596) );
  XOR U11049 ( .A(n10597), .B(n10560), .Z(n10685) );
  XNOR U11050 ( .A(n10599), .B(n11005), .Z(n10593) );
  XOR U11051 ( .A(n11006), .B(n10553), .Z(n11005) );
  OR U11052 ( .A(n11007), .B(n10694), .Z(n10553) );
  XOR U11053 ( .A(n10555), .B(n10690), .Z(n10694) );
  ANDN U11054 ( .B(n10690), .A(n11008), .Z(n11006) );
  XOR U11055 ( .A(n11009), .B(n10601), .Z(n10599) );
  OR U11056 ( .A(n10701), .B(n11010), .Z(n10601) );
  XOR U11057 ( .A(n11011), .B(n10603), .Z(n10701) );
  XNOR U11058 ( .A(n10690), .B(n10560), .Z(n10603) );
  XOR U11059 ( .A(n11012), .B(n11013), .Z(n10560) );
  NANDN U11060 ( .A(n11014), .B(n11015), .Z(n11013) );
  XOR U11061 ( .A(n11016), .B(n11017), .Z(n10690) );
  OR U11062 ( .A(n11014), .B(n11018), .Z(n11017) );
  ANDN U11063 ( .B(n11011), .A(n11019), .Z(n11009) );
  IV U11064 ( .A(n10704), .Z(n11011) );
  XOR U11065 ( .A(n10555), .B(n10597), .Z(n10704) );
  XNOR U11066 ( .A(n11020), .B(n11012), .Z(n10597) );
  NANDN U11067 ( .A(n11021), .B(n11022), .Z(n11012) );
  ANDN U11068 ( .B(n11023), .A(n11024), .Z(n11020) );
  NANDN U11069 ( .A(n11021), .B(n11026), .Z(n11016) );
  XOR U11070 ( .A(n11027), .B(n11014), .Z(n11021) );
  XNOR U11071 ( .A(n11028), .B(n11029), .Z(n11014) );
  XOR U11072 ( .A(n11030), .B(n11023), .Z(n11029) );
  XNOR U11073 ( .A(n11031), .B(n11032), .Z(n11028) );
  XNOR U11074 ( .A(n11033), .B(n11034), .Z(n11032) );
  ANDN U11075 ( .B(n11023), .A(n11035), .Z(n11033) );
  IV U11076 ( .A(n11036), .Z(n11023) );
  ANDN U11077 ( .B(n11027), .A(n11035), .Z(n11025) );
  IV U11078 ( .A(n11031), .Z(n11035) );
  IV U11079 ( .A(n11024), .Z(n11027) );
  XNOR U11080 ( .A(n11030), .B(n11037), .Z(n11024) );
  XOR U11081 ( .A(n11038), .B(n11034), .Z(n11037) );
  NAND U11082 ( .A(n11026), .B(n11022), .Z(n11034) );
  XNOR U11083 ( .A(n11015), .B(n11036), .Z(n11022) );
  XOR U11084 ( .A(n11039), .B(n11040), .Z(n11036) );
  XOR U11085 ( .A(n11041), .B(n11042), .Z(n11040) );
  XNOR U11086 ( .A(n10689), .B(n11043), .Z(n11042) );
  XNOR U11087 ( .A(n11044), .B(n11045), .Z(n11039) );
  XNOR U11088 ( .A(n11046), .B(n11047), .Z(n11045) );
  ANDN U11089 ( .B(n11048), .A(n10556), .Z(n11046) );
  XNOR U11090 ( .A(n11031), .B(n11018), .Z(n11026) );
  XOR U11091 ( .A(n11049), .B(n11050), .Z(n11031) );
  XNOR U11092 ( .A(n11051), .B(n11043), .Z(n11050) );
  XOR U11093 ( .A(n11052), .B(n11053), .Z(n11043) );
  XNOR U11094 ( .A(n11054), .B(n11055), .Z(n11053) );
  NAND U11095 ( .A(n10604), .B(n10699), .Z(n11055) );
  XNOR U11096 ( .A(n11056), .B(n11057), .Z(n11049) );
  ANDN U11097 ( .B(n11058), .A(n10598), .Z(n11056) );
  ANDN U11098 ( .B(n11015), .A(n11018), .Z(n11038) );
  XOR U11099 ( .A(n11018), .B(n11015), .Z(n11030) );
  XNOR U11100 ( .A(n11059), .B(n11060), .Z(n11015) );
  XNOR U11101 ( .A(n11052), .B(n11061), .Z(n11060) );
  XOR U11102 ( .A(n11051), .B(n10693), .Z(n11061) );
  XOR U11103 ( .A(n10556), .B(n11062), .Z(n11059) );
  XNOR U11104 ( .A(n11063), .B(n11047), .Z(n11062) );
  OR U11105 ( .A(n10695), .B(n11007), .Z(n11047) );
  XNOR U11106 ( .A(n10556), .B(n11008), .Z(n11007) );
  XOR U11107 ( .A(n10693), .B(n10689), .Z(n10695) );
  ANDN U11108 ( .B(n10689), .A(n11008), .Z(n11063) );
  XOR U11109 ( .A(n11064), .B(n11065), .Z(n11018) );
  XOR U11110 ( .A(n11052), .B(n11041), .Z(n11065) );
  XOR U11111 ( .A(n11003), .B(n10561), .Z(n11041) );
  XOR U11112 ( .A(n11066), .B(n11054), .Z(n11052) );
  NANDN U11113 ( .A(n11010), .B(n10702), .Z(n11054) );
  XOR U11114 ( .A(n10703), .B(n10699), .Z(n10702) );
  XNOR U11115 ( .A(n11058), .B(n11067), .Z(n10689) );
  XOR U11116 ( .A(n11068), .B(n11069), .Z(n11067) );
  XOR U11117 ( .A(n11019), .B(n10604), .Z(n11010) );
  XNOR U11118 ( .A(n11008), .B(n11003), .Z(n10604) );
  IV U11119 ( .A(n11044), .Z(n11008) );
  XOR U11120 ( .A(n11070), .B(n11071), .Z(n11044) );
  XOR U11121 ( .A(n11072), .B(n11073), .Z(n11071) );
  XNOR U11122 ( .A(n10556), .B(n11074), .Z(n11070) );
  ANDN U11123 ( .B(n10703), .A(n11019), .Z(n11066) );
  XNOR U11124 ( .A(n10556), .B(n10598), .Z(n11019) );
  XOR U11125 ( .A(n11058), .B(n11048), .Z(n10703) );
  IV U11126 ( .A(n10693), .Z(n11048) );
  XOR U11127 ( .A(n11075), .B(n11076), .Z(n10693) );
  XOR U11128 ( .A(n11077), .B(n11073), .Z(n11076) );
  XNOR U11129 ( .A(n11078), .B(n11079), .Z(n11073) );
  XOR U11130 ( .A(n11080), .B(n9932), .Z(n11079) );
  XOR U11131 ( .A(n9946), .B(n9954), .Z(n9932) );
  XNOR U11132 ( .A(n11081), .B(n11082), .Z(n11078) );
  XNOR U11133 ( .A(key[228]), .B(n9930), .Z(n11082) );
  IV U11134 ( .A(n10683), .Z(n11058) );
  XOR U11135 ( .A(n11051), .B(n11083), .Z(n11064) );
  XNOR U11136 ( .A(n11084), .B(n11057), .Z(n11083) );
  OR U11137 ( .A(n10684), .B(n11004), .Z(n11057) );
  XNOR U11138 ( .A(n11085), .B(n11003), .Z(n11004) );
  XNOR U11139 ( .A(n10683), .B(n10561), .Z(n10684) );
  ANDN U11140 ( .B(n11003), .A(n10561), .Z(n11084) );
  XOR U11141 ( .A(n11075), .B(n11086), .Z(n10561) );
  XNOR U11142 ( .A(n11069), .B(n11087), .Z(n11086) );
  XOR U11143 ( .A(n11077), .B(n11075), .Z(n11003) );
  XNOR U11144 ( .A(n10598), .B(n10683), .Z(n11051) );
  XOR U11145 ( .A(n11075), .B(n11088), .Z(n10683) );
  XNOR U11146 ( .A(n11077), .B(n11072), .Z(n11088) );
  XOR U11147 ( .A(n11089), .B(n11090), .Z(n11072) );
  XNOR U11148 ( .A(n11091), .B(n11092), .Z(n11090) );
  XNOR U11149 ( .A(key[231]), .B(n11093), .Z(n11089) );
  XNOR U11150 ( .A(n11094), .B(n11095), .Z(n11075) );
  XNOR U11151 ( .A(n11096), .B(n9937), .Z(n11095) );
  XOR U11152 ( .A(n9956), .B(n11097), .Z(n9937) );
  XNOR U11153 ( .A(key[229]), .B(n9953), .Z(n11094) );
  IV U11154 ( .A(n11085), .Z(n10598) );
  XOR U11155 ( .A(n11087), .B(n11098), .Z(n11085) );
  XNOR U11156 ( .A(n11068), .B(n11074), .Z(n11098) );
  XOR U11157 ( .A(n11099), .B(n11100), .Z(n11074) );
  XOR U11158 ( .A(n11069), .B(n11101), .Z(n11100) );
  XNOR U11159 ( .A(n11102), .B(n9910), .Z(n11101) );
  XNOR U11160 ( .A(n9946), .B(n9931), .Z(n9910) );
  XNOR U11161 ( .A(n11103), .B(n11104), .Z(n11069) );
  XNOR U11162 ( .A(n9150), .B(n9105), .Z(n11104) );
  XOR U11163 ( .A(n11105), .B(n9913), .Z(n9105) );
  XNOR U11164 ( .A(key[225]), .B(n11106), .Z(n11103) );
  XNOR U11165 ( .A(n11107), .B(n11108), .Z(n11099) );
  XNOR U11166 ( .A(key[227]), .B(n11109), .Z(n11108) );
  XOR U11167 ( .A(n11110), .B(n11111), .Z(n11068) );
  XOR U11168 ( .A(n11112), .B(n9137), .Z(n11111) );
  XOR U11169 ( .A(n9900), .B(n11102), .Z(n9137) );
  XNOR U11170 ( .A(key[226]), .B(n11105), .Z(n11110) );
  IV U11171 ( .A(n11077), .Z(n11087) );
  XOR U11172 ( .A(n11113), .B(n11114), .Z(n11077) );
  XOR U11173 ( .A(n10556), .B(n9947), .Z(n11114) );
  XNOR U11174 ( .A(n9946), .B(n9924), .Z(n9947) );
  XNOR U11175 ( .A(n11115), .B(n11116), .Z(n10556) );
  XOR U11176 ( .A(n11117), .B(n9142), .Z(n11116) );
  XOR U11177 ( .A(n11106), .B(n9944), .Z(n9142) );
  XNOR U11178 ( .A(key[224]), .B(n9938), .Z(n11115) );
  IV U11179 ( .A(n9916), .Z(n9938) );
  XNOR U11180 ( .A(key[230]), .B(n11119), .Z(n11118) );
  XOR U11181 ( .A(n11120), .B(n11121), .Z(n7953) );
  XOR U11182 ( .A(n10606), .B(n10564), .Z(n11121) );
  XNOR U11183 ( .A(n11122), .B(n11123), .Z(n10564) );
  XNOR U11184 ( .A(n11124), .B(n10498), .Z(n11123) );
  ANDN U11185 ( .B(n11125), .A(n11126), .Z(n10498) );
  ANDN U11186 ( .B(n11127), .A(n10716), .Z(n11124) );
  IV U11187 ( .A(n11128), .Z(n10716) );
  XOR U11188 ( .A(n10705), .B(n11129), .Z(n10606) );
  XOR U11189 ( .A(n10714), .B(n11130), .Z(n11129) );
  NANDN U11190 ( .A(n11131), .B(n10500), .Z(n11130) );
  XOR U11191 ( .A(n11128), .B(n10500), .Z(n11125) );
  XOR U11192 ( .A(n11133), .B(n10718), .Z(n10705) );
  OR U11193 ( .A(n11134), .B(n11135), .Z(n10718) );
  NOR U11194 ( .A(n11136), .B(n11137), .Z(n11133) );
  XNOR U11195 ( .A(n10608), .B(n10622), .Z(n11120) );
  XNOR U11196 ( .A(n10494), .B(n11138), .Z(n10622) );
  XNOR U11197 ( .A(n11139), .B(n11140), .Z(n11138) );
  NANDN U11198 ( .A(n11141), .B(n10710), .Z(n11140) );
  XNOR U11199 ( .A(n11139), .B(n11143), .Z(n11142) );
  NANDN U11200 ( .A(n11144), .B(n10620), .Z(n11143) );
  OR U11201 ( .A(n10709), .B(n11145), .Z(n11139) );
  XNOR U11202 ( .A(n10620), .B(n10710), .Z(n10709) );
  XNOR U11203 ( .A(n10494), .B(n11146), .Z(n11122) );
  XNOR U11204 ( .A(n11147), .B(n11148), .Z(n11146) );
  NANDN U11205 ( .A(n10720), .B(n11149), .Z(n11148) );
  XOR U11206 ( .A(n11150), .B(n11147), .Z(n10494) );
  NANDN U11207 ( .A(n11134), .B(n11151), .Z(n11147) );
  XNOR U11208 ( .A(n11136), .B(n10720), .Z(n11134) );
  XNOR U11209 ( .A(n10710), .B(n10500), .Z(n10720) );
  XOR U11210 ( .A(n11152), .B(n11153), .Z(n10500) );
  NANDN U11211 ( .A(n11154), .B(n11155), .Z(n11153) );
  XOR U11212 ( .A(n11156), .B(n11157), .Z(n10710) );
  NANDN U11213 ( .A(n11154), .B(n11158), .Z(n11157) );
  ANDN U11214 ( .B(n11159), .A(n11136), .Z(n11150) );
  XNOR U11215 ( .A(n11128), .B(n10620), .Z(n11136) );
  XNOR U11216 ( .A(n11160), .B(n11156), .Z(n10620) );
  NANDN U11217 ( .A(n11161), .B(n11162), .Z(n11156) );
  XOR U11218 ( .A(n11158), .B(n11163), .Z(n11162) );
  ANDN U11219 ( .B(n11163), .A(n11164), .Z(n11160) );
  XNOR U11220 ( .A(n11165), .B(n11152), .Z(n11128) );
  NANDN U11221 ( .A(n11161), .B(n11166), .Z(n11152) );
  XOR U11222 ( .A(n11167), .B(n11155), .Z(n11166) );
  XNOR U11223 ( .A(n11168), .B(n11169), .Z(n11154) );
  XOR U11224 ( .A(n11170), .B(n11171), .Z(n11169) );
  XNOR U11225 ( .A(n11172), .B(n11173), .Z(n11168) );
  XNOR U11226 ( .A(n11174), .B(n11175), .Z(n11173) );
  ANDN U11227 ( .B(n11167), .A(n11171), .Z(n11174) );
  ANDN U11228 ( .B(n11167), .A(n11164), .Z(n11165) );
  XNOR U11229 ( .A(n11170), .B(n11176), .Z(n11164) );
  XOR U11230 ( .A(n11177), .B(n11175), .Z(n11176) );
  NAND U11231 ( .A(n11178), .B(n11179), .Z(n11175) );
  XNOR U11232 ( .A(n11172), .B(n11155), .Z(n11179) );
  IV U11233 ( .A(n11167), .Z(n11172) );
  XNOR U11234 ( .A(n11158), .B(n11171), .Z(n11178) );
  IV U11235 ( .A(n11163), .Z(n11171) );
  XOR U11236 ( .A(n11180), .B(n11181), .Z(n11163) );
  XNOR U11237 ( .A(n11182), .B(n11183), .Z(n11181) );
  XNOR U11238 ( .A(n11184), .B(n11185), .Z(n11180) );
  ANDN U11239 ( .B(n10715), .A(n11186), .Z(n11184) );
  AND U11240 ( .A(n11155), .B(n11158), .Z(n11177) );
  XNOR U11241 ( .A(n11155), .B(n11158), .Z(n11170) );
  XNOR U11242 ( .A(n11187), .B(n11188), .Z(n11158) );
  XNOR U11243 ( .A(n11189), .B(n11183), .Z(n11188) );
  XOR U11244 ( .A(n11190), .B(n11191), .Z(n11187) );
  XNOR U11245 ( .A(n11192), .B(n11185), .Z(n11191) );
  OR U11246 ( .A(n11126), .B(n11132), .Z(n11185) );
  XNOR U11247 ( .A(n10715), .B(n11193), .Z(n11132) );
  XNOR U11248 ( .A(n11186), .B(n10501), .Z(n11126) );
  ANDN U11249 ( .B(n11194), .A(n11131), .Z(n11192) );
  XNOR U11250 ( .A(n11195), .B(n11196), .Z(n11155) );
  XNOR U11251 ( .A(n11183), .B(n11197), .Z(n11196) );
  XOR U11252 ( .A(n11144), .B(n11190), .Z(n11197) );
  XNOR U11253 ( .A(n10715), .B(n11186), .Z(n11183) );
  XOR U11254 ( .A(n10619), .B(n11198), .Z(n11195) );
  XNOR U11255 ( .A(n11199), .B(n11200), .Z(n11198) );
  ANDN U11256 ( .B(n11201), .A(n10711), .Z(n11199) );
  XNOR U11257 ( .A(n11202), .B(n11203), .Z(n11167) );
  XNOR U11258 ( .A(n11189), .B(n11204), .Z(n11203) );
  XNOR U11259 ( .A(n11141), .B(n11182), .Z(n11204) );
  XOR U11260 ( .A(n11190), .B(n11205), .Z(n11182) );
  XNOR U11261 ( .A(n11206), .B(n11207), .Z(n11205) );
  NAND U11262 ( .A(n10721), .B(n11149), .Z(n11207) );
  XNOR U11263 ( .A(n11208), .B(n11206), .Z(n11190) );
  NANDN U11264 ( .A(n11135), .B(n11151), .Z(n11206) );
  XOR U11265 ( .A(n11159), .B(n11149), .Z(n11151) );
  XNOR U11266 ( .A(n11201), .B(n10501), .Z(n11149) );
  XOR U11267 ( .A(n11137), .B(n10721), .Z(n11135) );
  XNOR U11268 ( .A(n10711), .B(n11193), .Z(n10721) );
  ANDN U11269 ( .B(n11159), .A(n11137), .Z(n11208) );
  XOR U11270 ( .A(n10619), .B(n10715), .Z(n11137) );
  XNOR U11271 ( .A(n11209), .B(n11210), .Z(n10715) );
  XNOR U11272 ( .A(n11211), .B(n11212), .Z(n11210) );
  XOR U11273 ( .A(n11193), .B(n11194), .Z(n11189) );
  IV U11274 ( .A(n10501), .Z(n11194) );
  XOR U11275 ( .A(n11213), .B(n11214), .Z(n10501) );
  XNOR U11276 ( .A(n11215), .B(n11212), .Z(n11214) );
  IV U11277 ( .A(n11131), .Z(n11193) );
  XOR U11278 ( .A(n11212), .B(n11216), .Z(n11131) );
  XNOR U11279 ( .A(n11217), .B(n11218), .Z(n11202) );
  XNOR U11280 ( .A(n11219), .B(n11200), .Z(n11218) );
  OR U11281 ( .A(n11145), .B(n10708), .Z(n11200) );
  XNOR U11282 ( .A(n10619), .B(n10711), .Z(n10708) );
  IV U11283 ( .A(n11217), .Z(n10711) );
  XOR U11284 ( .A(n11144), .B(n11201), .Z(n11145) );
  IV U11285 ( .A(n11141), .Z(n11201) );
  XOR U11286 ( .A(n11127), .B(n11220), .Z(n11141) );
  XNOR U11287 ( .A(n11215), .B(n11209), .Z(n11220) );
  XOR U11288 ( .A(n11221), .B(n11222), .Z(n11209) );
  XNOR U11289 ( .A(n9438), .B(n9443), .Z(n11222) );
  XNOR U11290 ( .A(n10365), .B(n11223), .Z(n11221) );
  XOR U11291 ( .A(key[218]), .B(n10370), .Z(n11223) );
  NOR U11292 ( .A(n11144), .B(n10619), .Z(n11219) );
  XOR U11293 ( .A(n11224), .B(n11225), .Z(n11217) );
  XNOR U11294 ( .A(n11226), .B(n11227), .Z(n11225) );
  XNOR U11295 ( .A(n10619), .B(n11211), .Z(n11224) );
  XOR U11296 ( .A(n11228), .B(n11229), .Z(n11211) );
  XNOR U11297 ( .A(n11215), .B(n11230), .Z(n11229) );
  XOR U11298 ( .A(n11231), .B(n10357), .Z(n11230) );
  XOR U11299 ( .A(n11232), .B(n10327), .Z(n10357) );
  XOR U11300 ( .A(n11233), .B(n11234), .Z(n11215) );
  XOR U11301 ( .A(n11235), .B(n10369), .Z(n11234) );
  XOR U11302 ( .A(key[217]), .B(n10361), .Z(n11236) );
  XNOR U11303 ( .A(n9399), .B(n11237), .Z(n11228) );
  XNOR U11304 ( .A(key[219]), .B(n11238), .Z(n11237) );
  IV U11305 ( .A(n11186), .Z(n11127) );
  XOR U11306 ( .A(n11213), .B(n11239), .Z(n11186) );
  XOR U11307 ( .A(n11212), .B(n11227), .Z(n11239) );
  XNOR U11308 ( .A(n11240), .B(n11241), .Z(n11227) );
  XNOR U11309 ( .A(n10337), .B(n9453), .Z(n11241) );
  XOR U11310 ( .A(n11242), .B(n11243), .Z(n9453) );
  XOR U11311 ( .A(n9425), .B(n11244), .Z(n10337) );
  XOR U11312 ( .A(key[223]), .B(n10346), .Z(n11240) );
  XOR U11313 ( .A(n11213), .B(n11245), .Z(n11144) );
  XOR U11314 ( .A(n11212), .B(n11226), .Z(n11245) );
  XNOR U11315 ( .A(n11246), .B(n11247), .Z(n11226) );
  XOR U11316 ( .A(n10325), .B(n10322), .Z(n11247) );
  XOR U11317 ( .A(n9434), .B(n11248), .Z(n10322) );
  XNOR U11318 ( .A(n11242), .B(n10340), .Z(n10325) );
  XOR U11319 ( .A(n10362), .B(n11249), .Z(n11246) );
  XNOR U11320 ( .A(key[220]), .B(n11250), .Z(n11249) );
  XOR U11321 ( .A(n11251), .B(n11252), .Z(n11212) );
  XNOR U11322 ( .A(n10619), .B(n10351), .Z(n11252) );
  XNOR U11323 ( .A(n11253), .B(n10336), .Z(n10351) );
  XOR U11324 ( .A(n11242), .B(n11254), .Z(n10336) );
  XNOR U11325 ( .A(n11255), .B(n11256), .Z(n10619) );
  XNOR U11326 ( .A(n11257), .B(n10360), .Z(n11256) );
  XNOR U11327 ( .A(n11258), .B(n11259), .Z(n11255) );
  XOR U11328 ( .A(key[216]), .B(n9427), .Z(n11259) );
  XNOR U11329 ( .A(n9418), .B(n11260), .Z(n11251) );
  XNOR U11330 ( .A(key[222]), .B(n11261), .Z(n11260) );
  IV U11331 ( .A(n11216), .Z(n11213) );
  XOR U11332 ( .A(n11262), .B(n11263), .Z(n11216) );
  XNOR U11333 ( .A(n10324), .B(n10341), .Z(n11263) );
  XOR U11334 ( .A(n9416), .B(n11264), .Z(n10341) );
  XNOR U11335 ( .A(n11265), .B(n11266), .Z(n11262) );
  XNOR U11336 ( .A(key[221]), .B(n10353), .Z(n11266) );
  XNOR U11337 ( .A(n8336), .B(n11267), .Z(n3947) );
  XOR U11338 ( .A(n8370), .B(n8338), .Z(n11267) );
  XOR U11339 ( .A(n8424), .B(n11268), .Z(n8338) );
  XOR U11340 ( .A(n11269), .B(n8514), .Z(n11268) );
  OR U11341 ( .A(n11270), .B(n11271), .Z(n8514) );
  AND U11342 ( .A(n11272), .B(n11273), .Z(n11269) );
  XNOR U11343 ( .A(n8508), .B(n11274), .Z(n8370) );
  XOR U11344 ( .A(n11275), .B(n8504), .Z(n11274) );
  OR U11345 ( .A(n11271), .B(n11276), .Z(n8504) );
  XOR U11346 ( .A(n8506), .B(n11273), .Z(n11271) );
  ANDN U11347 ( .B(n11273), .A(n11277), .Z(n11275) );
  XOR U11348 ( .A(n11278), .B(n8525), .Z(n8508) );
  OR U11349 ( .A(n11279), .B(n11280), .Z(n8525) );
  XNOR U11350 ( .A(n8517), .B(n11283), .Z(n8336) );
  XNOR U11351 ( .A(n8427), .B(n11284), .Z(n11283) );
  OR U11352 ( .A(n8523), .B(n11285), .Z(n11284) );
  NAND U11353 ( .A(n8521), .B(n11286), .Z(n8427) );
  XNOR U11354 ( .A(n8523), .B(n8428), .Z(n8521) );
  XNOR U11355 ( .A(n8424), .B(n11287), .Z(n8517) );
  XNOR U11356 ( .A(n11288), .B(n11289), .Z(n11287) );
  NAND U11357 ( .A(n11290), .B(n8527), .Z(n11289) );
  XOR U11358 ( .A(n11291), .B(n11288), .Z(n8424) );
  OR U11359 ( .A(n11279), .B(n11292), .Z(n11288) );
  XNOR U11360 ( .A(n11282), .B(n8527), .Z(n11279) );
  XOR U11361 ( .A(n11273), .B(n8428), .Z(n8527) );
  XOR U11362 ( .A(n11293), .B(n11294), .Z(n8428) );
  NANDN U11363 ( .A(n11295), .B(n11296), .Z(n11294) );
  XOR U11364 ( .A(n11297), .B(n11298), .Z(n11273) );
  OR U11365 ( .A(n11295), .B(n11299), .Z(n11298) );
  ANDN U11366 ( .B(n11282), .A(n11300), .Z(n11291) );
  XOR U11367 ( .A(n8506), .B(n8523), .Z(n11282) );
  XOR U11368 ( .A(n11301), .B(n11293), .Z(n8523) );
  NANDN U11369 ( .A(n11302), .B(n11303), .Z(n11293) );
  ANDN U11370 ( .B(n11304), .A(n11305), .Z(n11301) );
  NANDN U11371 ( .A(n11302), .B(n11307), .Z(n11297) );
  XOR U11372 ( .A(n11308), .B(n11295), .Z(n11302) );
  XNOR U11373 ( .A(n11309), .B(n11310), .Z(n11295) );
  XOR U11374 ( .A(n11311), .B(n11304), .Z(n11310) );
  XNOR U11375 ( .A(n11312), .B(n11313), .Z(n11309) );
  XNOR U11376 ( .A(n11314), .B(n11315), .Z(n11313) );
  ANDN U11377 ( .B(n11304), .A(n11316), .Z(n11314) );
  IV U11378 ( .A(n11317), .Z(n11304) );
  ANDN U11379 ( .B(n11308), .A(n11316), .Z(n11306) );
  IV U11380 ( .A(n11312), .Z(n11316) );
  IV U11381 ( .A(n11305), .Z(n11308) );
  XNOR U11382 ( .A(n11311), .B(n11318), .Z(n11305) );
  XOR U11383 ( .A(n11319), .B(n11315), .Z(n11318) );
  NAND U11384 ( .A(n11307), .B(n11303), .Z(n11315) );
  XNOR U11385 ( .A(n11296), .B(n11317), .Z(n11303) );
  XOR U11386 ( .A(n11320), .B(n11321), .Z(n11317) );
  XOR U11387 ( .A(n11322), .B(n11323), .Z(n11321) );
  XOR U11388 ( .A(n11324), .B(n11325), .Z(n11323) );
  XOR U11389 ( .A(n11272), .B(n11326), .Z(n11320) );
  XNOR U11390 ( .A(n11327), .B(n11328), .Z(n11326) );
  AND U11391 ( .A(n8516), .B(n8507), .Z(n11327) );
  XNOR U11392 ( .A(n11312), .B(n11299), .Z(n11307) );
  XOR U11393 ( .A(n11329), .B(n11330), .Z(n11312) );
  XNOR U11394 ( .A(n11331), .B(n11325), .Z(n11330) );
  XOR U11395 ( .A(n11332), .B(n11333), .Z(n11325) );
  XNOR U11396 ( .A(n11334), .B(n11335), .Z(n11333) );
  NAND U11397 ( .A(n8528), .B(n11290), .Z(n11335) );
  XNOR U11398 ( .A(n11336), .B(n11337), .Z(n11329) );
  ANDN U11399 ( .B(n8522), .A(n11285), .Z(n11336) );
  ANDN U11400 ( .B(n11296), .A(n11299), .Z(n11319) );
  XOR U11401 ( .A(n11299), .B(n11296), .Z(n11311) );
  XNOR U11402 ( .A(n11338), .B(n11339), .Z(n11296) );
  XNOR U11403 ( .A(n11332), .B(n11340), .Z(n11339) );
  XNOR U11404 ( .A(n8516), .B(n11331), .Z(n11340) );
  XNOR U11405 ( .A(n8507), .B(n11341), .Z(n11338) );
  XNOR U11406 ( .A(n11342), .B(n11328), .Z(n11341) );
  OR U11407 ( .A(n11270), .B(n11276), .Z(n11328) );
  XNOR U11408 ( .A(n8507), .B(n11324), .Z(n11276) );
  XNOR U11409 ( .A(n8516), .B(n11272), .Z(n11270) );
  ANDN U11410 ( .B(n11272), .A(n11277), .Z(n11342) );
  IV U11411 ( .A(n11324), .Z(n11277) );
  XOR U11412 ( .A(n11343), .B(n11344), .Z(n11299) );
  XOR U11413 ( .A(n11332), .B(n11322), .Z(n11344) );
  XOR U11414 ( .A(n11345), .B(n8512), .Z(n11322) );
  XOR U11415 ( .A(n11346), .B(n11334), .Z(n11332) );
  OR U11416 ( .A(n11280), .B(n11292), .Z(n11334) );
  XOR U11417 ( .A(n11300), .B(n11290), .Z(n11292) );
  XOR U11418 ( .A(n11345), .B(n11272), .Z(n11290) );
  XOR U11419 ( .A(n11347), .B(n11348), .Z(n11272) );
  XNOR U11420 ( .A(n11285), .B(n11349), .Z(n11348) );
  XNOR U11421 ( .A(n11281), .B(n8528), .Z(n11280) );
  XNOR U11422 ( .A(n8512), .B(n11324), .Z(n8528) );
  XOR U11423 ( .A(n11350), .B(n11351), .Z(n11324) );
  XNOR U11424 ( .A(n11352), .B(n11353), .Z(n11351) );
  XOR U11425 ( .A(n11354), .B(n8507), .Z(n11350) );
  ANDN U11426 ( .B(n11281), .A(n11300), .Z(n11346) );
  XNOR U11427 ( .A(n11355), .B(n8516), .Z(n11300) );
  XOR U11428 ( .A(n11352), .B(n11356), .Z(n8516) );
  XOR U11429 ( .A(n11357), .B(n11358), .Z(n11356) );
  XOR U11430 ( .A(n11359), .B(n6091), .Z(n11352) );
  XNOR U11431 ( .A(n11360), .B(n11361), .Z(n6091) );
  XOR U11432 ( .A(n6911), .B(n6916), .Z(n11361) );
  XNOR U11433 ( .A(n7752), .B(n11362), .Z(n6916) );
  IV U11434 ( .A(n6102), .Z(n7752) );
  XNOR U11435 ( .A(n11363), .B(n6883), .Z(n6911) );
  XOR U11436 ( .A(n6928), .B(n7768), .Z(n11360) );
  IV U11437 ( .A(n11364), .Z(n6928) );
  XNOR U11438 ( .A(n7780), .B(n11365), .Z(n11359) );
  XOR U11439 ( .A(key[356]), .B(n7781), .Z(n11365) );
  XNOR U11440 ( .A(n7777), .B(n6080), .Z(n7780) );
  XNOR U11441 ( .A(n11366), .B(n11367), .Z(n6080) );
  XNOR U11442 ( .A(n11368), .B(n11369), .Z(n11367) );
  XNOR U11443 ( .A(n11370), .B(n11371), .Z(n11366) );
  XOR U11444 ( .A(n11372), .B(n11373), .Z(n11371) );
  ANDN U11445 ( .B(n11374), .A(n11375), .Z(n11373) );
  XOR U11446 ( .A(n8507), .B(n8522), .Z(n11281) );
  XOR U11447 ( .A(n11331), .B(n11376), .Z(n11343) );
  XNOR U11448 ( .A(n11377), .B(n11337), .Z(n11376) );
  NANDN U11449 ( .A(n8520), .B(n11286), .Z(n11337) );
  XOR U11450 ( .A(n11285), .B(n8429), .Z(n11286) );
  XNOR U11451 ( .A(n8522), .B(n11378), .Z(n8520) );
  ANDN U11452 ( .B(n11345), .A(n8512), .Z(n11377) );
  IV U11453 ( .A(n11378), .Z(n8512) );
  IV U11454 ( .A(n8429), .Z(n11345) );
  XNOR U11455 ( .A(n11349), .B(n11378), .Z(n8429) );
  XNOR U11456 ( .A(n11379), .B(n11358), .Z(n11378) );
  XNOR U11457 ( .A(n11355), .B(n8522), .Z(n11331) );
  XNOR U11458 ( .A(n11353), .B(n11380), .Z(n8522) );
  XNOR U11459 ( .A(n11358), .B(n11347), .Z(n11380) );
  XOR U11460 ( .A(n11381), .B(n11382), .Z(n11347) );
  XOR U11461 ( .A(n7791), .B(n11383), .Z(n11382) );
  XOR U11462 ( .A(n6107), .B(n6063), .Z(n7791) );
  XOR U11463 ( .A(n11384), .B(n11385), .Z(n6107) );
  XNOR U11464 ( .A(n11386), .B(n11387), .Z(n11385) );
  XOR U11465 ( .A(n11388), .B(n11389), .Z(n11384) );
  XNOR U11466 ( .A(key[354]), .B(n6920), .Z(n11381) );
  XOR U11467 ( .A(n6883), .B(n6102), .Z(n6920) );
  XNOR U11468 ( .A(n11390), .B(n11391), .Z(n6102) );
  XOR U11469 ( .A(n11392), .B(n11393), .Z(n6883) );
  XOR U11470 ( .A(n11394), .B(n11395), .Z(n11353) );
  XNOR U11471 ( .A(n6099), .B(n11396), .Z(n11395) );
  XNOR U11472 ( .A(n7785), .B(n11349), .Z(n11396) );
  XOR U11473 ( .A(n11397), .B(n11398), .Z(n11349) );
  XOR U11474 ( .A(n6112), .B(n6881), .Z(n11398) );
  XNOR U11475 ( .A(n6061), .B(n11383), .Z(n6881) );
  XNOR U11476 ( .A(key[353]), .B(n6106), .Z(n11397) );
  XNOR U11477 ( .A(n7797), .B(n6116), .Z(n6106) );
  XOR U11478 ( .A(n11399), .B(n11400), .Z(n6116) );
  XOR U11479 ( .A(n11401), .B(n11402), .Z(n11400) );
  IV U11480 ( .A(n6921), .Z(n7797) );
  XOR U11481 ( .A(n11403), .B(n11404), .Z(n6921) );
  XOR U11482 ( .A(n11392), .B(n11405), .Z(n11404) );
  XOR U11483 ( .A(n7795), .B(n6094), .Z(n7785) );
  XOR U11484 ( .A(n11370), .B(n6061), .Z(n6094) );
  XOR U11485 ( .A(n11406), .B(n11407), .Z(n6061) );
  IV U11486 ( .A(n7777), .Z(n7795) );
  XNOR U11487 ( .A(n11364), .B(n7781), .Z(n6099) );
  XOR U11488 ( .A(n11408), .B(n11383), .Z(n7781) );
  IV U11489 ( .A(n6103), .Z(n11383) );
  XOR U11490 ( .A(n11409), .B(n11410), .Z(n6103) );
  XNOR U11491 ( .A(n6882), .B(n11411), .Z(n11394) );
  XNOR U11492 ( .A(key[355]), .B(n6063), .Z(n11411) );
  XOR U11493 ( .A(n11412), .B(n11413), .Z(n6063) );
  XNOR U11494 ( .A(n11410), .B(n11414), .Z(n11413) );
  XOR U11495 ( .A(n11415), .B(n11416), .Z(n11412) );
  IV U11496 ( .A(n6098), .Z(n6882) );
  XNOR U11497 ( .A(n6922), .B(n6062), .Z(n6098) );
  XNOR U11498 ( .A(n11417), .B(n11418), .Z(n6062) );
  XOR U11499 ( .A(n11419), .B(n11420), .Z(n11418) );
  XNOR U11500 ( .A(n11401), .B(n11402), .Z(n11417) );
  IV U11501 ( .A(n11390), .Z(n11401) );
  XOR U11502 ( .A(n11421), .B(n11422), .Z(n6922) );
  XNOR U11503 ( .A(n11423), .B(n11424), .Z(n11422) );
  IV U11504 ( .A(n11285), .Z(n11355) );
  XNOR U11505 ( .A(n11379), .B(n11354), .Z(n11425) );
  XOR U11506 ( .A(n11426), .B(n11427), .Z(n11354) );
  XNOR U11507 ( .A(n11428), .B(n6088), .Z(n11427) );
  XOR U11508 ( .A(n7765), .B(n6891), .Z(n6088) );
  XNOR U11509 ( .A(n11429), .B(n11430), .Z(n6891) );
  XNOR U11510 ( .A(n11399), .B(n11431), .Z(n11430) );
  XOR U11511 ( .A(n11390), .B(n11402), .Z(n11429) );
  XOR U11512 ( .A(n11432), .B(n11433), .Z(n11402) );
  XNOR U11513 ( .A(n11434), .B(n11435), .Z(n11433) );
  OR U11514 ( .A(n11436), .B(n11437), .Z(n11435) );
  XOR U11515 ( .A(n11438), .B(n11439), .Z(n11390) );
  XNOR U11516 ( .A(n11440), .B(n11441), .Z(n11439) );
  NAND U11517 ( .A(n11442), .B(n11443), .Z(n11441) );
  XOR U11518 ( .A(n11421), .B(n11444), .Z(n7765) );
  XOR U11519 ( .A(n11403), .B(n11445), .Z(n11444) );
  XNOR U11520 ( .A(n11392), .B(n11405), .Z(n11421) );
  XOR U11521 ( .A(n11446), .B(n11447), .Z(n11405) );
  XNOR U11522 ( .A(n11448), .B(n11449), .Z(n11447) );
  NANDN U11523 ( .A(n11450), .B(n11451), .Z(n11449) );
  XNOR U11524 ( .A(n11452), .B(n11453), .Z(n11392) );
  XNOR U11525 ( .A(n11454), .B(n11455), .Z(n11453) );
  NAND U11526 ( .A(n11456), .B(n11457), .Z(n11455) );
  XOR U11527 ( .A(key[359]), .B(n7777), .Z(n11426) );
  IV U11528 ( .A(n11357), .Z(n11379) );
  XNOR U11529 ( .A(n11458), .B(n11459), .Z(n11357) );
  XOR U11530 ( .A(n7768), .B(n6079), .Z(n11459) );
  XOR U11531 ( .A(n6898), .B(n6908), .Z(n6079) );
  XNOR U11532 ( .A(n11460), .B(n11461), .Z(n6908) );
  XOR U11533 ( .A(n11362), .B(n11431), .Z(n11461) );
  XNOR U11534 ( .A(n11462), .B(n11463), .Z(n11431) );
  XNOR U11535 ( .A(n11464), .B(n11465), .Z(n11463) );
  OR U11536 ( .A(n11436), .B(n11466), .Z(n11465) );
  XNOR U11537 ( .A(n11467), .B(n11468), .Z(n11460) );
  XNOR U11538 ( .A(n11469), .B(n11470), .Z(n11468) );
  ANDN U11539 ( .B(n11443), .A(n11471), .Z(n11470) );
  XOR U11540 ( .A(n11472), .B(n11473), .Z(n6898) );
  XNOR U11541 ( .A(n11363), .B(n11445), .Z(n11473) );
  XNOR U11542 ( .A(n11474), .B(n11475), .Z(n11445) );
  XNOR U11543 ( .A(n11476), .B(n11477), .Z(n11475) );
  OR U11544 ( .A(n11450), .B(n11478), .Z(n11477) );
  XNOR U11545 ( .A(n11479), .B(n11480), .Z(n11472) );
  XOR U11546 ( .A(n11481), .B(n11482), .Z(n11480) );
  ANDN U11547 ( .B(n11457), .A(n11483), .Z(n11482) );
  XNOR U11548 ( .A(n11484), .B(n11485), .Z(n7768) );
  XNOR U11549 ( .A(n11486), .B(n11487), .Z(n11485) );
  XNOR U11550 ( .A(n11408), .B(n11488), .Z(n11484) );
  XOR U11551 ( .A(n11489), .B(n11490), .Z(n11488) );
  ANDN U11552 ( .B(n11491), .A(n11492), .Z(n11490) );
  XNOR U11553 ( .A(key[357]), .B(n7763), .Z(n11458) );
  XOR U11554 ( .A(n6075), .B(n6082), .Z(n7763) );
  IV U11555 ( .A(n7770), .Z(n6075) );
  XOR U11556 ( .A(n11493), .B(n11387), .Z(n7770) );
  XNOR U11557 ( .A(n11494), .B(n11495), .Z(n11387) );
  XNOR U11558 ( .A(n11496), .B(n11372), .Z(n11495) );
  ANDN U11559 ( .B(n11497), .A(n11498), .Z(n11372) );
  ANDN U11560 ( .B(n11499), .A(n11500), .Z(n11496) );
  XOR U11561 ( .A(n11501), .B(n11502), .Z(n11358) );
  XOR U11562 ( .A(n8507), .B(n6072), .Z(n11502) );
  XOR U11563 ( .A(n6897), .B(n11428), .Z(n6072) );
  XNOR U11564 ( .A(n11364), .B(n7776), .Z(n11428) );
  XNOR U11565 ( .A(n11503), .B(n11504), .Z(n7776) );
  XNOR U11566 ( .A(n11410), .B(n11487), .Z(n11504) );
  XNOR U11567 ( .A(n11505), .B(n11506), .Z(n11487) );
  XNOR U11568 ( .A(n11507), .B(n11508), .Z(n11506) );
  NANDN U11569 ( .A(n11509), .B(n11510), .Z(n11508) );
  IV U11570 ( .A(n11511), .Z(n11410) );
  XOR U11571 ( .A(n11415), .B(n11512), .Z(n11503) );
  XOR U11572 ( .A(n6890), .B(n6078), .Z(n6897) );
  IV U11573 ( .A(n7761), .Z(n6078) );
  XOR U11574 ( .A(n11399), .B(n11420), .Z(n7761) );
  XOR U11575 ( .A(n11432), .B(n11513), .Z(n11420) );
  XOR U11576 ( .A(n11514), .B(n11469), .Z(n11513) );
  NANDN U11577 ( .A(n11515), .B(n11516), .Z(n11469) );
  ANDN U11578 ( .B(n11517), .A(n11518), .Z(n11514) );
  XNOR U11579 ( .A(n11467), .B(n11519), .Z(n11432) );
  XNOR U11580 ( .A(n11520), .B(n11521), .Z(n11519) );
  NAND U11581 ( .A(n11522), .B(n11523), .Z(n11521) );
  XOR U11582 ( .A(n11524), .B(n11419), .Z(n11399) );
  XNOR U11583 ( .A(n11467), .B(n11525), .Z(n11419) );
  XNOR U11584 ( .A(n11434), .B(n11526), .Z(n11525) );
  NANDN U11585 ( .A(n11527), .B(n11528), .Z(n11526) );
  OR U11586 ( .A(n11529), .B(n11530), .Z(n11434) );
  XOR U11587 ( .A(n11531), .B(n11520), .Z(n11467) );
  NANDN U11588 ( .A(n11532), .B(n11533), .Z(n11520) );
  ANDN U11589 ( .B(n11534), .A(n11535), .Z(n11531) );
  XOR U11590 ( .A(n11403), .B(n11424), .Z(n6890) );
  XNOR U11591 ( .A(n11446), .B(n11536), .Z(n11424) );
  XNOR U11592 ( .A(n11537), .B(n11481), .Z(n11536) );
  ANDN U11593 ( .B(n11538), .A(n11539), .Z(n11481) );
  ANDN U11594 ( .B(n11540), .A(n11541), .Z(n11537) );
  XNOR U11595 ( .A(n11479), .B(n11542), .Z(n11446) );
  XNOR U11596 ( .A(n11543), .B(n11544), .Z(n11542) );
  NAND U11597 ( .A(n11545), .B(n11546), .Z(n11544) );
  XNOR U11598 ( .A(n11423), .B(n11393), .Z(n11403) );
  XNOR U11599 ( .A(n11479), .B(n11547), .Z(n11423) );
  XNOR U11600 ( .A(n11448), .B(n11548), .Z(n11547) );
  NANDN U11601 ( .A(n11549), .B(n11550), .Z(n11548) );
  OR U11602 ( .A(n11551), .B(n11552), .Z(n11448) );
  XOR U11603 ( .A(n11553), .B(n11543), .Z(n11479) );
  NANDN U11604 ( .A(n11554), .B(n11555), .Z(n11543) );
  ANDN U11605 ( .B(n11556), .A(n11557), .Z(n11553) );
  XOR U11606 ( .A(n11558), .B(n11559), .Z(n8507) );
  XOR U11607 ( .A(n6919), .B(n6087), .Z(n11559) );
  XNOR U11608 ( .A(n11364), .B(n6113), .Z(n6087) );
  XNOR U11609 ( .A(n11524), .B(n11362), .Z(n6113) );
  XOR U11610 ( .A(n11462), .B(n11560), .Z(n11362) );
  XOR U11611 ( .A(n11561), .B(n11440), .Z(n11560) );
  NANDN U11612 ( .A(n11562), .B(n11516), .Z(n11440) );
  XOR U11613 ( .A(n11517), .B(n11443), .Z(n11516) );
  ANDN U11614 ( .B(n11517), .A(n11563), .Z(n11561) );
  XNOR U11615 ( .A(n11438), .B(n11564), .Z(n11462) );
  XNOR U11616 ( .A(n11565), .B(n11566), .Z(n11564) );
  NAND U11617 ( .A(n11523), .B(n11567), .Z(n11566) );
  IV U11618 ( .A(n11391), .Z(n11524) );
  XNOR U11619 ( .A(n11438), .B(n11568), .Z(n11391) );
  XOR U11620 ( .A(n11569), .B(n11464), .Z(n11568) );
  OR U11621 ( .A(n11570), .B(n11529), .Z(n11464) );
  XNOR U11622 ( .A(n11436), .B(n11527), .Z(n11529) );
  NOR U11623 ( .A(n11571), .B(n11527), .Z(n11569) );
  XOR U11624 ( .A(n11572), .B(n11565), .Z(n11438) );
  OR U11625 ( .A(n11532), .B(n11573), .Z(n11565) );
  XNOR U11626 ( .A(n11574), .B(n11523), .Z(n11532) );
  XNOR U11627 ( .A(n11527), .B(n11443), .Z(n11523) );
  XOR U11628 ( .A(n11575), .B(n11576), .Z(n11443) );
  NANDN U11629 ( .A(n11577), .B(n11578), .Z(n11576) );
  XNOR U11630 ( .A(n11579), .B(n11580), .Z(n11527) );
  OR U11631 ( .A(n11577), .B(n11581), .Z(n11580) );
  ANDN U11632 ( .B(n11574), .A(n11582), .Z(n11572) );
  IV U11633 ( .A(n11535), .Z(n11574) );
  XOR U11634 ( .A(n11436), .B(n11517), .Z(n11535) );
  XNOR U11635 ( .A(n11583), .B(n11575), .Z(n11517) );
  NANDN U11636 ( .A(n11584), .B(n11585), .Z(n11575) );
  ANDN U11637 ( .B(n11586), .A(n11587), .Z(n11583) );
  NANDN U11638 ( .A(n11584), .B(n11589), .Z(n11579) );
  XOR U11639 ( .A(n11590), .B(n11577), .Z(n11584) );
  XNOR U11640 ( .A(n11591), .B(n11592), .Z(n11577) );
  XOR U11641 ( .A(n11593), .B(n11586), .Z(n11592) );
  XNOR U11642 ( .A(n11594), .B(n11595), .Z(n11591) );
  XNOR U11643 ( .A(n11596), .B(n11597), .Z(n11595) );
  ANDN U11644 ( .B(n11586), .A(n11598), .Z(n11596) );
  IV U11645 ( .A(n11599), .Z(n11586) );
  ANDN U11646 ( .B(n11590), .A(n11598), .Z(n11588) );
  IV U11647 ( .A(n11594), .Z(n11598) );
  IV U11648 ( .A(n11587), .Z(n11590) );
  XNOR U11649 ( .A(n11593), .B(n11600), .Z(n11587) );
  XOR U11650 ( .A(n11601), .B(n11597), .Z(n11600) );
  NAND U11651 ( .A(n11589), .B(n11585), .Z(n11597) );
  XNOR U11652 ( .A(n11578), .B(n11599), .Z(n11585) );
  XOR U11653 ( .A(n11602), .B(n11603), .Z(n11599) );
  XOR U11654 ( .A(n11604), .B(n11605), .Z(n11603) );
  XNOR U11655 ( .A(n11528), .B(n11606), .Z(n11605) );
  XNOR U11656 ( .A(n11607), .B(n11608), .Z(n11602) );
  XNOR U11657 ( .A(n11609), .B(n11610), .Z(n11608) );
  ANDN U11658 ( .B(n11611), .A(n11466), .Z(n11609) );
  XNOR U11659 ( .A(n11594), .B(n11581), .Z(n11589) );
  XOR U11660 ( .A(n11612), .B(n11613), .Z(n11594) );
  XNOR U11661 ( .A(n11614), .B(n11606), .Z(n11613) );
  XOR U11662 ( .A(n11615), .B(n11616), .Z(n11606) );
  XNOR U11663 ( .A(n11617), .B(n11618), .Z(n11616) );
  NAND U11664 ( .A(n11567), .B(n11522), .Z(n11618) );
  XNOR U11665 ( .A(n11619), .B(n11620), .Z(n11612) );
  ANDN U11666 ( .B(n11621), .A(n11563), .Z(n11619) );
  ANDN U11667 ( .B(n11578), .A(n11581), .Z(n11601) );
  XOR U11668 ( .A(n11581), .B(n11578), .Z(n11593) );
  XNOR U11669 ( .A(n11622), .B(n11623), .Z(n11578) );
  XNOR U11670 ( .A(n11615), .B(n11624), .Z(n11623) );
  XOR U11671 ( .A(n11614), .B(n11437), .Z(n11624) );
  XOR U11672 ( .A(n11466), .B(n11625), .Z(n11622) );
  XNOR U11673 ( .A(n11626), .B(n11610), .Z(n11625) );
  OR U11674 ( .A(n11530), .B(n11570), .Z(n11610) );
  XNOR U11675 ( .A(n11466), .B(n11571), .Z(n11570) );
  XOR U11676 ( .A(n11437), .B(n11528), .Z(n11530) );
  ANDN U11677 ( .B(n11528), .A(n11571), .Z(n11626) );
  XOR U11678 ( .A(n11627), .B(n11628), .Z(n11581) );
  XOR U11679 ( .A(n11615), .B(n11604), .Z(n11628) );
  XOR U11680 ( .A(n11442), .B(n11471), .Z(n11604) );
  XOR U11681 ( .A(n11629), .B(n11617), .Z(n11615) );
  NANDN U11682 ( .A(n11573), .B(n11533), .Z(n11617) );
  XOR U11683 ( .A(n11534), .B(n11522), .Z(n11533) );
  XNOR U11684 ( .A(n11621), .B(n11630), .Z(n11528) );
  XNOR U11685 ( .A(n11631), .B(n11632), .Z(n11630) );
  XOR U11686 ( .A(n11582), .B(n11567), .Z(n11573) );
  XNOR U11687 ( .A(n11571), .B(n11442), .Z(n11567) );
  IV U11688 ( .A(n11607), .Z(n11571) );
  XOR U11689 ( .A(n11633), .B(n11634), .Z(n11607) );
  XOR U11690 ( .A(n11635), .B(n11636), .Z(n11634) );
  XNOR U11691 ( .A(n11466), .B(n11637), .Z(n11633) );
  ANDN U11692 ( .B(n11534), .A(n11582), .Z(n11629) );
  XNOR U11693 ( .A(n11466), .B(n11563), .Z(n11582) );
  XOR U11694 ( .A(n11621), .B(n11611), .Z(n11534) );
  IV U11695 ( .A(n11437), .Z(n11611) );
  XOR U11696 ( .A(n11638), .B(n11639), .Z(n11437) );
  XOR U11697 ( .A(n11640), .B(n11636), .Z(n11639) );
  XNOR U11698 ( .A(n11641), .B(n11642), .Z(n11636) );
  XOR U11699 ( .A(n9432), .B(n9430), .Z(n11642) );
  XOR U11700 ( .A(n10327), .B(n10362), .Z(n9430) );
  XOR U11701 ( .A(n11643), .B(n9443), .Z(n10362) );
  XNOR U11702 ( .A(n11644), .B(n10369), .Z(n10327) );
  XNOR U11703 ( .A(n10350), .B(n11264), .Z(n9432) );
  XNOR U11704 ( .A(n11250), .B(n11645), .Z(n11641) );
  XNOR U11705 ( .A(key[212]), .B(n11248), .Z(n11645) );
  XOR U11706 ( .A(n11243), .B(n9416), .Z(n11250) );
  XOR U11707 ( .A(n11646), .B(n11647), .Z(n9416) );
  XNOR U11708 ( .A(n11648), .B(n11649), .Z(n11647) );
  XNOR U11709 ( .A(n11650), .B(n11651), .Z(n11646) );
  XOR U11710 ( .A(n11652), .B(n11653), .Z(n11651) );
  ANDN U11711 ( .B(n11654), .A(n11655), .Z(n11653) );
  IV U11712 ( .A(n11518), .Z(n11621) );
  XOR U11713 ( .A(n11614), .B(n11656), .Z(n11627) );
  XNOR U11714 ( .A(n11657), .B(n11620), .Z(n11656) );
  OR U11715 ( .A(n11515), .B(n11562), .Z(n11620) );
  XNOR U11716 ( .A(n11658), .B(n11442), .Z(n11562) );
  XNOR U11717 ( .A(n11518), .B(n11471), .Z(n11515) );
  ANDN U11718 ( .B(n11442), .A(n11471), .Z(n11657) );
  XOR U11719 ( .A(n11638), .B(n11659), .Z(n11471) );
  XOR U11720 ( .A(n11631), .B(n11660), .Z(n11659) );
  XOR U11721 ( .A(n11640), .B(n11638), .Z(n11442) );
  XNOR U11722 ( .A(n11563), .B(n11518), .Z(n11614) );
  XOR U11723 ( .A(n11638), .B(n11661), .Z(n11518) );
  XNOR U11724 ( .A(n11640), .B(n11635), .Z(n11661) );
  XOR U11725 ( .A(n11662), .B(n11663), .Z(n11635) );
  XOR U11726 ( .A(n11664), .B(n9426), .Z(n11663) );
  XOR U11727 ( .A(n11254), .B(n10346), .Z(n9426) );
  XNOR U11728 ( .A(n11665), .B(n11666), .Z(n10346) );
  XOR U11729 ( .A(n11667), .B(n11668), .Z(n11666) );
  XNOR U11730 ( .A(n11669), .B(n11670), .Z(n11665) );
  XNOR U11731 ( .A(n11671), .B(n11672), .Z(n11254) );
  XNOR U11732 ( .A(n11673), .B(n11674), .Z(n11672) );
  XNOR U11733 ( .A(key[215]), .B(n11257), .Z(n11662) );
  XNOR U11734 ( .A(n11675), .B(n11676), .Z(n11638) );
  XNOR U11735 ( .A(n11253), .B(n9417), .Z(n11676) );
  XNOR U11736 ( .A(n11677), .B(n11678), .Z(n10324) );
  XNOR U11737 ( .A(n11679), .B(n11668), .Z(n11678) );
  XNOR U11738 ( .A(n11680), .B(n11681), .Z(n11668) );
  XNOR U11739 ( .A(n11682), .B(n11683), .Z(n11681) );
  NANDN U11740 ( .A(n11684), .B(n11685), .Z(n11683) );
  XNOR U11741 ( .A(n11643), .B(n11686), .Z(n11677) );
  XNOR U11742 ( .A(n11687), .B(n11688), .Z(n11686) );
  ANDN U11743 ( .B(n11689), .A(n11690), .Z(n11687) );
  XOR U11744 ( .A(n11691), .B(n11692), .Z(n10340) );
  XNOR U11745 ( .A(n11693), .B(n11674), .Z(n11692) );
  XNOR U11746 ( .A(n11694), .B(n11695), .Z(n11674) );
  XNOR U11747 ( .A(n11696), .B(n11697), .Z(n11695) );
  NANDN U11748 ( .A(n11698), .B(n11699), .Z(n11697) );
  XNOR U11749 ( .A(n11644), .B(n11700), .Z(n11691) );
  XOR U11750 ( .A(n11701), .B(n11702), .Z(n11700) );
  ANDN U11751 ( .B(n11703), .A(n11704), .Z(n11702) );
  XNOR U11752 ( .A(n9420), .B(n9411), .Z(n11253) );
  IV U11753 ( .A(n11265), .Z(n9411) );
  XOR U11754 ( .A(n11705), .B(n11706), .Z(n11265) );
  XNOR U11755 ( .A(key[213]), .B(n11264), .Z(n11675) );
  XOR U11756 ( .A(n11707), .B(n11708), .Z(n11264) );
  XNOR U11757 ( .A(n11709), .B(n11710), .Z(n11708) );
  XNOR U11758 ( .A(n11711), .B(n11712), .Z(n11707) );
  XOR U11759 ( .A(n11713), .B(n11714), .Z(n11712) );
  ANDN U11760 ( .B(n11715), .A(n11716), .Z(n11714) );
  IV U11761 ( .A(n11658), .Z(n11563) );
  XNOR U11762 ( .A(n11632), .B(n11717), .Z(n11658) );
  XOR U11763 ( .A(n11637), .B(n11660), .Z(n11717) );
  IV U11764 ( .A(n11640), .Z(n11660) );
  XOR U11765 ( .A(n11718), .B(n11719), .Z(n11640) );
  XNOR U11766 ( .A(n11261), .B(n9413), .Z(n11719) );
  XNOR U11767 ( .A(n10342), .B(n11664), .Z(n9413) );
  XNOR U11768 ( .A(n11720), .B(n11244), .Z(n11664) );
  XNOR U11769 ( .A(n11721), .B(n11722), .Z(n11244) );
  XNOR U11770 ( .A(n11723), .B(n11710), .Z(n11722) );
  XNOR U11771 ( .A(n11724), .B(n11725), .Z(n11710) );
  XNOR U11772 ( .A(n11726), .B(n11727), .Z(n11725) );
  NANDN U11773 ( .A(n11728), .B(n11729), .Z(n11727) );
  XNOR U11774 ( .A(n11730), .B(n11731), .Z(n11721) );
  XNOR U11775 ( .A(n9418), .B(n10353), .Z(n10342) );
  XNOR U11776 ( .A(n11673), .B(n11732), .Z(n10353) );
  XNOR U11777 ( .A(n11733), .B(n11669), .Z(n9418) );
  XOR U11778 ( .A(n11243), .B(n9425), .Z(n11261) );
  XOR U11779 ( .A(n11734), .B(n11735), .Z(n9425) );
  XOR U11780 ( .A(n11705), .B(n11649), .Z(n11735) );
  XNOR U11781 ( .A(n11736), .B(n11737), .Z(n11649) );
  XNOR U11782 ( .A(n11738), .B(n11739), .Z(n11737) );
  OR U11783 ( .A(n11740), .B(n11741), .Z(n11739) );
  XOR U11784 ( .A(n11742), .B(n11743), .Z(n11734) );
  XNOR U11785 ( .A(n9420), .B(n11744), .Z(n11718) );
  XOR U11786 ( .A(key[214]), .B(n11466), .Z(n11744) );
  XNOR U11787 ( .A(n11745), .B(n11746), .Z(n11466) );
  XOR U11788 ( .A(n11242), .B(n10361), .Z(n11746) );
  XOR U11789 ( .A(n9446), .B(n9454), .Z(n10361) );
  IV U11790 ( .A(n11258), .Z(n9446) );
  XOR U11791 ( .A(n11705), .B(n11747), .Z(n11258) );
  XOR U11792 ( .A(n11748), .B(n11743), .Z(n11747) );
  XOR U11793 ( .A(n11749), .B(n11750), .Z(n11705) );
  IV U11794 ( .A(n11232), .Z(n11242) );
  XOR U11795 ( .A(n11751), .B(n11644), .Z(n11232) );
  XNOR U11796 ( .A(n11694), .B(n11752), .Z(n11644) );
  XOR U11797 ( .A(n11753), .B(n11754), .Z(n11752) );
  NOR U11798 ( .A(n11755), .B(n11756), .Z(n11753) );
  XNOR U11799 ( .A(n11757), .B(n11758), .Z(n11694) );
  XNOR U11800 ( .A(n11759), .B(n11760), .Z(n11758) );
  NANDN U11801 ( .A(n11761), .B(n11762), .Z(n11760) );
  XOR U11802 ( .A(key[208]), .B(n9427), .Z(n11745) );
  XOR U11803 ( .A(n10323), .B(n11720), .Z(n9427) );
  IV U11804 ( .A(n10350), .Z(n11720) );
  XOR U11805 ( .A(n11763), .B(n11643), .Z(n10323) );
  XNOR U11806 ( .A(n11680), .B(n11764), .Z(n11643) );
  XOR U11807 ( .A(n11765), .B(n11766), .Z(n11764) );
  ANDN U11808 ( .B(n11767), .A(n11768), .Z(n11765) );
  XNOR U11809 ( .A(n11769), .B(n11770), .Z(n11680) );
  XNOR U11810 ( .A(n11771), .B(n11772), .Z(n11770) );
  NANDN U11811 ( .A(n11773), .B(n11774), .Z(n11772) );
  XNOR U11812 ( .A(n11775), .B(n11776), .Z(n9420) );
  XOR U11813 ( .A(n11777), .B(n11778), .Z(n11776) );
  XOR U11814 ( .A(n11779), .B(n11780), .Z(n11637) );
  XNOR U11815 ( .A(n9447), .B(n11781), .Z(n11780) );
  XNOR U11816 ( .A(n11631), .B(n9449), .Z(n11781) );
  IV U11817 ( .A(n10368), .Z(n9449) );
  XOR U11818 ( .A(n10365), .B(n9399), .Z(n10368) );
  XOR U11819 ( .A(n11782), .B(n11783), .Z(n9399) );
  XNOR U11820 ( .A(n11784), .B(n11733), .Z(n11783) );
  XNOR U11821 ( .A(n11785), .B(n11786), .Z(n11733) );
  XNOR U11822 ( .A(n11688), .B(n11787), .Z(n11786) );
  NAND U11823 ( .A(n11788), .B(n11767), .Z(n11787) );
  NANDN U11824 ( .A(n11789), .B(n11790), .Z(n11688) );
  XNOR U11825 ( .A(n11791), .B(n11670), .Z(n11782) );
  XOR U11826 ( .A(n11671), .B(n11792), .Z(n10365) );
  XNOR U11827 ( .A(n11793), .B(n11732), .Z(n11792) );
  XNOR U11828 ( .A(n11794), .B(n11795), .Z(n11732) );
  XNOR U11829 ( .A(n11796), .B(n11701), .Z(n11795) );
  NOR U11830 ( .A(n11797), .B(n11798), .Z(n11701) );
  NOR U11831 ( .A(n11799), .B(n11756), .Z(n11796) );
  XNOR U11832 ( .A(n11800), .B(n11801), .Z(n11671) );
  XOR U11833 ( .A(n11802), .B(n11803), .Z(n11631) );
  IV U11834 ( .A(n9442), .Z(n10349) );
  IV U11835 ( .A(n11235), .Z(n9452) );
  XOR U11836 ( .A(n11667), .B(n11804), .Z(n11235) );
  XOR U11837 ( .A(n11669), .B(n11670), .Z(n11804) );
  XNOR U11838 ( .A(n11763), .B(n11791), .Z(n11669) );
  XNOR U11839 ( .A(n11679), .B(n11805), .Z(n11791) );
  XOR U11840 ( .A(n11806), .B(n11807), .Z(n11805) );
  ANDN U11841 ( .B(n11808), .A(n11809), .Z(n11806) );
  IV U11842 ( .A(n11784), .Z(n11667) );
  XNOR U11843 ( .A(n11807), .B(n11811), .Z(n11810) );
  NANDN U11844 ( .A(n11684), .B(n11812), .Z(n11811) );
  OR U11845 ( .A(n11813), .B(n11814), .Z(n11807) );
  XNOR U11846 ( .A(n11679), .B(n11815), .Z(n11785) );
  XNOR U11847 ( .A(n11816), .B(n11817), .Z(n11815) );
  NANDN U11848 ( .A(n11773), .B(n11818), .Z(n11817) );
  XOR U11849 ( .A(n11819), .B(n11816), .Z(n11679) );
  NANDN U11850 ( .A(n11820), .B(n11821), .Z(n11816) );
  ANDN U11851 ( .B(n11822), .A(n11823), .Z(n11819) );
  XNOR U11852 ( .A(n11673), .B(n11824), .Z(n10360) );
  XOR U11853 ( .A(n11800), .B(n11801), .Z(n11824) );
  XOR U11854 ( .A(n11794), .B(n11825), .Z(n11801) );
  XNOR U11855 ( .A(n11826), .B(n11827), .Z(n11825) );
  NANDN U11856 ( .A(n11698), .B(n11828), .Z(n11827) );
  XNOR U11857 ( .A(n11693), .B(n11829), .Z(n11794) );
  XNOR U11858 ( .A(n11830), .B(n11831), .Z(n11829) );
  NANDN U11859 ( .A(n11761), .B(n11832), .Z(n11831) );
  XNOR U11860 ( .A(n11693), .B(n11833), .Z(n11793) );
  XNOR U11861 ( .A(n11826), .B(n11834), .Z(n11833) );
  OR U11862 ( .A(n11835), .B(n11836), .Z(n11834) );
  OR U11863 ( .A(n11837), .B(n11838), .Z(n11826) );
  XOR U11864 ( .A(n11839), .B(n11830), .Z(n11693) );
  NANDN U11865 ( .A(n11840), .B(n11841), .Z(n11830) );
  AND U11866 ( .A(n11842), .B(n11843), .Z(n11839) );
  XOR U11867 ( .A(n9401), .B(n9444), .Z(n10370) );
  XOR U11868 ( .A(key[209]), .B(n9454), .Z(n11802) );
  XOR U11869 ( .A(n11723), .B(n11844), .Z(n9454) );
  XOR U11870 ( .A(n11730), .B(n11731), .Z(n11844) );
  XNOR U11871 ( .A(n11845), .B(n11778), .Z(n11730) );
  XNOR U11872 ( .A(n10350), .B(n11248), .Z(n9447) );
  XOR U11873 ( .A(n11711), .B(n9444), .Z(n11248) );
  XOR U11874 ( .A(n11777), .B(n11711), .Z(n10350) );
  XNOR U11875 ( .A(n11724), .B(n11846), .Z(n11711) );
  XNOR U11876 ( .A(n11847), .B(n11848), .Z(n11846) );
  OR U11877 ( .A(n11849), .B(n11850), .Z(n11848) );
  XNOR U11878 ( .A(n11851), .B(n11852), .Z(n11724) );
  XNOR U11879 ( .A(n11853), .B(n11854), .Z(n11852) );
  NAND U11880 ( .A(n11855), .B(n11856), .Z(n11854) );
  XNOR U11881 ( .A(n11238), .B(n11857), .Z(n11779) );
  XNOR U11882 ( .A(key[211]), .B(n9403), .Z(n11857) );
  XOR U11883 ( .A(n11243), .B(n9434), .Z(n11238) );
  XOR U11884 ( .A(n11648), .B(n9401), .Z(n9434) );
  XNOR U11885 ( .A(n11742), .B(n11858), .Z(n9401) );
  IV U11886 ( .A(n11748), .Z(n11742) );
  IV U11887 ( .A(n11257), .Z(n11243) );
  XOR U11888 ( .A(n11749), .B(n11648), .Z(n11257) );
  XNOR U11889 ( .A(n11736), .B(n11859), .Z(n11648) );
  XOR U11890 ( .A(n11860), .B(n11861), .Z(n11859) );
  NOR U11891 ( .A(n11862), .B(n11863), .Z(n11860) );
  XNOR U11892 ( .A(n11864), .B(n11865), .Z(n11736) );
  XNOR U11893 ( .A(n11866), .B(n11867), .Z(n11865) );
  NANDN U11894 ( .A(n11868), .B(n11869), .Z(n11867) );
  IV U11895 ( .A(n11858), .Z(n11749) );
  XNOR U11896 ( .A(n11864), .B(n11870), .Z(n11858) );
  XOR U11897 ( .A(n11871), .B(n11738), .Z(n11870) );
  OR U11898 ( .A(n11872), .B(n11873), .Z(n11738) );
  ANDN U11899 ( .B(n11874), .A(n11875), .Z(n11871) );
  XOR U11900 ( .A(n11876), .B(n11877), .Z(n11632) );
  XNOR U11901 ( .A(n11231), .B(n9400), .Z(n11877) );
  XOR U11902 ( .A(n9443), .B(n10369), .Z(n9400) );
  XOR U11903 ( .A(n11751), .B(n11800), .Z(n10369) );
  XNOR U11904 ( .A(n11757), .B(n11878), .Z(n11800) );
  XNOR U11905 ( .A(n11754), .B(n11879), .Z(n11878) );
  NANDN U11906 ( .A(n11880), .B(n11881), .Z(n11879) );
  OR U11907 ( .A(n11882), .B(n11797), .Z(n11754) );
  XOR U11908 ( .A(n11756), .B(n11881), .Z(n11797) );
  XNOR U11909 ( .A(n11757), .B(n11883), .Z(n11751) );
  XOR U11910 ( .A(n11884), .B(n11696), .Z(n11883) );
  OR U11911 ( .A(n11885), .B(n11837), .Z(n11696) );
  XNOR U11912 ( .A(n11698), .B(n11835), .Z(n11837) );
  NOR U11913 ( .A(n11886), .B(n11835), .Z(n11884) );
  XOR U11914 ( .A(n11887), .B(n11759), .Z(n11757) );
  OR U11915 ( .A(n11840), .B(n11888), .Z(n11759) );
  XOR U11916 ( .A(n11835), .B(n11881), .Z(n11761) );
  IV U11917 ( .A(n11704), .Z(n11881) );
  XNOR U11918 ( .A(n11889), .B(n11890), .Z(n11704) );
  NANDN U11919 ( .A(n11891), .B(n11892), .Z(n11890) );
  XNOR U11920 ( .A(n11893), .B(n11894), .Z(n11835) );
  NANDN U11921 ( .A(n11891), .B(n11895), .Z(n11894) );
  ANDN U11922 ( .B(n11842), .A(n11896), .Z(n11887) );
  XOR U11923 ( .A(n11698), .B(n11756), .Z(n11842) );
  XOR U11924 ( .A(n11897), .B(n11889), .Z(n11756) );
  NANDN U11925 ( .A(n11898), .B(n11899), .Z(n11889) );
  XOR U11926 ( .A(n11892), .B(n11900), .Z(n11899) );
  ANDN U11927 ( .B(n11900), .A(n11901), .Z(n11897) );
  NANDN U11928 ( .A(n11898), .B(n11903), .Z(n11893) );
  XOR U11929 ( .A(n11904), .B(n11905), .Z(n11891) );
  XOR U11930 ( .A(n11906), .B(n11907), .Z(n11905) );
  XNOR U11931 ( .A(n11908), .B(n11909), .Z(n11904) );
  XNOR U11932 ( .A(n11910), .B(n11911), .Z(n11909) );
  ANDN U11933 ( .B(n11907), .A(n11906), .Z(n11910) );
  ANDN U11934 ( .B(n11907), .A(n11901), .Z(n11902) );
  XNOR U11935 ( .A(n11908), .B(n11912), .Z(n11901) );
  XOR U11936 ( .A(n11913), .B(n11911), .Z(n11912) );
  NAND U11937 ( .A(n11903), .B(n11914), .Z(n11911) );
  XNOR U11938 ( .A(n11892), .B(n11906), .Z(n11914) );
  IV U11939 ( .A(n11900), .Z(n11906) );
  XNOR U11940 ( .A(n11915), .B(n11916), .Z(n11900) );
  XNOR U11941 ( .A(n11917), .B(n11918), .Z(n11916) );
  XOR U11942 ( .A(n11836), .B(n11919), .Z(n11918) );
  XNOR U11943 ( .A(n11886), .B(n11920), .Z(n11915) );
  XNOR U11944 ( .A(n11921), .B(n11922), .Z(n11920) );
  AND U11945 ( .A(n11828), .B(n11699), .Z(n11921) );
  XOR U11946 ( .A(n11895), .B(n11907), .Z(n11903) );
  AND U11947 ( .A(n11892), .B(n11895), .Z(n11913) );
  XNOR U11948 ( .A(n11892), .B(n11895), .Z(n11908) );
  XNOR U11949 ( .A(n11923), .B(n11924), .Z(n11895) );
  XNOR U11950 ( .A(n11925), .B(n11919), .Z(n11924) );
  XOR U11951 ( .A(n11926), .B(n11927), .Z(n11923) );
  XNOR U11952 ( .A(n11928), .B(n11929), .Z(n11927) );
  ANDN U11953 ( .B(n11703), .A(n11880), .Z(n11928) );
  XNOR U11954 ( .A(n11930), .B(n11931), .Z(n11892) );
  XNOR U11955 ( .A(n11828), .B(n11926), .Z(n11932) );
  XOR U11956 ( .A(n11699), .B(n11933), .Z(n11930) );
  XNOR U11957 ( .A(n11934), .B(n11922), .Z(n11933) );
  OR U11958 ( .A(n11838), .B(n11885), .Z(n11922) );
  XOR U11959 ( .A(n11699), .B(n11886), .Z(n11885) );
  XNOR U11960 ( .A(n11828), .B(n11935), .Z(n11838) );
  ANDN U11961 ( .B(n11936), .A(n11836), .Z(n11934) );
  XNOR U11962 ( .A(n11937), .B(n11938), .Z(n11907) );
  XOR U11963 ( .A(n11925), .B(n11917), .Z(n11938) );
  XOR U11964 ( .A(n11926), .B(n11939), .Z(n11917) );
  XNOR U11965 ( .A(n11940), .B(n11941), .Z(n11939) );
  NAND U11966 ( .A(n11762), .B(n11832), .Z(n11941) );
  XNOR U11967 ( .A(n11942), .B(n11940), .Z(n11926) );
  NANDN U11968 ( .A(n11888), .B(n11841), .Z(n11940) );
  XOR U11969 ( .A(n11843), .B(n11832), .Z(n11841) );
  XOR U11970 ( .A(n11935), .B(n11703), .Z(n11832) );
  IV U11971 ( .A(n11836), .Z(n11935) );
  XOR U11972 ( .A(n11943), .B(n11944), .Z(n11836) );
  XNOR U11973 ( .A(n11945), .B(n11946), .Z(n11944) );
  XOR U11974 ( .A(n11896), .B(n11762), .Z(n11888) );
  XNOR U11975 ( .A(n11936), .B(n11880), .Z(n11762) );
  IV U11976 ( .A(n11886), .Z(n11936) );
  XOR U11977 ( .A(n11947), .B(n11948), .Z(n11886) );
  XOR U11978 ( .A(n11949), .B(n11950), .Z(n11948) );
  XNOR U11979 ( .A(n11699), .B(n11951), .Z(n11947) );
  ANDN U11980 ( .B(n11843), .A(n11896), .Z(n11942) );
  XNOR U11981 ( .A(n11699), .B(n11952), .Z(n11896) );
  XOR U11982 ( .A(n11828), .B(n11943), .Z(n11843) );
  XOR U11983 ( .A(n11953), .B(n11954), .Z(n11828) );
  XOR U11984 ( .A(n11955), .B(n11950), .Z(n11954) );
  XOR U11985 ( .A(state[92]), .B(key[92]), .Z(n11950) );
  XNOR U11986 ( .A(n11952), .B(n11799), .Z(n11925) );
  XNOR U11987 ( .A(n11956), .B(n11929), .Z(n11937) );
  OR U11988 ( .A(n11798), .B(n11882), .Z(n11929) );
  XNOR U11989 ( .A(n11755), .B(n11880), .Z(n11882) );
  XOR U11990 ( .A(n11957), .B(n11953), .Z(n11880) );
  XNOR U11991 ( .A(n11943), .B(n11703), .Z(n11798) );
  XOR U11992 ( .A(n11953), .B(n11958), .Z(n11703) );
  XOR U11993 ( .A(n11945), .B(n11957), .Z(n11958) );
  IV U11994 ( .A(n11799), .Z(n11943) );
  ANDN U11995 ( .B(n11952), .A(n11799), .Z(n11956) );
  XNOR U11996 ( .A(n11953), .B(n11959), .Z(n11799) );
  XNOR U11997 ( .A(n11955), .B(n11949), .Z(n11959) );
  XNOR U11998 ( .A(state[95]), .B(key[95]), .Z(n11949) );
  XNOR U11999 ( .A(state[93]), .B(key[93]), .Z(n11953) );
  IV U12000 ( .A(n11755), .Z(n11952) );
  XNOR U12001 ( .A(n11946), .B(n11960), .Z(n11755) );
  XOR U12002 ( .A(n11951), .B(n11957), .Z(n11960) );
  IV U12003 ( .A(n11955), .Z(n11957) );
  XOR U12004 ( .A(n11699), .B(n11961), .Z(n11955) );
  XNOR U12005 ( .A(state[94]), .B(key[94]), .Z(n11961) );
  XOR U12006 ( .A(state[88]), .B(key[88]), .Z(n11699) );
  XNOR U12007 ( .A(n11945), .B(n11962), .Z(n11951) );
  XNOR U12008 ( .A(state[91]), .B(key[91]), .Z(n11962) );
  XNOR U12009 ( .A(state[89]), .B(key[89]), .Z(n11945) );
  XNOR U12010 ( .A(state[90]), .B(key[90]), .Z(n11946) );
  XOR U12011 ( .A(n11763), .B(n11670), .Z(n9443) );
  XOR U12012 ( .A(n11769), .B(n11963), .Z(n11670) );
  XNOR U12013 ( .A(n11766), .B(n11964), .Z(n11963) );
  NANDN U12014 ( .A(n11966), .B(n11790), .Z(n11766) );
  XNOR U12015 ( .A(n11767), .B(n11690), .Z(n11790) );
  XNOR U12016 ( .A(n11769), .B(n11967), .Z(n11763) );
  XOR U12017 ( .A(n11968), .B(n11682), .Z(n11967) );
  OR U12018 ( .A(n11969), .B(n11813), .Z(n11682) );
  XOR U12019 ( .A(n11684), .B(n11970), .Z(n11813) );
  ANDN U12020 ( .B(n11971), .A(n11809), .Z(n11968) );
  IV U12021 ( .A(n11970), .Z(n11809) );
  XOR U12022 ( .A(n11972), .B(n11771), .Z(n11769) );
  OR U12023 ( .A(n11820), .B(n11973), .Z(n11771) );
  XNOR U12024 ( .A(n11823), .B(n11773), .Z(n11820) );
  XOR U12025 ( .A(n11970), .B(n11690), .Z(n11773) );
  XNOR U12026 ( .A(n11974), .B(n11975), .Z(n11690) );
  NANDN U12027 ( .A(n11976), .B(n11977), .Z(n11975) );
  XOR U12028 ( .A(n11978), .B(n11979), .Z(n11970) );
  NANDN U12029 ( .A(n11976), .B(n11980), .Z(n11979) );
  XOR U12030 ( .A(n11684), .B(n11767), .Z(n11823) );
  XNOR U12031 ( .A(n11982), .B(n11974), .Z(n11767) );
  NANDN U12032 ( .A(n11983), .B(n11984), .Z(n11974) );
  XOR U12033 ( .A(n11977), .B(n11985), .Z(n11984) );
  ANDN U12034 ( .B(n11985), .A(n11986), .Z(n11982) );
  NANDN U12035 ( .A(n11983), .B(n11988), .Z(n11978) );
  XOR U12036 ( .A(n11989), .B(n11990), .Z(n11976) );
  XOR U12037 ( .A(n11991), .B(n11992), .Z(n11990) );
  XNOR U12038 ( .A(n11993), .B(n11994), .Z(n11989) );
  XNOR U12039 ( .A(n11995), .B(n11996), .Z(n11994) );
  ANDN U12040 ( .B(n11992), .A(n11991), .Z(n11995) );
  ANDN U12041 ( .B(n11992), .A(n11986), .Z(n11987) );
  XNOR U12042 ( .A(n11993), .B(n11997), .Z(n11986) );
  XOR U12043 ( .A(n11998), .B(n11996), .Z(n11997) );
  NAND U12044 ( .A(n11988), .B(n11999), .Z(n11996) );
  XNOR U12045 ( .A(n11977), .B(n11991), .Z(n11999) );
  IV U12046 ( .A(n11985), .Z(n11991) );
  XNOR U12047 ( .A(n12000), .B(n12001), .Z(n11985) );
  XNOR U12048 ( .A(n12002), .B(n12003), .Z(n12001) );
  XOR U12049 ( .A(n12004), .B(n12005), .Z(n12003) );
  XNOR U12050 ( .A(n12006), .B(n12007), .Z(n12000) );
  XNOR U12051 ( .A(n12008), .B(n12009), .Z(n12007) );
  AND U12052 ( .A(n11812), .B(n11685), .Z(n12008) );
  XOR U12053 ( .A(n11980), .B(n11992), .Z(n11988) );
  AND U12054 ( .A(n11977), .B(n11980), .Z(n11998) );
  XNOR U12055 ( .A(n11977), .B(n11980), .Z(n11993) );
  XNOR U12056 ( .A(n12010), .B(n12011), .Z(n11980) );
  XNOR U12057 ( .A(n12012), .B(n12005), .Z(n12011) );
  XOR U12058 ( .A(n12013), .B(n12014), .Z(n12010) );
  XNOR U12059 ( .A(n12015), .B(n12016), .Z(n12014) );
  ANDN U12060 ( .B(n11689), .A(n11965), .Z(n12015) );
  XNOR U12061 ( .A(n12017), .B(n12018), .Z(n11977) );
  XNOR U12062 ( .A(n11812), .B(n12013), .Z(n12019) );
  XOR U12063 ( .A(n11685), .B(n12020), .Z(n12017) );
  XNOR U12064 ( .A(n12021), .B(n12009), .Z(n12020) );
  OR U12065 ( .A(n11814), .B(n11969), .Z(n12009) );
  XOR U12066 ( .A(n11685), .B(n12006), .Z(n11969) );
  XNOR U12067 ( .A(n11812), .B(n11808), .Z(n11814) );
  ANDN U12068 ( .B(n11971), .A(n12004), .Z(n12021) );
  XNOR U12069 ( .A(n12022), .B(n12023), .Z(n11992) );
  XOR U12070 ( .A(n12012), .B(n12002), .Z(n12023) );
  XOR U12071 ( .A(n12013), .B(n12024), .Z(n12002) );
  XNOR U12072 ( .A(n12025), .B(n12026), .Z(n12024) );
  NAND U12073 ( .A(n11774), .B(n11818), .Z(n12026) );
  XNOR U12074 ( .A(n12027), .B(n12025), .Z(n12013) );
  NANDN U12075 ( .A(n11973), .B(n11821), .Z(n12025) );
  XOR U12076 ( .A(n11822), .B(n11818), .Z(n11821) );
  XOR U12077 ( .A(n11808), .B(n11689), .Z(n11818) );
  IV U12078 ( .A(n12004), .Z(n11808) );
  XOR U12079 ( .A(n11788), .B(n12028), .Z(n12004) );
  XNOR U12080 ( .A(n12029), .B(n12030), .Z(n12028) );
  XOR U12081 ( .A(n11981), .B(n11774), .Z(n11973) );
  XNOR U12082 ( .A(n11971), .B(n11965), .Z(n11774) );
  IV U12083 ( .A(n12006), .Z(n11971) );
  XOR U12084 ( .A(n12031), .B(n12032), .Z(n12006) );
  XOR U12085 ( .A(n12033), .B(n12034), .Z(n12032) );
  XOR U12086 ( .A(n11685), .B(n12035), .Z(n12031) );
  ANDN U12087 ( .B(n11822), .A(n11981), .Z(n12027) );
  XNOR U12088 ( .A(n11685), .B(n12036), .Z(n11981) );
  XOR U12089 ( .A(n11812), .B(n11788), .Z(n11822) );
  XOR U12090 ( .A(n12037), .B(n12038), .Z(n11812) );
  XOR U12091 ( .A(n12039), .B(n12034), .Z(n12038) );
  XOR U12092 ( .A(state[100]), .B(key[100]), .Z(n12034) );
  XOR U12093 ( .A(n12036), .B(n11788), .Z(n12012) );
  IV U12094 ( .A(n11768), .Z(n12036) );
  XNOR U12095 ( .A(n12040), .B(n12016), .Z(n12022) );
  OR U12096 ( .A(n11789), .B(n11966), .Z(n12016) );
  XNOR U12097 ( .A(n11768), .B(n11965), .Z(n11966) );
  XOR U12098 ( .A(n12041), .B(n12037), .Z(n11965) );
  XNOR U12099 ( .A(n11788), .B(n11689), .Z(n11789) );
  XOR U12100 ( .A(n12037), .B(n12042), .Z(n11689) );
  XOR U12101 ( .A(n12030), .B(n12041), .Z(n12042) );
  ANDN U12102 ( .B(n11788), .A(n11768), .Z(n12040) );
  XOR U12103 ( .A(n12041), .B(n12043), .Z(n11768) );
  XOR U12104 ( .A(n12029), .B(n12035), .Z(n12043) );
  XOR U12105 ( .A(n12030), .B(n12044), .Z(n12035) );
  XNOR U12106 ( .A(state[99]), .B(key[99]), .Z(n12044) );
  XNOR U12107 ( .A(state[97]), .B(key[97]), .Z(n12030) );
  XNOR U12108 ( .A(state[98]), .B(key[98]), .Z(n12029) );
  IV U12109 ( .A(n12039), .Z(n12041) );
  XOR U12110 ( .A(n12037), .B(n12045), .Z(n11788) );
  XNOR U12111 ( .A(n12039), .B(n12033), .Z(n12045) );
  XNOR U12112 ( .A(state[103]), .B(key[103]), .Z(n12033) );
  XOR U12113 ( .A(n11685), .B(n12046), .Z(n12039) );
  XNOR U12114 ( .A(state[102]), .B(key[102]), .Z(n12046) );
  XOR U12115 ( .A(state[96]), .B(key[96]), .Z(n11685) );
  XNOR U12116 ( .A(state[101]), .B(key[101]), .Z(n12037) );
  IV U12117 ( .A(n10363), .Z(n11231) );
  XOR U12118 ( .A(n9403), .B(n9438), .Z(n10363) );
  XOR U12119 ( .A(n12047), .B(n12048), .Z(n9438) );
  XOR U12120 ( .A(n11750), .B(n11706), .Z(n12048) );
  XNOR U12121 ( .A(n12049), .B(n12050), .Z(n11706) );
  XNOR U12122 ( .A(n12051), .B(n11652), .Z(n12050) );
  NOR U12123 ( .A(n12052), .B(n12053), .Z(n11652) );
  NOR U12124 ( .A(n12054), .B(n11863), .Z(n12051) );
  XOR U12125 ( .A(n11650), .B(n12055), .Z(n11750) );
  XNOR U12126 ( .A(n12056), .B(n12057), .Z(n12055) );
  NANDN U12127 ( .A(n11875), .B(n12058), .Z(n12057) );
  XNOR U12128 ( .A(n11748), .B(n11743), .Z(n12047) );
  XNOR U12129 ( .A(n12056), .B(n12060), .Z(n12059) );
  OR U12130 ( .A(n11740), .B(n12061), .Z(n12060) );
  OR U12131 ( .A(n11872), .B(n12062), .Z(n12056) );
  XOR U12132 ( .A(n11740), .B(n12063), .Z(n11872) );
  XNOR U12133 ( .A(n11650), .B(n12064), .Z(n12049) );
  XNOR U12134 ( .A(n12065), .B(n12066), .Z(n12064) );
  OR U12135 ( .A(n11868), .B(n12067), .Z(n12066) );
  XOR U12136 ( .A(n12068), .B(n12065), .Z(n11650) );
  NANDN U12137 ( .A(n12069), .B(n12070), .Z(n12065) );
  AND U12138 ( .A(n12071), .B(n12072), .Z(n12068) );
  XNOR U12139 ( .A(n11864), .B(n12073), .Z(n11748) );
  XNOR U12140 ( .A(n11861), .B(n12074), .Z(n12073) );
  NANDN U12141 ( .A(n12075), .B(n11654), .Z(n12074) );
  OR U12142 ( .A(n12076), .B(n12052), .Z(n11861) );
  XOR U12143 ( .A(n11863), .B(n11654), .Z(n12052) );
  XOR U12144 ( .A(n12077), .B(n11866), .Z(n11864) );
  OR U12145 ( .A(n12069), .B(n12078), .Z(n11866) );
  XOR U12146 ( .A(n12071), .B(n11868), .Z(n12069) );
  XNOR U12147 ( .A(n12063), .B(n11654), .Z(n11868) );
  XOR U12148 ( .A(n12079), .B(n12080), .Z(n11654) );
  NANDN U12149 ( .A(n12081), .B(n12082), .Z(n12080) );
  IV U12150 ( .A(n11875), .Z(n12063) );
  XNOR U12151 ( .A(n12083), .B(n12084), .Z(n11875) );
  NANDN U12152 ( .A(n12081), .B(n12085), .Z(n12084) );
  ANDN U12153 ( .B(n12071), .A(n12086), .Z(n12077) );
  XOR U12154 ( .A(n11863), .B(n11740), .Z(n12071) );
  XOR U12155 ( .A(n12087), .B(n12083), .Z(n11740) );
  NANDN U12156 ( .A(n12088), .B(n12089), .Z(n12083) );
  NANDN U12157 ( .A(n12088), .B(n12093), .Z(n12079) );
  XOR U12158 ( .A(n12094), .B(n12095), .Z(n12081) );
  XOR U12159 ( .A(n12096), .B(n12091), .Z(n12095) );
  XNOR U12160 ( .A(n12097), .B(n12098), .Z(n12094) );
  XNOR U12161 ( .A(n12099), .B(n12100), .Z(n12098) );
  ANDN U12162 ( .B(n12096), .A(n12091), .Z(n12099) );
  ANDN U12163 ( .B(n12096), .A(n12090), .Z(n12092) );
  XNOR U12164 ( .A(n12097), .B(n12101), .Z(n12090) );
  XOR U12165 ( .A(n12102), .B(n12100), .Z(n12101) );
  NAND U12166 ( .A(n12089), .B(n12093), .Z(n12100) );
  XNOR U12167 ( .A(n12085), .B(n12091), .Z(n12089) );
  XOR U12168 ( .A(n12103), .B(n12104), .Z(n12091) );
  XOR U12169 ( .A(n12105), .B(n12106), .Z(n12104) );
  XNOR U12170 ( .A(n12107), .B(n12108), .Z(n12103) );
  ANDN U12171 ( .B(n12109), .A(n12054), .Z(n12107) );
  AND U12172 ( .A(n12082), .B(n12085), .Z(n12102) );
  XNOR U12173 ( .A(n12082), .B(n12085), .Z(n12097) );
  XNOR U12174 ( .A(n12110), .B(n12111), .Z(n12085) );
  XNOR U12175 ( .A(n12112), .B(n12113), .Z(n12111) );
  XOR U12176 ( .A(n12105), .B(n12114), .Z(n12110) );
  XNOR U12177 ( .A(n12115), .B(n12108), .Z(n12114) );
  OR U12178 ( .A(n12053), .B(n12076), .Z(n12108) );
  XNOR U12179 ( .A(n11862), .B(n12075), .Z(n12076) );
  XNOR U12180 ( .A(n12054), .B(n11655), .Z(n12053) );
  NOR U12181 ( .A(n11655), .B(n12075), .Z(n12115) );
  XNOR U12182 ( .A(n12116), .B(n12117), .Z(n12082) );
  XNOR U12183 ( .A(n12118), .B(n12119), .Z(n12117) );
  XOR U12184 ( .A(n12061), .B(n12105), .Z(n12119) );
  XOR U12185 ( .A(n12109), .B(n12120), .Z(n12105) );
  XNOR U12186 ( .A(n11741), .B(n12121), .Z(n12116) );
  XNOR U12187 ( .A(n12122), .B(n12123), .Z(n12121) );
  ANDN U12188 ( .B(n12058), .A(n12124), .Z(n12122) );
  XNOR U12189 ( .A(n12125), .B(n12126), .Z(n12096) );
  XNOR U12190 ( .A(n12106), .B(n12127), .Z(n12126) );
  XNOR U12191 ( .A(n12058), .B(n12113), .Z(n12127) );
  XOR U12192 ( .A(n12075), .B(n11655), .Z(n12113) );
  XNOR U12193 ( .A(n12118), .B(n12128), .Z(n12106) );
  XNOR U12194 ( .A(n12129), .B(n12130), .Z(n12128) );
  NANDN U12195 ( .A(n12067), .B(n11869), .Z(n12130) );
  IV U12196 ( .A(n12112), .Z(n12118) );
  XNOR U12197 ( .A(n12131), .B(n12129), .Z(n12112) );
  NANDN U12198 ( .A(n12078), .B(n12070), .Z(n12129) );
  XOR U12199 ( .A(n12058), .B(n11655), .Z(n12067) );
  XOR U12200 ( .A(n12132), .B(n12133), .Z(n11655) );
  XNOR U12201 ( .A(n12134), .B(n12135), .Z(n12133) );
  XOR U12202 ( .A(n12086), .B(n11869), .Z(n12078) );
  XNOR U12203 ( .A(n11874), .B(n12075), .Z(n11869) );
  XNOR U12204 ( .A(n12135), .B(n12136), .Z(n12075) );
  ANDN U12205 ( .B(n12072), .A(n12086), .Z(n12131) );
  XNOR U12206 ( .A(n12137), .B(n12109), .Z(n12086) );
  IV U12207 ( .A(n11862), .Z(n12109) );
  XNOR U12208 ( .A(n12138), .B(n12139), .Z(n11862) );
  XNOR U12209 ( .A(n12140), .B(n12135), .Z(n12139) );
  XOR U12210 ( .A(n12141), .B(n12120), .Z(n12072) );
  XNOR U12211 ( .A(n12124), .B(n12142), .Z(n12125) );
  XNOR U12212 ( .A(n12143), .B(n12123), .Z(n12142) );
  OR U12213 ( .A(n12062), .B(n11873), .Z(n12123) );
  XOR U12214 ( .A(n11741), .B(n11874), .Z(n11873) );
  IV U12215 ( .A(n12124), .Z(n11874) );
  XOR U12216 ( .A(n12061), .B(n12058), .Z(n12062) );
  XNOR U12217 ( .A(n12120), .B(n12144), .Z(n12058) );
  XNOR U12218 ( .A(n12134), .B(n12138), .Z(n12144) );
  XNOR U12219 ( .A(state[50]), .B(key[50]), .Z(n12138) );
  IV U12220 ( .A(n12054), .Z(n12120) );
  XOR U12221 ( .A(n12132), .B(n12145), .Z(n12054) );
  XOR U12222 ( .A(n12135), .B(n12146), .Z(n12145) );
  IV U12223 ( .A(n12141), .Z(n12061) );
  ANDN U12224 ( .B(n12141), .A(n11741), .Z(n12143) );
  XOR U12225 ( .A(n12136), .B(n12147), .Z(n12141) );
  XNOR U12226 ( .A(n12135), .B(n12148), .Z(n12147) );
  XOR U12227 ( .A(n12137), .B(n12149), .Z(n12135) );
  XNOR U12228 ( .A(state[54]), .B(key[54]), .Z(n12149) );
  IV U12229 ( .A(n12132), .Z(n12136) );
  XOR U12230 ( .A(state[53]), .B(key[53]), .Z(n12132) );
  XOR U12231 ( .A(n12150), .B(n12151), .Z(n12124) );
  XOR U12232 ( .A(n12148), .B(n12146), .Z(n12151) );
  XOR U12233 ( .A(state[55]), .B(key[55]), .Z(n12146) );
  XNOR U12234 ( .A(state[52]), .B(key[52]), .Z(n12148) );
  XOR U12235 ( .A(n11741), .B(n12140), .Z(n12150) );
  XNOR U12236 ( .A(n12134), .B(n12152), .Z(n12140) );
  XNOR U12237 ( .A(state[51]), .B(key[51]), .Z(n12152) );
  XNOR U12238 ( .A(state[49]), .B(key[49]), .Z(n12134) );
  IV U12239 ( .A(n12137), .Z(n11741) );
  XOR U12240 ( .A(state[48]), .B(key[48]), .Z(n12137) );
  XOR U12241 ( .A(n12153), .B(n12154), .Z(n9403) );
  XNOR U12242 ( .A(n11723), .B(n11775), .Z(n12154) );
  XNOR U12243 ( .A(n12155), .B(n12156), .Z(n11775) );
  XNOR U12244 ( .A(n12157), .B(n11713), .Z(n12156) );
  NOR U12245 ( .A(n12158), .B(n12159), .Z(n11713) );
  NOR U12246 ( .A(n12160), .B(n11849), .Z(n12157) );
  XNOR U12247 ( .A(n12155), .B(n12161), .Z(n11723) );
  XOR U12248 ( .A(n12162), .B(n12163), .Z(n12161) );
  ANDN U12249 ( .B(n12164), .A(n11728), .Z(n12162) );
  XNOR U12250 ( .A(n11709), .B(n12165), .Z(n12155) );
  XNOR U12251 ( .A(n12166), .B(n12167), .Z(n12165) );
  NAND U12252 ( .A(n12168), .B(n11855), .Z(n12167) );
  XNOR U12253 ( .A(n11778), .B(n11731), .Z(n12153) );
  XNOR U12254 ( .A(n11709), .B(n12169), .Z(n11778) );
  XNOR U12255 ( .A(n12163), .B(n12170), .Z(n12169) );
  NANDN U12256 ( .A(n12171), .B(n12172), .Z(n12170) );
  OR U12257 ( .A(n12173), .B(n12174), .Z(n12163) );
  XOR U12258 ( .A(n12175), .B(n12166), .Z(n11709) );
  NANDN U12259 ( .A(n12176), .B(n12177), .Z(n12166) );
  AND U12260 ( .A(n12178), .B(n12179), .Z(n12175) );
  XOR U12261 ( .A(key[210]), .B(n9444), .Z(n11876) );
  XOR U12262 ( .A(n11777), .B(n11731), .Z(n9444) );
  XOR U12263 ( .A(n11851), .B(n12180), .Z(n11731) );
  XNOR U12264 ( .A(n11847), .B(n12181), .Z(n12180) );
  NANDN U12265 ( .A(n12182), .B(n12183), .Z(n12181) );
  OR U12266 ( .A(n12184), .B(n12158), .Z(n11847) );
  XOR U12267 ( .A(n11849), .B(n12183), .Z(n12158) );
  IV U12268 ( .A(n11845), .Z(n11777) );
  XNOR U12269 ( .A(n11851), .B(n12185), .Z(n11845) );
  XOR U12270 ( .A(n12186), .B(n11726), .Z(n12185) );
  OR U12271 ( .A(n12187), .B(n12173), .Z(n11726) );
  XNOR U12272 ( .A(n11728), .B(n12171), .Z(n12173) );
  NOR U12273 ( .A(n12188), .B(n12171), .Z(n12186) );
  XOR U12274 ( .A(n12189), .B(n11853), .Z(n11851) );
  OR U12275 ( .A(n12176), .B(n12190), .Z(n11853) );
  XNOR U12276 ( .A(n12178), .B(n11855), .Z(n12176) );
  XOR U12277 ( .A(n12171), .B(n11716), .Z(n11855) );
  IV U12278 ( .A(n12183), .Z(n11716) );
  XOR U12279 ( .A(n12191), .B(n12192), .Z(n12183) );
  NAND U12280 ( .A(n12193), .B(n12194), .Z(n12192) );
  XNOR U12281 ( .A(n12195), .B(n12196), .Z(n12171) );
  NANDN U12282 ( .A(n12197), .B(n12193), .Z(n12196) );
  ANDN U12283 ( .B(n12178), .A(n12198), .Z(n12189) );
  XOR U12284 ( .A(n11728), .B(n11849), .Z(n12178) );
  XNOR U12285 ( .A(n12191), .B(n12199), .Z(n11849) );
  NANDN U12286 ( .A(n12200), .B(n12201), .Z(n12199) );
  NAND U12287 ( .A(n12202), .B(n12203), .Z(n12191) );
  NANDN U12288 ( .A(n12205), .B(n12203), .Z(n12195) );
  XNOR U12289 ( .A(n12200), .B(n12193), .Z(n12203) );
  XNOR U12290 ( .A(n12206), .B(n12207), .Z(n12193) );
  XOR U12291 ( .A(n12208), .B(n12201), .Z(n12207) );
  IV U12292 ( .A(n12209), .Z(n12201) );
  XNOR U12293 ( .A(n12210), .B(n12211), .Z(n12206) );
  XNOR U12294 ( .A(n12212), .B(n12213), .Z(n12211) );
  NOR U12295 ( .A(n12209), .B(n12210), .Z(n12212) );
  NOR U12296 ( .A(n12200), .B(n12210), .Z(n12204) );
  XNOR U12297 ( .A(n12208), .B(n12214), .Z(n12200) );
  XNOR U12298 ( .A(n12213), .B(n12215), .Z(n12214) );
  NANDN U12299 ( .A(n12197), .B(n12194), .Z(n12215) );
  NANDN U12300 ( .A(n12205), .B(n12202), .Z(n12213) );
  XNOR U12301 ( .A(n12194), .B(n12209), .Z(n12202) );
  XOR U12302 ( .A(n12216), .B(n12217), .Z(n12209) );
  XOR U12303 ( .A(n12218), .B(n12219), .Z(n12217) );
  XOR U12304 ( .A(n12172), .B(n12220), .Z(n12219) );
  XNOR U12305 ( .A(n12188), .B(n12221), .Z(n12216) );
  XNOR U12306 ( .A(n12222), .B(n12223), .Z(n12221) );
  AND U12307 ( .A(n11729), .B(n12164), .Z(n12222) );
  XOR U12308 ( .A(n12224), .B(n12225), .Z(n12210) );
  XNOR U12309 ( .A(n12226), .B(n12220), .Z(n12225) );
  XNOR U12310 ( .A(n12227), .B(n12228), .Z(n12220) );
  XNOR U12311 ( .A(n12229), .B(n12230), .Z(n12228) );
  NAND U12312 ( .A(n11856), .B(n12168), .Z(n12230) );
  XNOR U12313 ( .A(n12231), .B(n12232), .Z(n12224) );
  ANDN U12314 ( .B(n12233), .A(n12160), .Z(n12231) );
  XOR U12315 ( .A(n12197), .B(n12194), .Z(n12208) );
  XNOR U12316 ( .A(n12234), .B(n12235), .Z(n12194) );
  XOR U12317 ( .A(n12236), .B(n12237), .Z(n12235) );
  XOR U12318 ( .A(n12226), .B(n12164), .Z(n12237) );
  XOR U12319 ( .A(n11729), .B(n12238), .Z(n12234) );
  XNOR U12320 ( .A(n12239), .B(n12223), .Z(n12238) );
  OR U12321 ( .A(n12174), .B(n12187), .Z(n12223) );
  XNOR U12322 ( .A(n11729), .B(n12240), .Z(n12187) );
  XNOR U12323 ( .A(n12164), .B(n12172), .Z(n12174) );
  ANDN U12324 ( .B(n12172), .A(n12188), .Z(n12239) );
  XOR U12325 ( .A(n12241), .B(n12242), .Z(n12197) );
  XOR U12326 ( .A(n12227), .B(n12218), .Z(n12242) );
  XOR U12327 ( .A(n12243), .B(n11715), .Z(n12218) );
  IV U12328 ( .A(n12236), .Z(n12227) );
  XNOR U12329 ( .A(n12244), .B(n12229), .Z(n12236) );
  NANDN U12330 ( .A(n12190), .B(n12177), .Z(n12229) );
  XOR U12331 ( .A(n12179), .B(n12168), .Z(n12177) );
  XOR U12332 ( .A(n11715), .B(n12172), .Z(n12168) );
  XNOR U12333 ( .A(n12245), .B(n12246), .Z(n12172) );
  XNOR U12334 ( .A(n12247), .B(n12248), .Z(n12246) );
  IV U12335 ( .A(n12249), .Z(n11715) );
  XOR U12336 ( .A(n12198), .B(n11856), .Z(n12190) );
  XNOR U12337 ( .A(n12240), .B(n12182), .Z(n11856) );
  IV U12338 ( .A(n12188), .Z(n12240) );
  XOR U12339 ( .A(n12250), .B(n12251), .Z(n12188) );
  XOR U12340 ( .A(n12252), .B(n12253), .Z(n12251) );
  XNOR U12341 ( .A(n11729), .B(n12254), .Z(n12250) );
  ANDN U12342 ( .B(n12179), .A(n12198), .Z(n12244) );
  XNOR U12343 ( .A(n11729), .B(n12233), .Z(n12198) );
  XOR U12344 ( .A(n12245), .B(n12164), .Z(n12179) );
  XNOR U12345 ( .A(n12255), .B(n12256), .Z(n12164) );
  XOR U12346 ( .A(n12257), .B(n12253), .Z(n12256) );
  XOR U12347 ( .A(state[12]), .B(key[12]), .Z(n12253) );
  IV U12348 ( .A(n12160), .Z(n12245) );
  XNOR U12349 ( .A(n12226), .B(n12258), .Z(n12241) );
  XNOR U12350 ( .A(n12259), .B(n12232), .Z(n12258) );
  OR U12351 ( .A(n12159), .B(n12184), .Z(n12232) );
  XNOR U12352 ( .A(n11850), .B(n12182), .Z(n12184) );
  IV U12353 ( .A(n12243), .Z(n12182) );
  XNOR U12354 ( .A(n12160), .B(n12249), .Z(n12159) );
  ANDN U12355 ( .B(n12243), .A(n12249), .Z(n12259) );
  XOR U12356 ( .A(n12255), .B(n12260), .Z(n12249) );
  XOR U12357 ( .A(n12248), .B(n12261), .Z(n12260) );
  XOR U12358 ( .A(n12233), .B(n12160), .Z(n12226) );
  XOR U12359 ( .A(n12255), .B(n12262), .Z(n12160) );
  XNOR U12360 ( .A(n12257), .B(n12252), .Z(n12262) );
  XNOR U12361 ( .A(state[15]), .B(key[15]), .Z(n12252) );
  XOR U12362 ( .A(state[13]), .B(key[13]), .Z(n12255) );
  IV U12363 ( .A(n11850), .Z(n12233) );
  XOR U12364 ( .A(n12261), .B(n12263), .Z(n11850) );
  XNOR U12365 ( .A(n12247), .B(n12254), .Z(n12263) );
  XNOR U12366 ( .A(n12248), .B(n12264), .Z(n12254) );
  XNOR U12367 ( .A(state[11]), .B(key[11]), .Z(n12264) );
  XNOR U12368 ( .A(state[9]), .B(key[9]), .Z(n12248) );
  XNOR U12369 ( .A(state[10]), .B(key[10]), .Z(n12247) );
  IV U12370 ( .A(n12257), .Z(n12261) );
  XOR U12371 ( .A(n11729), .B(n12265), .Z(n12257) );
  XNOR U12372 ( .A(state[14]), .B(key[14]), .Z(n12265) );
  XOR U12373 ( .A(state[8]), .B(key[8]), .Z(n11729) );
  XOR U12374 ( .A(n11408), .B(n11409), .Z(n11364) );
  XNOR U12375 ( .A(n11505), .B(n12266), .Z(n11408) );
  XNOR U12376 ( .A(n12267), .B(n12268), .Z(n12266) );
  ANDN U12377 ( .B(n12269), .A(n12270), .Z(n12267) );
  XNOR U12378 ( .A(n12271), .B(n12272), .Z(n11505) );
  XNOR U12379 ( .A(n12273), .B(n12274), .Z(n12272) );
  NANDN U12380 ( .A(n12275), .B(n12276), .Z(n12274) );
  XNOR U12381 ( .A(n6104), .B(n6112), .Z(n6919) );
  XNOR U12382 ( .A(n11511), .B(n12277), .Z(n6112) );
  XNOR U12383 ( .A(n11415), .B(n11512), .Z(n12277) );
  XNOR U12384 ( .A(n12279), .B(n12280), .Z(n12278) );
  NANDN U12385 ( .A(n12281), .B(n11510), .Z(n12280) );
  XOR U12386 ( .A(n12271), .B(n12283), .Z(n11511) );
  XOR U12387 ( .A(n12268), .B(n12284), .Z(n12283) );
  NANDN U12388 ( .A(n12285), .B(n11491), .Z(n12284) );
  IV U12389 ( .A(n7794), .Z(n6104) );
  XOR U12390 ( .A(n11407), .B(n12288), .Z(n7794) );
  XNOR U12391 ( .A(n11388), .B(n11493), .Z(n12288) );
  XNOR U12392 ( .A(key[352]), .B(n7764), .Z(n11558) );
  XOR U12393 ( .A(n11393), .B(n11363), .Z(n7764) );
  XNOR U12394 ( .A(n11474), .B(n12289), .Z(n11363) );
  XOR U12395 ( .A(n12290), .B(n11454), .Z(n12289) );
  XOR U12396 ( .A(n11540), .B(n11457), .Z(n11538) );
  ANDN U12397 ( .B(n11540), .A(n12292), .Z(n12290) );
  XNOR U12398 ( .A(n11452), .B(n12293), .Z(n11474) );
  XNOR U12399 ( .A(n12294), .B(n12295), .Z(n12293) );
  NAND U12400 ( .A(n11546), .B(n12296), .Z(n12295) );
  XOR U12401 ( .A(n11452), .B(n12297), .Z(n11393) );
  XOR U12402 ( .A(n12298), .B(n11476), .Z(n12297) );
  OR U12403 ( .A(n11551), .B(n12299), .Z(n11476) );
  XNOR U12404 ( .A(n11450), .B(n11549), .Z(n11551) );
  NOR U12405 ( .A(n12300), .B(n11549), .Z(n12298) );
  XOR U12406 ( .A(n12301), .B(n12294), .Z(n11452) );
  OR U12407 ( .A(n11554), .B(n12302), .Z(n12294) );
  XOR U12408 ( .A(n11557), .B(n11546), .Z(n11554) );
  XNOR U12409 ( .A(n11549), .B(n11457), .Z(n11546) );
  XOR U12410 ( .A(n12303), .B(n12304), .Z(n11457) );
  NANDN U12411 ( .A(n12305), .B(n12306), .Z(n12304) );
  XNOR U12412 ( .A(n12307), .B(n12308), .Z(n11549) );
  OR U12413 ( .A(n12305), .B(n12309), .Z(n12308) );
  ANDN U12414 ( .B(n12310), .A(n11557), .Z(n12301) );
  XOR U12415 ( .A(n11450), .B(n11540), .Z(n11557) );
  XNOR U12416 ( .A(n12311), .B(n12303), .Z(n11540) );
  NANDN U12417 ( .A(n12312), .B(n12313), .Z(n12303) );
  ANDN U12418 ( .B(n12314), .A(n12315), .Z(n12311) );
  NANDN U12419 ( .A(n12312), .B(n12317), .Z(n12307) );
  XOR U12420 ( .A(n12318), .B(n12305), .Z(n12312) );
  XNOR U12421 ( .A(n12319), .B(n12320), .Z(n12305) );
  XOR U12422 ( .A(n12321), .B(n12314), .Z(n12320) );
  XNOR U12423 ( .A(n12322), .B(n12323), .Z(n12319) );
  XNOR U12424 ( .A(n12324), .B(n12325), .Z(n12323) );
  ANDN U12425 ( .B(n12314), .A(n12326), .Z(n12324) );
  IV U12426 ( .A(n12327), .Z(n12314) );
  ANDN U12427 ( .B(n12318), .A(n12326), .Z(n12316) );
  IV U12428 ( .A(n12322), .Z(n12326) );
  IV U12429 ( .A(n12315), .Z(n12318) );
  XNOR U12430 ( .A(n12321), .B(n12328), .Z(n12315) );
  XOR U12431 ( .A(n12329), .B(n12325), .Z(n12328) );
  NAND U12432 ( .A(n12317), .B(n12313), .Z(n12325) );
  XNOR U12433 ( .A(n12306), .B(n12327), .Z(n12313) );
  XOR U12434 ( .A(n12330), .B(n12331), .Z(n12327) );
  XOR U12435 ( .A(n12332), .B(n12333), .Z(n12331) );
  XNOR U12436 ( .A(n11550), .B(n12334), .Z(n12333) );
  XNOR U12437 ( .A(n12335), .B(n12336), .Z(n12330) );
  XNOR U12438 ( .A(n12337), .B(n12338), .Z(n12336) );
  ANDN U12439 ( .B(n11451), .A(n11478), .Z(n12337) );
  XNOR U12440 ( .A(n12322), .B(n12309), .Z(n12317) );
  XOR U12441 ( .A(n12339), .B(n12340), .Z(n12322) );
  XNOR U12442 ( .A(n12341), .B(n12334), .Z(n12340) );
  XOR U12443 ( .A(n12342), .B(n12343), .Z(n12334) );
  XNOR U12444 ( .A(n12344), .B(n12345), .Z(n12343) );
  NAND U12445 ( .A(n12296), .B(n11545), .Z(n12345) );
  XNOR U12446 ( .A(n12346), .B(n12347), .Z(n12339) );
  ANDN U12447 ( .B(n12348), .A(n12292), .Z(n12346) );
  ANDN U12448 ( .B(n12306), .A(n12309), .Z(n12329) );
  XOR U12449 ( .A(n12309), .B(n12306), .Z(n12321) );
  XNOR U12450 ( .A(n12349), .B(n12350), .Z(n12306) );
  XNOR U12451 ( .A(n12342), .B(n12351), .Z(n12350) );
  XNOR U12452 ( .A(n12341), .B(n11451), .Z(n12351) );
  XNOR U12453 ( .A(n12352), .B(n12353), .Z(n12349) );
  XNOR U12454 ( .A(n12354), .B(n12338), .Z(n12353) );
  OR U12455 ( .A(n11552), .B(n12299), .Z(n12338) );
  XNOR U12456 ( .A(n12352), .B(n12335), .Z(n12299) );
  XNOR U12457 ( .A(n11451), .B(n11550), .Z(n11552) );
  ANDN U12458 ( .B(n11550), .A(n12300), .Z(n12354) );
  XOR U12459 ( .A(n12355), .B(n12356), .Z(n12309) );
  XOR U12460 ( .A(n12342), .B(n12332), .Z(n12356) );
  XOR U12461 ( .A(n11456), .B(n11483), .Z(n12332) );
  XOR U12462 ( .A(n12357), .B(n12344), .Z(n12342) );
  NANDN U12463 ( .A(n12302), .B(n11555), .Z(n12344) );
  XOR U12464 ( .A(n11556), .B(n11545), .Z(n11555) );
  XNOR U12465 ( .A(n12348), .B(n12358), .Z(n11550) );
  XNOR U12466 ( .A(n12359), .B(n12360), .Z(n12358) );
  XNOR U12467 ( .A(n12310), .B(n12296), .Z(n12302) );
  XNOR U12468 ( .A(n12300), .B(n11456), .Z(n12296) );
  IV U12469 ( .A(n12335), .Z(n12300) );
  XOR U12470 ( .A(n12361), .B(n12362), .Z(n12335) );
  XOR U12471 ( .A(n12363), .B(n12364), .Z(n12362) );
  XOR U12472 ( .A(n12352), .B(n12365), .Z(n12361) );
  AND U12473 ( .A(n11556), .B(n12310), .Z(n12357) );
  XOR U12474 ( .A(n12348), .B(n11451), .Z(n11556) );
  XNOR U12475 ( .A(n12366), .B(n12367), .Z(n11451) );
  XOR U12476 ( .A(n12368), .B(n12364), .Z(n12367) );
  XNOR U12477 ( .A(n12369), .B(n12370), .Z(n12364) );
  XNOR U12478 ( .A(n10986), .B(n9279), .Z(n12370) );
  XOR U12479 ( .A(n12371), .B(n12372), .Z(n9279) );
  XNOR U12480 ( .A(n10191), .B(n9281), .Z(n10986) );
  XOR U12481 ( .A(n12373), .B(n9252), .Z(n9281) );
  XNOR U12482 ( .A(n10187), .B(n12374), .Z(n12369) );
  XNOR U12483 ( .A(key[172]), .B(n10987), .Z(n12374) );
  XOR U12484 ( .A(n12375), .B(n10206), .Z(n10987) );
  XOR U12485 ( .A(n12376), .B(n12377), .Z(n10206) );
  XOR U12486 ( .A(n12378), .B(n12379), .Z(n12377) );
  XNOR U12487 ( .A(n12380), .B(n12381), .Z(n12376) );
  XOR U12488 ( .A(n12382), .B(n12383), .Z(n12381) );
  ANDN U12489 ( .B(n12384), .A(n12385), .Z(n12383) );
  XOR U12490 ( .A(n12386), .B(n10225), .Z(n10187) );
  IV U12491 ( .A(n11541), .Z(n12348) );
  XOR U12492 ( .A(n12341), .B(n12387), .Z(n12355) );
  XNOR U12493 ( .A(n12388), .B(n12347), .Z(n12387) );
  OR U12494 ( .A(n11539), .B(n12291), .Z(n12347) );
  XNOR U12495 ( .A(n12389), .B(n11456), .Z(n12291) );
  XNOR U12496 ( .A(n11541), .B(n11483), .Z(n11539) );
  ANDN U12497 ( .B(n11456), .A(n11483), .Z(n12388) );
  XOR U12498 ( .A(n12366), .B(n12390), .Z(n11483) );
  XOR U12499 ( .A(n12359), .B(n12391), .Z(n12390) );
  XOR U12500 ( .A(n12368), .B(n12366), .Z(n11456) );
  XNOR U12501 ( .A(n12292), .B(n11541), .Z(n12341) );
  XOR U12502 ( .A(n12366), .B(n12392), .Z(n11541) );
  XNOR U12503 ( .A(n12368), .B(n12363), .Z(n12392) );
  XOR U12504 ( .A(n12393), .B(n12394), .Z(n12363) );
  XOR U12505 ( .A(n10201), .B(n10982), .Z(n12394) );
  XOR U12506 ( .A(n10199), .B(n10215), .Z(n10982) );
  XNOR U12507 ( .A(n12395), .B(n12396), .Z(n10215) );
  XOR U12508 ( .A(n12397), .B(n12398), .Z(n12396) );
  XOR U12509 ( .A(n12399), .B(n12400), .Z(n12395) );
  XNOR U12510 ( .A(n12401), .B(n12402), .Z(n10201) );
  XOR U12511 ( .A(n12403), .B(n12404), .Z(n12402) );
  XOR U12512 ( .A(n12405), .B(n12406), .Z(n12401) );
  XNOR U12513 ( .A(key[175]), .B(n10239), .Z(n12393) );
  IV U12514 ( .A(n10993), .Z(n10239) );
  XNOR U12515 ( .A(n9276), .B(n9298), .Z(n10993) );
  IV U12516 ( .A(n12375), .Z(n9298) );
  XNOR U12517 ( .A(n12407), .B(n12408), .Z(n12366) );
  XOR U12518 ( .A(n10207), .B(n10999), .Z(n12408) );
  XNOR U12519 ( .A(n12372), .B(n9267), .Z(n10999) );
  XNOR U12520 ( .A(n12409), .B(n12410), .Z(n9267) );
  XNOR U12521 ( .A(n12411), .B(n12398), .Z(n12410) );
  XNOR U12522 ( .A(n12412), .B(n12413), .Z(n12398) );
  XNOR U12523 ( .A(n12414), .B(n12415), .Z(n12413) );
  OR U12524 ( .A(n12416), .B(n12417), .Z(n12415) );
  XNOR U12525 ( .A(n12373), .B(n12418), .Z(n12409) );
  XOR U12526 ( .A(n12419), .B(n12420), .Z(n12418) );
  ANDN U12527 ( .B(n12421), .A(n12422), .Z(n12420) );
  IV U12528 ( .A(n10205), .Z(n12372) );
  XOR U12529 ( .A(n12423), .B(n12424), .Z(n10205) );
  XNOR U12530 ( .A(n12425), .B(n12426), .Z(n12424) );
  XNOR U12531 ( .A(n12427), .B(n12428), .Z(n12423) );
  XOR U12532 ( .A(n12429), .B(n12430), .Z(n12428) );
  ANDN U12533 ( .B(n12431), .A(n12432), .Z(n12430) );
  XNOR U12534 ( .A(n12433), .B(n12434), .Z(n10207) );
  XNOR U12535 ( .A(n12435), .B(n12404), .Z(n12434) );
  XNOR U12536 ( .A(n12436), .B(n12437), .Z(n12404) );
  XNOR U12537 ( .A(n12438), .B(n12439), .Z(n12437) );
  NANDN U12538 ( .A(n12440), .B(n12441), .Z(n12439) );
  XNOR U12539 ( .A(n12386), .B(n12442), .Z(n12433) );
  XOR U12540 ( .A(n12443), .B(n12444), .Z(n12442) );
  ANDN U12541 ( .B(n12445), .A(n12446), .Z(n12444) );
  XOR U12542 ( .A(n10994), .B(n12447), .Z(n12407) );
  XNOR U12543 ( .A(key[173]), .B(n10218), .Z(n12447) );
  XOR U12544 ( .A(n12448), .B(n12449), .Z(n10994) );
  XOR U12545 ( .A(n11478), .B(n12292), .Z(n12310) );
  IV U12546 ( .A(n12389), .Z(n12292) );
  XNOR U12547 ( .A(n12360), .B(n12450), .Z(n12389) );
  XOR U12548 ( .A(n12365), .B(n12391), .Z(n12450) );
  IV U12549 ( .A(n12368), .Z(n12391) );
  XOR U12550 ( .A(n12451), .B(n12452), .Z(n12368) );
  XNOR U12551 ( .A(n10996), .B(n9262), .Z(n12452) );
  XOR U12552 ( .A(n9276), .B(n10199), .Z(n9262) );
  XOR U12553 ( .A(n12453), .B(n12454), .Z(n10199) );
  XOR U12554 ( .A(n12455), .B(n12426), .Z(n12454) );
  XNOR U12555 ( .A(n12456), .B(n12457), .Z(n12426) );
  XNOR U12556 ( .A(n12458), .B(n12459), .Z(n12457) );
  OR U12557 ( .A(n12460), .B(n12461), .Z(n12459) );
  XOR U12558 ( .A(n12462), .B(n12463), .Z(n12453) );
  XNOR U12559 ( .A(n9269), .B(n10981), .Z(n10996) );
  XOR U12560 ( .A(n12375), .B(n10200), .Z(n10981) );
  XOR U12561 ( .A(n12464), .B(n12465), .Z(n10200) );
  XNOR U12562 ( .A(n12448), .B(n12379), .Z(n12465) );
  XNOR U12563 ( .A(n12466), .B(n12467), .Z(n12379) );
  XNOR U12564 ( .A(n12468), .B(n12469), .Z(n12467) );
  NANDN U12565 ( .A(n12470), .B(n12471), .Z(n12469) );
  XOR U12566 ( .A(n12472), .B(n12473), .Z(n12464) );
  XNOR U12567 ( .A(n10218), .B(n9264), .Z(n9269) );
  XOR U12568 ( .A(n12474), .B(n12397), .Z(n9264) );
  XOR U12569 ( .A(n12463), .B(n12475), .Z(n10218) );
  XNOR U12570 ( .A(n10209), .B(n12476), .Z(n12451) );
  XNOR U12571 ( .A(key[174]), .B(n12352), .Z(n12476) );
  XOR U12572 ( .A(n12477), .B(n12403), .Z(n10209) );
  XOR U12573 ( .A(n12478), .B(n12479), .Z(n12365) );
  XNOR U12574 ( .A(n9292), .B(n12480), .Z(n12479) );
  XNOR U12575 ( .A(n12359), .B(n10976), .Z(n12480) );
  XOR U12576 ( .A(n12375), .B(n10186), .Z(n10976) );
  XOR U12577 ( .A(n10963), .B(n12378), .Z(n10186) );
  XNOR U12578 ( .A(n12481), .B(n12378), .Z(n12375) );
  XOR U12579 ( .A(n12466), .B(n12482), .Z(n12378) );
  XOR U12580 ( .A(n12483), .B(n12484), .Z(n12482) );
  NOR U12581 ( .A(n12485), .B(n12486), .Z(n12483) );
  XNOR U12582 ( .A(n12487), .B(n12488), .Z(n12466) );
  XNOR U12583 ( .A(n12489), .B(n12490), .Z(n12488) );
  NANDN U12584 ( .A(n12491), .B(n12492), .Z(n12490) );
  XOR U12585 ( .A(n12493), .B(n12494), .Z(n12359) );
  XOR U12586 ( .A(n10963), .B(n9297), .Z(n12494) );
  IV U12587 ( .A(n10973), .Z(n9297) );
  XNOR U12588 ( .A(n10227), .B(n10238), .Z(n10973) );
  IV U12589 ( .A(n9291), .Z(n10238) );
  XOR U12590 ( .A(n12397), .B(n12495), .Z(n9291) );
  IV U12591 ( .A(n12498), .Z(n10227) );
  XOR U12592 ( .A(n12472), .B(n12481), .Z(n10963) );
  IV U12593 ( .A(n12499), .Z(n12472) );
  XOR U12594 ( .A(n10240), .B(n12500), .Z(n12493) );
  XOR U12595 ( .A(key[169]), .B(n10233), .Z(n12500) );
  XNOR U12596 ( .A(n12403), .B(n12501), .Z(n10240) );
  XNOR U12597 ( .A(n12405), .B(n12406), .Z(n12501) );
  XOR U12598 ( .A(n12502), .B(n12503), .Z(n12403) );
  XOR U12599 ( .A(n9276), .B(n10191), .Z(n9292) );
  XOR U12600 ( .A(n12427), .B(n10233), .Z(n10191) );
  XNOR U12601 ( .A(n10234), .B(n12504), .Z(n12478) );
  XOR U12602 ( .A(key[171]), .B(n9254), .Z(n12504) );
  XOR U12603 ( .A(n10230), .B(n9294), .Z(n9254) );
  XOR U12604 ( .A(n12505), .B(n12506), .Z(n9294) );
  XNOR U12605 ( .A(n12399), .B(n12400), .Z(n12506) );
  XOR U12606 ( .A(n12507), .B(n12508), .Z(n12400) );
  XNOR U12607 ( .A(n12509), .B(n12510), .Z(n12508) );
  OR U12608 ( .A(n12416), .B(n12511), .Z(n12510) );
  XNOR U12609 ( .A(n12496), .B(n12474), .Z(n12505) );
  XNOR U12610 ( .A(n12507), .B(n12512), .Z(n12474) );
  XNOR U12611 ( .A(n12513), .B(n12419), .Z(n12512) );
  NOR U12612 ( .A(n12514), .B(n12515), .Z(n12419) );
  NOR U12613 ( .A(n12516), .B(n12517), .Z(n12513) );
  XNOR U12614 ( .A(n12411), .B(n12518), .Z(n12507) );
  XNOR U12615 ( .A(n12519), .B(n12520), .Z(n12518) );
  OR U12616 ( .A(n12521), .B(n12522), .Z(n12520) );
  XOR U12617 ( .A(n12411), .B(n12523), .Z(n12496) );
  XNOR U12618 ( .A(n12509), .B(n12524), .Z(n12523) );
  NANDN U12619 ( .A(n12525), .B(n12526), .Z(n12524) );
  OR U12620 ( .A(n12527), .B(n12528), .Z(n12509) );
  XOR U12621 ( .A(n12529), .B(n12519), .Z(n12411) );
  NANDN U12622 ( .A(n12530), .B(n12531), .Z(n12519) );
  AND U12623 ( .A(n12532), .B(n12533), .Z(n12529) );
  XOR U12624 ( .A(n12534), .B(n12535), .Z(n10234) );
  XOR U12625 ( .A(n12406), .B(n12477), .Z(n12535) );
  XNOR U12626 ( .A(n12536), .B(n12537), .Z(n12477) );
  XNOR U12627 ( .A(n12538), .B(n12443), .Z(n12537) );
  NOR U12628 ( .A(n12539), .B(n12540), .Z(n12443) );
  NOR U12629 ( .A(n12541), .B(n12542), .Z(n12538) );
  XOR U12630 ( .A(n12405), .B(n12503), .Z(n12534) );
  XOR U12631 ( .A(n12435), .B(n12543), .Z(n12503) );
  XNOR U12632 ( .A(n12544), .B(n12545), .Z(n12543) );
  OR U12633 ( .A(n12546), .B(n12547), .Z(n12545) );
  XNOR U12634 ( .A(n12544), .B(n12549), .Z(n12548) );
  NANDN U12635 ( .A(n12440), .B(n12550), .Z(n12549) );
  OR U12636 ( .A(n12551), .B(n12552), .Z(n12544) );
  XNOR U12637 ( .A(n12435), .B(n12553), .Z(n12536) );
  XNOR U12638 ( .A(n12554), .B(n12555), .Z(n12553) );
  NANDN U12639 ( .A(n12556), .B(n12557), .Z(n12555) );
  XOR U12640 ( .A(n12558), .B(n12554), .Z(n12435) );
  NANDN U12641 ( .A(n12559), .B(n12560), .Z(n12554) );
  AND U12642 ( .A(n12561), .B(n12562), .Z(n12558) );
  XOR U12643 ( .A(n12563), .B(n12564), .Z(n12360) );
  XOR U12644 ( .A(n9289), .B(n10225), .Z(n12564) );
  XOR U12645 ( .A(n12502), .B(n12406), .Z(n10225) );
  XOR U12646 ( .A(n12565), .B(n12566), .Z(n12406) );
  XNOR U12647 ( .A(n12567), .B(n12568), .Z(n12566) );
  NANDN U12648 ( .A(n12569), .B(n12570), .Z(n12568) );
  IV U12649 ( .A(n12571), .Z(n12502) );
  XNOR U12650 ( .A(n10233), .B(n9252), .Z(n9289) );
  XNOR U12651 ( .A(n12497), .B(n12399), .Z(n9252) );
  XOR U12652 ( .A(n12572), .B(n12573), .Z(n12399) );
  XNOR U12653 ( .A(n12574), .B(n12575), .Z(n12573) );
  NANDN U12654 ( .A(n12576), .B(n12421), .Z(n12575) );
  XOR U12655 ( .A(n12577), .B(n12455), .Z(n10233) );
  XOR U12656 ( .A(n10962), .B(n12578), .Z(n12563) );
  XNOR U12657 ( .A(key[170]), .B(n10230), .Z(n12578) );
  XOR U12658 ( .A(n12579), .B(n12580), .Z(n10230) );
  XOR U12659 ( .A(n12455), .B(n12475), .Z(n12580) );
  XNOR U12660 ( .A(n12581), .B(n12582), .Z(n12475) );
  XNOR U12661 ( .A(n12583), .B(n12429), .Z(n12582) );
  NOR U12662 ( .A(n12584), .B(n12585), .Z(n12429) );
  NOR U12663 ( .A(n12586), .B(n12587), .Z(n12583) );
  XOR U12664 ( .A(n12462), .B(n12588), .Z(n12579) );
  XNOR U12665 ( .A(n12589), .B(n12590), .Z(n10962) );
  XOR U12666 ( .A(n12591), .B(n12449), .Z(n12590) );
  XNOR U12667 ( .A(n12592), .B(n12593), .Z(n12449) );
  XNOR U12668 ( .A(n12594), .B(n12382), .Z(n12593) );
  NOR U12669 ( .A(n12595), .B(n12596), .Z(n12382) );
  NOR U12670 ( .A(n12597), .B(n12486), .Z(n12594) );
  XNOR U12671 ( .A(n12499), .B(n12473), .Z(n12589) );
  IV U12672 ( .A(n12352), .Z(n11478) );
  XOR U12673 ( .A(n12598), .B(n12599), .Z(n12352) );
  XOR U12674 ( .A(n12498), .B(n10202), .Z(n12599) );
  IV U12675 ( .A(n9299), .Z(n10202) );
  XNOR U12676 ( .A(n10214), .B(n10242), .Z(n9299) );
  XOR U12677 ( .A(n12571), .B(n12386), .Z(n10242) );
  XNOR U12678 ( .A(n12436), .B(n12600), .Z(n12386) );
  XOR U12679 ( .A(n12601), .B(n12567), .Z(n12600) );
  OR U12680 ( .A(n12602), .B(n12539), .Z(n12567) );
  XOR U12681 ( .A(n12542), .B(n12570), .Z(n12539) );
  NOR U12682 ( .A(n12603), .B(n12542), .Z(n12601) );
  XNOR U12683 ( .A(n12565), .B(n12604), .Z(n12436) );
  XNOR U12684 ( .A(n12605), .B(n12606), .Z(n12604) );
  NANDN U12685 ( .A(n12556), .B(n12607), .Z(n12606) );
  XNOR U12686 ( .A(n12565), .B(n12608), .Z(n12571) );
  XOR U12687 ( .A(n12609), .B(n12438), .Z(n12608) );
  OR U12688 ( .A(n12610), .B(n12551), .Z(n12438) );
  XNOR U12689 ( .A(n12440), .B(n12546), .Z(n12551) );
  NOR U12690 ( .A(n12611), .B(n12546), .Z(n12609) );
  XOR U12691 ( .A(n12612), .B(n12605), .Z(n12565) );
  OR U12692 ( .A(n12559), .B(n12613), .Z(n12605) );
  XOR U12693 ( .A(n12546), .B(n12570), .Z(n12556) );
  IV U12694 ( .A(n12446), .Z(n12570) );
  XNOR U12695 ( .A(n12614), .B(n12615), .Z(n12446) );
  NANDN U12696 ( .A(n12616), .B(n12617), .Z(n12615) );
  XNOR U12697 ( .A(n12618), .B(n12619), .Z(n12546) );
  NANDN U12698 ( .A(n12616), .B(n12620), .Z(n12619) );
  ANDN U12699 ( .B(n12561), .A(n12621), .Z(n12612) );
  XOR U12700 ( .A(n12440), .B(n12542), .Z(n12561) );
  XOR U12701 ( .A(n12622), .B(n12614), .Z(n12542) );
  NANDN U12702 ( .A(n12623), .B(n12624), .Z(n12614) );
  XOR U12703 ( .A(n12617), .B(n12625), .Z(n12624) );
  ANDN U12704 ( .B(n12625), .A(n12626), .Z(n12622) );
  NANDN U12705 ( .A(n12623), .B(n12628), .Z(n12618) );
  XOR U12706 ( .A(n12629), .B(n12630), .Z(n12616) );
  XOR U12707 ( .A(n12631), .B(n12632), .Z(n12630) );
  XNOR U12708 ( .A(n12633), .B(n12634), .Z(n12629) );
  XNOR U12709 ( .A(n12635), .B(n12636), .Z(n12634) );
  ANDN U12710 ( .B(n12632), .A(n12631), .Z(n12635) );
  ANDN U12711 ( .B(n12632), .A(n12626), .Z(n12627) );
  XNOR U12712 ( .A(n12633), .B(n12637), .Z(n12626) );
  XOR U12713 ( .A(n12638), .B(n12636), .Z(n12637) );
  NAND U12714 ( .A(n12628), .B(n12639), .Z(n12636) );
  XNOR U12715 ( .A(n12617), .B(n12631), .Z(n12639) );
  IV U12716 ( .A(n12625), .Z(n12631) );
  XNOR U12717 ( .A(n12640), .B(n12641), .Z(n12625) );
  XNOR U12718 ( .A(n12642), .B(n12643), .Z(n12641) );
  XOR U12719 ( .A(n12547), .B(n12644), .Z(n12643) );
  XNOR U12720 ( .A(n12611), .B(n12645), .Z(n12640) );
  XNOR U12721 ( .A(n12646), .B(n12647), .Z(n12645) );
  AND U12722 ( .A(n12550), .B(n12441), .Z(n12646) );
  XOR U12723 ( .A(n12620), .B(n12632), .Z(n12628) );
  AND U12724 ( .A(n12617), .B(n12620), .Z(n12638) );
  XNOR U12725 ( .A(n12617), .B(n12620), .Z(n12633) );
  XNOR U12726 ( .A(n12648), .B(n12649), .Z(n12620) );
  XNOR U12727 ( .A(n12650), .B(n12644), .Z(n12649) );
  XOR U12728 ( .A(n12651), .B(n12652), .Z(n12648) );
  XNOR U12729 ( .A(n12653), .B(n12654), .Z(n12652) );
  ANDN U12730 ( .B(n12445), .A(n12569), .Z(n12653) );
  XNOR U12731 ( .A(n12655), .B(n12656), .Z(n12617) );
  XNOR U12732 ( .A(n12550), .B(n12651), .Z(n12657) );
  XOR U12733 ( .A(n12441), .B(n12658), .Z(n12655) );
  XNOR U12734 ( .A(n12659), .B(n12647), .Z(n12658) );
  OR U12735 ( .A(n12552), .B(n12610), .Z(n12647) );
  XOR U12736 ( .A(n12441), .B(n12611), .Z(n12610) );
  XNOR U12737 ( .A(n12550), .B(n12660), .Z(n12552) );
  ANDN U12738 ( .B(n12661), .A(n12547), .Z(n12659) );
  XNOR U12739 ( .A(n12662), .B(n12663), .Z(n12632) );
  XOR U12740 ( .A(n12650), .B(n12642), .Z(n12663) );
  XOR U12741 ( .A(n12651), .B(n12664), .Z(n12642) );
  XNOR U12742 ( .A(n12665), .B(n12666), .Z(n12664) );
  NAND U12743 ( .A(n12607), .B(n12557), .Z(n12666) );
  XNOR U12744 ( .A(n12667), .B(n12665), .Z(n12651) );
  NANDN U12745 ( .A(n12613), .B(n12560), .Z(n12665) );
  XOR U12746 ( .A(n12562), .B(n12557), .Z(n12560) );
  XOR U12747 ( .A(n12660), .B(n12445), .Z(n12557) );
  IV U12748 ( .A(n12547), .Z(n12660) );
  XOR U12749 ( .A(n12668), .B(n12669), .Z(n12547) );
  XNOR U12750 ( .A(n12670), .B(n12671), .Z(n12669) );
  XOR U12751 ( .A(n12621), .B(n12607), .Z(n12613) );
  XNOR U12752 ( .A(n12661), .B(n12569), .Z(n12607) );
  IV U12753 ( .A(n12611), .Z(n12661) );
  XOR U12754 ( .A(n12672), .B(n12673), .Z(n12611) );
  XOR U12755 ( .A(n12674), .B(n12675), .Z(n12673) );
  XNOR U12756 ( .A(n12441), .B(n12676), .Z(n12672) );
  ANDN U12757 ( .B(n12562), .A(n12621), .Z(n12667) );
  XNOR U12758 ( .A(n12441), .B(n12677), .Z(n12621) );
  XOR U12759 ( .A(n12550), .B(n12668), .Z(n12562) );
  XOR U12760 ( .A(n12678), .B(n12679), .Z(n12550) );
  XOR U12761 ( .A(n12680), .B(n12675), .Z(n12679) );
  XOR U12762 ( .A(state[20]), .B(key[20]), .Z(n12675) );
  XNOR U12763 ( .A(n12677), .B(n12541), .Z(n12650) );
  XNOR U12764 ( .A(n12681), .B(n12654), .Z(n12662) );
  OR U12765 ( .A(n12540), .B(n12602), .Z(n12654) );
  XNOR U12766 ( .A(n12603), .B(n12569), .Z(n12602) );
  XOR U12767 ( .A(n12682), .B(n12678), .Z(n12569) );
  XNOR U12768 ( .A(n12668), .B(n12445), .Z(n12540) );
  XOR U12769 ( .A(n12678), .B(n12683), .Z(n12445) );
  XOR U12770 ( .A(n12670), .B(n12682), .Z(n12683) );
  IV U12771 ( .A(n12541), .Z(n12668) );
  ANDN U12772 ( .B(n12677), .A(n12541), .Z(n12681) );
  XNOR U12773 ( .A(n12678), .B(n12684), .Z(n12541) );
  XNOR U12774 ( .A(n12680), .B(n12674), .Z(n12684) );
  XNOR U12775 ( .A(state[23]), .B(key[23]), .Z(n12674) );
  XNOR U12776 ( .A(state[21]), .B(key[21]), .Z(n12678) );
  IV U12777 ( .A(n12603), .Z(n12677) );
  XNOR U12778 ( .A(n12671), .B(n12685), .Z(n12603) );
  XOR U12779 ( .A(n12676), .B(n12682), .Z(n12685) );
  IV U12780 ( .A(n12680), .Z(n12682) );
  XOR U12781 ( .A(n12441), .B(n12686), .Z(n12680) );
  XNOR U12782 ( .A(state[22]), .B(key[22]), .Z(n12686) );
  XOR U12783 ( .A(state[16]), .B(key[16]), .Z(n12441) );
  XNOR U12784 ( .A(n12670), .B(n12687), .Z(n12676) );
  XNOR U12785 ( .A(state[19]), .B(key[19]), .Z(n12687) );
  XNOR U12786 ( .A(state[17]), .B(key[17]), .Z(n12670) );
  XNOR U12787 ( .A(state[18]), .B(key[18]), .Z(n12671) );
  XOR U12788 ( .A(n12373), .B(n12497), .Z(n10214) );
  XNOR U12789 ( .A(n12572), .B(n12688), .Z(n12497) );
  XOR U12790 ( .A(n12689), .B(n12414), .Z(n12688) );
  OR U12791 ( .A(n12690), .B(n12527), .Z(n12414) );
  XOR U12792 ( .A(n12416), .B(n12691), .Z(n12527) );
  ANDN U12793 ( .B(n12692), .A(n12525), .Z(n12689) );
  XNOR U12794 ( .A(n12412), .B(n12693), .Z(n12373) );
  XOR U12795 ( .A(n12694), .B(n12574), .Z(n12693) );
  OR U12796 ( .A(n12695), .B(n12514), .Z(n12574) );
  XOR U12797 ( .A(n12517), .B(n12421), .Z(n12514) );
  NOR U12798 ( .A(n12696), .B(n12517), .Z(n12694) );
  XNOR U12799 ( .A(n12572), .B(n12697), .Z(n12412) );
  XNOR U12800 ( .A(n12698), .B(n12699), .Z(n12697) );
  NANDN U12801 ( .A(n12521), .B(n12700), .Z(n12699) );
  XOR U12802 ( .A(n12701), .B(n12698), .Z(n12572) );
  OR U12803 ( .A(n12530), .B(n12702), .Z(n12698) );
  XOR U12804 ( .A(n12532), .B(n12521), .Z(n12530) );
  XNOR U12805 ( .A(n12691), .B(n12421), .Z(n12521) );
  XOR U12806 ( .A(n12703), .B(n12704), .Z(n12421) );
  NANDN U12807 ( .A(n12705), .B(n12706), .Z(n12704) );
  IV U12808 ( .A(n12525), .Z(n12691) );
  XNOR U12809 ( .A(n12707), .B(n12708), .Z(n12525) );
  NANDN U12810 ( .A(n12705), .B(n12709), .Z(n12708) );
  ANDN U12811 ( .B(n12532), .A(n12710), .Z(n12701) );
  XOR U12812 ( .A(n12517), .B(n12416), .Z(n12532) );
  XOR U12813 ( .A(n12711), .B(n12707), .Z(n12416) );
  NANDN U12814 ( .A(n12712), .B(n12713), .Z(n12707) );
  NANDN U12815 ( .A(n12712), .B(n12717), .Z(n12703) );
  XOR U12816 ( .A(n12718), .B(n12719), .Z(n12705) );
  XOR U12817 ( .A(n12720), .B(n12715), .Z(n12719) );
  XNOR U12818 ( .A(n12721), .B(n12722), .Z(n12718) );
  XNOR U12819 ( .A(n12723), .B(n12724), .Z(n12722) );
  ANDN U12820 ( .B(n12720), .A(n12715), .Z(n12723) );
  ANDN U12821 ( .B(n12720), .A(n12714), .Z(n12716) );
  XNOR U12822 ( .A(n12721), .B(n12725), .Z(n12714) );
  XOR U12823 ( .A(n12726), .B(n12724), .Z(n12725) );
  NAND U12824 ( .A(n12713), .B(n12717), .Z(n12724) );
  XNOR U12825 ( .A(n12709), .B(n12715), .Z(n12713) );
  XOR U12826 ( .A(n12727), .B(n12728), .Z(n12715) );
  XOR U12827 ( .A(n12729), .B(n12730), .Z(n12728) );
  XNOR U12828 ( .A(n12731), .B(n12732), .Z(n12727) );
  ANDN U12829 ( .B(n12733), .A(n12516), .Z(n12731) );
  AND U12830 ( .A(n12706), .B(n12709), .Z(n12726) );
  XNOR U12831 ( .A(n12706), .B(n12709), .Z(n12721) );
  XNOR U12832 ( .A(n12734), .B(n12735), .Z(n12709) );
  XNOR U12833 ( .A(n12736), .B(n12737), .Z(n12735) );
  XOR U12834 ( .A(n12729), .B(n12738), .Z(n12734) );
  XNOR U12835 ( .A(n12739), .B(n12732), .Z(n12738) );
  OR U12836 ( .A(n12515), .B(n12695), .Z(n12732) );
  XNOR U12837 ( .A(n12696), .B(n12576), .Z(n12695) );
  XNOR U12838 ( .A(n12516), .B(n12422), .Z(n12515) );
  NOR U12839 ( .A(n12422), .B(n12576), .Z(n12739) );
  XNOR U12840 ( .A(n12740), .B(n12741), .Z(n12706) );
  XNOR U12841 ( .A(n12742), .B(n12743), .Z(n12741) );
  XOR U12842 ( .A(n12511), .B(n12729), .Z(n12743) );
  XOR U12843 ( .A(n12733), .B(n12744), .Z(n12729) );
  XNOR U12844 ( .A(n12417), .B(n12745), .Z(n12740) );
  XNOR U12845 ( .A(n12746), .B(n12747), .Z(n12745) );
  ANDN U12846 ( .B(n12526), .A(n12748), .Z(n12746) );
  XNOR U12847 ( .A(n12749), .B(n12750), .Z(n12720) );
  XNOR U12848 ( .A(n12730), .B(n12751), .Z(n12750) );
  XNOR U12849 ( .A(n12526), .B(n12737), .Z(n12751) );
  XOR U12850 ( .A(n12576), .B(n12422), .Z(n12737) );
  XNOR U12851 ( .A(n12742), .B(n12752), .Z(n12730) );
  XNOR U12852 ( .A(n12753), .B(n12754), .Z(n12752) );
  NANDN U12853 ( .A(n12522), .B(n12700), .Z(n12754) );
  IV U12854 ( .A(n12736), .Z(n12742) );
  XNOR U12855 ( .A(n12755), .B(n12753), .Z(n12736) );
  NANDN U12856 ( .A(n12702), .B(n12531), .Z(n12753) );
  XOR U12857 ( .A(n12526), .B(n12422), .Z(n12522) );
  XOR U12858 ( .A(n12756), .B(n12757), .Z(n12422) );
  XNOR U12859 ( .A(n12758), .B(n12759), .Z(n12757) );
  XOR U12860 ( .A(n12710), .B(n12700), .Z(n12702) );
  XNOR U12861 ( .A(n12692), .B(n12576), .Z(n12700) );
  XNOR U12862 ( .A(n12759), .B(n12760), .Z(n12576) );
  ANDN U12863 ( .B(n12533), .A(n12710), .Z(n12755) );
  XNOR U12864 ( .A(n12761), .B(n12733), .Z(n12710) );
  IV U12865 ( .A(n12696), .Z(n12733) );
  XNOR U12866 ( .A(n12762), .B(n12763), .Z(n12696) );
  XNOR U12867 ( .A(n12764), .B(n12759), .Z(n12763) );
  XOR U12868 ( .A(n12765), .B(n12744), .Z(n12533) );
  XNOR U12869 ( .A(n12748), .B(n12766), .Z(n12749) );
  XNOR U12870 ( .A(n12767), .B(n12747), .Z(n12766) );
  OR U12871 ( .A(n12528), .B(n12690), .Z(n12747) );
  XOR U12872 ( .A(n12417), .B(n12692), .Z(n12690) );
  IV U12873 ( .A(n12748), .Z(n12692) );
  XOR U12874 ( .A(n12511), .B(n12526), .Z(n12528) );
  XNOR U12875 ( .A(n12744), .B(n12768), .Z(n12526) );
  XNOR U12876 ( .A(n12758), .B(n12762), .Z(n12768) );
  XNOR U12877 ( .A(state[58]), .B(key[58]), .Z(n12762) );
  IV U12878 ( .A(n12516), .Z(n12744) );
  XOR U12879 ( .A(n12756), .B(n12769), .Z(n12516) );
  XOR U12880 ( .A(n12759), .B(n12770), .Z(n12769) );
  IV U12881 ( .A(n12765), .Z(n12511) );
  ANDN U12882 ( .B(n12765), .A(n12417), .Z(n12767) );
  XOR U12883 ( .A(n12760), .B(n12771), .Z(n12765) );
  XNOR U12884 ( .A(n12759), .B(n12772), .Z(n12771) );
  XOR U12885 ( .A(n12761), .B(n12773), .Z(n12759) );
  XNOR U12886 ( .A(state[62]), .B(key[62]), .Z(n12773) );
  IV U12887 ( .A(n12756), .Z(n12760) );
  XOR U12888 ( .A(state[61]), .B(key[61]), .Z(n12756) );
  XOR U12889 ( .A(n12774), .B(n12775), .Z(n12748) );
  XOR U12890 ( .A(n12772), .B(n12770), .Z(n12775) );
  XOR U12891 ( .A(state[63]), .B(key[63]), .Z(n12770) );
  XNOR U12892 ( .A(state[60]), .B(key[60]), .Z(n12772) );
  XOR U12893 ( .A(n12417), .B(n12764), .Z(n12774) );
  XNOR U12894 ( .A(n12758), .B(n12776), .Z(n12764) );
  XNOR U12895 ( .A(state[59]), .B(key[59]), .Z(n12776) );
  XNOR U12896 ( .A(state[57]), .B(key[57]), .Z(n12758) );
  IV U12897 ( .A(n12761), .Z(n12417) );
  XOR U12898 ( .A(state[56]), .B(key[56]), .Z(n12761) );
  XOR U12899 ( .A(n12455), .B(n12777), .Z(n12498) );
  XOR U12900 ( .A(n12577), .B(n12588), .Z(n12463) );
  XOR U12901 ( .A(n12425), .B(n12778), .Z(n12588) );
  XNOR U12902 ( .A(n12779), .B(n12780), .Z(n12778) );
  NANDN U12903 ( .A(n12781), .B(n12782), .Z(n12780) );
  IV U12904 ( .A(n12783), .Z(n12577) );
  XNOR U12905 ( .A(n12779), .B(n12785), .Z(n12784) );
  OR U12906 ( .A(n12460), .B(n12786), .Z(n12785) );
  OR U12907 ( .A(n12787), .B(n12788), .Z(n12779) );
  XNOR U12908 ( .A(n12425), .B(n12789), .Z(n12581) );
  XNOR U12909 ( .A(n12790), .B(n12791), .Z(n12789) );
  OR U12910 ( .A(n12792), .B(n12793), .Z(n12791) );
  XOR U12911 ( .A(n12794), .B(n12790), .Z(n12425) );
  NANDN U12912 ( .A(n12795), .B(n12796), .Z(n12790) );
  XOR U12913 ( .A(n12799), .B(n12800), .Z(n12455) );
  XNOR U12914 ( .A(n12801), .B(n12802), .Z(n12800) );
  NANDN U12915 ( .A(n12803), .B(n12431), .Z(n12802) );
  XNOR U12916 ( .A(n10974), .B(n12804), .Z(n12598) );
  XNOR U12917 ( .A(key[168]), .B(n12371), .Z(n12804) );
  IV U12918 ( .A(n9276), .Z(n12371) );
  XOR U12919 ( .A(n12427), .B(n12783), .Z(n9276) );
  XNOR U12920 ( .A(n12799), .B(n12805), .Z(n12783) );
  XOR U12921 ( .A(n12806), .B(n12458), .Z(n12805) );
  OR U12922 ( .A(n12787), .B(n12807), .Z(n12458) );
  XOR U12923 ( .A(n12460), .B(n12808), .Z(n12787) );
  ANDN U12924 ( .B(n12809), .A(n12781), .Z(n12806) );
  XNOR U12925 ( .A(n12456), .B(n12810), .Z(n12427) );
  XOR U12926 ( .A(n12811), .B(n12801), .Z(n12810) );
  OR U12927 ( .A(n12812), .B(n12584), .Z(n12801) );
  XOR U12928 ( .A(n12587), .B(n12431), .Z(n12584) );
  NOR U12929 ( .A(n12813), .B(n12587), .Z(n12811) );
  XNOR U12930 ( .A(n12799), .B(n12814), .Z(n12456) );
  XNOR U12931 ( .A(n12815), .B(n12816), .Z(n12814) );
  NANDN U12932 ( .A(n12792), .B(n12817), .Z(n12816) );
  XOR U12933 ( .A(n12818), .B(n12815), .Z(n12799) );
  OR U12934 ( .A(n12795), .B(n12819), .Z(n12815) );
  XOR U12935 ( .A(n12798), .B(n12792), .Z(n12795) );
  XNOR U12936 ( .A(n12808), .B(n12431), .Z(n12792) );
  XOR U12937 ( .A(n12820), .B(n12821), .Z(n12431) );
  NANDN U12938 ( .A(n12822), .B(n12823), .Z(n12821) );
  IV U12939 ( .A(n12781), .Z(n12808) );
  XNOR U12940 ( .A(n12824), .B(n12825), .Z(n12781) );
  NANDN U12941 ( .A(n12822), .B(n12826), .Z(n12825) );
  ANDN U12942 ( .B(n12798), .A(n12827), .Z(n12818) );
  XOR U12943 ( .A(n12587), .B(n12460), .Z(n12798) );
  XOR U12944 ( .A(n12828), .B(n12824), .Z(n12460) );
  NANDN U12945 ( .A(n12829), .B(n12830), .Z(n12824) );
  NANDN U12946 ( .A(n12829), .B(n12834), .Z(n12820) );
  XOR U12947 ( .A(n12835), .B(n12836), .Z(n12822) );
  XOR U12948 ( .A(n12837), .B(n12832), .Z(n12836) );
  XNOR U12949 ( .A(n12838), .B(n12839), .Z(n12835) );
  XNOR U12950 ( .A(n12840), .B(n12841), .Z(n12839) );
  ANDN U12951 ( .B(n12837), .A(n12832), .Z(n12840) );
  ANDN U12952 ( .B(n12837), .A(n12831), .Z(n12833) );
  XNOR U12953 ( .A(n12838), .B(n12842), .Z(n12831) );
  XOR U12954 ( .A(n12843), .B(n12841), .Z(n12842) );
  NAND U12955 ( .A(n12830), .B(n12834), .Z(n12841) );
  XNOR U12956 ( .A(n12826), .B(n12832), .Z(n12830) );
  XOR U12957 ( .A(n12844), .B(n12845), .Z(n12832) );
  XOR U12958 ( .A(n12846), .B(n12847), .Z(n12845) );
  XNOR U12959 ( .A(n12848), .B(n12849), .Z(n12844) );
  ANDN U12960 ( .B(n12850), .A(n12586), .Z(n12848) );
  AND U12961 ( .A(n12823), .B(n12826), .Z(n12843) );
  XNOR U12962 ( .A(n12823), .B(n12826), .Z(n12838) );
  XNOR U12963 ( .A(n12851), .B(n12852), .Z(n12826) );
  XNOR U12964 ( .A(n12853), .B(n12854), .Z(n12852) );
  XOR U12965 ( .A(n12846), .B(n12855), .Z(n12851) );
  XNOR U12966 ( .A(n12856), .B(n12849), .Z(n12855) );
  OR U12967 ( .A(n12585), .B(n12812), .Z(n12849) );
  XNOR U12968 ( .A(n12813), .B(n12803), .Z(n12812) );
  XNOR U12969 ( .A(n12586), .B(n12432), .Z(n12585) );
  NOR U12970 ( .A(n12432), .B(n12803), .Z(n12856) );
  XNOR U12971 ( .A(n12857), .B(n12858), .Z(n12823) );
  XNOR U12972 ( .A(n12859), .B(n12860), .Z(n12858) );
  XOR U12973 ( .A(n12786), .B(n12846), .Z(n12860) );
  XOR U12974 ( .A(n12850), .B(n12861), .Z(n12846) );
  XNOR U12975 ( .A(n12461), .B(n12862), .Z(n12857) );
  XNOR U12976 ( .A(n12863), .B(n12864), .Z(n12862) );
  ANDN U12977 ( .B(n12782), .A(n12865), .Z(n12863) );
  XNOR U12978 ( .A(n12866), .B(n12867), .Z(n12837) );
  XNOR U12979 ( .A(n12847), .B(n12868), .Z(n12867) );
  XNOR U12980 ( .A(n12782), .B(n12854), .Z(n12868) );
  XOR U12981 ( .A(n12803), .B(n12432), .Z(n12854) );
  XNOR U12982 ( .A(n12859), .B(n12869), .Z(n12847) );
  XNOR U12983 ( .A(n12870), .B(n12871), .Z(n12869) );
  NANDN U12984 ( .A(n12793), .B(n12817), .Z(n12871) );
  IV U12985 ( .A(n12853), .Z(n12859) );
  XNOR U12986 ( .A(n12872), .B(n12870), .Z(n12853) );
  NANDN U12987 ( .A(n12819), .B(n12796), .Z(n12870) );
  XOR U12988 ( .A(n12782), .B(n12432), .Z(n12793) );
  XOR U12989 ( .A(n12873), .B(n12874), .Z(n12432) );
  XNOR U12990 ( .A(n12875), .B(n12876), .Z(n12874) );
  XOR U12991 ( .A(n12827), .B(n12817), .Z(n12819) );
  XNOR U12992 ( .A(n12809), .B(n12803), .Z(n12817) );
  XNOR U12993 ( .A(n12876), .B(n12877), .Z(n12803) );
  ANDN U12994 ( .B(n12797), .A(n12827), .Z(n12872) );
  XNOR U12995 ( .A(n12878), .B(n12850), .Z(n12827) );
  IV U12996 ( .A(n12813), .Z(n12850) );
  XNOR U12997 ( .A(n12879), .B(n12880), .Z(n12813) );
  XNOR U12998 ( .A(n12881), .B(n12876), .Z(n12880) );
  XOR U12999 ( .A(n12882), .B(n12861), .Z(n12797) );
  XNOR U13000 ( .A(n12865), .B(n12883), .Z(n12866) );
  XNOR U13001 ( .A(n12884), .B(n12864), .Z(n12883) );
  OR U13002 ( .A(n12788), .B(n12807), .Z(n12864) );
  XOR U13003 ( .A(n12461), .B(n12809), .Z(n12807) );
  IV U13004 ( .A(n12865), .Z(n12809) );
  XOR U13005 ( .A(n12786), .B(n12782), .Z(n12788) );
  XNOR U13006 ( .A(n12861), .B(n12885), .Z(n12782) );
  XNOR U13007 ( .A(n12875), .B(n12879), .Z(n12885) );
  XNOR U13008 ( .A(state[66]), .B(key[66]), .Z(n12879) );
  IV U13009 ( .A(n12586), .Z(n12861) );
  XOR U13010 ( .A(n12873), .B(n12886), .Z(n12586) );
  XOR U13011 ( .A(n12876), .B(n12887), .Z(n12886) );
  IV U13012 ( .A(n12882), .Z(n12786) );
  ANDN U13013 ( .B(n12882), .A(n12461), .Z(n12884) );
  XOR U13014 ( .A(n12877), .B(n12888), .Z(n12882) );
  XNOR U13015 ( .A(n12876), .B(n12889), .Z(n12888) );
  XOR U13016 ( .A(n12878), .B(n12890), .Z(n12876) );
  XNOR U13017 ( .A(state[70]), .B(key[70]), .Z(n12890) );
  IV U13018 ( .A(n12873), .Z(n12877) );
  XOR U13019 ( .A(state[69]), .B(key[69]), .Z(n12873) );
  XOR U13020 ( .A(n12891), .B(n12892), .Z(n12865) );
  XOR U13021 ( .A(n12889), .B(n12887), .Z(n12892) );
  XOR U13022 ( .A(state[71]), .B(key[71]), .Z(n12887) );
  XNOR U13023 ( .A(state[68]), .B(key[68]), .Z(n12889) );
  XOR U13024 ( .A(n12461), .B(n12881), .Z(n12891) );
  XNOR U13025 ( .A(n12875), .B(n12893), .Z(n12881) );
  XNOR U13026 ( .A(state[67]), .B(key[67]), .Z(n12893) );
  XNOR U13027 ( .A(state[65]), .B(key[65]), .Z(n12875) );
  IV U13028 ( .A(n12878), .Z(n12461) );
  XOR U13029 ( .A(state[64]), .B(key[64]), .Z(n12878) );
  XNOR U13030 ( .A(n12448), .B(n12894), .Z(n10974) );
  XOR U13031 ( .A(n12499), .B(n12473), .Z(n12894) );
  XNOR U13032 ( .A(n12896), .B(n12897), .Z(n12895) );
  NANDN U13033 ( .A(n12470), .B(n12898), .Z(n12897) );
  XNOR U13034 ( .A(n12380), .B(n12899), .Z(n12592) );
  XNOR U13035 ( .A(n12900), .B(n12901), .Z(n12899) );
  NANDN U13036 ( .A(n12491), .B(n12902), .Z(n12901) );
  XNOR U13037 ( .A(n12487), .B(n12903), .Z(n12499) );
  XNOR U13038 ( .A(n12484), .B(n12904), .Z(n12903) );
  NANDN U13039 ( .A(n12905), .B(n12906), .Z(n12904) );
  OR U13040 ( .A(n12907), .B(n12595), .Z(n12484) );
  XOR U13041 ( .A(n12486), .B(n12906), .Z(n12595) );
  XOR U13042 ( .A(n12481), .B(n12591), .Z(n12448) );
  XOR U13043 ( .A(n12380), .B(n12908), .Z(n12591) );
  XNOR U13044 ( .A(n12896), .B(n12909), .Z(n12908) );
  NANDN U13045 ( .A(n12910), .B(n12911), .Z(n12909) );
  OR U13046 ( .A(n12912), .B(n12913), .Z(n12896) );
  XOR U13047 ( .A(n12914), .B(n12900), .Z(n12380) );
  NANDN U13048 ( .A(n12915), .B(n12916), .Z(n12900) );
  AND U13049 ( .A(n12917), .B(n12918), .Z(n12914) );
  XNOR U13050 ( .A(n12487), .B(n12919), .Z(n12481) );
  XOR U13051 ( .A(n12920), .B(n12468), .Z(n12919) );
  OR U13052 ( .A(n12912), .B(n12921), .Z(n12468) );
  XOR U13053 ( .A(n12470), .B(n12911), .Z(n12912) );
  ANDN U13054 ( .B(n12911), .A(n12922), .Z(n12920) );
  XOR U13055 ( .A(n12923), .B(n12489), .Z(n12487) );
  OR U13056 ( .A(n12915), .B(n12924), .Z(n12489) );
  XOR U13057 ( .A(n12917), .B(n12491), .Z(n12915) );
  XNOR U13058 ( .A(n12911), .B(n12906), .Z(n12491) );
  IV U13059 ( .A(n12385), .Z(n12906) );
  XNOR U13060 ( .A(n12925), .B(n12926), .Z(n12385) );
  NANDN U13061 ( .A(n12927), .B(n12928), .Z(n12926) );
  XOR U13062 ( .A(n12929), .B(n12930), .Z(n12911) );
  NANDN U13063 ( .A(n12927), .B(n12931), .Z(n12930) );
  ANDN U13064 ( .B(n12917), .A(n12932), .Z(n12923) );
  XOR U13065 ( .A(n12470), .B(n12486), .Z(n12917) );
  XOR U13066 ( .A(n12933), .B(n12925), .Z(n12486) );
  NANDN U13067 ( .A(n12934), .B(n12935), .Z(n12925) );
  XOR U13068 ( .A(n12928), .B(n12936), .Z(n12935) );
  ANDN U13069 ( .B(n12936), .A(n12937), .Z(n12933) );
  NANDN U13070 ( .A(n12934), .B(n12939), .Z(n12929) );
  XOR U13071 ( .A(n12940), .B(n12941), .Z(n12927) );
  XOR U13072 ( .A(n12942), .B(n12943), .Z(n12941) );
  XNOR U13073 ( .A(n12944), .B(n12945), .Z(n12940) );
  XNOR U13074 ( .A(n12946), .B(n12947), .Z(n12945) );
  ANDN U13075 ( .B(n12943), .A(n12942), .Z(n12946) );
  ANDN U13076 ( .B(n12943), .A(n12937), .Z(n12938) );
  XNOR U13077 ( .A(n12944), .B(n12948), .Z(n12937) );
  XOR U13078 ( .A(n12949), .B(n12947), .Z(n12948) );
  NAND U13079 ( .A(n12939), .B(n12950), .Z(n12947) );
  XNOR U13080 ( .A(n12928), .B(n12942), .Z(n12950) );
  IV U13081 ( .A(n12936), .Z(n12942) );
  XNOR U13082 ( .A(n12951), .B(n12952), .Z(n12936) );
  XNOR U13083 ( .A(n12953), .B(n12954), .Z(n12952) );
  XOR U13084 ( .A(n12910), .B(n12955), .Z(n12954) );
  XNOR U13085 ( .A(n12922), .B(n12956), .Z(n12951) );
  XNOR U13086 ( .A(n12957), .B(n12958), .Z(n12956) );
  AND U13087 ( .A(n12898), .B(n12471), .Z(n12957) );
  XOR U13088 ( .A(n12931), .B(n12943), .Z(n12939) );
  AND U13089 ( .A(n12928), .B(n12931), .Z(n12949) );
  XNOR U13090 ( .A(n12928), .B(n12931), .Z(n12944) );
  XNOR U13091 ( .A(n12959), .B(n12960), .Z(n12931) );
  XNOR U13092 ( .A(n12961), .B(n12955), .Z(n12960) );
  XOR U13093 ( .A(n12962), .B(n12963), .Z(n12959) );
  XNOR U13094 ( .A(n12964), .B(n12965), .Z(n12963) );
  ANDN U13095 ( .B(n12384), .A(n12905), .Z(n12964) );
  XNOR U13096 ( .A(n12966), .B(n12967), .Z(n12928) );
  XNOR U13097 ( .A(n12898), .B(n12962), .Z(n12968) );
  XOR U13098 ( .A(n12471), .B(n12969), .Z(n12966) );
  XNOR U13099 ( .A(n12970), .B(n12958), .Z(n12969) );
  OR U13100 ( .A(n12913), .B(n12921), .Z(n12958) );
  XOR U13101 ( .A(n12471), .B(n12922), .Z(n12921) );
  XNOR U13102 ( .A(n12898), .B(n12971), .Z(n12913) );
  ANDN U13103 ( .B(n12972), .A(n12910), .Z(n12970) );
  XNOR U13104 ( .A(n12973), .B(n12974), .Z(n12943) );
  XOR U13105 ( .A(n12961), .B(n12953), .Z(n12974) );
  XOR U13106 ( .A(n12962), .B(n12975), .Z(n12953) );
  XNOR U13107 ( .A(n12976), .B(n12977), .Z(n12975) );
  NAND U13108 ( .A(n12492), .B(n12902), .Z(n12977) );
  XNOR U13109 ( .A(n12978), .B(n12976), .Z(n12962) );
  NANDN U13110 ( .A(n12924), .B(n12916), .Z(n12976) );
  XOR U13111 ( .A(n12918), .B(n12902), .Z(n12916) );
  XOR U13112 ( .A(n12971), .B(n12384), .Z(n12902) );
  IV U13113 ( .A(n12910), .Z(n12971) );
  XOR U13114 ( .A(n12979), .B(n12980), .Z(n12910) );
  XNOR U13115 ( .A(n12981), .B(n12982), .Z(n12980) );
  XOR U13116 ( .A(n12932), .B(n12492), .Z(n12924) );
  XNOR U13117 ( .A(n12972), .B(n12905), .Z(n12492) );
  IV U13118 ( .A(n12922), .Z(n12972) );
  XOR U13119 ( .A(n12983), .B(n12984), .Z(n12922) );
  XOR U13120 ( .A(n12985), .B(n12986), .Z(n12984) );
  XNOR U13121 ( .A(n12471), .B(n12987), .Z(n12983) );
  ANDN U13122 ( .B(n12918), .A(n12932), .Z(n12978) );
  XNOR U13123 ( .A(n12471), .B(n12988), .Z(n12932) );
  XOR U13124 ( .A(n12898), .B(n12979), .Z(n12918) );
  XOR U13125 ( .A(n12989), .B(n12990), .Z(n12898) );
  XOR U13126 ( .A(n12991), .B(n12986), .Z(n12990) );
  XOR U13127 ( .A(state[108]), .B(key[108]), .Z(n12986) );
  XNOR U13128 ( .A(n12988), .B(n12597), .Z(n12961) );
  XNOR U13129 ( .A(n12992), .B(n12965), .Z(n12973) );
  OR U13130 ( .A(n12596), .B(n12907), .Z(n12965) );
  XNOR U13131 ( .A(n12485), .B(n12905), .Z(n12907) );
  XOR U13132 ( .A(n12993), .B(n12989), .Z(n12905) );
  XNOR U13133 ( .A(n12979), .B(n12384), .Z(n12596) );
  XOR U13134 ( .A(n12989), .B(n12994), .Z(n12384) );
  XOR U13135 ( .A(n12981), .B(n12993), .Z(n12994) );
  IV U13136 ( .A(n12597), .Z(n12979) );
  ANDN U13137 ( .B(n12988), .A(n12597), .Z(n12992) );
  XNOR U13138 ( .A(n12989), .B(n12995), .Z(n12597) );
  XNOR U13139 ( .A(n12991), .B(n12985), .Z(n12995) );
  XNOR U13140 ( .A(state[111]), .B(key[111]), .Z(n12985) );
  XNOR U13141 ( .A(state[109]), .B(key[109]), .Z(n12989) );
  IV U13142 ( .A(n12485), .Z(n12988) );
  XNOR U13143 ( .A(n12982), .B(n12996), .Z(n12485) );
  XOR U13144 ( .A(n12987), .B(n12993), .Z(n12996) );
  IV U13145 ( .A(n12991), .Z(n12993) );
  XOR U13146 ( .A(n12471), .B(n12997), .Z(n12991) );
  XNOR U13147 ( .A(state[110]), .B(key[110]), .Z(n12997) );
  XOR U13148 ( .A(state[104]), .B(key[104]), .Z(n12471) );
  XNOR U13149 ( .A(n12981), .B(n12998), .Z(n12987) );
  XNOR U13150 ( .A(state[107]), .B(key[107]), .Z(n12998) );
  XNOR U13151 ( .A(state[105]), .B(key[105]), .Z(n12981) );
  XNOR U13152 ( .A(state[106]), .B(key[106]), .Z(n12982) );
  XOR U13153 ( .A(n7760), .B(n12999), .Z(n11501) );
  XNOR U13154 ( .A(key[358]), .B(n6082), .Z(n12999) );
  XOR U13155 ( .A(n11512), .B(n11414), .Z(n6082) );
  XNOR U13156 ( .A(n12282), .B(n13000), .Z(n11414) );
  XNOR U13157 ( .A(n13001), .B(n11489), .Z(n13000) );
  ANDN U13158 ( .B(n12287), .A(n13002), .Z(n11489) );
  XOR U13159 ( .A(n13003), .B(n11491), .Z(n12287) );
  ANDN U13160 ( .B(n13004), .A(n12270), .Z(n13001) );
  IV U13161 ( .A(n13003), .Z(n12270) );
  XNOR U13162 ( .A(n11486), .B(n13005), .Z(n12282) );
  XNOR U13163 ( .A(n13006), .B(n13007), .Z(n13005) );
  NANDN U13164 ( .A(n12275), .B(n13008), .Z(n13007) );
  XNOR U13165 ( .A(n11409), .B(n11416), .Z(n11512) );
  XOR U13166 ( .A(n11486), .B(n13009), .Z(n11416) );
  XNOR U13167 ( .A(n12279), .B(n13010), .Z(n13009) );
  NANDN U13168 ( .A(n13011), .B(n13012), .Z(n13010) );
  OR U13169 ( .A(n13013), .B(n13014), .Z(n12279) );
  XOR U13170 ( .A(n13015), .B(n13006), .Z(n11486) );
  NANDN U13171 ( .A(n13016), .B(n13017), .Z(n13006) );
  ANDN U13172 ( .B(n13018), .A(n13019), .Z(n13015) );
  XNOR U13173 ( .A(n12271), .B(n13020), .Z(n11409) );
  XOR U13174 ( .A(n13021), .B(n11507), .Z(n13020) );
  OR U13175 ( .A(n13022), .B(n13013), .Z(n11507) );
  XNOR U13176 ( .A(n11510), .B(n13012), .Z(n13013) );
  ANDN U13177 ( .B(n13012), .A(n13023), .Z(n13021) );
  XOR U13178 ( .A(n13024), .B(n12273), .Z(n12271) );
  OR U13179 ( .A(n13016), .B(n13025), .Z(n12273) );
  XNOR U13180 ( .A(n13019), .B(n12275), .Z(n13016) );
  XNOR U13181 ( .A(n13012), .B(n11491), .Z(n12275) );
  XOR U13182 ( .A(n13026), .B(n13027), .Z(n11491) );
  NANDN U13183 ( .A(n13028), .B(n13029), .Z(n13027) );
  XOR U13184 ( .A(n13030), .B(n13031), .Z(n13012) );
  NANDN U13185 ( .A(n13028), .B(n13032), .Z(n13031) );
  NOR U13186 ( .A(n13019), .B(n13033), .Z(n13024) );
  XNOR U13187 ( .A(n13003), .B(n11510), .Z(n13019) );
  XNOR U13188 ( .A(n13034), .B(n13030), .Z(n11510) );
  NANDN U13189 ( .A(n13035), .B(n13036), .Z(n13030) );
  XOR U13190 ( .A(n13032), .B(n13037), .Z(n13036) );
  ANDN U13191 ( .B(n13037), .A(n13038), .Z(n13034) );
  XNOR U13192 ( .A(n13039), .B(n13026), .Z(n13003) );
  NANDN U13193 ( .A(n13035), .B(n13040), .Z(n13026) );
  XOR U13194 ( .A(n13041), .B(n13029), .Z(n13040) );
  XNOR U13195 ( .A(n13042), .B(n13043), .Z(n13028) );
  XOR U13196 ( .A(n13044), .B(n13045), .Z(n13043) );
  XNOR U13197 ( .A(n13046), .B(n13047), .Z(n13042) );
  XNOR U13198 ( .A(n13048), .B(n13049), .Z(n13047) );
  ANDN U13199 ( .B(n13041), .A(n13045), .Z(n13048) );
  ANDN U13200 ( .B(n13041), .A(n13038), .Z(n13039) );
  XNOR U13201 ( .A(n13044), .B(n13050), .Z(n13038) );
  XOR U13202 ( .A(n13051), .B(n13049), .Z(n13050) );
  NAND U13203 ( .A(n13052), .B(n13053), .Z(n13049) );
  XNOR U13204 ( .A(n13046), .B(n13029), .Z(n13053) );
  IV U13205 ( .A(n13041), .Z(n13046) );
  XNOR U13206 ( .A(n13032), .B(n13045), .Z(n13052) );
  IV U13207 ( .A(n13037), .Z(n13045) );
  XOR U13208 ( .A(n13054), .B(n13055), .Z(n13037) );
  XNOR U13209 ( .A(n13056), .B(n13057), .Z(n13055) );
  XNOR U13210 ( .A(n13058), .B(n13059), .Z(n13054) );
  ANDN U13211 ( .B(n12269), .A(n13060), .Z(n13058) );
  AND U13212 ( .A(n13029), .B(n13032), .Z(n13051) );
  XNOR U13213 ( .A(n13029), .B(n13032), .Z(n13044) );
  XNOR U13214 ( .A(n13061), .B(n13062), .Z(n13032) );
  XNOR U13215 ( .A(n13063), .B(n13057), .Z(n13062) );
  XOR U13216 ( .A(n13064), .B(n13065), .Z(n13061) );
  XNOR U13217 ( .A(n13066), .B(n13059), .Z(n13065) );
  OR U13218 ( .A(n13002), .B(n12286), .Z(n13059) );
  XNOR U13219 ( .A(n12269), .B(n13067), .Z(n12286) );
  XNOR U13220 ( .A(n13060), .B(n11492), .Z(n13002) );
  ANDN U13221 ( .B(n13068), .A(n12285), .Z(n13066) );
  XNOR U13222 ( .A(n13069), .B(n13070), .Z(n13029) );
  XNOR U13223 ( .A(n13057), .B(n13071), .Z(n13070) );
  XOR U13224 ( .A(n12281), .B(n13064), .Z(n13071) );
  XNOR U13225 ( .A(n12269), .B(n13060), .Z(n13057) );
  XOR U13226 ( .A(n11509), .B(n13072), .Z(n13069) );
  XNOR U13227 ( .A(n13073), .B(n13074), .Z(n13072) );
  ANDN U13228 ( .B(n13075), .A(n13023), .Z(n13073) );
  XNOR U13229 ( .A(n13076), .B(n13077), .Z(n13041) );
  XNOR U13230 ( .A(n13063), .B(n13078), .Z(n13077) );
  XNOR U13231 ( .A(n13011), .B(n13056), .Z(n13078) );
  XOR U13232 ( .A(n13064), .B(n13079), .Z(n13056) );
  XNOR U13233 ( .A(n13080), .B(n13081), .Z(n13079) );
  NAND U13234 ( .A(n12276), .B(n13008), .Z(n13081) );
  XNOR U13235 ( .A(n13082), .B(n13080), .Z(n13064) );
  NANDN U13236 ( .A(n13025), .B(n13017), .Z(n13080) );
  XOR U13237 ( .A(n13018), .B(n13008), .Z(n13017) );
  XNOR U13238 ( .A(n13075), .B(n11492), .Z(n13008) );
  XOR U13239 ( .A(n13033), .B(n12276), .Z(n13025) );
  XNOR U13240 ( .A(n13023), .B(n13067), .Z(n12276) );
  ANDN U13241 ( .B(n13018), .A(n13033), .Z(n13082) );
  XOR U13242 ( .A(n11509), .B(n12269), .Z(n13033) );
  XNOR U13243 ( .A(n13083), .B(n13084), .Z(n12269) );
  XNOR U13244 ( .A(n13085), .B(n13086), .Z(n13084) );
  XOR U13245 ( .A(n13067), .B(n13068), .Z(n13063) );
  IV U13246 ( .A(n11492), .Z(n13068) );
  XOR U13247 ( .A(n13087), .B(n13088), .Z(n11492) );
  XNOR U13248 ( .A(n13089), .B(n13086), .Z(n13088) );
  IV U13249 ( .A(n12285), .Z(n13067) );
  XOR U13250 ( .A(n13086), .B(n13090), .Z(n12285) );
  XNOR U13251 ( .A(n13091), .B(n13092), .Z(n13076) );
  XNOR U13252 ( .A(n13093), .B(n13074), .Z(n13092) );
  OR U13253 ( .A(n13014), .B(n13022), .Z(n13074) );
  XNOR U13254 ( .A(n11509), .B(n13023), .Z(n13022) );
  IV U13255 ( .A(n13091), .Z(n13023) );
  XOR U13256 ( .A(n12281), .B(n13075), .Z(n13014) );
  IV U13257 ( .A(n13011), .Z(n13075) );
  XOR U13258 ( .A(n13004), .B(n13094), .Z(n13011) );
  XNOR U13259 ( .A(n13089), .B(n13083), .Z(n13094) );
  XOR U13260 ( .A(n13095), .B(n13096), .Z(n13083) );
  XOR U13261 ( .A(n9913), .B(n11112), .Z(n13096) );
  IV U13262 ( .A(n9141), .Z(n11112) );
  XOR U13263 ( .A(n9901), .B(n9104), .Z(n9141) );
  XOR U13264 ( .A(n11102), .B(n13097), .Z(n13095) );
  XNOR U13265 ( .A(key[250]), .B(n9918), .Z(n13097) );
  XNOR U13266 ( .A(n13098), .B(n13099), .Z(n11102) );
  XNOR U13267 ( .A(n13100), .B(n13101), .Z(n13099) );
  XNOR U13268 ( .A(n13102), .B(n13103), .Z(n13098) );
  IV U13269 ( .A(n13060), .Z(n13004) );
  XOR U13270 ( .A(n13087), .B(n13104), .Z(n13060) );
  XOR U13271 ( .A(n13086), .B(n13105), .Z(n13104) );
  NOR U13272 ( .A(n12281), .B(n11509), .Z(n13093) );
  XOR U13273 ( .A(n13087), .B(n13106), .Z(n12281) );
  XOR U13274 ( .A(n13086), .B(n13107), .Z(n13106) );
  XOR U13275 ( .A(n13108), .B(n13109), .Z(n13086) );
  XOR U13276 ( .A(n11119), .B(n9114), .Z(n13109) );
  XNOR U13277 ( .A(n9128), .B(n9922), .Z(n9114) );
  XNOR U13278 ( .A(n11091), .B(n9121), .Z(n11119) );
  XOR U13279 ( .A(n9949), .B(n9116), .Z(n9121) );
  XNOR U13280 ( .A(n13110), .B(n13111), .Z(n9116) );
  XOR U13281 ( .A(n13112), .B(n9923), .Z(n11091) );
  XOR U13282 ( .A(n13113), .B(n13114), .Z(n9923) );
  XNOR U13283 ( .A(n13115), .B(n13116), .Z(n13114) );
  XNOR U13284 ( .A(n13117), .B(n13103), .Z(n13113) );
  XOR U13285 ( .A(n9956), .B(n13118), .Z(n13108) );
  XOR U13286 ( .A(key[254]), .B(n11509), .Z(n13118) );
  XOR U13287 ( .A(n13119), .B(n13120), .Z(n9956) );
  IV U13288 ( .A(n13090), .Z(n13087) );
  XOR U13289 ( .A(n13121), .B(n13122), .Z(n13090) );
  XNOR U13290 ( .A(n11097), .B(n11096), .Z(n13122) );
  XOR U13291 ( .A(n9952), .B(n9119), .Z(n11096) );
  XNOR U13292 ( .A(n13123), .B(n13124), .Z(n9119) );
  XNOR U13293 ( .A(n13125), .B(n13126), .Z(n13124) );
  XNOR U13294 ( .A(n13127), .B(n13128), .Z(n13123) );
  XNOR U13295 ( .A(n13129), .B(n13130), .Z(n13128) );
  ANDN U13296 ( .B(n13131), .A(n13132), .Z(n13130) );
  XOR U13297 ( .A(n13117), .B(n13101), .Z(n11097) );
  XNOR U13298 ( .A(n13133), .B(n13134), .Z(n13101) );
  XOR U13299 ( .A(n13135), .B(n13136), .Z(n13134) );
  NOR U13300 ( .A(n13137), .B(n13138), .Z(n13135) );
  XOR U13301 ( .A(n9954), .B(n13139), .Z(n13121) );
  XOR U13302 ( .A(key[253]), .B(n9949), .Z(n13139) );
  XNOR U13303 ( .A(n13140), .B(n13141), .Z(n9949) );
  XNOR U13304 ( .A(n13142), .B(n13143), .Z(n9954) );
  XNOR U13305 ( .A(n13144), .B(n13145), .Z(n13143) );
  XOR U13306 ( .A(n13146), .B(n13147), .Z(n13142) );
  XNOR U13307 ( .A(n13148), .B(n13149), .Z(n13147) );
  ANDN U13308 ( .B(n13150), .A(n13151), .Z(n13149) );
  XOR U13309 ( .A(n13152), .B(n13153), .Z(n13091) );
  XNOR U13310 ( .A(n13107), .B(n13105), .Z(n13153) );
  XNOR U13311 ( .A(n13154), .B(n13155), .Z(n13105) );
  XOR U13312 ( .A(n9943), .B(n9924), .Z(n13155) );
  XNOR U13313 ( .A(n13156), .B(n13157), .Z(n9924) );
  XNOR U13314 ( .A(n13119), .B(n13145), .Z(n13157) );
  XOR U13315 ( .A(n13158), .B(n13159), .Z(n13145) );
  XNOR U13316 ( .A(n13160), .B(n13161), .Z(n13159) );
  OR U13317 ( .A(n13162), .B(n13163), .Z(n13161) );
  XOR U13318 ( .A(n13164), .B(n13165), .Z(n13156) );
  IV U13319 ( .A(n11117), .Z(n9943) );
  XOR U13320 ( .A(n9128), .B(n9149), .Z(n11117) );
  XNOR U13321 ( .A(key[255]), .B(n11092), .Z(n13154) );
  XNOR U13322 ( .A(n9922), .B(n9939), .Z(n11092) );
  XNOR U13323 ( .A(n13166), .B(n13167), .Z(n9939) );
  XOR U13324 ( .A(n13168), .B(n13126), .Z(n13167) );
  XNOR U13325 ( .A(n13169), .B(n13170), .Z(n13126) );
  XNOR U13326 ( .A(n13171), .B(n13172), .Z(n13170) );
  OR U13327 ( .A(n13173), .B(n13174), .Z(n13172) );
  XNOR U13328 ( .A(n13175), .B(n13176), .Z(n13166) );
  XNOR U13329 ( .A(n13177), .B(n13178), .Z(n9922) );
  XOR U13330 ( .A(n13179), .B(n13180), .Z(n13178) );
  XOR U13331 ( .A(n13140), .B(n13181), .Z(n13177) );
  XNOR U13332 ( .A(n13182), .B(n13183), .Z(n13107) );
  XNOR U13333 ( .A(n9931), .B(n9131), .Z(n13183) );
  XNOR U13334 ( .A(n9128), .B(n9952), .Z(n9131) );
  XOR U13335 ( .A(n13184), .B(n13185), .Z(n9952) );
  XNOR U13336 ( .A(n13186), .B(n13180), .Z(n13185) );
  XNOR U13337 ( .A(n13187), .B(n13188), .Z(n13180) );
  XNOR U13338 ( .A(n13189), .B(n13190), .Z(n13188) );
  OR U13339 ( .A(n13191), .B(n13192), .Z(n13190) );
  XNOR U13340 ( .A(n13193), .B(n13194), .Z(n13184) );
  XNOR U13341 ( .A(n13195), .B(n13196), .Z(n13194) );
  ANDN U13342 ( .B(n13197), .A(n13198), .Z(n13196) );
  XNOR U13343 ( .A(n13146), .B(n9913), .Z(n9931) );
  XNOR U13344 ( .A(n13199), .B(n13164), .Z(n9913) );
  XNOR U13345 ( .A(n11080), .B(n13200), .Z(n13182) );
  XNOR U13346 ( .A(key[252]), .B(n11081), .Z(n13200) );
  XNOR U13347 ( .A(n9934), .B(n9133), .Z(n11081) );
  XOR U13348 ( .A(n13127), .B(n9104), .Z(n9133) );
  XNOR U13349 ( .A(n13201), .B(n13202), .Z(n9104) );
  XOR U13350 ( .A(n13112), .B(n9953), .Z(n11080) );
  XOR U13351 ( .A(n13203), .B(n13204), .Z(n9953) );
  XNOR U13352 ( .A(n13205), .B(n13116), .Z(n13204) );
  XNOR U13353 ( .A(n13206), .B(n13207), .Z(n13116) );
  XNOR U13354 ( .A(n13208), .B(n13209), .Z(n13207) );
  OR U13355 ( .A(n13210), .B(n13211), .Z(n13209) );
  XNOR U13356 ( .A(n13212), .B(n13213), .Z(n13203) );
  XNOR U13357 ( .A(n13136), .B(n13214), .Z(n13213) );
  ANDN U13358 ( .B(n13215), .A(n13216), .Z(n13214) );
  NANDN U13359 ( .A(n13217), .B(n13218), .Z(n13136) );
  XNOR U13360 ( .A(n11509), .B(n13085), .Z(n13152) );
  XOR U13361 ( .A(n13219), .B(n13220), .Z(n13085) );
  XNOR U13362 ( .A(n9144), .B(n13221), .Z(n13220) );
  XNOR U13363 ( .A(n13222), .B(n13223), .Z(n9900) );
  XNOR U13364 ( .A(n13224), .B(n13120), .Z(n13223) );
  XNOR U13365 ( .A(n13225), .B(n13226), .Z(n13120) );
  XOR U13366 ( .A(n13227), .B(n13148), .Z(n13226) );
  NANDN U13367 ( .A(n13228), .B(n13229), .Z(n13148) );
  NOR U13368 ( .A(n13230), .B(n13231), .Z(n13227) );
  XNOR U13369 ( .A(n13164), .B(n13232), .Z(n13222) );
  XOR U13370 ( .A(n13233), .B(n13234), .Z(n13089) );
  XNOR U13371 ( .A(n13235), .B(n9150), .Z(n13234) );
  XOR U13372 ( .A(n9915), .B(n9942), .Z(n9150) );
  IV U13373 ( .A(n9143), .Z(n9942) );
  XOR U13374 ( .A(n13168), .B(n13236), .Z(n9143) );
  XOR U13375 ( .A(n13175), .B(n13176), .Z(n13236) );
  IV U13376 ( .A(n13111), .Z(n13168) );
  XOR U13377 ( .A(n13201), .B(n13237), .Z(n13111) );
  XOR U13378 ( .A(n9944), .B(n13238), .Z(n13233) );
  XNOR U13379 ( .A(key[249]), .B(n11105), .Z(n13238) );
  XOR U13380 ( .A(n13119), .B(n13239), .Z(n9944) );
  XOR U13381 ( .A(n13164), .B(n13232), .Z(n13239) );
  IV U13382 ( .A(n13165), .Z(n13232) );
  XOR U13383 ( .A(n13225), .B(n13240), .Z(n13165) );
  XNOR U13384 ( .A(n13241), .B(n13242), .Z(n13240) );
  OR U13385 ( .A(n13162), .B(n13243), .Z(n13242) );
  XNOR U13386 ( .A(n13144), .B(n13244), .Z(n13225) );
  XNOR U13387 ( .A(n13245), .B(n13246), .Z(n13244) );
  OR U13388 ( .A(n13247), .B(n13248), .Z(n13246) );
  XOR U13389 ( .A(n13249), .B(n13250), .Z(n13164) );
  XOR U13390 ( .A(n13251), .B(n13252), .Z(n13250) );
  OR U13391 ( .A(n13253), .B(n13151), .Z(n13252) );
  XNOR U13392 ( .A(n13199), .B(n13224), .Z(n13119) );
  XNOR U13393 ( .A(n13144), .B(n13254), .Z(n13224) );
  XNOR U13394 ( .A(n13241), .B(n13255), .Z(n13254) );
  NANDN U13395 ( .A(n13256), .B(n13257), .Z(n13255) );
  OR U13396 ( .A(n13258), .B(n13259), .Z(n13241) );
  XOR U13397 ( .A(n13260), .B(n13245), .Z(n13144) );
  NANDN U13398 ( .A(n13261), .B(n13262), .Z(n13245) );
  AND U13399 ( .A(n13263), .B(n13264), .Z(n13260) );
  XNOR U13400 ( .A(n9128), .B(n9934), .Z(n9144) );
  XOR U13401 ( .A(n13193), .B(n9901), .Z(n9934) );
  IV U13402 ( .A(n13235), .Z(n9901) );
  XOR U13403 ( .A(n13265), .B(n13181), .Z(n13235) );
  XNOR U13404 ( .A(n11107), .B(n13266), .Z(n13219) );
  XNOR U13405 ( .A(key[251]), .B(n11109), .Z(n13266) );
  IV U13406 ( .A(n9106), .Z(n11109) );
  XOR U13407 ( .A(n9146), .B(n9918), .Z(n9106) );
  XOR U13408 ( .A(n13267), .B(n13268), .Z(n9918) );
  XNOR U13409 ( .A(n13269), .B(n13141), .Z(n13268) );
  XNOR U13410 ( .A(n13270), .B(n13271), .Z(n13141) );
  XOR U13411 ( .A(n13272), .B(n13195), .Z(n13271) );
  NANDN U13412 ( .A(n13273), .B(n13274), .Z(n13195) );
  NOR U13413 ( .A(n13275), .B(n13276), .Z(n13272) );
  XNOR U13414 ( .A(n13277), .B(n13181), .Z(n13267) );
  XOR U13415 ( .A(n13278), .B(n13279), .Z(n9146) );
  XOR U13416 ( .A(n13176), .B(n13110), .Z(n13279) );
  XNOR U13417 ( .A(n13280), .B(n13281), .Z(n13110) );
  XOR U13418 ( .A(n13282), .B(n13129), .Z(n13281) );
  NANDN U13419 ( .A(n13283), .B(n13284), .Z(n13129) );
  NOR U13420 ( .A(n13285), .B(n13286), .Z(n13282) );
  XOR U13421 ( .A(n13280), .B(n13287), .Z(n13176) );
  XNOR U13422 ( .A(n13288), .B(n13289), .Z(n13287) );
  OR U13423 ( .A(n13173), .B(n13290), .Z(n13289) );
  XNOR U13424 ( .A(n13125), .B(n13291), .Z(n13280) );
  XNOR U13425 ( .A(n13292), .B(n13293), .Z(n13291) );
  OR U13426 ( .A(n13294), .B(n13295), .Z(n13293) );
  XNOR U13427 ( .A(n13175), .B(n13237), .Z(n13278) );
  XOR U13428 ( .A(n13125), .B(n13296), .Z(n13237) );
  XNOR U13429 ( .A(n13288), .B(n13297), .Z(n13296) );
  NANDN U13430 ( .A(n13298), .B(n13299), .Z(n13297) );
  OR U13431 ( .A(n13300), .B(n13301), .Z(n13288) );
  XOR U13432 ( .A(n13302), .B(n13292), .Z(n13125) );
  NANDN U13433 ( .A(n13303), .B(n13304), .Z(n13292) );
  AND U13434 ( .A(n13305), .B(n13306), .Z(n13302) );
  IV U13435 ( .A(n13202), .Z(n13175) );
  XOR U13436 ( .A(n13307), .B(n13308), .Z(n13202) );
  XOR U13437 ( .A(n13309), .B(n13310), .Z(n13308) );
  OR U13438 ( .A(n13311), .B(n13132), .Z(n13310) );
  XOR U13439 ( .A(n13112), .B(n9930), .Z(n11107) );
  XOR U13440 ( .A(n13312), .B(n13103), .Z(n11105) );
  IV U13441 ( .A(n9149), .Z(n13112) );
  XOR U13442 ( .A(n13313), .B(n13205), .Z(n9149) );
  XNOR U13443 ( .A(n13206), .B(n13314), .Z(n13205) );
  XOR U13444 ( .A(n13315), .B(n13316), .Z(n13314) );
  NOR U13445 ( .A(n13317), .B(n13138), .Z(n13315) );
  XNOR U13446 ( .A(n13318), .B(n13319), .Z(n13206) );
  XNOR U13447 ( .A(n13320), .B(n13321), .Z(n13319) );
  NANDN U13448 ( .A(n13322), .B(n13323), .Z(n13321) );
  XNOR U13449 ( .A(n13324), .B(n13325), .Z(n11509) );
  XOR U13450 ( .A(n9915), .B(n9925), .Z(n13325) );
  IV U13451 ( .A(n9151), .Z(n9925) );
  XNOR U13452 ( .A(n9946), .B(n9916), .Z(n9151) );
  XOR U13453 ( .A(n13201), .B(n13127), .Z(n9916) );
  XNOR U13454 ( .A(n13169), .B(n13326), .Z(n13127) );
  XNOR U13455 ( .A(n13327), .B(n13309), .Z(n13326) );
  ANDN U13456 ( .B(n13284), .A(n13328), .Z(n13309) );
  XOR U13457 ( .A(n13286), .B(n13132), .Z(n13284) );
  NOR U13458 ( .A(n13329), .B(n13286), .Z(n13327) );
  XNOR U13459 ( .A(n13307), .B(n13330), .Z(n13169) );
  XNOR U13460 ( .A(n13331), .B(n13332), .Z(n13330) );
  NANDN U13461 ( .A(n13294), .B(n13333), .Z(n13332) );
  XNOR U13462 ( .A(n13307), .B(n13334), .Z(n13201) );
  XOR U13463 ( .A(n13335), .B(n13171), .Z(n13334) );
  OR U13464 ( .A(n13336), .B(n13300), .Z(n13171) );
  XOR U13465 ( .A(n13173), .B(n13337), .Z(n13300) );
  ANDN U13466 ( .B(n13338), .A(n13298), .Z(n13335) );
  XOR U13467 ( .A(n13339), .B(n13331), .Z(n13307) );
  OR U13468 ( .A(n13303), .B(n13340), .Z(n13331) );
  XOR U13469 ( .A(n13305), .B(n13294), .Z(n13303) );
  XOR U13470 ( .A(n13337), .B(n13132), .Z(n13294) );
  XNOR U13471 ( .A(n13341), .B(n13342), .Z(n13132) );
  NANDN U13472 ( .A(n13343), .B(n13344), .Z(n13342) );
  IV U13473 ( .A(n13298), .Z(n13337) );
  XNOR U13474 ( .A(n13345), .B(n13346), .Z(n13298) );
  NANDN U13475 ( .A(n13343), .B(n13347), .Z(n13346) );
  ANDN U13476 ( .B(n13305), .A(n13348), .Z(n13339) );
  XOR U13477 ( .A(n13286), .B(n13173), .Z(n13305) );
  XOR U13478 ( .A(n13349), .B(n13345), .Z(n13173) );
  NANDN U13479 ( .A(n13350), .B(n13351), .Z(n13345) );
  NANDN U13480 ( .A(n13350), .B(n13355), .Z(n13341) );
  XOR U13481 ( .A(n13356), .B(n13357), .Z(n13343) );
  XOR U13482 ( .A(n13358), .B(n13353), .Z(n13357) );
  XNOR U13483 ( .A(n13359), .B(n13360), .Z(n13356) );
  XNOR U13484 ( .A(n13361), .B(n13362), .Z(n13360) );
  ANDN U13485 ( .B(n13358), .A(n13353), .Z(n13361) );
  ANDN U13486 ( .B(n13358), .A(n13352), .Z(n13354) );
  XNOR U13487 ( .A(n13359), .B(n13363), .Z(n13352) );
  XOR U13488 ( .A(n13364), .B(n13362), .Z(n13363) );
  NAND U13489 ( .A(n13351), .B(n13355), .Z(n13362) );
  XNOR U13490 ( .A(n13347), .B(n13353), .Z(n13351) );
  XOR U13491 ( .A(n13365), .B(n13366), .Z(n13353) );
  XOR U13492 ( .A(n13367), .B(n13368), .Z(n13366) );
  XNOR U13493 ( .A(n13369), .B(n13370), .Z(n13365) );
  ANDN U13494 ( .B(n13371), .A(n13285), .Z(n13369) );
  AND U13495 ( .A(n13344), .B(n13347), .Z(n13364) );
  XNOR U13496 ( .A(n13344), .B(n13347), .Z(n13359) );
  XNOR U13497 ( .A(n13372), .B(n13373), .Z(n13347) );
  XNOR U13498 ( .A(n13374), .B(n13375), .Z(n13373) );
  XOR U13499 ( .A(n13367), .B(n13376), .Z(n13372) );
  XNOR U13500 ( .A(n13377), .B(n13370), .Z(n13376) );
  OR U13501 ( .A(n13283), .B(n13328), .Z(n13370) );
  XNOR U13502 ( .A(n13329), .B(n13311), .Z(n13328) );
  XNOR U13503 ( .A(n13285), .B(n13378), .Z(n13283) );
  NOR U13504 ( .A(n13378), .B(n13311), .Z(n13377) );
  XNOR U13505 ( .A(n13379), .B(n13380), .Z(n13344) );
  XNOR U13506 ( .A(n13381), .B(n13382), .Z(n13380) );
  XOR U13507 ( .A(n13290), .B(n13367), .Z(n13382) );
  XOR U13508 ( .A(n13371), .B(n13383), .Z(n13367) );
  XNOR U13509 ( .A(n13174), .B(n13384), .Z(n13379) );
  XNOR U13510 ( .A(n13385), .B(n13386), .Z(n13384) );
  ANDN U13511 ( .B(n13299), .A(n13387), .Z(n13385) );
  XNOR U13512 ( .A(n13388), .B(n13389), .Z(n13358) );
  XNOR U13513 ( .A(n13368), .B(n13390), .Z(n13389) );
  XNOR U13514 ( .A(n13299), .B(n13375), .Z(n13390) );
  XOR U13515 ( .A(n13311), .B(n13378), .Z(n13375) );
  XNOR U13516 ( .A(n13381), .B(n13391), .Z(n13368) );
  XNOR U13517 ( .A(n13392), .B(n13393), .Z(n13391) );
  NANDN U13518 ( .A(n13295), .B(n13333), .Z(n13393) );
  IV U13519 ( .A(n13374), .Z(n13381) );
  XNOR U13520 ( .A(n13394), .B(n13392), .Z(n13374) );
  NANDN U13521 ( .A(n13340), .B(n13304), .Z(n13392) );
  XOR U13522 ( .A(n13299), .B(n13378), .Z(n13295) );
  IV U13523 ( .A(n13131), .Z(n13378) );
  XOR U13524 ( .A(n13395), .B(n13396), .Z(n13131) );
  XNOR U13525 ( .A(n13397), .B(n13398), .Z(n13396) );
  XOR U13526 ( .A(n13348), .B(n13333), .Z(n13340) );
  XNOR U13527 ( .A(n13338), .B(n13311), .Z(n13333) );
  XNOR U13528 ( .A(n13398), .B(n13395), .Z(n13311) );
  ANDN U13529 ( .B(n13306), .A(n13348), .Z(n13394) );
  XNOR U13530 ( .A(n13399), .B(n13371), .Z(n13348) );
  IV U13531 ( .A(n13329), .Z(n13371) );
  XNOR U13532 ( .A(n13400), .B(n13401), .Z(n13329) );
  XNOR U13533 ( .A(n13402), .B(n13398), .Z(n13401) );
  XOR U13534 ( .A(n13403), .B(n13383), .Z(n13306) );
  XNOR U13535 ( .A(n13387), .B(n13404), .Z(n13388) );
  XNOR U13536 ( .A(n13405), .B(n13386), .Z(n13404) );
  OR U13537 ( .A(n13301), .B(n13336), .Z(n13386) );
  XOR U13538 ( .A(n13174), .B(n13338), .Z(n13336) );
  IV U13539 ( .A(n13387), .Z(n13338) );
  XOR U13540 ( .A(n13290), .B(n13299), .Z(n13301) );
  XNOR U13541 ( .A(n13383), .B(n13406), .Z(n13299) );
  XNOR U13542 ( .A(n13397), .B(n13400), .Z(n13406) );
  XNOR U13543 ( .A(state[42]), .B(key[42]), .Z(n13400) );
  IV U13544 ( .A(n13285), .Z(n13383) );
  XOR U13545 ( .A(n13407), .B(n13408), .Z(n13285) );
  XOR U13546 ( .A(n13398), .B(n13409), .Z(n13408) );
  IV U13547 ( .A(n13403), .Z(n13290) );
  ANDN U13548 ( .B(n13403), .A(n13174), .Z(n13405) );
  XOR U13549 ( .A(n13395), .B(n13410), .Z(n13403) );
  XNOR U13550 ( .A(n13398), .B(n13411), .Z(n13410) );
  XOR U13551 ( .A(n13399), .B(n13412), .Z(n13398) );
  XNOR U13552 ( .A(state[46]), .B(key[46]), .Z(n13412) );
  IV U13553 ( .A(n13407), .Z(n13395) );
  XOR U13554 ( .A(state[45]), .B(key[45]), .Z(n13407) );
  XOR U13555 ( .A(n13413), .B(n13414), .Z(n13387) );
  XOR U13556 ( .A(n13411), .B(n13409), .Z(n13414) );
  XOR U13557 ( .A(state[47]), .B(key[47]), .Z(n13409) );
  XNOR U13558 ( .A(state[44]), .B(key[44]), .Z(n13411) );
  XOR U13559 ( .A(n13174), .B(n13402), .Z(n13413) );
  XNOR U13560 ( .A(n13397), .B(n13415), .Z(n13402) );
  XNOR U13561 ( .A(state[43]), .B(key[43]), .Z(n13415) );
  XNOR U13562 ( .A(state[41]), .B(key[41]), .Z(n13397) );
  IV U13563 ( .A(n13399), .Z(n13174) );
  XOR U13564 ( .A(state[40]), .B(key[40]), .Z(n13399) );
  IV U13565 ( .A(n11093), .Z(n9946) );
  XOR U13566 ( .A(n13146), .B(n13199), .Z(n11093) );
  XNOR U13567 ( .A(n13249), .B(n13416), .Z(n13199) );
  XOR U13568 ( .A(n13417), .B(n13160), .Z(n13416) );
  OR U13569 ( .A(n13418), .B(n13258), .Z(n13160) );
  XOR U13570 ( .A(n13162), .B(n13419), .Z(n13258) );
  ANDN U13571 ( .B(n13420), .A(n13256), .Z(n13417) );
  XNOR U13572 ( .A(n13158), .B(n13421), .Z(n13146) );
  XNOR U13573 ( .A(n13422), .B(n13251), .Z(n13421) );
  ANDN U13574 ( .B(n13229), .A(n13423), .Z(n13251) );
  XOR U13575 ( .A(n13231), .B(n13151), .Z(n13229) );
  NOR U13576 ( .A(n13424), .B(n13231), .Z(n13422) );
  XOR U13577 ( .A(n13249), .B(n13425), .Z(n13158) );
  XNOR U13578 ( .A(n13426), .B(n13427), .Z(n13425) );
  NANDN U13579 ( .A(n13247), .B(n13428), .Z(n13427) );
  XOR U13580 ( .A(n13429), .B(n13426), .Z(n13249) );
  OR U13581 ( .A(n13261), .B(n13430), .Z(n13426) );
  XOR U13582 ( .A(n13263), .B(n13247), .Z(n13261) );
  XOR U13583 ( .A(n13419), .B(n13151), .Z(n13247) );
  XNOR U13584 ( .A(n13431), .B(n13432), .Z(n13151) );
  NANDN U13585 ( .A(n13433), .B(n13434), .Z(n13432) );
  IV U13586 ( .A(n13256), .Z(n13419) );
  XNOR U13587 ( .A(n13435), .B(n13436), .Z(n13256) );
  NANDN U13588 ( .A(n13433), .B(n13437), .Z(n13436) );
  ANDN U13589 ( .B(n13263), .A(n13438), .Z(n13429) );
  XOR U13590 ( .A(n13231), .B(n13162), .Z(n13263) );
  XOR U13591 ( .A(n13439), .B(n13435), .Z(n13162) );
  NANDN U13592 ( .A(n13440), .B(n13441), .Z(n13435) );
  NANDN U13593 ( .A(n13440), .B(n13445), .Z(n13431) );
  XOR U13594 ( .A(n13446), .B(n13447), .Z(n13433) );
  XOR U13595 ( .A(n13448), .B(n13443), .Z(n13447) );
  XNOR U13596 ( .A(n13449), .B(n13450), .Z(n13446) );
  XNOR U13597 ( .A(n13451), .B(n13452), .Z(n13450) );
  ANDN U13598 ( .B(n13448), .A(n13443), .Z(n13451) );
  ANDN U13599 ( .B(n13448), .A(n13442), .Z(n13444) );
  XNOR U13600 ( .A(n13449), .B(n13453), .Z(n13442) );
  XOR U13601 ( .A(n13454), .B(n13452), .Z(n13453) );
  NAND U13602 ( .A(n13441), .B(n13445), .Z(n13452) );
  XNOR U13603 ( .A(n13437), .B(n13443), .Z(n13441) );
  XOR U13604 ( .A(n13455), .B(n13456), .Z(n13443) );
  XOR U13605 ( .A(n13457), .B(n13458), .Z(n13456) );
  XNOR U13606 ( .A(n13459), .B(n13460), .Z(n13455) );
  ANDN U13607 ( .B(n13461), .A(n13230), .Z(n13459) );
  AND U13608 ( .A(n13434), .B(n13437), .Z(n13454) );
  XNOR U13609 ( .A(n13434), .B(n13437), .Z(n13449) );
  XNOR U13610 ( .A(n13462), .B(n13463), .Z(n13437) );
  XNOR U13611 ( .A(n13464), .B(n13465), .Z(n13463) );
  XOR U13612 ( .A(n13457), .B(n13466), .Z(n13462) );
  XNOR U13613 ( .A(n13467), .B(n13460), .Z(n13466) );
  OR U13614 ( .A(n13228), .B(n13423), .Z(n13460) );
  XNOR U13615 ( .A(n13424), .B(n13253), .Z(n13423) );
  XNOR U13616 ( .A(n13230), .B(n13468), .Z(n13228) );
  NOR U13617 ( .A(n13468), .B(n13253), .Z(n13467) );
  XNOR U13618 ( .A(n13469), .B(n13470), .Z(n13434) );
  XNOR U13619 ( .A(n13471), .B(n13472), .Z(n13470) );
  XOR U13620 ( .A(n13243), .B(n13457), .Z(n13472) );
  XOR U13621 ( .A(n13461), .B(n13473), .Z(n13457) );
  XNOR U13622 ( .A(n13163), .B(n13474), .Z(n13469) );
  XNOR U13623 ( .A(n13475), .B(n13476), .Z(n13474) );
  ANDN U13624 ( .B(n13257), .A(n13477), .Z(n13475) );
  XNOR U13625 ( .A(n13478), .B(n13479), .Z(n13448) );
  XNOR U13626 ( .A(n13458), .B(n13480), .Z(n13479) );
  XNOR U13627 ( .A(n13257), .B(n13465), .Z(n13480) );
  XOR U13628 ( .A(n13253), .B(n13468), .Z(n13465) );
  XNOR U13629 ( .A(n13471), .B(n13481), .Z(n13458) );
  XNOR U13630 ( .A(n13482), .B(n13483), .Z(n13481) );
  NANDN U13631 ( .A(n13248), .B(n13428), .Z(n13483) );
  IV U13632 ( .A(n13464), .Z(n13471) );
  XNOR U13633 ( .A(n13484), .B(n13482), .Z(n13464) );
  NANDN U13634 ( .A(n13430), .B(n13262), .Z(n13482) );
  XOR U13635 ( .A(n13257), .B(n13468), .Z(n13248) );
  IV U13636 ( .A(n13150), .Z(n13468) );
  XOR U13637 ( .A(n13485), .B(n13486), .Z(n13150) );
  XNOR U13638 ( .A(n13487), .B(n13488), .Z(n13486) );
  XOR U13639 ( .A(n13438), .B(n13428), .Z(n13430) );
  XNOR U13640 ( .A(n13420), .B(n13253), .Z(n13428) );
  XNOR U13641 ( .A(n13488), .B(n13485), .Z(n13253) );
  ANDN U13642 ( .B(n13264), .A(n13438), .Z(n13484) );
  XNOR U13643 ( .A(n13489), .B(n13461), .Z(n13438) );
  IV U13644 ( .A(n13424), .Z(n13461) );
  XNOR U13645 ( .A(n13490), .B(n13491), .Z(n13424) );
  XNOR U13646 ( .A(n13492), .B(n13488), .Z(n13491) );
  XOR U13647 ( .A(n13493), .B(n13473), .Z(n13264) );
  XNOR U13648 ( .A(n13477), .B(n13494), .Z(n13478) );
  XNOR U13649 ( .A(n13495), .B(n13476), .Z(n13494) );
  OR U13650 ( .A(n13259), .B(n13418), .Z(n13476) );
  XOR U13651 ( .A(n13163), .B(n13420), .Z(n13418) );
  IV U13652 ( .A(n13477), .Z(n13420) );
  XOR U13653 ( .A(n13243), .B(n13257), .Z(n13259) );
  XNOR U13654 ( .A(n13473), .B(n13496), .Z(n13257) );
  XNOR U13655 ( .A(n13487), .B(n13490), .Z(n13496) );
  XNOR U13656 ( .A(state[2]), .B(key[2]), .Z(n13490) );
  IV U13657 ( .A(n13230), .Z(n13473) );
  XOR U13658 ( .A(n13497), .B(n13498), .Z(n13230) );
  XOR U13659 ( .A(n13488), .B(n13499), .Z(n13498) );
  IV U13660 ( .A(n13493), .Z(n13243) );
  ANDN U13661 ( .B(n13493), .A(n13163), .Z(n13495) );
  XOR U13662 ( .A(n13485), .B(n13500), .Z(n13493) );
  XNOR U13663 ( .A(n13488), .B(n13501), .Z(n13500) );
  XOR U13664 ( .A(n13489), .B(n13502), .Z(n13488) );
  XNOR U13665 ( .A(state[6]), .B(key[6]), .Z(n13502) );
  IV U13666 ( .A(n13497), .Z(n13485) );
  XOR U13667 ( .A(state[5]), .B(key[5]), .Z(n13497) );
  XOR U13668 ( .A(n13503), .B(n13504), .Z(n13477) );
  XOR U13669 ( .A(n13501), .B(n13499), .Z(n13504) );
  XOR U13670 ( .A(state[7]), .B(key[7]), .Z(n13499) );
  XNOR U13671 ( .A(state[4]), .B(key[4]), .Z(n13501) );
  XOR U13672 ( .A(n13163), .B(n13492), .Z(n13503) );
  XNOR U13673 ( .A(n13487), .B(n13505), .Z(n13492) );
  XNOR U13674 ( .A(state[3]), .B(key[3]), .Z(n13505) );
  XNOR U13675 ( .A(state[1]), .B(key[1]), .Z(n13487) );
  IV U13676 ( .A(n13489), .Z(n13163) );
  XOR U13677 ( .A(state[0]), .B(key[0]), .Z(n13489) );
  XOR U13678 ( .A(n13179), .B(n13506), .Z(n9915) );
  XNOR U13679 ( .A(n13140), .B(n13181), .Z(n13506) );
  XOR U13680 ( .A(n13507), .B(n13508), .Z(n13181) );
  XOR U13681 ( .A(n13509), .B(n13510), .Z(n13508) );
  OR U13682 ( .A(n13511), .B(n13198), .Z(n13510) );
  XOR U13683 ( .A(n13265), .B(n13277), .Z(n13140) );
  XNOR U13684 ( .A(n13186), .B(n13512), .Z(n13277) );
  XNOR U13685 ( .A(n13513), .B(n13514), .Z(n13512) );
  NANDN U13686 ( .A(n13515), .B(n13516), .Z(n13514) );
  IV U13687 ( .A(n13269), .Z(n13179) );
  XNOR U13688 ( .A(n13513), .B(n13518), .Z(n13517) );
  OR U13689 ( .A(n13191), .B(n13519), .Z(n13518) );
  OR U13690 ( .A(n13520), .B(n13521), .Z(n13513) );
  XNOR U13691 ( .A(n13186), .B(n13522), .Z(n13270) );
  XNOR U13692 ( .A(n13523), .B(n13524), .Z(n13522) );
  OR U13693 ( .A(n13525), .B(n13526), .Z(n13524) );
  XOR U13694 ( .A(n13527), .B(n13523), .Z(n13186) );
  NANDN U13695 ( .A(n13528), .B(n13529), .Z(n13523) );
  AND U13696 ( .A(n13530), .B(n13531), .Z(n13527) );
  XNOR U13697 ( .A(n11106), .B(n13532), .Z(n13324) );
  XNOR U13698 ( .A(key[248]), .B(n9128), .Z(n13532) );
  XNOR U13699 ( .A(n13187), .B(n13533), .Z(n13193) );
  XNOR U13700 ( .A(n13534), .B(n13509), .Z(n13533) );
  ANDN U13701 ( .B(n13274), .A(n13535), .Z(n13509) );
  XOR U13702 ( .A(n13276), .B(n13198), .Z(n13274) );
  NOR U13703 ( .A(n13536), .B(n13276), .Z(n13534) );
  XNOR U13704 ( .A(n13507), .B(n13537), .Z(n13187) );
  XNOR U13705 ( .A(n13538), .B(n13539), .Z(n13537) );
  NANDN U13706 ( .A(n13525), .B(n13540), .Z(n13539) );
  XNOR U13707 ( .A(n13507), .B(n13541), .Z(n13265) );
  XOR U13708 ( .A(n13542), .B(n13189), .Z(n13541) );
  OR U13709 ( .A(n13543), .B(n13520), .Z(n13189) );
  XOR U13710 ( .A(n13191), .B(n13544), .Z(n13520) );
  ANDN U13711 ( .B(n13545), .A(n13515), .Z(n13542) );
  XOR U13712 ( .A(n13546), .B(n13538), .Z(n13507) );
  OR U13713 ( .A(n13528), .B(n13547), .Z(n13538) );
  XOR U13714 ( .A(n13530), .B(n13525), .Z(n13528) );
  XOR U13715 ( .A(n13544), .B(n13198), .Z(n13525) );
  XNOR U13716 ( .A(n13548), .B(n13549), .Z(n13198) );
  NANDN U13717 ( .A(n13550), .B(n13551), .Z(n13549) );
  IV U13718 ( .A(n13515), .Z(n13544) );
  XNOR U13719 ( .A(n13552), .B(n13553), .Z(n13515) );
  NANDN U13720 ( .A(n13550), .B(n13554), .Z(n13553) );
  ANDN U13721 ( .B(n13530), .A(n13555), .Z(n13546) );
  XOR U13722 ( .A(n13276), .B(n13191), .Z(n13530) );
  XOR U13723 ( .A(n13556), .B(n13552), .Z(n13191) );
  NANDN U13724 ( .A(n13557), .B(n13558), .Z(n13552) );
  NANDN U13725 ( .A(n13557), .B(n13562), .Z(n13548) );
  XOR U13726 ( .A(n13563), .B(n13564), .Z(n13550) );
  XOR U13727 ( .A(n13565), .B(n13560), .Z(n13564) );
  XNOR U13728 ( .A(n13566), .B(n13567), .Z(n13563) );
  XNOR U13729 ( .A(n13568), .B(n13569), .Z(n13567) );
  ANDN U13730 ( .B(n13565), .A(n13560), .Z(n13568) );
  ANDN U13731 ( .B(n13565), .A(n13559), .Z(n13561) );
  XNOR U13732 ( .A(n13566), .B(n13570), .Z(n13559) );
  XOR U13733 ( .A(n13571), .B(n13569), .Z(n13570) );
  NAND U13734 ( .A(n13558), .B(n13562), .Z(n13569) );
  XNOR U13735 ( .A(n13554), .B(n13560), .Z(n13558) );
  XOR U13736 ( .A(n13572), .B(n13573), .Z(n13560) );
  XOR U13737 ( .A(n13574), .B(n13575), .Z(n13573) );
  XNOR U13738 ( .A(n13576), .B(n13577), .Z(n13572) );
  ANDN U13739 ( .B(n13578), .A(n13275), .Z(n13576) );
  AND U13740 ( .A(n13551), .B(n13554), .Z(n13571) );
  XNOR U13741 ( .A(n13551), .B(n13554), .Z(n13566) );
  XNOR U13742 ( .A(n13579), .B(n13580), .Z(n13554) );
  XNOR U13743 ( .A(n13581), .B(n13582), .Z(n13580) );
  XOR U13744 ( .A(n13574), .B(n13583), .Z(n13579) );
  XNOR U13745 ( .A(n13584), .B(n13577), .Z(n13583) );
  OR U13746 ( .A(n13273), .B(n13535), .Z(n13577) );
  XNOR U13747 ( .A(n13536), .B(n13511), .Z(n13535) );
  XNOR U13748 ( .A(n13275), .B(n13585), .Z(n13273) );
  NOR U13749 ( .A(n13585), .B(n13511), .Z(n13584) );
  XNOR U13750 ( .A(n13586), .B(n13587), .Z(n13551) );
  XNOR U13751 ( .A(n13588), .B(n13589), .Z(n13587) );
  XOR U13752 ( .A(n13519), .B(n13574), .Z(n13589) );
  XOR U13753 ( .A(n13578), .B(n13590), .Z(n13574) );
  XNOR U13754 ( .A(n13192), .B(n13591), .Z(n13586) );
  XNOR U13755 ( .A(n13592), .B(n13593), .Z(n13591) );
  ANDN U13756 ( .B(n13516), .A(n13594), .Z(n13592) );
  XNOR U13757 ( .A(n13595), .B(n13596), .Z(n13565) );
  XNOR U13758 ( .A(n13575), .B(n13597), .Z(n13596) );
  XNOR U13759 ( .A(n13516), .B(n13582), .Z(n13597) );
  XOR U13760 ( .A(n13511), .B(n13585), .Z(n13582) );
  XNOR U13761 ( .A(n13588), .B(n13598), .Z(n13575) );
  XNOR U13762 ( .A(n13599), .B(n13600), .Z(n13598) );
  NANDN U13763 ( .A(n13526), .B(n13540), .Z(n13600) );
  IV U13764 ( .A(n13581), .Z(n13588) );
  XNOR U13765 ( .A(n13601), .B(n13599), .Z(n13581) );
  NANDN U13766 ( .A(n13547), .B(n13529), .Z(n13599) );
  XOR U13767 ( .A(n13516), .B(n13585), .Z(n13526) );
  IV U13768 ( .A(n13197), .Z(n13585) );
  XOR U13769 ( .A(n13602), .B(n13603), .Z(n13197) );
  XNOR U13770 ( .A(n13604), .B(n13605), .Z(n13603) );
  XOR U13771 ( .A(n13555), .B(n13540), .Z(n13547) );
  XNOR U13772 ( .A(n13545), .B(n13511), .Z(n13540) );
  XNOR U13773 ( .A(n13605), .B(n13602), .Z(n13511) );
  ANDN U13774 ( .B(n13531), .A(n13555), .Z(n13601) );
  XNOR U13775 ( .A(n13606), .B(n13578), .Z(n13555) );
  IV U13776 ( .A(n13536), .Z(n13578) );
  XNOR U13777 ( .A(n13607), .B(n13608), .Z(n13536) );
  XNOR U13778 ( .A(n13609), .B(n13605), .Z(n13608) );
  XOR U13779 ( .A(n13610), .B(n13590), .Z(n13531) );
  XNOR U13780 ( .A(n13594), .B(n13611), .Z(n13595) );
  XNOR U13781 ( .A(n13612), .B(n13593), .Z(n13611) );
  OR U13782 ( .A(n13521), .B(n13543), .Z(n13593) );
  XOR U13783 ( .A(n13192), .B(n13545), .Z(n13543) );
  IV U13784 ( .A(n13594), .Z(n13545) );
  XOR U13785 ( .A(n13519), .B(n13516), .Z(n13521) );
  XNOR U13786 ( .A(n13590), .B(n13613), .Z(n13516) );
  XNOR U13787 ( .A(n13604), .B(n13607), .Z(n13613) );
  XNOR U13788 ( .A(state[82]), .B(key[82]), .Z(n13607) );
  IV U13789 ( .A(n13275), .Z(n13590) );
  XOR U13790 ( .A(n13614), .B(n13615), .Z(n13275) );
  XOR U13791 ( .A(n13605), .B(n13616), .Z(n13615) );
  IV U13792 ( .A(n13610), .Z(n13519) );
  ANDN U13793 ( .B(n13610), .A(n13192), .Z(n13612) );
  XOR U13794 ( .A(n13602), .B(n13617), .Z(n13610) );
  XNOR U13795 ( .A(n13605), .B(n13618), .Z(n13617) );
  XOR U13796 ( .A(n13606), .B(n13619), .Z(n13605) );
  XNOR U13797 ( .A(state[86]), .B(key[86]), .Z(n13619) );
  IV U13798 ( .A(n13614), .Z(n13602) );
  XOR U13799 ( .A(state[85]), .B(key[85]), .Z(n13614) );
  XOR U13800 ( .A(n13620), .B(n13621), .Z(n13594) );
  XOR U13801 ( .A(n13618), .B(n13616), .Z(n13621) );
  XOR U13802 ( .A(state[87]), .B(key[87]), .Z(n13616) );
  XNOR U13803 ( .A(state[84]), .B(key[84]), .Z(n13618) );
  XOR U13804 ( .A(n13192), .B(n13609), .Z(n13620) );
  XNOR U13805 ( .A(n13604), .B(n13622), .Z(n13609) );
  XNOR U13806 ( .A(state[83]), .B(key[83]), .Z(n13622) );
  XNOR U13807 ( .A(state[81]), .B(key[81]), .Z(n13604) );
  IV U13808 ( .A(n13606), .Z(n13192) );
  XOR U13809 ( .A(state[80]), .B(key[80]), .Z(n13606) );
  XOR U13810 ( .A(n13100), .B(n13623), .Z(n11106) );
  XOR U13811 ( .A(n13117), .B(n13103), .Z(n13623) );
  XOR U13812 ( .A(n13318), .B(n13624), .Z(n13103) );
  XNOR U13813 ( .A(n13316), .B(n13625), .Z(n13624) );
  NANDN U13814 ( .A(n13626), .B(n13215), .Z(n13625) );
  NANDN U13815 ( .A(n13627), .B(n13218), .Z(n13316) );
  XNOR U13816 ( .A(n13138), .B(n13215), .Z(n13218) );
  XOR U13817 ( .A(n13313), .B(n13102), .Z(n13117) );
  XNOR U13818 ( .A(n13212), .B(n13628), .Z(n13102) );
  XNOR U13819 ( .A(n13629), .B(n13630), .Z(n13628) );
  NANDN U13820 ( .A(n13631), .B(n13632), .Z(n13630) );
  IV U13821 ( .A(n13312), .Z(n13313) );
  XNOR U13822 ( .A(n13318), .B(n13633), .Z(n13312) );
  XOR U13823 ( .A(n13634), .B(n13208), .Z(n13633) );
  OR U13824 ( .A(n13635), .B(n13636), .Z(n13208) );
  ANDN U13825 ( .B(n13637), .A(n13631), .Z(n13634) );
  XOR U13826 ( .A(n13638), .B(n13320), .Z(n13318) );
  OR U13827 ( .A(n13639), .B(n13640), .Z(n13320) );
  ANDN U13828 ( .B(n13641), .A(n13642), .Z(n13638) );
  IV U13829 ( .A(n13115), .Z(n13100) );
  XOR U13830 ( .A(n13133), .B(n13643), .Z(n13115) );
  XNOR U13831 ( .A(n13629), .B(n13644), .Z(n13643) );
  OR U13832 ( .A(n13210), .B(n13645), .Z(n13644) );
  OR U13833 ( .A(n13635), .B(n13646), .Z(n13629) );
  XOR U13834 ( .A(n13210), .B(n13647), .Z(n13635) );
  XOR U13835 ( .A(n13212), .B(n13648), .Z(n13133) );
  XNOR U13836 ( .A(n13649), .B(n13650), .Z(n13648) );
  OR U13837 ( .A(n13322), .B(n13651), .Z(n13650) );
  XOR U13838 ( .A(n13652), .B(n13649), .Z(n13212) );
  NANDN U13839 ( .A(n13639), .B(n13653), .Z(n13649) );
  XOR U13840 ( .A(n13641), .B(n13322), .Z(n13639) );
  XNOR U13841 ( .A(n13647), .B(n13215), .Z(n13322) );
  XOR U13842 ( .A(n13654), .B(n13655), .Z(n13215) );
  NANDN U13843 ( .A(n13656), .B(n13657), .Z(n13655) );
  IV U13844 ( .A(n13631), .Z(n13647) );
  XNOR U13845 ( .A(n13658), .B(n13659), .Z(n13631) );
  NANDN U13846 ( .A(n13656), .B(n13660), .Z(n13659) );
  XOR U13847 ( .A(n13138), .B(n13210), .Z(n13641) );
  XOR U13848 ( .A(n13662), .B(n13658), .Z(n13210) );
  NANDN U13849 ( .A(n13663), .B(n13664), .Z(n13658) );
  NANDN U13850 ( .A(n13663), .B(n13668), .Z(n13654) );
  XOR U13851 ( .A(n13669), .B(n13670), .Z(n13656) );
  XOR U13852 ( .A(n13671), .B(n13666), .Z(n13670) );
  XNOR U13853 ( .A(n13672), .B(n13673), .Z(n13669) );
  XNOR U13854 ( .A(n13674), .B(n13675), .Z(n13673) );
  ANDN U13855 ( .B(n13671), .A(n13666), .Z(n13674) );
  ANDN U13856 ( .B(n13671), .A(n13665), .Z(n13667) );
  XNOR U13857 ( .A(n13672), .B(n13676), .Z(n13665) );
  XOR U13858 ( .A(n13677), .B(n13675), .Z(n13676) );
  NAND U13859 ( .A(n13664), .B(n13668), .Z(n13675) );
  XNOR U13860 ( .A(n13660), .B(n13666), .Z(n13664) );
  XOR U13861 ( .A(n13678), .B(n13679), .Z(n13666) );
  XOR U13862 ( .A(n13680), .B(n13681), .Z(n13679) );
  XNOR U13863 ( .A(n13682), .B(n13683), .Z(n13678) );
  ANDN U13864 ( .B(n13684), .A(n13137), .Z(n13682) );
  AND U13865 ( .A(n13657), .B(n13660), .Z(n13677) );
  XNOR U13866 ( .A(n13657), .B(n13660), .Z(n13672) );
  XNOR U13867 ( .A(n13685), .B(n13686), .Z(n13660) );
  XNOR U13868 ( .A(n13687), .B(n13688), .Z(n13686) );
  XOR U13869 ( .A(n13680), .B(n13689), .Z(n13685) );
  XNOR U13870 ( .A(n13690), .B(n13683), .Z(n13689) );
  OR U13871 ( .A(n13217), .B(n13627), .Z(n13683) );
  XNOR U13872 ( .A(n13317), .B(n13626), .Z(n13627) );
  XNOR U13873 ( .A(n13137), .B(n13216), .Z(n13217) );
  NOR U13874 ( .A(n13216), .B(n13626), .Z(n13690) );
  XNOR U13875 ( .A(n13691), .B(n13692), .Z(n13657) );
  XNOR U13876 ( .A(n13693), .B(n13694), .Z(n13692) );
  XOR U13877 ( .A(n13645), .B(n13680), .Z(n13694) );
  XOR U13878 ( .A(n13684), .B(n13695), .Z(n13680) );
  XNOR U13879 ( .A(n13211), .B(n13696), .Z(n13691) );
  XNOR U13880 ( .A(n13697), .B(n13698), .Z(n13696) );
  ANDN U13881 ( .B(n13632), .A(n13699), .Z(n13697) );
  XNOR U13882 ( .A(n13700), .B(n13701), .Z(n13671) );
  XNOR U13883 ( .A(n13681), .B(n13702), .Z(n13701) );
  XNOR U13884 ( .A(n13632), .B(n13688), .Z(n13702) );
  XOR U13885 ( .A(n13626), .B(n13216), .Z(n13688) );
  XNOR U13886 ( .A(n13693), .B(n13703), .Z(n13681) );
  XNOR U13887 ( .A(n13704), .B(n13705), .Z(n13703) );
  NANDN U13888 ( .A(n13651), .B(n13323), .Z(n13705) );
  IV U13889 ( .A(n13687), .Z(n13693) );
  XNOR U13890 ( .A(n13706), .B(n13704), .Z(n13687) );
  NANDN U13891 ( .A(n13640), .B(n13653), .Z(n13704) );
  XOR U13892 ( .A(n13632), .B(n13216), .Z(n13651) );
  XOR U13893 ( .A(n13707), .B(n13708), .Z(n13216) );
  XNOR U13894 ( .A(n13709), .B(n13710), .Z(n13708) );
  XOR U13895 ( .A(n13642), .B(n13323), .Z(n13640) );
  XNOR U13896 ( .A(n13637), .B(n13626), .Z(n13323) );
  XNOR U13897 ( .A(n13710), .B(n13711), .Z(n13626) );
  ANDN U13898 ( .B(n13661), .A(n13642), .Z(n13706) );
  XNOR U13899 ( .A(n13712), .B(n13684), .Z(n13642) );
  IV U13900 ( .A(n13317), .Z(n13684) );
  XNOR U13901 ( .A(n13713), .B(n13714), .Z(n13317) );
  XNOR U13902 ( .A(n13715), .B(n13710), .Z(n13714) );
  XNOR U13903 ( .A(n13699), .B(n13716), .Z(n13700) );
  XNOR U13904 ( .A(n13717), .B(n13698), .Z(n13716) );
  OR U13905 ( .A(n13646), .B(n13636), .Z(n13698) );
  XOR U13906 ( .A(n13211), .B(n13637), .Z(n13636) );
  IV U13907 ( .A(n13699), .Z(n13637) );
  XOR U13908 ( .A(n13645), .B(n13632), .Z(n13646) );
  XNOR U13909 ( .A(n13695), .B(n13718), .Z(n13632) );
  XNOR U13910 ( .A(n13709), .B(n13713), .Z(n13718) );
  XNOR U13911 ( .A(state[122]), .B(key[122]), .Z(n13713) );
  IV U13912 ( .A(n13719), .Z(n13645) );
  ANDN U13913 ( .B(n13719), .A(n13211), .Z(n13717) );
  XOR U13914 ( .A(n13720), .B(n13721), .Z(n13699) );
  XOR U13915 ( .A(n13722), .B(n13723), .Z(n13721) );
  XOR U13916 ( .A(n13211), .B(n13715), .Z(n13720) );
  XNOR U13917 ( .A(n13709), .B(n13724), .Z(n13715) );
  XNOR U13918 ( .A(state[123]), .B(key[123]), .Z(n13724) );
  XNOR U13919 ( .A(state[121]), .B(key[121]), .Z(n13709) );
  IV U13920 ( .A(n13712), .Z(n13211) );
  XOR U13921 ( .A(n13719), .B(n13695), .Z(n13661) );
  IV U13922 ( .A(n13137), .Z(n13695) );
  XOR U13923 ( .A(n13707), .B(n13725), .Z(n13137) );
  XOR U13924 ( .A(n13710), .B(n13723), .Z(n13725) );
  XOR U13925 ( .A(state[127]), .B(key[127]), .Z(n13723) );
  XOR U13926 ( .A(n13711), .B(n13726), .Z(n13719) );
  XNOR U13927 ( .A(n13710), .B(n13722), .Z(n13726) );
  XNOR U13928 ( .A(state[124]), .B(key[124]), .Z(n13722) );
  XOR U13929 ( .A(n13712), .B(n13727), .Z(n13710) );
  XNOR U13930 ( .A(state[126]), .B(key[126]), .Z(n13727) );
  XOR U13931 ( .A(state[120]), .B(key[120]), .Z(n13712) );
  IV U13932 ( .A(n13707), .Z(n13711) );
  XOR U13933 ( .A(state[125]), .B(key[125]), .Z(n13707) );
  XOR U13934 ( .A(n7777), .B(n7775), .Z(n7760) );
  IV U13935 ( .A(n6089), .Z(n7775) );
  XOR U13936 ( .A(n13728), .B(n13729), .Z(n6089) );
  XNOR U13937 ( .A(n11386), .B(n11369), .Z(n13729) );
  XNOR U13938 ( .A(n13730), .B(n13731), .Z(n11369) );
  XNOR U13939 ( .A(n13732), .B(n13733), .Z(n13731) );
  NANDN U13940 ( .A(n13734), .B(n13735), .Z(n13733) );
  IV U13941 ( .A(n11407), .Z(n11386) );
  XOR U13942 ( .A(n13736), .B(n13737), .Z(n11407) );
  XOR U13943 ( .A(n13738), .B(n13739), .Z(n13737) );
  NANDN U13944 ( .A(n13740), .B(n11374), .Z(n13739) );
  XOR U13945 ( .A(n11388), .B(n11493), .Z(n13728) );
  XNOR U13946 ( .A(n11406), .B(n11389), .Z(n11493) );
  XOR U13947 ( .A(n11368), .B(n13741), .Z(n11389) );
  XNOR U13948 ( .A(n13742), .B(n13743), .Z(n13741) );
  NANDN U13949 ( .A(n13744), .B(n13745), .Z(n13743) );
  XNOR U13950 ( .A(n13742), .B(n13747), .Z(n13746) );
  NANDN U13951 ( .A(n13748), .B(n13735), .Z(n13747) );
  OR U13952 ( .A(n13749), .B(n13750), .Z(n13742) );
  XNOR U13953 ( .A(n11368), .B(n13751), .Z(n11494) );
  XNOR U13954 ( .A(n13752), .B(n13753), .Z(n13751) );
  NANDN U13955 ( .A(n13754), .B(n13755), .Z(n13753) );
  XOR U13956 ( .A(n13756), .B(n13752), .Z(n11368) );
  NANDN U13957 ( .A(n13757), .B(n13758), .Z(n13752) );
  ANDN U13958 ( .B(n13759), .A(n13760), .Z(n13756) );
  XOR U13959 ( .A(n11370), .B(n11406), .Z(n7777) );
  XNOR U13960 ( .A(n13736), .B(n13761), .Z(n11406) );
  XOR U13961 ( .A(n13762), .B(n13732), .Z(n13761) );
  OR U13962 ( .A(n13763), .B(n13749), .Z(n13732) );
  XNOR U13963 ( .A(n13735), .B(n13745), .Z(n13749) );
  ANDN U13964 ( .B(n13745), .A(n13764), .Z(n13762) );
  XNOR U13965 ( .A(n13730), .B(n13765), .Z(n11370) );
  XNOR U13966 ( .A(n13766), .B(n13738), .Z(n13765) );
  XOR U13967 ( .A(n13768), .B(n11374), .Z(n11497) );
  ANDN U13968 ( .B(n13769), .A(n11500), .Z(n13766) );
  IV U13969 ( .A(n13768), .Z(n11500) );
  XNOR U13970 ( .A(n13736), .B(n13770), .Z(n13730) );
  XNOR U13971 ( .A(n13771), .B(n13772), .Z(n13770) );
  NANDN U13972 ( .A(n13754), .B(n13773), .Z(n13772) );
  XOR U13973 ( .A(n13774), .B(n13771), .Z(n13736) );
  OR U13974 ( .A(n13757), .B(n13775), .Z(n13771) );
  XNOR U13975 ( .A(n13760), .B(n13754), .Z(n13757) );
  XNOR U13976 ( .A(n13745), .B(n11374), .Z(n13754) );
  XOR U13977 ( .A(n13776), .B(n13777), .Z(n11374) );
  NANDN U13978 ( .A(n13778), .B(n13779), .Z(n13777) );
  XOR U13979 ( .A(n13780), .B(n13781), .Z(n13745) );
  NANDN U13980 ( .A(n13778), .B(n13782), .Z(n13781) );
  NOR U13981 ( .A(n13760), .B(n13783), .Z(n13774) );
  XNOR U13982 ( .A(n13768), .B(n13735), .Z(n13760) );
  XNOR U13983 ( .A(n13784), .B(n13780), .Z(n13735) );
  NANDN U13984 ( .A(n13785), .B(n13786), .Z(n13780) );
  XOR U13985 ( .A(n13782), .B(n13787), .Z(n13786) );
  ANDN U13986 ( .B(n13787), .A(n13788), .Z(n13784) );
  XNOR U13987 ( .A(n13789), .B(n13776), .Z(n13768) );
  NANDN U13988 ( .A(n13785), .B(n13790), .Z(n13776) );
  XOR U13989 ( .A(n13791), .B(n13779), .Z(n13790) );
  XNOR U13990 ( .A(n13792), .B(n13793), .Z(n13778) );
  XOR U13991 ( .A(n13794), .B(n13795), .Z(n13793) );
  XNOR U13992 ( .A(n13796), .B(n13797), .Z(n13792) );
  XNOR U13993 ( .A(n13798), .B(n13799), .Z(n13797) );
  ANDN U13994 ( .B(n13791), .A(n13795), .Z(n13798) );
  ANDN U13995 ( .B(n13791), .A(n13788), .Z(n13789) );
  XNOR U13996 ( .A(n13794), .B(n13800), .Z(n13788) );
  XOR U13997 ( .A(n13801), .B(n13799), .Z(n13800) );
  NAND U13998 ( .A(n13802), .B(n13803), .Z(n13799) );
  XNOR U13999 ( .A(n13796), .B(n13779), .Z(n13803) );
  IV U14000 ( .A(n13791), .Z(n13796) );
  XNOR U14001 ( .A(n13782), .B(n13795), .Z(n13802) );
  IV U14002 ( .A(n13787), .Z(n13795) );
  XOR U14003 ( .A(n13804), .B(n13805), .Z(n13787) );
  XNOR U14004 ( .A(n13806), .B(n13807), .Z(n13805) );
  XNOR U14005 ( .A(n13808), .B(n13809), .Z(n13804) );
  ANDN U14006 ( .B(n13769), .A(n13810), .Z(n13808) );
  AND U14007 ( .A(n13779), .B(n13782), .Z(n13801) );
  XNOR U14008 ( .A(n13779), .B(n13782), .Z(n13794) );
  XNOR U14009 ( .A(n13811), .B(n13812), .Z(n13782) );
  XNOR U14010 ( .A(n13813), .B(n13807), .Z(n13812) );
  XOR U14011 ( .A(n13814), .B(n13815), .Z(n13811) );
  XNOR U14012 ( .A(n13816), .B(n13809), .Z(n13815) );
  OR U14013 ( .A(n11498), .B(n13767), .Z(n13809) );
  XNOR U14014 ( .A(n13769), .B(n13817), .Z(n13767) );
  XNOR U14015 ( .A(n13810), .B(n11375), .Z(n11498) );
  ANDN U14016 ( .B(n13818), .A(n13740), .Z(n13816) );
  XNOR U14017 ( .A(n13819), .B(n13820), .Z(n13779) );
  XNOR U14018 ( .A(n13807), .B(n13821), .Z(n13820) );
  XOR U14019 ( .A(n13748), .B(n13814), .Z(n13821) );
  XNOR U14020 ( .A(n13769), .B(n13810), .Z(n13807) );
  XOR U14021 ( .A(n13734), .B(n13822), .Z(n13819) );
  XNOR U14022 ( .A(n13823), .B(n13824), .Z(n13822) );
  ANDN U14023 ( .B(n13825), .A(n13764), .Z(n13823) );
  XNOR U14024 ( .A(n13826), .B(n13827), .Z(n13791) );
  XNOR U14025 ( .A(n13813), .B(n13828), .Z(n13827) );
  XNOR U14026 ( .A(n13744), .B(n13806), .Z(n13828) );
  XOR U14027 ( .A(n13814), .B(n13829), .Z(n13806) );
  XNOR U14028 ( .A(n13830), .B(n13831), .Z(n13829) );
  NAND U14029 ( .A(n13773), .B(n13755), .Z(n13831) );
  XNOR U14030 ( .A(n13832), .B(n13830), .Z(n13814) );
  NANDN U14031 ( .A(n13775), .B(n13758), .Z(n13830) );
  XOR U14032 ( .A(n13759), .B(n13755), .Z(n13758) );
  XNOR U14033 ( .A(n13825), .B(n11375), .Z(n13755) );
  XOR U14034 ( .A(n13783), .B(n13773), .Z(n13775) );
  XNOR U14035 ( .A(n13764), .B(n13817), .Z(n13773) );
  ANDN U14036 ( .B(n13759), .A(n13783), .Z(n13832) );
  XOR U14037 ( .A(n13734), .B(n13769), .Z(n13783) );
  XNOR U14038 ( .A(n13833), .B(n13834), .Z(n13769) );
  XNOR U14039 ( .A(n13835), .B(n13836), .Z(n13834) );
  XOR U14040 ( .A(n13817), .B(n13818), .Z(n13813) );
  IV U14041 ( .A(n11375), .Z(n13818) );
  XOR U14042 ( .A(n13837), .B(n13838), .Z(n11375) );
  XNOR U14043 ( .A(n13839), .B(n13836), .Z(n13838) );
  IV U14044 ( .A(n13740), .Z(n13817) );
  XOR U14045 ( .A(n13836), .B(n13840), .Z(n13740) );
  XNOR U14046 ( .A(n13841), .B(n13842), .Z(n13826) );
  XNOR U14047 ( .A(n13843), .B(n13824), .Z(n13842) );
  OR U14048 ( .A(n13750), .B(n13763), .Z(n13824) );
  XNOR U14049 ( .A(n13734), .B(n13764), .Z(n13763) );
  IV U14050 ( .A(n13841), .Z(n13764) );
  XOR U14051 ( .A(n13748), .B(n13825), .Z(n13750) );
  IV U14052 ( .A(n13744), .Z(n13825) );
  XOR U14053 ( .A(n11499), .B(n13844), .Z(n13744) );
  XNOR U14054 ( .A(n13839), .B(n13833), .Z(n13844) );
  XOR U14055 ( .A(n13845), .B(n13846), .Z(n13833) );
  XNOR U14056 ( .A(n10078), .B(n9000), .Z(n13846) );
  XOR U14057 ( .A(n8990), .B(n10838), .Z(n9000) );
  XOR U14058 ( .A(n9001), .B(n8985), .Z(n10078) );
  XOR U14059 ( .A(n13847), .B(n13848), .Z(n8985) );
  XNOR U14060 ( .A(n13849), .B(n13850), .Z(n13848) );
  XNOR U14061 ( .A(n13851), .B(n13852), .Z(n13847) );
  XOR U14062 ( .A(key[130]), .B(n8991), .Z(n13845) );
  IV U14063 ( .A(n13810), .Z(n11499) );
  XOR U14064 ( .A(n13837), .B(n13853), .Z(n13810) );
  XOR U14065 ( .A(n13836), .B(n13854), .Z(n13853) );
  NOR U14066 ( .A(n13748), .B(n13734), .Z(n13843) );
  XOR U14067 ( .A(n13837), .B(n13855), .Z(n13748) );
  XOR U14068 ( .A(n13836), .B(n13856), .Z(n13855) );
  XOR U14069 ( .A(n13857), .B(n13858), .Z(n13836) );
  XOR U14070 ( .A(n10857), .B(n8981), .Z(n13858) );
  XOR U14071 ( .A(n10106), .B(n13859), .Z(n8981) );
  XOR U14072 ( .A(n8965), .B(n10101), .Z(n10106) );
  IV U14073 ( .A(n10831), .Z(n10101) );
  XNOR U14074 ( .A(n13860), .B(n13861), .Z(n10831) );
  XNOR U14075 ( .A(n13862), .B(n13863), .Z(n8965) );
  XOR U14076 ( .A(n13864), .B(n8958), .Z(n10857) );
  XOR U14077 ( .A(n13865), .B(n13866), .Z(n8958) );
  XNOR U14078 ( .A(n13867), .B(n13868), .Z(n13866) );
  XNOR U14079 ( .A(n13869), .B(n13852), .Z(n13865) );
  XNOR U14080 ( .A(n8967), .B(n13870), .Z(n13857) );
  XOR U14081 ( .A(key[134]), .B(n13734), .Z(n13870) );
  IV U14082 ( .A(n13840), .Z(n13837) );
  XOR U14083 ( .A(n13871), .B(n13872), .Z(n13840) );
  XOR U14084 ( .A(n10850), .B(n8964), .Z(n13872) );
  XOR U14085 ( .A(n10812), .B(n10090), .Z(n8964) );
  XNOR U14086 ( .A(n13873), .B(n13874), .Z(n10090) );
  XNOR U14087 ( .A(n13875), .B(n13876), .Z(n13874) );
  XNOR U14088 ( .A(n13877), .B(n13878), .Z(n13873) );
  XNOR U14089 ( .A(n13879), .B(n13880), .Z(n13878) );
  ANDN U14090 ( .B(n13881), .A(n13882), .Z(n13880) );
  IV U14091 ( .A(n10104), .Z(n10812) );
  XOR U14092 ( .A(n13883), .B(n13884), .Z(n10104) );
  XNOR U14093 ( .A(n13885), .B(n13886), .Z(n13884) );
  XNOR U14094 ( .A(n13887), .B(n13888), .Z(n13883) );
  XNOR U14095 ( .A(n13889), .B(n13890), .Z(n13888) );
  ANDN U14096 ( .B(n13891), .A(n13892), .Z(n13890) );
  XOR U14097 ( .A(n8967), .B(n8979), .Z(n10850) );
  IV U14098 ( .A(n10829), .Z(n8979) );
  XOR U14099 ( .A(n13869), .B(n13850), .Z(n10829) );
  XNOR U14100 ( .A(n13893), .B(n13894), .Z(n13850) );
  XOR U14101 ( .A(n13895), .B(n13896), .Z(n13894) );
  NOR U14102 ( .A(n13897), .B(n13898), .Z(n13895) );
  XOR U14103 ( .A(n13899), .B(n13900), .Z(n8967) );
  XNOR U14104 ( .A(key[133]), .B(n10828), .Z(n13871) );
  XOR U14105 ( .A(n13901), .B(n13902), .Z(n13841) );
  XNOR U14106 ( .A(n13856), .B(n13854), .Z(n13902) );
  XNOR U14107 ( .A(n13903), .B(n13904), .Z(n13854) );
  XNOR U14108 ( .A(n13859), .B(n8959), .Z(n13904) );
  XNOR U14109 ( .A(n13905), .B(n13906), .Z(n10851) );
  XNOR U14110 ( .A(n13860), .B(n13886), .Z(n13906) );
  XNOR U14111 ( .A(n13907), .B(n13908), .Z(n13886) );
  XNOR U14112 ( .A(n13909), .B(n13910), .Z(n13908) );
  OR U14113 ( .A(n13911), .B(n13912), .Z(n13910) );
  XOR U14114 ( .A(n13913), .B(n13914), .Z(n13905) );
  XOR U14115 ( .A(n13915), .B(n13916), .Z(n10094) );
  XNOR U14116 ( .A(n13862), .B(n13876), .Z(n13916) );
  XNOR U14117 ( .A(n13917), .B(n13918), .Z(n13876) );
  XNOR U14118 ( .A(n13919), .B(n13920), .Z(n13918) );
  OR U14119 ( .A(n13921), .B(n13922), .Z(n13920) );
  XOR U14120 ( .A(n13923), .B(n10825), .Z(n13859) );
  XNOR U14121 ( .A(n13924), .B(n13925), .Z(n10825) );
  XOR U14122 ( .A(n13926), .B(n13927), .Z(n13925) );
  XNOR U14123 ( .A(n13899), .B(n13928), .Z(n13924) );
  XNOR U14124 ( .A(key[135]), .B(n10824), .Z(n13903) );
  XNOR U14125 ( .A(n13929), .B(n13930), .Z(n13856) );
  XOR U14126 ( .A(n8948), .B(n8946), .Z(n13930) );
  XOR U14127 ( .A(n10077), .B(n10091), .Z(n8946) );
  XOR U14128 ( .A(n13887), .B(n10838), .Z(n10091) );
  IV U14129 ( .A(n10062), .Z(n10838) );
  XNOR U14130 ( .A(n13931), .B(n13913), .Z(n10062) );
  XOR U14131 ( .A(n13877), .B(n8990), .Z(n10077) );
  XOR U14132 ( .A(n13932), .B(n13933), .Z(n8990) );
  XNOR U14133 ( .A(n13923), .B(n10828), .Z(n8948) );
  XOR U14134 ( .A(n13934), .B(n13935), .Z(n10828) );
  XNOR U14135 ( .A(n13936), .B(n13927), .Z(n13935) );
  XNOR U14136 ( .A(n13937), .B(n13938), .Z(n13927) );
  XNOR U14137 ( .A(n13939), .B(n13940), .Z(n13938) );
  OR U14138 ( .A(n13941), .B(n13942), .Z(n13940) );
  XNOR U14139 ( .A(n13943), .B(n13944), .Z(n13934) );
  XNOR U14140 ( .A(n13945), .B(n13946), .Z(n13944) );
  ANDN U14141 ( .B(n13947), .A(n13948), .Z(n13946) );
  IV U14142 ( .A(n10098), .Z(n13923) );
  XNOR U14143 ( .A(n10814), .B(n13949), .Z(n13929) );
  XNOR U14144 ( .A(key[132]), .B(n10811), .Z(n13949) );
  XOR U14145 ( .A(n13864), .B(n8963), .Z(n10814) );
  XOR U14146 ( .A(n13950), .B(n13951), .Z(n8963) );
  XNOR U14147 ( .A(n13952), .B(n13868), .Z(n13951) );
  XNOR U14148 ( .A(n13953), .B(n13954), .Z(n13868) );
  XNOR U14149 ( .A(n13955), .B(n13956), .Z(n13954) );
  OR U14150 ( .A(n13957), .B(n13958), .Z(n13956) );
  XNOR U14151 ( .A(n13959), .B(n13960), .Z(n13950) );
  XNOR U14152 ( .A(n13896), .B(n13961), .Z(n13960) );
  ANDN U14153 ( .B(n13962), .A(n13963), .Z(n13961) );
  NANDN U14154 ( .A(n13964), .B(n13965), .Z(n13896) );
  XNOR U14155 ( .A(n13734), .B(n13835), .Z(n13901) );
  XOR U14156 ( .A(n13966), .B(n13967), .Z(n13835) );
  XNOR U14157 ( .A(n8994), .B(n13968), .Z(n13967) );
  XNOR U14158 ( .A(n13839), .B(n8996), .Z(n13968) );
  IV U14159 ( .A(n10061), .Z(n8996) );
  XOR U14160 ( .A(n8999), .B(n10080), .Z(n10061) );
  XOR U14161 ( .A(n13969), .B(n13970), .Z(n10080) );
  XNOR U14162 ( .A(n13971), .B(n13861), .Z(n13970) );
  XNOR U14163 ( .A(n13972), .B(n13973), .Z(n13861) );
  XOR U14164 ( .A(n13974), .B(n13889), .Z(n13973) );
  NANDN U14165 ( .A(n13975), .B(n13976), .Z(n13889) );
  NOR U14166 ( .A(n13977), .B(n13978), .Z(n13974) );
  XNOR U14167 ( .A(n13913), .B(n13979), .Z(n13969) );
  XOR U14168 ( .A(n13915), .B(n13980), .Z(n8999) );
  XNOR U14169 ( .A(n13981), .B(n13863), .Z(n13980) );
  XNOR U14170 ( .A(n13982), .B(n13983), .Z(n13863) );
  XOR U14171 ( .A(n13984), .B(n13879), .Z(n13983) );
  NANDN U14172 ( .A(n13985), .B(n13986), .Z(n13879) );
  NOR U14173 ( .A(n13987), .B(n13988), .Z(n13984) );
  XNOR U14174 ( .A(n13989), .B(n13933), .Z(n13915) );
  XOR U14175 ( .A(n13990), .B(n13991), .Z(n13839) );
  XOR U14176 ( .A(n10847), .B(n10097), .Z(n13991) );
  IV U14177 ( .A(n8989), .Z(n10097) );
  XNOR U14178 ( .A(n13862), .B(n13992), .Z(n8974) );
  XOR U14179 ( .A(n13989), .B(n13933), .Z(n13992) );
  XOR U14180 ( .A(n13993), .B(n13994), .Z(n13933) );
  XOR U14181 ( .A(n13995), .B(n13996), .Z(n13994) );
  OR U14182 ( .A(n13997), .B(n13882), .Z(n13996) );
  XNOR U14183 ( .A(n13982), .B(n13998), .Z(n13989) );
  XNOR U14184 ( .A(n13999), .B(n14000), .Z(n13998) );
  OR U14185 ( .A(n13921), .B(n14001), .Z(n14000) );
  XNOR U14186 ( .A(n13875), .B(n14002), .Z(n13982) );
  XNOR U14187 ( .A(n14003), .B(n14004), .Z(n14002) );
  OR U14188 ( .A(n14005), .B(n14006), .Z(n14004) );
  XOR U14189 ( .A(n14007), .B(n13981), .Z(n13862) );
  XNOR U14190 ( .A(n13875), .B(n14008), .Z(n13981) );
  XNOR U14191 ( .A(n13999), .B(n14009), .Z(n14008) );
  NANDN U14192 ( .A(n14010), .B(n14011), .Z(n14009) );
  OR U14193 ( .A(n14012), .B(n14013), .Z(n13999) );
  XOR U14194 ( .A(n14014), .B(n14003), .Z(n13875) );
  NANDN U14195 ( .A(n14015), .B(n14016), .Z(n14003) );
  AND U14196 ( .A(n14017), .B(n14018), .Z(n14014) );
  XNOR U14197 ( .A(n13860), .B(n14019), .Z(n10074) );
  XOR U14198 ( .A(n13913), .B(n13979), .Z(n14019) );
  IV U14199 ( .A(n13914), .Z(n13979) );
  XOR U14200 ( .A(n13972), .B(n14020), .Z(n13914) );
  XNOR U14201 ( .A(n14021), .B(n14022), .Z(n14020) );
  OR U14202 ( .A(n13911), .B(n14023), .Z(n14022) );
  XNOR U14203 ( .A(n13885), .B(n14024), .Z(n13972) );
  XNOR U14204 ( .A(n14025), .B(n14026), .Z(n14024) );
  OR U14205 ( .A(n14027), .B(n14028), .Z(n14026) );
  XOR U14206 ( .A(n14029), .B(n14030), .Z(n13913) );
  XOR U14207 ( .A(n14031), .B(n14032), .Z(n14030) );
  OR U14208 ( .A(n14033), .B(n13892), .Z(n14032) );
  XNOR U14209 ( .A(n13931), .B(n13971), .Z(n13860) );
  XNOR U14210 ( .A(n13885), .B(n14034), .Z(n13971) );
  XNOR U14211 ( .A(n14021), .B(n14035), .Z(n14034) );
  NANDN U14212 ( .A(n14036), .B(n14037), .Z(n14035) );
  OR U14213 ( .A(n14038), .B(n14039), .Z(n14021) );
  XOR U14214 ( .A(n14040), .B(n14025), .Z(n13885) );
  NANDN U14215 ( .A(n14041), .B(n14042), .Z(n14025) );
  AND U14216 ( .A(n14043), .B(n14044), .Z(n14040) );
  IV U14217 ( .A(n10063), .Z(n10847) );
  XOR U14218 ( .A(n9003), .B(n8991), .Z(n10063) );
  XNOR U14219 ( .A(key[129]), .B(n14045), .Z(n13990) );
  XOR U14220 ( .A(n10098), .B(n10811), .Z(n8994) );
  XOR U14221 ( .A(n13943), .B(n8991), .Z(n10811) );
  XNOR U14222 ( .A(n14046), .B(n14047), .Z(n8991) );
  XNOR U14223 ( .A(n9001), .B(n14048), .Z(n13966) );
  XNOR U14224 ( .A(key[131]), .B(n10843), .Z(n14048) );
  XOR U14225 ( .A(n13864), .B(n8950), .Z(n10843) );
  XOR U14226 ( .A(n13952), .B(n9003), .Z(n8950) );
  IV U14227 ( .A(n10839), .Z(n9003) );
  XOR U14228 ( .A(n14049), .B(n13852), .Z(n10839) );
  IV U14229 ( .A(n10824), .Z(n13864) );
  XOR U14230 ( .A(n14050), .B(n13952), .Z(n10824) );
  XNOR U14231 ( .A(n13953), .B(n14051), .Z(n13952) );
  XOR U14232 ( .A(n14052), .B(n14053), .Z(n14051) );
  NOR U14233 ( .A(n14054), .B(n13898), .Z(n14052) );
  XNOR U14234 ( .A(n14055), .B(n14056), .Z(n13953) );
  XNOR U14235 ( .A(n14057), .B(n14058), .Z(n14056) );
  NANDN U14236 ( .A(n14059), .B(n14060), .Z(n14058) );
  XOR U14237 ( .A(n14061), .B(n14062), .Z(n9001) );
  XNOR U14238 ( .A(n14063), .B(n13900), .Z(n14062) );
  XNOR U14239 ( .A(n14064), .B(n14065), .Z(n13900) );
  XOR U14240 ( .A(n14066), .B(n13945), .Z(n14065) );
  NANDN U14241 ( .A(n14067), .B(n14068), .Z(n13945) );
  NOR U14242 ( .A(n14069), .B(n14070), .Z(n14066) );
  XOR U14243 ( .A(n14071), .B(n13928), .Z(n14061) );
  IV U14244 ( .A(n14047), .Z(n13928) );
  XNOR U14245 ( .A(n14072), .B(n14073), .Z(n13734) );
  XOR U14246 ( .A(n8960), .B(n10075), .Z(n14073) );
  IV U14247 ( .A(n10841), .Z(n10075) );
  XNOR U14248 ( .A(n8993), .B(n8976), .Z(n10841) );
  IV U14249 ( .A(n14045), .Z(n8976) );
  XOR U14250 ( .A(n13926), .B(n14074), .Z(n14045) );
  XNOR U14251 ( .A(n13899), .B(n14047), .Z(n14074) );
  XOR U14252 ( .A(n14075), .B(n14076), .Z(n14047) );
  XOR U14253 ( .A(n14077), .B(n14078), .Z(n14076) );
  OR U14254 ( .A(n14079), .B(n13948), .Z(n14078) );
  XOR U14255 ( .A(n14046), .B(n14071), .Z(n13899) );
  XNOR U14256 ( .A(n13936), .B(n14080), .Z(n14071) );
  XNOR U14257 ( .A(n14081), .B(n14082), .Z(n14080) );
  NANDN U14258 ( .A(n14083), .B(n14084), .Z(n14082) );
  IV U14259 ( .A(n14063), .Z(n13926) );
  XNOR U14260 ( .A(n14081), .B(n14086), .Z(n14085) );
  OR U14261 ( .A(n13941), .B(n14087), .Z(n14086) );
  OR U14262 ( .A(n14088), .B(n14089), .Z(n14081) );
  XNOR U14263 ( .A(n13936), .B(n14090), .Z(n14064) );
  XNOR U14264 ( .A(n14091), .B(n14092), .Z(n14090) );
  OR U14265 ( .A(n14093), .B(n14094), .Z(n14092) );
  XOR U14266 ( .A(n14095), .B(n14091), .Z(n13936) );
  NANDN U14267 ( .A(n14096), .B(n14097), .Z(n14091) );
  AND U14268 ( .A(n14098), .B(n14099), .Z(n14095) );
  IV U14269 ( .A(n10854), .Z(n8993) );
  XOR U14270 ( .A(n13849), .B(n14100), .Z(n10854) );
  XOR U14271 ( .A(n13869), .B(n13852), .Z(n14100) );
  XOR U14272 ( .A(n14055), .B(n14101), .Z(n13852) );
  XNOR U14273 ( .A(n14053), .B(n14102), .Z(n14101) );
  NANDN U14274 ( .A(n14103), .B(n13962), .Z(n14102) );
  NANDN U14275 ( .A(n14104), .B(n13965), .Z(n14053) );
  XNOR U14276 ( .A(n13898), .B(n13962), .Z(n13965) );
  XOR U14277 ( .A(n14050), .B(n13851), .Z(n13869) );
  XNOR U14278 ( .A(n13959), .B(n14105), .Z(n13851) );
  XNOR U14279 ( .A(n14106), .B(n14107), .Z(n14105) );
  NANDN U14280 ( .A(n14108), .B(n14109), .Z(n14107) );
  IV U14281 ( .A(n14049), .Z(n14050) );
  XNOR U14282 ( .A(n14055), .B(n14110), .Z(n14049) );
  XOR U14283 ( .A(n14111), .B(n13955), .Z(n14110) );
  OR U14284 ( .A(n14112), .B(n14113), .Z(n13955) );
  ANDN U14285 ( .B(n14114), .A(n14108), .Z(n14111) );
  XOR U14286 ( .A(n14115), .B(n14057), .Z(n14055) );
  OR U14287 ( .A(n14116), .B(n14117), .Z(n14057) );
  ANDN U14288 ( .B(n14118), .A(n14119), .Z(n14115) );
  IV U14289 ( .A(n13867), .Z(n13849) );
  XOR U14290 ( .A(n13893), .B(n14120), .Z(n13867) );
  XNOR U14291 ( .A(n14106), .B(n14121), .Z(n14120) );
  OR U14292 ( .A(n13957), .B(n14122), .Z(n14121) );
  OR U14293 ( .A(n14112), .B(n14123), .Z(n14106) );
  XOR U14294 ( .A(n13957), .B(n14124), .Z(n14112) );
  XOR U14295 ( .A(n13959), .B(n14125), .Z(n13893) );
  XNOR U14296 ( .A(n14126), .B(n14127), .Z(n14125) );
  OR U14297 ( .A(n14059), .B(n14128), .Z(n14127) );
  XOR U14298 ( .A(n14129), .B(n14126), .Z(n13959) );
  NANDN U14299 ( .A(n14116), .B(n14130), .Z(n14126) );
  XOR U14300 ( .A(n14118), .B(n14059), .Z(n14116) );
  XNOR U14301 ( .A(n14124), .B(n13962), .Z(n14059) );
  XOR U14302 ( .A(n14131), .B(n14132), .Z(n13962) );
  NANDN U14303 ( .A(n14133), .B(n14134), .Z(n14132) );
  IV U14304 ( .A(n14108), .Z(n14124) );
  XNOR U14305 ( .A(n14135), .B(n14136), .Z(n14108) );
  NANDN U14306 ( .A(n14133), .B(n14137), .Z(n14136) );
  XOR U14307 ( .A(n13898), .B(n13957), .Z(n14118) );
  XOR U14308 ( .A(n14139), .B(n14135), .Z(n13957) );
  NANDN U14309 ( .A(n14140), .B(n14141), .Z(n14135) );
  NANDN U14310 ( .A(n14140), .B(n14145), .Z(n14131) );
  XOR U14311 ( .A(n14146), .B(n14147), .Z(n14133) );
  XOR U14312 ( .A(n14148), .B(n14143), .Z(n14147) );
  XNOR U14313 ( .A(n14149), .B(n14150), .Z(n14146) );
  XNOR U14314 ( .A(n14151), .B(n14152), .Z(n14150) );
  ANDN U14315 ( .B(n14148), .A(n14143), .Z(n14151) );
  ANDN U14316 ( .B(n14148), .A(n14142), .Z(n14144) );
  XNOR U14317 ( .A(n14149), .B(n14153), .Z(n14142) );
  XOR U14318 ( .A(n14154), .B(n14152), .Z(n14153) );
  NAND U14319 ( .A(n14141), .B(n14145), .Z(n14152) );
  XNOR U14320 ( .A(n14137), .B(n14143), .Z(n14141) );
  XOR U14321 ( .A(n14155), .B(n14156), .Z(n14143) );
  XOR U14322 ( .A(n14157), .B(n14158), .Z(n14156) );
  XNOR U14323 ( .A(n14159), .B(n14160), .Z(n14155) );
  ANDN U14324 ( .B(n14161), .A(n13897), .Z(n14159) );
  AND U14325 ( .A(n14134), .B(n14137), .Z(n14154) );
  XNOR U14326 ( .A(n14134), .B(n14137), .Z(n14149) );
  XNOR U14327 ( .A(n14162), .B(n14163), .Z(n14137) );
  XNOR U14328 ( .A(n14164), .B(n14165), .Z(n14163) );
  XOR U14329 ( .A(n14157), .B(n14166), .Z(n14162) );
  XNOR U14330 ( .A(n14167), .B(n14160), .Z(n14166) );
  OR U14331 ( .A(n13964), .B(n14104), .Z(n14160) );
  XNOR U14332 ( .A(n14054), .B(n14103), .Z(n14104) );
  XNOR U14333 ( .A(n13897), .B(n13963), .Z(n13964) );
  NOR U14334 ( .A(n13963), .B(n14103), .Z(n14167) );
  XNOR U14335 ( .A(n14168), .B(n14169), .Z(n14134) );
  XNOR U14336 ( .A(n14170), .B(n14171), .Z(n14169) );
  XOR U14337 ( .A(n14122), .B(n14157), .Z(n14171) );
  XOR U14338 ( .A(n14161), .B(n14172), .Z(n14157) );
  XNOR U14339 ( .A(n13958), .B(n14173), .Z(n14168) );
  XNOR U14340 ( .A(n14174), .B(n14175), .Z(n14173) );
  ANDN U14341 ( .B(n14109), .A(n14176), .Z(n14174) );
  XNOR U14342 ( .A(n14177), .B(n14178), .Z(n14148) );
  XNOR U14343 ( .A(n14158), .B(n14179), .Z(n14178) );
  XNOR U14344 ( .A(n14109), .B(n14165), .Z(n14179) );
  XOR U14345 ( .A(n14103), .B(n13963), .Z(n14165) );
  XNOR U14346 ( .A(n14170), .B(n14180), .Z(n14158) );
  XNOR U14347 ( .A(n14181), .B(n14182), .Z(n14180) );
  NANDN U14348 ( .A(n14128), .B(n14060), .Z(n14182) );
  IV U14349 ( .A(n14164), .Z(n14170) );
  XNOR U14350 ( .A(n14183), .B(n14181), .Z(n14164) );
  NANDN U14351 ( .A(n14117), .B(n14130), .Z(n14181) );
  XOR U14352 ( .A(n14109), .B(n13963), .Z(n14128) );
  XOR U14353 ( .A(n14184), .B(n14185), .Z(n13963) );
  XNOR U14354 ( .A(n14186), .B(n14187), .Z(n14185) );
  XOR U14355 ( .A(n14119), .B(n14060), .Z(n14117) );
  XNOR U14356 ( .A(n14114), .B(n14103), .Z(n14060) );
  XNOR U14357 ( .A(n14187), .B(n14188), .Z(n14103) );
  ANDN U14358 ( .B(n14138), .A(n14119), .Z(n14183) );
  XNOR U14359 ( .A(n14189), .B(n14161), .Z(n14119) );
  IV U14360 ( .A(n14054), .Z(n14161) );
  XNOR U14361 ( .A(n14190), .B(n14191), .Z(n14054) );
  XNOR U14362 ( .A(n14192), .B(n14187), .Z(n14191) );
  XNOR U14363 ( .A(n14176), .B(n14193), .Z(n14177) );
  XNOR U14364 ( .A(n14194), .B(n14175), .Z(n14193) );
  OR U14365 ( .A(n14123), .B(n14113), .Z(n14175) );
  XOR U14366 ( .A(n13958), .B(n14114), .Z(n14113) );
  IV U14367 ( .A(n14176), .Z(n14114) );
  XOR U14368 ( .A(n14122), .B(n14109), .Z(n14123) );
  XNOR U14369 ( .A(n14172), .B(n14195), .Z(n14109) );
  XNOR U14370 ( .A(n14186), .B(n14190), .Z(n14195) );
  XNOR U14371 ( .A(state[34]), .B(key[34]), .Z(n14190) );
  IV U14372 ( .A(n14196), .Z(n14122) );
  ANDN U14373 ( .B(n14196), .A(n13958), .Z(n14194) );
  XOR U14374 ( .A(n14197), .B(n14198), .Z(n14176) );
  XOR U14375 ( .A(n14199), .B(n14200), .Z(n14198) );
  XOR U14376 ( .A(n13958), .B(n14192), .Z(n14197) );
  XNOR U14377 ( .A(n14186), .B(n14201), .Z(n14192) );
  XNOR U14378 ( .A(state[35]), .B(key[35]), .Z(n14201) );
  XNOR U14379 ( .A(state[33]), .B(key[33]), .Z(n14186) );
  IV U14380 ( .A(n14189), .Z(n13958) );
  XOR U14381 ( .A(n14196), .B(n14172), .Z(n14138) );
  IV U14382 ( .A(n13897), .Z(n14172) );
  XOR U14383 ( .A(n14184), .B(n14202), .Z(n13897) );
  XOR U14384 ( .A(n14187), .B(n14200), .Z(n14202) );
  XOR U14385 ( .A(state[39]), .B(key[39]), .Z(n14200) );
  XOR U14386 ( .A(n14188), .B(n14203), .Z(n14196) );
  XNOR U14387 ( .A(n14187), .B(n14199), .Z(n14203) );
  XNOR U14388 ( .A(state[36]), .B(key[36]), .Z(n14199) );
  XOR U14389 ( .A(n14189), .B(n14204), .Z(n14187) );
  XNOR U14390 ( .A(state[38]), .B(key[38]), .Z(n14204) );
  XOR U14391 ( .A(state[32]), .B(key[32]), .Z(n14189) );
  IV U14392 ( .A(n14184), .Z(n14188) );
  XOR U14393 ( .A(state[37]), .B(key[37]), .Z(n14184) );
  XNOR U14394 ( .A(n10076), .B(n10098), .Z(n8960) );
  XOR U14395 ( .A(n14046), .B(n13943), .Z(n10098) );
  XNOR U14396 ( .A(n13937), .B(n14205), .Z(n13943) );
  XNOR U14397 ( .A(n14206), .B(n14077), .Z(n14205) );
  ANDN U14398 ( .B(n14068), .A(n14207), .Z(n14077) );
  XOR U14399 ( .A(n14070), .B(n13948), .Z(n14068) );
  NOR U14400 ( .A(n14208), .B(n14070), .Z(n14206) );
  XNOR U14401 ( .A(n14075), .B(n14209), .Z(n13937) );
  XNOR U14402 ( .A(n14210), .B(n14211), .Z(n14209) );
  NANDN U14403 ( .A(n14093), .B(n14212), .Z(n14211) );
  XNOR U14404 ( .A(n14075), .B(n14213), .Z(n14046) );
  XOR U14405 ( .A(n14214), .B(n13939), .Z(n14213) );
  OR U14406 ( .A(n14215), .B(n14088), .Z(n13939) );
  XOR U14407 ( .A(n13941), .B(n14216), .Z(n14088) );
  ANDN U14408 ( .B(n14217), .A(n14083), .Z(n14214) );
  XOR U14409 ( .A(n14218), .B(n14210), .Z(n14075) );
  OR U14410 ( .A(n14096), .B(n14219), .Z(n14210) );
  XOR U14411 ( .A(n14098), .B(n14093), .Z(n14096) );
  XOR U14412 ( .A(n14216), .B(n13948), .Z(n14093) );
  XNOR U14413 ( .A(n14220), .B(n14221), .Z(n13948) );
  NANDN U14414 ( .A(n14222), .B(n14223), .Z(n14221) );
  IV U14415 ( .A(n14083), .Z(n14216) );
  XNOR U14416 ( .A(n14224), .B(n14225), .Z(n14083) );
  NANDN U14417 ( .A(n14222), .B(n14226), .Z(n14225) );
  ANDN U14418 ( .B(n14098), .A(n14227), .Z(n14218) );
  XOR U14419 ( .A(n14070), .B(n13941), .Z(n14098) );
  XOR U14420 ( .A(n14228), .B(n14224), .Z(n13941) );
  NANDN U14421 ( .A(n14229), .B(n14230), .Z(n14224) );
  NANDN U14422 ( .A(n14229), .B(n14234), .Z(n14220) );
  XOR U14423 ( .A(n14235), .B(n14236), .Z(n14222) );
  XOR U14424 ( .A(n14237), .B(n14232), .Z(n14236) );
  XNOR U14425 ( .A(n14238), .B(n14239), .Z(n14235) );
  XNOR U14426 ( .A(n14240), .B(n14241), .Z(n14239) );
  ANDN U14427 ( .B(n14237), .A(n14232), .Z(n14240) );
  ANDN U14428 ( .B(n14237), .A(n14231), .Z(n14233) );
  XNOR U14429 ( .A(n14238), .B(n14242), .Z(n14231) );
  XOR U14430 ( .A(n14243), .B(n14241), .Z(n14242) );
  NAND U14431 ( .A(n14230), .B(n14234), .Z(n14241) );
  XNOR U14432 ( .A(n14226), .B(n14232), .Z(n14230) );
  XOR U14433 ( .A(n14244), .B(n14245), .Z(n14232) );
  XOR U14434 ( .A(n14246), .B(n14247), .Z(n14245) );
  XNOR U14435 ( .A(n14248), .B(n14249), .Z(n14244) );
  ANDN U14436 ( .B(n14250), .A(n14069), .Z(n14248) );
  AND U14437 ( .A(n14223), .B(n14226), .Z(n14243) );
  XNOR U14438 ( .A(n14223), .B(n14226), .Z(n14238) );
  XNOR U14439 ( .A(n14251), .B(n14252), .Z(n14226) );
  XNOR U14440 ( .A(n14253), .B(n14254), .Z(n14252) );
  XOR U14441 ( .A(n14246), .B(n14255), .Z(n14251) );
  XNOR U14442 ( .A(n14256), .B(n14249), .Z(n14255) );
  OR U14443 ( .A(n14067), .B(n14207), .Z(n14249) );
  XNOR U14444 ( .A(n14208), .B(n14079), .Z(n14207) );
  XNOR U14445 ( .A(n14069), .B(n14257), .Z(n14067) );
  NOR U14446 ( .A(n14257), .B(n14079), .Z(n14256) );
  XNOR U14447 ( .A(n14258), .B(n14259), .Z(n14223) );
  XNOR U14448 ( .A(n14260), .B(n14261), .Z(n14259) );
  XOR U14449 ( .A(n14087), .B(n14246), .Z(n14261) );
  XOR U14450 ( .A(n14250), .B(n14262), .Z(n14246) );
  XNOR U14451 ( .A(n13942), .B(n14263), .Z(n14258) );
  XNOR U14452 ( .A(n14264), .B(n14265), .Z(n14263) );
  ANDN U14453 ( .B(n14084), .A(n14266), .Z(n14264) );
  XNOR U14454 ( .A(n14267), .B(n14268), .Z(n14237) );
  XNOR U14455 ( .A(n14247), .B(n14269), .Z(n14268) );
  XNOR U14456 ( .A(n14084), .B(n14254), .Z(n14269) );
  XOR U14457 ( .A(n14079), .B(n14257), .Z(n14254) );
  XNOR U14458 ( .A(n14260), .B(n14270), .Z(n14247) );
  XNOR U14459 ( .A(n14271), .B(n14272), .Z(n14270) );
  NANDN U14460 ( .A(n14094), .B(n14212), .Z(n14272) );
  IV U14461 ( .A(n14253), .Z(n14260) );
  XNOR U14462 ( .A(n14273), .B(n14271), .Z(n14253) );
  NANDN U14463 ( .A(n14219), .B(n14097), .Z(n14271) );
  XOR U14464 ( .A(n14084), .B(n14257), .Z(n14094) );
  IV U14465 ( .A(n13947), .Z(n14257) );
  XOR U14466 ( .A(n14274), .B(n14275), .Z(n13947) );
  XNOR U14467 ( .A(n14276), .B(n14277), .Z(n14275) );
  XOR U14468 ( .A(n14227), .B(n14212), .Z(n14219) );
  XNOR U14469 ( .A(n14217), .B(n14079), .Z(n14212) );
  XNOR U14470 ( .A(n14277), .B(n14274), .Z(n14079) );
  ANDN U14471 ( .B(n14099), .A(n14227), .Z(n14273) );
  XNOR U14472 ( .A(n14278), .B(n14250), .Z(n14227) );
  IV U14473 ( .A(n14208), .Z(n14250) );
  XNOR U14474 ( .A(n14279), .B(n14280), .Z(n14208) );
  XNOR U14475 ( .A(n14281), .B(n14277), .Z(n14280) );
  XOR U14476 ( .A(n14282), .B(n14262), .Z(n14099) );
  XNOR U14477 ( .A(n14266), .B(n14283), .Z(n14267) );
  XNOR U14478 ( .A(n14284), .B(n14265), .Z(n14283) );
  OR U14479 ( .A(n14089), .B(n14215), .Z(n14265) );
  XOR U14480 ( .A(n13942), .B(n14217), .Z(n14215) );
  IV U14481 ( .A(n14266), .Z(n14217) );
  XOR U14482 ( .A(n14087), .B(n14084), .Z(n14089) );
  XNOR U14483 ( .A(n14262), .B(n14285), .Z(n14084) );
  XNOR U14484 ( .A(n14276), .B(n14279), .Z(n14285) );
  XNOR U14485 ( .A(state[26]), .B(key[26]), .Z(n14279) );
  IV U14486 ( .A(n14069), .Z(n14262) );
  XOR U14487 ( .A(n14286), .B(n14287), .Z(n14069) );
  XOR U14488 ( .A(n14277), .B(n14288), .Z(n14287) );
  IV U14489 ( .A(n14282), .Z(n14087) );
  ANDN U14490 ( .B(n14282), .A(n13942), .Z(n14284) );
  XOR U14491 ( .A(n14274), .B(n14289), .Z(n14282) );
  XNOR U14492 ( .A(n14277), .B(n14290), .Z(n14289) );
  XOR U14493 ( .A(n14278), .B(n14291), .Z(n14277) );
  XNOR U14494 ( .A(state[30]), .B(key[30]), .Z(n14291) );
  IV U14495 ( .A(n14286), .Z(n14274) );
  XOR U14496 ( .A(state[29]), .B(key[29]), .Z(n14286) );
  XOR U14497 ( .A(n14292), .B(n14293), .Z(n14266) );
  XOR U14498 ( .A(n14290), .B(n14288), .Z(n14293) );
  XOR U14499 ( .A(state[31]), .B(key[31]), .Z(n14288) );
  XNOR U14500 ( .A(state[28]), .B(key[28]), .Z(n14290) );
  XOR U14501 ( .A(n13942), .B(n14281), .Z(n14292) );
  XNOR U14502 ( .A(n14276), .B(n14294), .Z(n14281) );
  XNOR U14503 ( .A(state[27]), .B(key[27]), .Z(n14294) );
  XNOR U14504 ( .A(state[25]), .B(key[25]), .Z(n14276) );
  IV U14505 ( .A(n14278), .Z(n13942) );
  XOR U14506 ( .A(state[24]), .B(key[24]), .Z(n14278) );
  IV U14507 ( .A(n8978), .Z(n10076) );
  XOR U14508 ( .A(n14007), .B(n13877), .Z(n8978) );
  XNOR U14509 ( .A(n13917), .B(n14295), .Z(n13877) );
  XNOR U14510 ( .A(n14296), .B(n13995), .Z(n14295) );
  ANDN U14511 ( .B(n13986), .A(n14297), .Z(n13995) );
  XOR U14512 ( .A(n13988), .B(n13882), .Z(n13986) );
  NOR U14513 ( .A(n14298), .B(n13988), .Z(n14296) );
  XNOR U14514 ( .A(n13993), .B(n14299), .Z(n13917) );
  XNOR U14515 ( .A(n14300), .B(n14301), .Z(n14299) );
  NANDN U14516 ( .A(n14005), .B(n14302), .Z(n14301) );
  IV U14517 ( .A(n13932), .Z(n14007) );
  XNOR U14518 ( .A(n13993), .B(n14303), .Z(n13932) );
  XOR U14519 ( .A(n14304), .B(n13919), .Z(n14303) );
  OR U14520 ( .A(n14305), .B(n14012), .Z(n13919) );
  XOR U14521 ( .A(n13921), .B(n14306), .Z(n14012) );
  ANDN U14522 ( .B(n14307), .A(n14010), .Z(n14304) );
  XOR U14523 ( .A(n14308), .B(n14300), .Z(n13993) );
  OR U14524 ( .A(n14015), .B(n14309), .Z(n14300) );
  XOR U14525 ( .A(n14017), .B(n14005), .Z(n14015) );
  XOR U14526 ( .A(n14306), .B(n13882), .Z(n14005) );
  XNOR U14527 ( .A(n14310), .B(n14311), .Z(n13882) );
  NANDN U14528 ( .A(n14312), .B(n14313), .Z(n14311) );
  IV U14529 ( .A(n14010), .Z(n14306) );
  XNOR U14530 ( .A(n14314), .B(n14315), .Z(n14010) );
  NANDN U14531 ( .A(n14312), .B(n14316), .Z(n14315) );
  ANDN U14532 ( .B(n14017), .A(n14317), .Z(n14308) );
  XOR U14533 ( .A(n13988), .B(n13921), .Z(n14017) );
  XOR U14534 ( .A(n14318), .B(n14314), .Z(n13921) );
  NANDN U14535 ( .A(n14319), .B(n14320), .Z(n14314) );
  NANDN U14536 ( .A(n14319), .B(n14324), .Z(n14310) );
  XOR U14537 ( .A(n14325), .B(n14326), .Z(n14312) );
  XOR U14538 ( .A(n14327), .B(n14322), .Z(n14326) );
  XNOR U14539 ( .A(n14328), .B(n14329), .Z(n14325) );
  XNOR U14540 ( .A(n14330), .B(n14331), .Z(n14329) );
  ANDN U14541 ( .B(n14327), .A(n14322), .Z(n14330) );
  ANDN U14542 ( .B(n14327), .A(n14321), .Z(n14323) );
  XNOR U14543 ( .A(n14328), .B(n14332), .Z(n14321) );
  XOR U14544 ( .A(n14333), .B(n14331), .Z(n14332) );
  NAND U14545 ( .A(n14320), .B(n14324), .Z(n14331) );
  XNOR U14546 ( .A(n14316), .B(n14322), .Z(n14320) );
  XOR U14547 ( .A(n14334), .B(n14335), .Z(n14322) );
  XOR U14548 ( .A(n14336), .B(n14337), .Z(n14335) );
  XNOR U14549 ( .A(n14338), .B(n14339), .Z(n14334) );
  ANDN U14550 ( .B(n14340), .A(n13987), .Z(n14338) );
  AND U14551 ( .A(n14313), .B(n14316), .Z(n14333) );
  XNOR U14552 ( .A(n14313), .B(n14316), .Z(n14328) );
  XNOR U14553 ( .A(n14341), .B(n14342), .Z(n14316) );
  XNOR U14554 ( .A(n14343), .B(n14344), .Z(n14342) );
  XOR U14555 ( .A(n14336), .B(n14345), .Z(n14341) );
  XNOR U14556 ( .A(n14346), .B(n14339), .Z(n14345) );
  OR U14557 ( .A(n13985), .B(n14297), .Z(n14339) );
  XNOR U14558 ( .A(n14298), .B(n13997), .Z(n14297) );
  XNOR U14559 ( .A(n13987), .B(n14347), .Z(n13985) );
  NOR U14560 ( .A(n14347), .B(n13997), .Z(n14346) );
  XNOR U14561 ( .A(n14348), .B(n14349), .Z(n14313) );
  XNOR U14562 ( .A(n14350), .B(n14351), .Z(n14349) );
  XOR U14563 ( .A(n14001), .B(n14336), .Z(n14351) );
  XOR U14564 ( .A(n14340), .B(n14352), .Z(n14336) );
  XNOR U14565 ( .A(n13922), .B(n14353), .Z(n14348) );
  XNOR U14566 ( .A(n14354), .B(n14355), .Z(n14353) );
  ANDN U14567 ( .B(n14011), .A(n14356), .Z(n14354) );
  XNOR U14568 ( .A(n14357), .B(n14358), .Z(n14327) );
  XNOR U14569 ( .A(n14337), .B(n14359), .Z(n14358) );
  XNOR U14570 ( .A(n14011), .B(n14344), .Z(n14359) );
  XOR U14571 ( .A(n13997), .B(n14347), .Z(n14344) );
  XNOR U14572 ( .A(n14350), .B(n14360), .Z(n14337) );
  XNOR U14573 ( .A(n14361), .B(n14362), .Z(n14360) );
  NANDN U14574 ( .A(n14006), .B(n14302), .Z(n14362) );
  IV U14575 ( .A(n14343), .Z(n14350) );
  XNOR U14576 ( .A(n14363), .B(n14361), .Z(n14343) );
  NANDN U14577 ( .A(n14309), .B(n14016), .Z(n14361) );
  XOR U14578 ( .A(n14011), .B(n14347), .Z(n14006) );
  IV U14579 ( .A(n13881), .Z(n14347) );
  XOR U14580 ( .A(n14364), .B(n14365), .Z(n13881) );
  XNOR U14581 ( .A(n14366), .B(n14367), .Z(n14365) );
  XOR U14582 ( .A(n14317), .B(n14302), .Z(n14309) );
  XNOR U14583 ( .A(n14307), .B(n13997), .Z(n14302) );
  XNOR U14584 ( .A(n14367), .B(n14364), .Z(n13997) );
  ANDN U14585 ( .B(n14018), .A(n14317), .Z(n14363) );
  XNOR U14586 ( .A(n14368), .B(n14340), .Z(n14317) );
  IV U14587 ( .A(n14298), .Z(n14340) );
  XNOR U14588 ( .A(n14369), .B(n14370), .Z(n14298) );
  XNOR U14589 ( .A(n14371), .B(n14367), .Z(n14370) );
  XOR U14590 ( .A(n14372), .B(n14352), .Z(n14018) );
  XNOR U14591 ( .A(n14356), .B(n14373), .Z(n14357) );
  XNOR U14592 ( .A(n14374), .B(n14355), .Z(n14373) );
  OR U14593 ( .A(n14013), .B(n14305), .Z(n14355) );
  XOR U14594 ( .A(n13922), .B(n14307), .Z(n14305) );
  IV U14595 ( .A(n14356), .Z(n14307) );
  XOR U14596 ( .A(n14001), .B(n14011), .Z(n14013) );
  XNOR U14597 ( .A(n14352), .B(n14375), .Z(n14011) );
  XNOR U14598 ( .A(n14366), .B(n14369), .Z(n14375) );
  XNOR U14599 ( .A(state[114]), .B(key[114]), .Z(n14369) );
  IV U14600 ( .A(n13987), .Z(n14352) );
  XOR U14601 ( .A(n14376), .B(n14377), .Z(n13987) );
  XOR U14602 ( .A(n14367), .B(n14378), .Z(n14377) );
  IV U14603 ( .A(n14372), .Z(n14001) );
  ANDN U14604 ( .B(n14372), .A(n13922), .Z(n14374) );
  XOR U14605 ( .A(n14364), .B(n14379), .Z(n14372) );
  XNOR U14606 ( .A(n14367), .B(n14380), .Z(n14379) );
  XOR U14607 ( .A(n14368), .B(n14381), .Z(n14367) );
  XNOR U14608 ( .A(state[118]), .B(key[118]), .Z(n14381) );
  IV U14609 ( .A(n14376), .Z(n14364) );
  XOR U14610 ( .A(state[117]), .B(key[117]), .Z(n14376) );
  XOR U14611 ( .A(n14382), .B(n14383), .Z(n14356) );
  XOR U14612 ( .A(n14380), .B(n14378), .Z(n14383) );
  XOR U14613 ( .A(state[119]), .B(key[119]), .Z(n14378) );
  XNOR U14614 ( .A(state[116]), .B(key[116]), .Z(n14380) );
  XOR U14615 ( .A(n13922), .B(n14371), .Z(n14382) );
  XNOR U14616 ( .A(n14366), .B(n14384), .Z(n14371) );
  XNOR U14617 ( .A(state[115]), .B(key[115]), .Z(n14384) );
  XNOR U14618 ( .A(state[113]), .B(key[113]), .Z(n14366) );
  IV U14619 ( .A(n14368), .Z(n13922) );
  XOR U14620 ( .A(state[112]), .B(key[112]), .Z(n14368) );
  XOR U14621 ( .A(n13887), .B(n13931), .Z(n10813) );
  XNOR U14622 ( .A(n14029), .B(n14385), .Z(n13931) );
  XOR U14623 ( .A(n14386), .B(n13909), .Z(n14385) );
  OR U14624 ( .A(n14387), .B(n14038), .Z(n13909) );
  XOR U14625 ( .A(n13911), .B(n14388), .Z(n14038) );
  ANDN U14626 ( .B(n14389), .A(n14036), .Z(n14386) );
  XNOR U14627 ( .A(n13907), .B(n14390), .Z(n13887) );
  XNOR U14628 ( .A(n14391), .B(n14031), .Z(n14390) );
  ANDN U14629 ( .B(n13976), .A(n14392), .Z(n14031) );
  XOR U14630 ( .A(n13978), .B(n13892), .Z(n13976) );
  NOR U14631 ( .A(n14393), .B(n13978), .Z(n14391) );
  XNOR U14632 ( .A(n14029), .B(n14394), .Z(n13907) );
  XNOR U14633 ( .A(n14395), .B(n14396), .Z(n14394) );
  NANDN U14634 ( .A(n14027), .B(n14397), .Z(n14396) );
  XOR U14635 ( .A(n14398), .B(n14395), .Z(n14029) );
  OR U14636 ( .A(n14041), .B(n14399), .Z(n14395) );
  XOR U14637 ( .A(n14043), .B(n14027), .Z(n14041) );
  XOR U14638 ( .A(n14388), .B(n13892), .Z(n14027) );
  XNOR U14639 ( .A(n14400), .B(n14401), .Z(n13892) );
  NANDN U14640 ( .A(n14402), .B(n14403), .Z(n14401) );
  IV U14641 ( .A(n14036), .Z(n14388) );
  XNOR U14642 ( .A(n14404), .B(n14405), .Z(n14036) );
  NANDN U14643 ( .A(n14402), .B(n14406), .Z(n14405) );
  ANDN U14644 ( .B(n14043), .A(n14407), .Z(n14398) );
  XOR U14645 ( .A(n13978), .B(n13911), .Z(n14043) );
  XOR U14646 ( .A(n14408), .B(n14404), .Z(n13911) );
  NANDN U14647 ( .A(n14409), .B(n14410), .Z(n14404) );
  NANDN U14648 ( .A(n14409), .B(n14414), .Z(n14400) );
  XOR U14649 ( .A(n14415), .B(n14416), .Z(n14402) );
  XOR U14650 ( .A(n14417), .B(n14412), .Z(n14416) );
  XNOR U14651 ( .A(n14418), .B(n14419), .Z(n14415) );
  XNOR U14652 ( .A(n14420), .B(n14421), .Z(n14419) );
  ANDN U14653 ( .B(n14417), .A(n14412), .Z(n14420) );
  ANDN U14654 ( .B(n14417), .A(n14411), .Z(n14413) );
  XNOR U14655 ( .A(n14418), .B(n14422), .Z(n14411) );
  XOR U14656 ( .A(n14423), .B(n14421), .Z(n14422) );
  NAND U14657 ( .A(n14410), .B(n14414), .Z(n14421) );
  XNOR U14658 ( .A(n14406), .B(n14412), .Z(n14410) );
  XOR U14659 ( .A(n14424), .B(n14425), .Z(n14412) );
  XOR U14660 ( .A(n14426), .B(n14427), .Z(n14425) );
  XNOR U14661 ( .A(n14428), .B(n14429), .Z(n14424) );
  ANDN U14662 ( .B(n14430), .A(n13977), .Z(n14428) );
  AND U14663 ( .A(n14403), .B(n14406), .Z(n14423) );
  XNOR U14664 ( .A(n14403), .B(n14406), .Z(n14418) );
  XNOR U14665 ( .A(n14431), .B(n14432), .Z(n14406) );
  XNOR U14666 ( .A(n14433), .B(n14434), .Z(n14432) );
  XOR U14667 ( .A(n14426), .B(n14435), .Z(n14431) );
  XNOR U14668 ( .A(n14436), .B(n14429), .Z(n14435) );
  OR U14669 ( .A(n13975), .B(n14392), .Z(n14429) );
  XNOR U14670 ( .A(n14393), .B(n14033), .Z(n14392) );
  XNOR U14671 ( .A(n13977), .B(n14437), .Z(n13975) );
  NOR U14672 ( .A(n14437), .B(n14033), .Z(n14436) );
  XNOR U14673 ( .A(n14438), .B(n14439), .Z(n14403) );
  XNOR U14674 ( .A(n14440), .B(n14441), .Z(n14439) );
  XOR U14675 ( .A(n14023), .B(n14426), .Z(n14441) );
  XOR U14676 ( .A(n14430), .B(n14442), .Z(n14426) );
  XNOR U14677 ( .A(n13912), .B(n14443), .Z(n14438) );
  XNOR U14678 ( .A(n14444), .B(n14445), .Z(n14443) );
  ANDN U14679 ( .B(n14037), .A(n14446), .Z(n14444) );
  XNOR U14680 ( .A(n14447), .B(n14448), .Z(n14417) );
  XNOR U14681 ( .A(n14427), .B(n14449), .Z(n14448) );
  XNOR U14682 ( .A(n14037), .B(n14434), .Z(n14449) );
  XOR U14683 ( .A(n14033), .B(n14437), .Z(n14434) );
  XNOR U14684 ( .A(n14440), .B(n14450), .Z(n14427) );
  XNOR U14685 ( .A(n14451), .B(n14452), .Z(n14450) );
  NANDN U14686 ( .A(n14028), .B(n14397), .Z(n14452) );
  IV U14687 ( .A(n14433), .Z(n14440) );
  XNOR U14688 ( .A(n14453), .B(n14451), .Z(n14433) );
  NANDN U14689 ( .A(n14399), .B(n14042), .Z(n14451) );
  XOR U14690 ( .A(n14037), .B(n14437), .Z(n14028) );
  IV U14691 ( .A(n13891), .Z(n14437) );
  XOR U14692 ( .A(n14454), .B(n14455), .Z(n13891) );
  XNOR U14693 ( .A(n14456), .B(n14457), .Z(n14455) );
  XOR U14694 ( .A(n14407), .B(n14397), .Z(n14399) );
  XNOR U14695 ( .A(n14389), .B(n14033), .Z(n14397) );
  XNOR U14696 ( .A(n14457), .B(n14454), .Z(n14033) );
  ANDN U14697 ( .B(n14044), .A(n14407), .Z(n14453) );
  XNOR U14698 ( .A(n14458), .B(n14430), .Z(n14407) );
  IV U14699 ( .A(n14393), .Z(n14430) );
  XNOR U14700 ( .A(n14459), .B(n14460), .Z(n14393) );
  XNOR U14701 ( .A(n14461), .B(n14457), .Z(n14460) );
  XOR U14702 ( .A(n14462), .B(n14442), .Z(n14044) );
  XNOR U14703 ( .A(n14446), .B(n14463), .Z(n14447) );
  XNOR U14704 ( .A(n14464), .B(n14445), .Z(n14463) );
  OR U14705 ( .A(n14039), .B(n14387), .Z(n14445) );
  XOR U14706 ( .A(n13912), .B(n14389), .Z(n14387) );
  IV U14707 ( .A(n14446), .Z(n14389) );
  XOR U14708 ( .A(n14023), .B(n14037), .Z(n14039) );
  XNOR U14709 ( .A(n14442), .B(n14465), .Z(n14037) );
  XNOR U14710 ( .A(n14456), .B(n14459), .Z(n14465) );
  XNOR U14711 ( .A(state[74]), .B(key[74]), .Z(n14459) );
  IV U14712 ( .A(n13977), .Z(n14442) );
  XOR U14713 ( .A(n14466), .B(n14467), .Z(n13977) );
  XOR U14714 ( .A(n14457), .B(n14468), .Z(n14467) );
  IV U14715 ( .A(n14462), .Z(n14023) );
  ANDN U14716 ( .B(n14462), .A(n13912), .Z(n14464) );
  XOR U14717 ( .A(n14454), .B(n14469), .Z(n14462) );
  XNOR U14718 ( .A(n14457), .B(n14470), .Z(n14469) );
  XOR U14719 ( .A(n14458), .B(n14471), .Z(n14457) );
  XNOR U14720 ( .A(state[78]), .B(key[78]), .Z(n14471) );
  IV U14721 ( .A(n14466), .Z(n14454) );
  XOR U14722 ( .A(state[77]), .B(key[77]), .Z(n14466) );
  XOR U14723 ( .A(n14472), .B(n14473), .Z(n14446) );
  XOR U14724 ( .A(n14470), .B(n14468), .Z(n14473) );
  XOR U14725 ( .A(state[79]), .B(key[79]), .Z(n14468) );
  XNOR U14726 ( .A(state[76]), .B(key[76]), .Z(n14470) );
  XOR U14727 ( .A(n13912), .B(n14461), .Z(n14472) );
  XNOR U14728 ( .A(n14456), .B(n14474), .Z(n14461) );
  XNOR U14729 ( .A(state[75]), .B(key[75]), .Z(n14474) );
  XNOR U14730 ( .A(state[73]), .B(key[73]), .Z(n14456) );
  IV U14731 ( .A(n14458), .Z(n13912) );
  XOR U14732 ( .A(state[72]), .B(key[72]), .Z(n14458) );
endmodule

