
module mult_N64_CC64 ( clk, rst, a, b, c );
  input [63:0] a;
  input [0:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317;
  wire   [127:0] sreg;

  DFF \sreg_reg[126]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(sreg[63]) );
  DFF \sreg_reg[62]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[1]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U4 ( .A(b[0]), .B(a[0]), .Z(n1) );
  XNOR U5 ( .A(n1), .B(sreg[63]), .Z(c[63]) );
  NAND U6 ( .A(b[0]), .B(a[1]), .Z(n2) );
  XOR U7 ( .A(sreg[64]), .B(n2), .Z(n4) );
  NANDN U8 ( .A(n1), .B(sreg[63]), .Z(n3) );
  XOR U9 ( .A(n4), .B(n3), .Z(c[64]) );
  NAND U10 ( .A(b[0]), .B(a[2]), .Z(n7) );
  XOR U11 ( .A(sreg[65]), .B(n7), .Z(n9) );
  NANDN U12 ( .A(n2), .B(sreg[64]), .Z(n6) );
  OR U13 ( .A(n4), .B(n3), .Z(n5) );
  AND U14 ( .A(n6), .B(n5), .Z(n8) );
  XOR U15 ( .A(n9), .B(n8), .Z(c[65]) );
  NAND U16 ( .A(b[0]), .B(a[3]), .Z(n12) );
  XOR U17 ( .A(sreg[66]), .B(n12), .Z(n14) );
  NANDN U18 ( .A(n7), .B(sreg[65]), .Z(n11) );
  OR U19 ( .A(n9), .B(n8), .Z(n10) );
  AND U20 ( .A(n11), .B(n10), .Z(n13) );
  XOR U21 ( .A(n14), .B(n13), .Z(c[66]) );
  NAND U22 ( .A(b[0]), .B(a[4]), .Z(n17) );
  XOR U23 ( .A(sreg[67]), .B(n17), .Z(n19) );
  NANDN U24 ( .A(n12), .B(sreg[66]), .Z(n16) );
  OR U25 ( .A(n14), .B(n13), .Z(n15) );
  AND U26 ( .A(n16), .B(n15), .Z(n18) );
  XOR U27 ( .A(n19), .B(n18), .Z(c[67]) );
  NAND U28 ( .A(b[0]), .B(a[5]), .Z(n22) );
  XOR U29 ( .A(sreg[68]), .B(n22), .Z(n24) );
  NANDN U30 ( .A(n17), .B(sreg[67]), .Z(n21) );
  OR U31 ( .A(n19), .B(n18), .Z(n20) );
  AND U32 ( .A(n21), .B(n20), .Z(n23) );
  XOR U33 ( .A(n24), .B(n23), .Z(c[68]) );
  NAND U34 ( .A(b[0]), .B(a[6]), .Z(n27) );
  XOR U35 ( .A(sreg[69]), .B(n27), .Z(n29) );
  NANDN U36 ( .A(n22), .B(sreg[68]), .Z(n26) );
  OR U37 ( .A(n24), .B(n23), .Z(n25) );
  AND U38 ( .A(n26), .B(n25), .Z(n28) );
  XOR U39 ( .A(n29), .B(n28), .Z(c[69]) );
  NAND U40 ( .A(b[0]), .B(a[7]), .Z(n32) );
  XOR U41 ( .A(sreg[70]), .B(n32), .Z(n34) );
  NANDN U42 ( .A(n27), .B(sreg[69]), .Z(n31) );
  OR U43 ( .A(n29), .B(n28), .Z(n30) );
  AND U44 ( .A(n31), .B(n30), .Z(n33) );
  XOR U45 ( .A(n34), .B(n33), .Z(c[70]) );
  NAND U46 ( .A(b[0]), .B(a[8]), .Z(n37) );
  XOR U47 ( .A(sreg[71]), .B(n37), .Z(n39) );
  NANDN U48 ( .A(n32), .B(sreg[70]), .Z(n36) );
  OR U49 ( .A(n34), .B(n33), .Z(n35) );
  AND U50 ( .A(n36), .B(n35), .Z(n38) );
  XOR U51 ( .A(n39), .B(n38), .Z(c[71]) );
  NAND U52 ( .A(b[0]), .B(a[9]), .Z(n42) );
  XOR U53 ( .A(sreg[72]), .B(n42), .Z(n44) );
  NANDN U54 ( .A(n37), .B(sreg[71]), .Z(n41) );
  OR U55 ( .A(n39), .B(n38), .Z(n40) );
  AND U56 ( .A(n41), .B(n40), .Z(n43) );
  XOR U57 ( .A(n44), .B(n43), .Z(c[72]) );
  NAND U58 ( .A(b[0]), .B(a[10]), .Z(n47) );
  XOR U59 ( .A(sreg[73]), .B(n47), .Z(n49) );
  NANDN U60 ( .A(n42), .B(sreg[72]), .Z(n46) );
  OR U61 ( .A(n44), .B(n43), .Z(n45) );
  AND U62 ( .A(n46), .B(n45), .Z(n48) );
  XOR U63 ( .A(n49), .B(n48), .Z(c[73]) );
  NAND U64 ( .A(b[0]), .B(a[11]), .Z(n52) );
  XOR U65 ( .A(sreg[74]), .B(n52), .Z(n54) );
  NANDN U66 ( .A(n47), .B(sreg[73]), .Z(n51) );
  OR U67 ( .A(n49), .B(n48), .Z(n50) );
  AND U68 ( .A(n51), .B(n50), .Z(n53) );
  XOR U69 ( .A(n54), .B(n53), .Z(c[74]) );
  NAND U70 ( .A(b[0]), .B(a[12]), .Z(n57) );
  XOR U71 ( .A(sreg[75]), .B(n57), .Z(n59) );
  NANDN U72 ( .A(n52), .B(sreg[74]), .Z(n56) );
  OR U73 ( .A(n54), .B(n53), .Z(n55) );
  AND U74 ( .A(n56), .B(n55), .Z(n58) );
  XOR U75 ( .A(n59), .B(n58), .Z(c[75]) );
  NAND U76 ( .A(b[0]), .B(a[13]), .Z(n62) );
  XOR U77 ( .A(sreg[76]), .B(n62), .Z(n64) );
  NANDN U78 ( .A(n57), .B(sreg[75]), .Z(n61) );
  OR U79 ( .A(n59), .B(n58), .Z(n60) );
  AND U80 ( .A(n61), .B(n60), .Z(n63) );
  XOR U81 ( .A(n64), .B(n63), .Z(c[76]) );
  NAND U82 ( .A(b[0]), .B(a[14]), .Z(n67) );
  XOR U83 ( .A(sreg[77]), .B(n67), .Z(n69) );
  NANDN U84 ( .A(n62), .B(sreg[76]), .Z(n66) );
  OR U85 ( .A(n64), .B(n63), .Z(n65) );
  AND U86 ( .A(n66), .B(n65), .Z(n68) );
  XOR U87 ( .A(n69), .B(n68), .Z(c[77]) );
  NAND U88 ( .A(b[0]), .B(a[15]), .Z(n72) );
  XOR U89 ( .A(sreg[78]), .B(n72), .Z(n74) );
  NANDN U90 ( .A(n67), .B(sreg[77]), .Z(n71) );
  OR U91 ( .A(n69), .B(n68), .Z(n70) );
  AND U92 ( .A(n71), .B(n70), .Z(n73) );
  XOR U93 ( .A(n74), .B(n73), .Z(c[78]) );
  NAND U94 ( .A(b[0]), .B(a[16]), .Z(n77) );
  XOR U95 ( .A(sreg[79]), .B(n77), .Z(n79) );
  NANDN U96 ( .A(n72), .B(sreg[78]), .Z(n76) );
  OR U97 ( .A(n74), .B(n73), .Z(n75) );
  AND U98 ( .A(n76), .B(n75), .Z(n78) );
  XOR U99 ( .A(n79), .B(n78), .Z(c[79]) );
  NAND U100 ( .A(b[0]), .B(a[17]), .Z(n82) );
  XOR U101 ( .A(sreg[80]), .B(n82), .Z(n84) );
  NANDN U102 ( .A(n77), .B(sreg[79]), .Z(n81) );
  OR U103 ( .A(n79), .B(n78), .Z(n80) );
  AND U104 ( .A(n81), .B(n80), .Z(n83) );
  XOR U105 ( .A(n84), .B(n83), .Z(c[80]) );
  NAND U106 ( .A(b[0]), .B(a[18]), .Z(n87) );
  XOR U107 ( .A(sreg[81]), .B(n87), .Z(n89) );
  NANDN U108 ( .A(n82), .B(sreg[80]), .Z(n86) );
  OR U109 ( .A(n84), .B(n83), .Z(n85) );
  AND U110 ( .A(n86), .B(n85), .Z(n88) );
  XOR U111 ( .A(n89), .B(n88), .Z(c[81]) );
  NAND U112 ( .A(b[0]), .B(a[19]), .Z(n92) );
  XOR U113 ( .A(sreg[82]), .B(n92), .Z(n94) );
  NANDN U114 ( .A(n87), .B(sreg[81]), .Z(n91) );
  OR U115 ( .A(n89), .B(n88), .Z(n90) );
  AND U116 ( .A(n91), .B(n90), .Z(n93) );
  XOR U117 ( .A(n94), .B(n93), .Z(c[82]) );
  NAND U118 ( .A(b[0]), .B(a[20]), .Z(n97) );
  XOR U119 ( .A(sreg[83]), .B(n97), .Z(n99) );
  NANDN U120 ( .A(n92), .B(sreg[82]), .Z(n96) );
  OR U121 ( .A(n94), .B(n93), .Z(n95) );
  AND U122 ( .A(n96), .B(n95), .Z(n98) );
  XOR U123 ( .A(n99), .B(n98), .Z(c[83]) );
  NAND U124 ( .A(b[0]), .B(a[21]), .Z(n102) );
  XOR U125 ( .A(sreg[84]), .B(n102), .Z(n104) );
  NANDN U126 ( .A(n97), .B(sreg[83]), .Z(n101) );
  OR U127 ( .A(n99), .B(n98), .Z(n100) );
  AND U128 ( .A(n101), .B(n100), .Z(n103) );
  XOR U129 ( .A(n104), .B(n103), .Z(c[84]) );
  NAND U130 ( .A(b[0]), .B(a[22]), .Z(n107) );
  XOR U131 ( .A(sreg[85]), .B(n107), .Z(n109) );
  NANDN U132 ( .A(n102), .B(sreg[84]), .Z(n106) );
  OR U133 ( .A(n104), .B(n103), .Z(n105) );
  AND U134 ( .A(n106), .B(n105), .Z(n108) );
  XOR U135 ( .A(n109), .B(n108), .Z(c[85]) );
  NAND U136 ( .A(b[0]), .B(a[23]), .Z(n112) );
  XOR U137 ( .A(sreg[86]), .B(n112), .Z(n114) );
  NANDN U138 ( .A(n107), .B(sreg[85]), .Z(n111) );
  OR U139 ( .A(n109), .B(n108), .Z(n110) );
  AND U140 ( .A(n111), .B(n110), .Z(n113) );
  XOR U141 ( .A(n114), .B(n113), .Z(c[86]) );
  NAND U142 ( .A(b[0]), .B(a[24]), .Z(n117) );
  XOR U143 ( .A(sreg[87]), .B(n117), .Z(n119) );
  NANDN U144 ( .A(n112), .B(sreg[86]), .Z(n116) );
  OR U145 ( .A(n114), .B(n113), .Z(n115) );
  AND U146 ( .A(n116), .B(n115), .Z(n118) );
  XOR U147 ( .A(n119), .B(n118), .Z(c[87]) );
  NAND U148 ( .A(b[0]), .B(a[25]), .Z(n122) );
  XOR U149 ( .A(sreg[88]), .B(n122), .Z(n124) );
  NANDN U150 ( .A(n117), .B(sreg[87]), .Z(n121) );
  OR U151 ( .A(n119), .B(n118), .Z(n120) );
  AND U152 ( .A(n121), .B(n120), .Z(n123) );
  XOR U153 ( .A(n124), .B(n123), .Z(c[88]) );
  NAND U154 ( .A(b[0]), .B(a[26]), .Z(n127) );
  XOR U155 ( .A(sreg[89]), .B(n127), .Z(n129) );
  NANDN U156 ( .A(n122), .B(sreg[88]), .Z(n126) );
  OR U157 ( .A(n124), .B(n123), .Z(n125) );
  AND U158 ( .A(n126), .B(n125), .Z(n128) );
  XOR U159 ( .A(n129), .B(n128), .Z(c[89]) );
  NAND U160 ( .A(b[0]), .B(a[27]), .Z(n132) );
  XOR U161 ( .A(sreg[90]), .B(n132), .Z(n134) );
  NANDN U162 ( .A(n127), .B(sreg[89]), .Z(n131) );
  OR U163 ( .A(n129), .B(n128), .Z(n130) );
  AND U164 ( .A(n131), .B(n130), .Z(n133) );
  XOR U165 ( .A(n134), .B(n133), .Z(c[90]) );
  NAND U166 ( .A(b[0]), .B(a[28]), .Z(n137) );
  XOR U167 ( .A(sreg[91]), .B(n137), .Z(n139) );
  NANDN U168 ( .A(n132), .B(sreg[90]), .Z(n136) );
  OR U169 ( .A(n134), .B(n133), .Z(n135) );
  AND U170 ( .A(n136), .B(n135), .Z(n138) );
  XOR U171 ( .A(n139), .B(n138), .Z(c[91]) );
  NAND U172 ( .A(b[0]), .B(a[29]), .Z(n142) );
  XOR U173 ( .A(sreg[92]), .B(n142), .Z(n144) );
  NANDN U174 ( .A(n137), .B(sreg[91]), .Z(n141) );
  OR U175 ( .A(n139), .B(n138), .Z(n140) );
  AND U176 ( .A(n141), .B(n140), .Z(n143) );
  XOR U177 ( .A(n144), .B(n143), .Z(c[92]) );
  NAND U178 ( .A(b[0]), .B(a[30]), .Z(n147) );
  XOR U179 ( .A(sreg[93]), .B(n147), .Z(n149) );
  NANDN U180 ( .A(n142), .B(sreg[92]), .Z(n146) );
  OR U181 ( .A(n144), .B(n143), .Z(n145) );
  AND U182 ( .A(n146), .B(n145), .Z(n148) );
  XOR U183 ( .A(n149), .B(n148), .Z(c[93]) );
  NAND U184 ( .A(b[0]), .B(a[31]), .Z(n152) );
  XOR U185 ( .A(sreg[94]), .B(n152), .Z(n154) );
  NANDN U186 ( .A(n147), .B(sreg[93]), .Z(n151) );
  OR U187 ( .A(n149), .B(n148), .Z(n150) );
  AND U188 ( .A(n151), .B(n150), .Z(n153) );
  XOR U189 ( .A(n154), .B(n153), .Z(c[94]) );
  NAND U190 ( .A(b[0]), .B(a[32]), .Z(n157) );
  XOR U191 ( .A(sreg[95]), .B(n157), .Z(n159) );
  NANDN U192 ( .A(n152), .B(sreg[94]), .Z(n156) );
  OR U193 ( .A(n154), .B(n153), .Z(n155) );
  AND U194 ( .A(n156), .B(n155), .Z(n158) );
  XOR U195 ( .A(n159), .B(n158), .Z(c[95]) );
  NAND U196 ( .A(b[0]), .B(a[33]), .Z(n162) );
  XOR U197 ( .A(sreg[96]), .B(n162), .Z(n164) );
  NANDN U198 ( .A(n157), .B(sreg[95]), .Z(n161) );
  OR U199 ( .A(n159), .B(n158), .Z(n160) );
  AND U200 ( .A(n161), .B(n160), .Z(n163) );
  XOR U201 ( .A(n164), .B(n163), .Z(c[96]) );
  NAND U202 ( .A(b[0]), .B(a[34]), .Z(n167) );
  XOR U203 ( .A(sreg[97]), .B(n167), .Z(n169) );
  NANDN U204 ( .A(n162), .B(sreg[96]), .Z(n166) );
  OR U205 ( .A(n164), .B(n163), .Z(n165) );
  AND U206 ( .A(n166), .B(n165), .Z(n168) );
  XOR U207 ( .A(n169), .B(n168), .Z(c[97]) );
  NAND U208 ( .A(b[0]), .B(a[35]), .Z(n172) );
  XOR U209 ( .A(sreg[98]), .B(n172), .Z(n174) );
  NANDN U210 ( .A(n167), .B(sreg[97]), .Z(n171) );
  OR U211 ( .A(n169), .B(n168), .Z(n170) );
  AND U212 ( .A(n171), .B(n170), .Z(n173) );
  XOR U213 ( .A(n174), .B(n173), .Z(c[98]) );
  NAND U214 ( .A(b[0]), .B(a[36]), .Z(n177) );
  XOR U215 ( .A(sreg[99]), .B(n177), .Z(n179) );
  NANDN U216 ( .A(n172), .B(sreg[98]), .Z(n176) );
  OR U217 ( .A(n174), .B(n173), .Z(n175) );
  AND U218 ( .A(n176), .B(n175), .Z(n178) );
  XOR U219 ( .A(n179), .B(n178), .Z(c[99]) );
  NAND U220 ( .A(b[0]), .B(a[37]), .Z(n182) );
  XOR U221 ( .A(sreg[100]), .B(n182), .Z(n184) );
  NANDN U222 ( .A(n177), .B(sreg[99]), .Z(n181) );
  OR U223 ( .A(n179), .B(n178), .Z(n180) );
  AND U224 ( .A(n181), .B(n180), .Z(n183) );
  XOR U225 ( .A(n184), .B(n183), .Z(c[100]) );
  NAND U226 ( .A(b[0]), .B(a[38]), .Z(n187) );
  XOR U227 ( .A(sreg[101]), .B(n187), .Z(n189) );
  NANDN U228 ( .A(n182), .B(sreg[100]), .Z(n186) );
  OR U229 ( .A(n184), .B(n183), .Z(n185) );
  AND U230 ( .A(n186), .B(n185), .Z(n188) );
  XOR U231 ( .A(n189), .B(n188), .Z(c[101]) );
  NAND U232 ( .A(b[0]), .B(a[39]), .Z(n192) );
  XOR U233 ( .A(sreg[102]), .B(n192), .Z(n194) );
  NANDN U234 ( .A(n187), .B(sreg[101]), .Z(n191) );
  OR U235 ( .A(n189), .B(n188), .Z(n190) );
  AND U236 ( .A(n191), .B(n190), .Z(n193) );
  XOR U237 ( .A(n194), .B(n193), .Z(c[102]) );
  NAND U238 ( .A(b[0]), .B(a[40]), .Z(n197) );
  XOR U239 ( .A(sreg[103]), .B(n197), .Z(n199) );
  NANDN U240 ( .A(n192), .B(sreg[102]), .Z(n196) );
  OR U241 ( .A(n194), .B(n193), .Z(n195) );
  AND U242 ( .A(n196), .B(n195), .Z(n198) );
  XOR U243 ( .A(n199), .B(n198), .Z(c[103]) );
  NAND U244 ( .A(b[0]), .B(a[41]), .Z(n202) );
  XOR U245 ( .A(sreg[104]), .B(n202), .Z(n204) );
  NANDN U246 ( .A(n197), .B(sreg[103]), .Z(n201) );
  OR U247 ( .A(n199), .B(n198), .Z(n200) );
  AND U248 ( .A(n201), .B(n200), .Z(n203) );
  XOR U249 ( .A(n204), .B(n203), .Z(c[104]) );
  NAND U250 ( .A(b[0]), .B(a[42]), .Z(n207) );
  XOR U251 ( .A(sreg[105]), .B(n207), .Z(n209) );
  NANDN U252 ( .A(n202), .B(sreg[104]), .Z(n206) );
  OR U253 ( .A(n204), .B(n203), .Z(n205) );
  AND U254 ( .A(n206), .B(n205), .Z(n208) );
  XOR U255 ( .A(n209), .B(n208), .Z(c[105]) );
  NAND U256 ( .A(b[0]), .B(a[43]), .Z(n212) );
  XOR U257 ( .A(sreg[106]), .B(n212), .Z(n214) );
  NANDN U258 ( .A(n207), .B(sreg[105]), .Z(n211) );
  OR U259 ( .A(n209), .B(n208), .Z(n210) );
  AND U260 ( .A(n211), .B(n210), .Z(n213) );
  XOR U261 ( .A(n214), .B(n213), .Z(c[106]) );
  NAND U262 ( .A(b[0]), .B(a[44]), .Z(n217) );
  XOR U263 ( .A(sreg[107]), .B(n217), .Z(n219) );
  NANDN U264 ( .A(n212), .B(sreg[106]), .Z(n216) );
  OR U265 ( .A(n214), .B(n213), .Z(n215) );
  AND U266 ( .A(n216), .B(n215), .Z(n218) );
  XOR U267 ( .A(n219), .B(n218), .Z(c[107]) );
  NAND U268 ( .A(b[0]), .B(a[45]), .Z(n222) );
  XOR U269 ( .A(sreg[108]), .B(n222), .Z(n224) );
  NANDN U270 ( .A(n217), .B(sreg[107]), .Z(n221) );
  OR U271 ( .A(n219), .B(n218), .Z(n220) );
  AND U272 ( .A(n221), .B(n220), .Z(n223) );
  XOR U273 ( .A(n224), .B(n223), .Z(c[108]) );
  NAND U274 ( .A(b[0]), .B(a[46]), .Z(n227) );
  XOR U275 ( .A(sreg[109]), .B(n227), .Z(n229) );
  NANDN U276 ( .A(n222), .B(sreg[108]), .Z(n226) );
  OR U277 ( .A(n224), .B(n223), .Z(n225) );
  AND U278 ( .A(n226), .B(n225), .Z(n228) );
  XOR U279 ( .A(n229), .B(n228), .Z(c[109]) );
  NAND U280 ( .A(b[0]), .B(a[47]), .Z(n232) );
  XOR U281 ( .A(sreg[110]), .B(n232), .Z(n234) );
  NANDN U282 ( .A(n227), .B(sreg[109]), .Z(n231) );
  OR U283 ( .A(n229), .B(n228), .Z(n230) );
  AND U284 ( .A(n231), .B(n230), .Z(n233) );
  XOR U285 ( .A(n234), .B(n233), .Z(c[110]) );
  NAND U286 ( .A(b[0]), .B(a[48]), .Z(n237) );
  XOR U287 ( .A(sreg[111]), .B(n237), .Z(n239) );
  NANDN U288 ( .A(n232), .B(sreg[110]), .Z(n236) );
  OR U289 ( .A(n234), .B(n233), .Z(n235) );
  AND U290 ( .A(n236), .B(n235), .Z(n238) );
  XOR U291 ( .A(n239), .B(n238), .Z(c[111]) );
  NAND U292 ( .A(b[0]), .B(a[49]), .Z(n242) );
  XOR U293 ( .A(sreg[112]), .B(n242), .Z(n244) );
  NANDN U294 ( .A(n237), .B(sreg[111]), .Z(n241) );
  OR U295 ( .A(n239), .B(n238), .Z(n240) );
  AND U296 ( .A(n241), .B(n240), .Z(n243) );
  XOR U297 ( .A(n244), .B(n243), .Z(c[112]) );
  NAND U298 ( .A(b[0]), .B(a[50]), .Z(n247) );
  XOR U299 ( .A(sreg[113]), .B(n247), .Z(n249) );
  NANDN U300 ( .A(n242), .B(sreg[112]), .Z(n246) );
  OR U301 ( .A(n244), .B(n243), .Z(n245) );
  AND U302 ( .A(n246), .B(n245), .Z(n248) );
  XOR U303 ( .A(n249), .B(n248), .Z(c[113]) );
  NAND U304 ( .A(b[0]), .B(a[51]), .Z(n252) );
  XOR U305 ( .A(sreg[114]), .B(n252), .Z(n254) );
  NANDN U306 ( .A(n247), .B(sreg[113]), .Z(n251) );
  OR U307 ( .A(n249), .B(n248), .Z(n250) );
  AND U308 ( .A(n251), .B(n250), .Z(n253) );
  XOR U309 ( .A(n254), .B(n253), .Z(c[114]) );
  NAND U310 ( .A(b[0]), .B(a[52]), .Z(n257) );
  XOR U311 ( .A(sreg[115]), .B(n257), .Z(n259) );
  NANDN U312 ( .A(n252), .B(sreg[114]), .Z(n256) );
  OR U313 ( .A(n254), .B(n253), .Z(n255) );
  AND U314 ( .A(n256), .B(n255), .Z(n258) );
  XOR U315 ( .A(n259), .B(n258), .Z(c[115]) );
  NAND U316 ( .A(b[0]), .B(a[53]), .Z(n262) );
  XOR U317 ( .A(sreg[116]), .B(n262), .Z(n264) );
  NANDN U318 ( .A(n257), .B(sreg[115]), .Z(n261) );
  OR U319 ( .A(n259), .B(n258), .Z(n260) );
  AND U320 ( .A(n261), .B(n260), .Z(n263) );
  XOR U321 ( .A(n264), .B(n263), .Z(c[116]) );
  NAND U322 ( .A(b[0]), .B(a[54]), .Z(n267) );
  XOR U323 ( .A(sreg[117]), .B(n267), .Z(n269) );
  NANDN U324 ( .A(n262), .B(sreg[116]), .Z(n266) );
  OR U325 ( .A(n264), .B(n263), .Z(n265) );
  AND U326 ( .A(n266), .B(n265), .Z(n268) );
  XOR U327 ( .A(n269), .B(n268), .Z(c[117]) );
  NAND U328 ( .A(b[0]), .B(a[55]), .Z(n272) );
  XOR U329 ( .A(sreg[118]), .B(n272), .Z(n274) );
  NANDN U330 ( .A(n267), .B(sreg[117]), .Z(n271) );
  OR U331 ( .A(n269), .B(n268), .Z(n270) );
  AND U332 ( .A(n271), .B(n270), .Z(n273) );
  XOR U333 ( .A(n274), .B(n273), .Z(c[118]) );
  NAND U334 ( .A(b[0]), .B(a[56]), .Z(n277) );
  XOR U335 ( .A(sreg[119]), .B(n277), .Z(n279) );
  NANDN U336 ( .A(n272), .B(sreg[118]), .Z(n276) );
  OR U337 ( .A(n274), .B(n273), .Z(n275) );
  AND U338 ( .A(n276), .B(n275), .Z(n278) );
  XOR U339 ( .A(n279), .B(n278), .Z(c[119]) );
  NAND U340 ( .A(b[0]), .B(a[57]), .Z(n282) );
  XOR U341 ( .A(sreg[120]), .B(n282), .Z(n284) );
  NANDN U342 ( .A(n277), .B(sreg[119]), .Z(n281) );
  OR U343 ( .A(n279), .B(n278), .Z(n280) );
  AND U344 ( .A(n281), .B(n280), .Z(n283) );
  XOR U345 ( .A(n284), .B(n283), .Z(c[120]) );
  NAND U346 ( .A(b[0]), .B(a[58]), .Z(n287) );
  XOR U347 ( .A(sreg[121]), .B(n287), .Z(n289) );
  NANDN U348 ( .A(n282), .B(sreg[120]), .Z(n286) );
  OR U349 ( .A(n284), .B(n283), .Z(n285) );
  AND U350 ( .A(n286), .B(n285), .Z(n288) );
  XOR U351 ( .A(n289), .B(n288), .Z(c[121]) );
  NAND U352 ( .A(b[0]), .B(a[59]), .Z(n292) );
  XOR U353 ( .A(sreg[122]), .B(n292), .Z(n294) );
  NANDN U354 ( .A(n287), .B(sreg[121]), .Z(n291) );
  OR U355 ( .A(n289), .B(n288), .Z(n290) );
  AND U356 ( .A(n291), .B(n290), .Z(n293) );
  XOR U357 ( .A(n294), .B(n293), .Z(c[122]) );
  NAND U358 ( .A(b[0]), .B(a[60]), .Z(n297) );
  XOR U359 ( .A(sreg[123]), .B(n297), .Z(n299) );
  NANDN U360 ( .A(n292), .B(sreg[122]), .Z(n296) );
  OR U361 ( .A(n294), .B(n293), .Z(n295) );
  AND U362 ( .A(n296), .B(n295), .Z(n298) );
  XOR U363 ( .A(n299), .B(n298), .Z(c[123]) );
  NAND U364 ( .A(b[0]), .B(a[61]), .Z(n302) );
  XOR U365 ( .A(sreg[124]), .B(n302), .Z(n304) );
  NANDN U366 ( .A(n297), .B(sreg[123]), .Z(n301) );
  OR U367 ( .A(n299), .B(n298), .Z(n300) );
  AND U368 ( .A(n301), .B(n300), .Z(n303) );
  XOR U369 ( .A(n304), .B(n303), .Z(c[124]) );
  NAND U370 ( .A(b[0]), .B(a[62]), .Z(n307) );
  XOR U371 ( .A(sreg[125]), .B(n307), .Z(n309) );
  NANDN U372 ( .A(n302), .B(sreg[124]), .Z(n306) );
  OR U373 ( .A(n304), .B(n303), .Z(n305) );
  AND U374 ( .A(n306), .B(n305), .Z(n308) );
  XOR U375 ( .A(n309), .B(n308), .Z(c[125]) );
  NANDN U376 ( .A(n307), .B(sreg[125]), .Z(n311) );
  OR U377 ( .A(n309), .B(n308), .Z(n310) );
  AND U378 ( .A(n311), .B(n310), .Z(n315) );
  AND U379 ( .A(a[63]), .B(b[0]), .Z(n313) );
  XNOR U380 ( .A(sreg[126]), .B(n313), .Z(n312) );
  XOR U381 ( .A(n315), .B(n312), .Z(c[126]) );
  NAND U382 ( .A(sreg[126]), .B(n313), .Z(n317) );
  XOR U383 ( .A(n313), .B(sreg[126]), .Z(n314) );
  NANDN U384 ( .A(n315), .B(n314), .Z(n316) );
  NAND U385 ( .A(n317), .B(n316), .Z(c[127]) );
endmodule

