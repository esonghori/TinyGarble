
module sum_N256_CC1 ( clk, rst, a, b, c );
  input [255:0] a;
  input [255:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274;

  XOR U2 ( .A(a[24]), .B(b[24]), .Z(n2) );
  NANDN U3 ( .A(n1096), .B(n2), .Z(n3) );
  NAND U4 ( .A(a[24]), .B(b[24]), .Z(n4) );
  AND U5 ( .A(n3), .B(n4), .Z(n763) );
  XOR U6 ( .A(a[3]), .B(b[3]), .Z(n5) );
  NANDN U7 ( .A(n1141), .B(n5), .Z(n6) );
  NAND U8 ( .A(a[3]), .B(b[3]), .Z(n7) );
  AND U9 ( .A(n6), .B(n7), .Z(n1163) );
  XOR U10 ( .A(a[6]), .B(b[6]), .Z(n8) );
  NANDN U11 ( .A(n1207), .B(n8), .Z(n9) );
  NAND U12 ( .A(a[6]), .B(b[6]), .Z(n10) );
  AND U13 ( .A(n9), .B(n10), .Z(n1229) );
  XOR U14 ( .A(b[9]), .B(a[9]), .Z(n11) );
  NANDN U15 ( .A(n1273), .B(n11), .Z(n12) );
  NAND U16 ( .A(b[9]), .B(a[9]), .Z(n13) );
  AND U17 ( .A(n12), .B(n13), .Z(n786) );
  XOR U18 ( .A(a[12]), .B(b[12]), .Z(n14) );
  NANDN U19 ( .A(n830), .B(n14), .Z(n15) );
  NAND U20 ( .A(a[12]), .B(b[12]), .Z(n16) );
  AND U21 ( .A(n15), .B(n16), .Z(n852) );
  XOR U22 ( .A(a[15]), .B(b[15]), .Z(n17) );
  NANDN U23 ( .A(n896), .B(n17), .Z(n18) );
  NAND U24 ( .A(a[15]), .B(b[15]), .Z(n19) );
  AND U25 ( .A(n18), .B(n19), .Z(n918) );
  XOR U26 ( .A(a[18]), .B(b[18]), .Z(n20) );
  NANDN U27 ( .A(n962), .B(n20), .Z(n21) );
  NAND U28 ( .A(a[18]), .B(b[18]), .Z(n22) );
  AND U29 ( .A(n21), .B(n22), .Z(n984) );
  XOR U30 ( .A(a[21]), .B(b[21]), .Z(n23) );
  NANDN U31 ( .A(n1030), .B(n23), .Z(n24) );
  NAND U32 ( .A(a[21]), .B(b[21]), .Z(n25) );
  AND U33 ( .A(n24), .B(n25), .Z(n1052) );
  XOR U34 ( .A(a[27]), .B(b[27]), .Z(n26) );
  NANDN U35 ( .A(n1113), .B(n26), .Z(n27) );
  NAND U36 ( .A(a[27]), .B(b[27]), .Z(n28) );
  AND U37 ( .A(n27), .B(n28), .Z(n1115) );
  XOR U38 ( .A(a[30]), .B(b[30]), .Z(n29) );
  NANDN U39 ( .A(n1121), .B(n29), .Z(n30) );
  NAND U40 ( .A(a[30]), .B(b[30]), .Z(n31) );
  AND U41 ( .A(n30), .B(n31), .Z(n1123) );
  XOR U42 ( .A(a[33]), .B(b[33]), .Z(n32) );
  NANDN U43 ( .A(n1127), .B(n32), .Z(n33) );
  NAND U44 ( .A(a[33]), .B(b[33]), .Z(n34) );
  AND U45 ( .A(n33), .B(n34), .Z(n1129) );
  XOR U46 ( .A(a[36]), .B(b[36]), .Z(n35) );
  NANDN U47 ( .A(n1133), .B(n35), .Z(n36) );
  NAND U48 ( .A(a[36]), .B(b[36]), .Z(n37) );
  AND U49 ( .A(n36), .B(n37), .Z(n1135) );
  XOR U50 ( .A(a[39]), .B(b[39]), .Z(n38) );
  NANDN U51 ( .A(n1139), .B(n38), .Z(n39) );
  NAND U52 ( .A(a[39]), .B(b[39]), .Z(n40) );
  AND U53 ( .A(n39), .B(n40), .Z(n1143) );
  XOR U54 ( .A(a[42]), .B(b[42]), .Z(n41) );
  NANDN U55 ( .A(n1147), .B(n41), .Z(n42) );
  NAND U56 ( .A(a[42]), .B(b[42]), .Z(n43) );
  AND U57 ( .A(n42), .B(n43), .Z(n1149) );
  XOR U58 ( .A(a[45]), .B(b[45]), .Z(n44) );
  NANDN U59 ( .A(n1153), .B(n44), .Z(n45) );
  NAND U60 ( .A(a[45]), .B(b[45]), .Z(n46) );
  AND U61 ( .A(n45), .B(n46), .Z(n1155) );
  XOR U62 ( .A(a[48]), .B(b[48]), .Z(n47) );
  NANDN U63 ( .A(n1159), .B(n47), .Z(n48) );
  NAND U64 ( .A(a[48]), .B(b[48]), .Z(n49) );
  AND U65 ( .A(n48), .B(n49), .Z(n1161) );
  XOR U66 ( .A(a[51]), .B(b[51]), .Z(n50) );
  NANDN U67 ( .A(n1167), .B(n50), .Z(n51) );
  NAND U68 ( .A(a[51]), .B(b[51]), .Z(n52) );
  AND U69 ( .A(n51), .B(n52), .Z(n1169) );
  XOR U70 ( .A(a[54]), .B(b[54]), .Z(n53) );
  NANDN U71 ( .A(n1173), .B(n53), .Z(n54) );
  NAND U72 ( .A(a[54]), .B(b[54]), .Z(n55) );
  AND U73 ( .A(n54), .B(n55), .Z(n1175) );
  XOR U74 ( .A(a[57]), .B(b[57]), .Z(n56) );
  NANDN U75 ( .A(n1179), .B(n56), .Z(n57) );
  NAND U76 ( .A(a[57]), .B(b[57]), .Z(n58) );
  AND U77 ( .A(n57), .B(n58), .Z(n1181) );
  XOR U78 ( .A(a[60]), .B(b[60]), .Z(n59) );
  NANDN U79 ( .A(n1187), .B(n59), .Z(n60) );
  NAND U80 ( .A(a[60]), .B(b[60]), .Z(n61) );
  AND U81 ( .A(n60), .B(n61), .Z(n1189) );
  XOR U82 ( .A(a[63]), .B(b[63]), .Z(n62) );
  NANDN U83 ( .A(n1193), .B(n62), .Z(n63) );
  NAND U84 ( .A(a[63]), .B(b[63]), .Z(n64) );
  AND U85 ( .A(n63), .B(n64), .Z(n1195) );
  XOR U86 ( .A(a[66]), .B(b[66]), .Z(n65) );
  NANDN U87 ( .A(n1199), .B(n65), .Z(n66) );
  NAND U88 ( .A(a[66]), .B(b[66]), .Z(n67) );
  AND U89 ( .A(n66), .B(n67), .Z(n1201) );
  XOR U90 ( .A(a[69]), .B(b[69]), .Z(n68) );
  NANDN U91 ( .A(n1205), .B(n68), .Z(n69) );
  NAND U92 ( .A(a[69]), .B(b[69]), .Z(n70) );
  AND U93 ( .A(n69), .B(n70), .Z(n1209) );
  XOR U94 ( .A(a[72]), .B(b[72]), .Z(n71) );
  NANDN U95 ( .A(n1213), .B(n71), .Z(n72) );
  NAND U96 ( .A(a[72]), .B(b[72]), .Z(n73) );
  AND U97 ( .A(n72), .B(n73), .Z(n1215) );
  XOR U98 ( .A(a[75]), .B(b[75]), .Z(n74) );
  NANDN U99 ( .A(n1219), .B(n74), .Z(n75) );
  NAND U100 ( .A(a[75]), .B(b[75]), .Z(n76) );
  AND U101 ( .A(n75), .B(n76), .Z(n1221) );
  XOR U102 ( .A(a[78]), .B(b[78]), .Z(n77) );
  NANDN U103 ( .A(n1225), .B(n77), .Z(n78) );
  NAND U104 ( .A(a[78]), .B(b[78]), .Z(n79) );
  AND U105 ( .A(n78), .B(n79), .Z(n1227) );
  XOR U106 ( .A(a[81]), .B(b[81]), .Z(n80) );
  NANDN U107 ( .A(n1233), .B(n80), .Z(n81) );
  NAND U108 ( .A(a[81]), .B(b[81]), .Z(n82) );
  AND U109 ( .A(n81), .B(n82), .Z(n1235) );
  XOR U110 ( .A(a[84]), .B(b[84]), .Z(n83) );
  NANDN U111 ( .A(n1239), .B(n83), .Z(n84) );
  NAND U112 ( .A(a[84]), .B(b[84]), .Z(n85) );
  AND U113 ( .A(n84), .B(n85), .Z(n1241) );
  XOR U114 ( .A(a[87]), .B(b[87]), .Z(n86) );
  NANDN U115 ( .A(n1245), .B(n86), .Z(n87) );
  NAND U116 ( .A(a[87]), .B(b[87]), .Z(n88) );
  AND U117 ( .A(n87), .B(n88), .Z(n1247) );
  XOR U118 ( .A(a[90]), .B(b[90]), .Z(n89) );
  NANDN U119 ( .A(n1253), .B(n89), .Z(n90) );
  NAND U120 ( .A(a[90]), .B(b[90]), .Z(n91) );
  AND U121 ( .A(n90), .B(n91), .Z(n1255) );
  XOR U122 ( .A(a[93]), .B(b[93]), .Z(n92) );
  NANDN U123 ( .A(n1259), .B(n92), .Z(n93) );
  NAND U124 ( .A(a[93]), .B(b[93]), .Z(n94) );
  AND U125 ( .A(n93), .B(n94), .Z(n1261) );
  XOR U126 ( .A(a[96]), .B(b[96]), .Z(n95) );
  NANDN U127 ( .A(n1265), .B(n95), .Z(n96) );
  NAND U128 ( .A(a[96]), .B(b[96]), .Z(n97) );
  AND U129 ( .A(n96), .B(n97), .Z(n1267) );
  XOR U130 ( .A(b[99]), .B(a[99]), .Z(n98) );
  NANDN U131 ( .A(n1271), .B(n98), .Z(n99) );
  NAND U132 ( .A(b[99]), .B(a[99]), .Z(n100) );
  AND U133 ( .A(n99), .B(n100), .Z(n768) );
  XOR U134 ( .A(b[102]), .B(a[102]), .Z(n101) );
  NANDN U135 ( .A(n772), .B(n101), .Z(n102) );
  NAND U136 ( .A(b[102]), .B(a[102]), .Z(n103) );
  AND U137 ( .A(n102), .B(n103), .Z(n774) );
  XOR U138 ( .A(b[105]), .B(a[105]), .Z(n104) );
  NANDN U139 ( .A(n778), .B(n104), .Z(n105) );
  NAND U140 ( .A(b[105]), .B(a[105]), .Z(n106) );
  AND U141 ( .A(n105), .B(n106), .Z(n780) );
  XOR U142 ( .A(b[108]), .B(a[108]), .Z(n107) );
  NANDN U143 ( .A(n784), .B(n107), .Z(n108) );
  NAND U144 ( .A(b[108]), .B(a[108]), .Z(n109) );
  AND U145 ( .A(n108), .B(n109), .Z(n788) );
  XOR U146 ( .A(b[111]), .B(a[111]), .Z(n110) );
  NANDN U147 ( .A(n792), .B(n110), .Z(n111) );
  NAND U148 ( .A(b[111]), .B(a[111]), .Z(n112) );
  AND U149 ( .A(n111), .B(n112), .Z(n794) );
  XOR U150 ( .A(b[114]), .B(a[114]), .Z(n113) );
  NANDN U151 ( .A(n798), .B(n113), .Z(n114) );
  NAND U152 ( .A(b[114]), .B(a[114]), .Z(n115) );
  AND U153 ( .A(n114), .B(n115), .Z(n800) );
  XOR U154 ( .A(b[117]), .B(a[117]), .Z(n116) );
  NANDN U155 ( .A(n804), .B(n116), .Z(n117) );
  NAND U156 ( .A(b[117]), .B(a[117]), .Z(n118) );
  AND U157 ( .A(n117), .B(n118), .Z(n806) );
  XOR U158 ( .A(b[120]), .B(a[120]), .Z(n119) );
  NANDN U159 ( .A(n812), .B(n119), .Z(n120) );
  NAND U160 ( .A(b[120]), .B(a[120]), .Z(n121) );
  AND U161 ( .A(n120), .B(n121), .Z(n814) );
  XOR U162 ( .A(b[123]), .B(a[123]), .Z(n122) );
  NANDN U163 ( .A(n818), .B(n122), .Z(n123) );
  NAND U164 ( .A(b[123]), .B(a[123]), .Z(n124) );
  AND U165 ( .A(n123), .B(n124), .Z(n820) );
  XOR U166 ( .A(b[126]), .B(a[126]), .Z(n125) );
  NANDN U167 ( .A(n824), .B(n125), .Z(n126) );
  NAND U168 ( .A(b[126]), .B(a[126]), .Z(n127) );
  AND U169 ( .A(n126), .B(n127), .Z(n826) );
  XOR U170 ( .A(b[129]), .B(a[129]), .Z(n128) );
  NANDN U171 ( .A(n832), .B(n128), .Z(n129) );
  NAND U172 ( .A(b[129]), .B(a[129]), .Z(n130) );
  AND U173 ( .A(n129), .B(n130), .Z(n834) );
  XOR U174 ( .A(b[132]), .B(a[132]), .Z(n131) );
  NANDN U175 ( .A(n838), .B(n131), .Z(n132) );
  NAND U176 ( .A(b[132]), .B(a[132]), .Z(n133) );
  AND U177 ( .A(n132), .B(n133), .Z(n840) );
  XOR U178 ( .A(b[135]), .B(a[135]), .Z(n134) );
  NANDN U179 ( .A(n844), .B(n134), .Z(n135) );
  NAND U180 ( .A(b[135]), .B(a[135]), .Z(n136) );
  AND U181 ( .A(n135), .B(n136), .Z(n846) );
  XOR U182 ( .A(b[138]), .B(a[138]), .Z(n137) );
  NANDN U183 ( .A(n850), .B(n137), .Z(n138) );
  NAND U184 ( .A(b[138]), .B(a[138]), .Z(n139) );
  AND U185 ( .A(n138), .B(n139), .Z(n854) );
  XOR U186 ( .A(b[141]), .B(a[141]), .Z(n140) );
  NANDN U187 ( .A(n858), .B(n140), .Z(n141) );
  NAND U188 ( .A(b[141]), .B(a[141]), .Z(n142) );
  AND U189 ( .A(n141), .B(n142), .Z(n860) );
  XOR U190 ( .A(b[144]), .B(a[144]), .Z(n143) );
  NANDN U191 ( .A(n864), .B(n143), .Z(n144) );
  NAND U192 ( .A(b[144]), .B(a[144]), .Z(n145) );
  AND U193 ( .A(n144), .B(n145), .Z(n866) );
  XOR U194 ( .A(b[147]), .B(a[147]), .Z(n146) );
  NANDN U195 ( .A(n870), .B(n146), .Z(n147) );
  NAND U196 ( .A(b[147]), .B(a[147]), .Z(n148) );
  AND U197 ( .A(n147), .B(n148), .Z(n872) );
  XOR U198 ( .A(b[150]), .B(a[150]), .Z(n149) );
  NANDN U199 ( .A(n878), .B(n149), .Z(n150) );
  NAND U200 ( .A(b[150]), .B(a[150]), .Z(n151) );
  AND U201 ( .A(n150), .B(n151), .Z(n880) );
  XOR U202 ( .A(b[153]), .B(a[153]), .Z(n152) );
  NANDN U203 ( .A(n884), .B(n152), .Z(n153) );
  NAND U204 ( .A(b[153]), .B(a[153]), .Z(n154) );
  AND U205 ( .A(n153), .B(n154), .Z(n886) );
  XOR U206 ( .A(b[156]), .B(a[156]), .Z(n155) );
  NANDN U207 ( .A(n890), .B(n155), .Z(n156) );
  NAND U208 ( .A(b[156]), .B(a[156]), .Z(n157) );
  AND U209 ( .A(n156), .B(n157), .Z(n892) );
  XOR U210 ( .A(b[159]), .B(a[159]), .Z(n158) );
  NANDN U211 ( .A(n898), .B(n158), .Z(n159) );
  NAND U212 ( .A(b[159]), .B(a[159]), .Z(n160) );
  AND U213 ( .A(n159), .B(n160), .Z(n900) );
  XOR U214 ( .A(b[162]), .B(a[162]), .Z(n161) );
  NANDN U215 ( .A(n904), .B(n161), .Z(n162) );
  NAND U216 ( .A(b[162]), .B(a[162]), .Z(n163) );
  AND U217 ( .A(n162), .B(n163), .Z(n906) );
  XOR U218 ( .A(b[165]), .B(a[165]), .Z(n164) );
  NANDN U219 ( .A(n910), .B(n164), .Z(n165) );
  NAND U220 ( .A(b[165]), .B(a[165]), .Z(n166) );
  AND U221 ( .A(n165), .B(n166), .Z(n912) );
  XOR U222 ( .A(b[168]), .B(a[168]), .Z(n167) );
  NANDN U223 ( .A(n916), .B(n167), .Z(n168) );
  NAND U224 ( .A(b[168]), .B(a[168]), .Z(n169) );
  AND U225 ( .A(n168), .B(n169), .Z(n920) );
  XOR U226 ( .A(b[171]), .B(a[171]), .Z(n170) );
  NANDN U227 ( .A(n924), .B(n170), .Z(n171) );
  NAND U228 ( .A(b[171]), .B(a[171]), .Z(n172) );
  AND U229 ( .A(n171), .B(n172), .Z(n926) );
  XOR U230 ( .A(b[174]), .B(a[174]), .Z(n173) );
  NANDN U231 ( .A(n930), .B(n173), .Z(n174) );
  NAND U232 ( .A(b[174]), .B(a[174]), .Z(n175) );
  AND U233 ( .A(n174), .B(n175), .Z(n932) );
  XOR U234 ( .A(b[177]), .B(a[177]), .Z(n176) );
  NANDN U235 ( .A(n936), .B(n176), .Z(n177) );
  NAND U236 ( .A(b[177]), .B(a[177]), .Z(n178) );
  AND U237 ( .A(n177), .B(n178), .Z(n938) );
  XOR U238 ( .A(b[180]), .B(a[180]), .Z(n179) );
  NANDN U239 ( .A(n944), .B(n179), .Z(n180) );
  NAND U240 ( .A(b[180]), .B(a[180]), .Z(n181) );
  AND U241 ( .A(n180), .B(n181), .Z(n946) );
  XOR U242 ( .A(b[183]), .B(a[183]), .Z(n182) );
  NANDN U243 ( .A(n950), .B(n182), .Z(n183) );
  NAND U244 ( .A(b[183]), .B(a[183]), .Z(n184) );
  AND U245 ( .A(n183), .B(n184), .Z(n952) );
  XOR U246 ( .A(b[186]), .B(a[186]), .Z(n185) );
  NANDN U247 ( .A(n956), .B(n185), .Z(n186) );
  NAND U248 ( .A(b[186]), .B(a[186]), .Z(n187) );
  AND U249 ( .A(n186), .B(n187), .Z(n958) );
  XOR U250 ( .A(b[189]), .B(a[189]), .Z(n188) );
  NANDN U251 ( .A(n964), .B(n188), .Z(n189) );
  NAND U252 ( .A(b[189]), .B(a[189]), .Z(n190) );
  AND U253 ( .A(n189), .B(n190), .Z(n966) );
  XOR U254 ( .A(b[192]), .B(a[192]), .Z(n191) );
  NANDN U255 ( .A(n970), .B(n191), .Z(n192) );
  NAND U256 ( .A(b[192]), .B(a[192]), .Z(n193) );
  AND U257 ( .A(n192), .B(n193), .Z(n972) );
  XOR U258 ( .A(b[195]), .B(a[195]), .Z(n194) );
  NANDN U259 ( .A(n976), .B(n194), .Z(n195) );
  NAND U260 ( .A(b[195]), .B(a[195]), .Z(n196) );
  AND U261 ( .A(n195), .B(n196), .Z(n978) );
  XOR U262 ( .A(b[198]), .B(a[198]), .Z(n197) );
  NANDN U263 ( .A(n982), .B(n197), .Z(n198) );
  NAND U264 ( .A(b[198]), .B(a[198]), .Z(n199) );
  AND U265 ( .A(n198), .B(n199), .Z(n988) );
  XOR U266 ( .A(b[201]), .B(a[201]), .Z(n200) );
  NANDN U267 ( .A(n992), .B(n200), .Z(n201) );
  NAND U268 ( .A(b[201]), .B(a[201]), .Z(n202) );
  AND U269 ( .A(n201), .B(n202), .Z(n994) );
  XOR U270 ( .A(b[204]), .B(a[204]), .Z(n203) );
  NANDN U271 ( .A(n998), .B(n203), .Z(n204) );
  NAND U272 ( .A(b[204]), .B(a[204]), .Z(n205) );
  AND U273 ( .A(n204), .B(n205), .Z(n1000) );
  XOR U274 ( .A(b[207]), .B(a[207]), .Z(n206) );
  NANDN U275 ( .A(n1004), .B(n206), .Z(n207) );
  NAND U276 ( .A(b[207]), .B(a[207]), .Z(n208) );
  AND U277 ( .A(n207), .B(n208), .Z(n1006) );
  XOR U278 ( .A(b[210]), .B(a[210]), .Z(n209) );
  NANDN U279 ( .A(n1012), .B(n209), .Z(n210) );
  NAND U280 ( .A(b[210]), .B(a[210]), .Z(n211) );
  AND U281 ( .A(n210), .B(n211), .Z(n1014) );
  XOR U282 ( .A(b[213]), .B(a[213]), .Z(n212) );
  NANDN U283 ( .A(n1018), .B(n212), .Z(n213) );
  NAND U284 ( .A(b[213]), .B(a[213]), .Z(n214) );
  AND U285 ( .A(n213), .B(n214), .Z(n1020) );
  XOR U286 ( .A(b[216]), .B(a[216]), .Z(n215) );
  NANDN U287 ( .A(n1024), .B(n215), .Z(n216) );
  NAND U288 ( .A(b[216]), .B(a[216]), .Z(n217) );
  AND U289 ( .A(n216), .B(n217), .Z(n1026) );
  XOR U290 ( .A(b[219]), .B(a[219]), .Z(n218) );
  NANDN U291 ( .A(n1032), .B(n218), .Z(n219) );
  NAND U292 ( .A(b[219]), .B(a[219]), .Z(n220) );
  AND U293 ( .A(n219), .B(n220), .Z(n1034) );
  XOR U294 ( .A(b[222]), .B(a[222]), .Z(n221) );
  NANDN U295 ( .A(n1038), .B(n221), .Z(n222) );
  NAND U296 ( .A(b[222]), .B(a[222]), .Z(n223) );
  AND U297 ( .A(n222), .B(n223), .Z(n1040) );
  XOR U298 ( .A(b[225]), .B(a[225]), .Z(n224) );
  NANDN U299 ( .A(n1044), .B(n224), .Z(n225) );
  NAND U300 ( .A(b[225]), .B(a[225]), .Z(n226) );
  AND U301 ( .A(n225), .B(n226), .Z(n1046) );
  XOR U302 ( .A(b[228]), .B(a[228]), .Z(n227) );
  NANDN U303 ( .A(n1050), .B(n227), .Z(n228) );
  NAND U304 ( .A(b[228]), .B(a[228]), .Z(n229) );
  AND U305 ( .A(n228), .B(n229), .Z(n1054) );
  XOR U306 ( .A(b[231]), .B(a[231]), .Z(n230) );
  NANDN U307 ( .A(n1058), .B(n230), .Z(n231) );
  NAND U308 ( .A(b[231]), .B(a[231]), .Z(n232) );
  AND U309 ( .A(n231), .B(n232), .Z(n1060) );
  XOR U310 ( .A(b[234]), .B(a[234]), .Z(n233) );
  NANDN U311 ( .A(n1064), .B(n233), .Z(n234) );
  NAND U312 ( .A(b[234]), .B(a[234]), .Z(n235) );
  AND U313 ( .A(n234), .B(n235), .Z(n1066) );
  XOR U314 ( .A(b[237]), .B(a[237]), .Z(n236) );
  NANDN U315 ( .A(n1070), .B(n236), .Z(n237) );
  NAND U316 ( .A(b[237]), .B(a[237]), .Z(n238) );
  AND U317 ( .A(n237), .B(n238), .Z(n1072) );
  XOR U318 ( .A(b[240]), .B(a[240]), .Z(n239) );
  NANDN U319 ( .A(n1078), .B(n239), .Z(n240) );
  NAND U320 ( .A(b[240]), .B(a[240]), .Z(n241) );
  AND U321 ( .A(n240), .B(n241), .Z(n1080) );
  XOR U322 ( .A(b[243]), .B(a[243]), .Z(n242) );
  NANDN U323 ( .A(n1084), .B(n242), .Z(n243) );
  NAND U324 ( .A(b[243]), .B(a[243]), .Z(n244) );
  AND U325 ( .A(n243), .B(n244), .Z(n1086) );
  XOR U326 ( .A(b[246]), .B(a[246]), .Z(n245) );
  NANDN U327 ( .A(n1090), .B(n245), .Z(n246) );
  NAND U328 ( .A(b[246]), .B(a[246]), .Z(n247) );
  AND U329 ( .A(n246), .B(n247), .Z(n1092) );
  XOR U330 ( .A(b[249]), .B(a[249]), .Z(n248) );
  NANDN U331 ( .A(n1098), .B(n248), .Z(n249) );
  NAND U332 ( .A(b[249]), .B(a[249]), .Z(n250) );
  AND U333 ( .A(n249), .B(n250), .Z(n1100) );
  XOR U334 ( .A(b[252]), .B(a[252]), .Z(n251) );
  NANDN U335 ( .A(n1104), .B(n251), .Z(n252) );
  NAND U336 ( .A(b[252]), .B(a[252]), .Z(n253) );
  AND U337 ( .A(n252), .B(n253), .Z(n1106) );
  XOR U338 ( .A(b[1]), .B(a[1]), .Z(n254) );
  NANDN U339 ( .A(n987), .B(n254), .Z(n255) );
  NAND U340 ( .A(b[1]), .B(a[1]), .Z(n256) );
  AND U341 ( .A(n255), .B(n256), .Z(n1119) );
  XOR U342 ( .A(a[4]), .B(b[4]), .Z(n257) );
  NANDN U343 ( .A(n1163), .B(n257), .Z(n258) );
  NAND U344 ( .A(a[4]), .B(b[4]), .Z(n259) );
  AND U345 ( .A(n258), .B(n259), .Z(n1185) );
  XOR U346 ( .A(a[7]), .B(b[7]), .Z(n260) );
  NANDN U347 ( .A(n1229), .B(n260), .Z(n261) );
  NAND U348 ( .A(a[7]), .B(b[7]), .Z(n262) );
  AND U349 ( .A(n261), .B(n262), .Z(n1251) );
  XOR U350 ( .A(a[10]), .B(b[10]), .Z(n263) );
  NANDN U351 ( .A(n786), .B(n263), .Z(n264) );
  NAND U352 ( .A(a[10]), .B(b[10]), .Z(n265) );
  AND U353 ( .A(n264), .B(n265), .Z(n808) );
  XOR U354 ( .A(a[13]), .B(b[13]), .Z(n266) );
  NANDN U355 ( .A(n852), .B(n266), .Z(n267) );
  NAND U356 ( .A(a[13]), .B(b[13]), .Z(n268) );
  AND U357 ( .A(n267), .B(n268), .Z(n874) );
  XOR U358 ( .A(a[16]), .B(b[16]), .Z(n269) );
  NANDN U359 ( .A(n918), .B(n269), .Z(n270) );
  NAND U360 ( .A(a[16]), .B(b[16]), .Z(n271) );
  AND U361 ( .A(n270), .B(n271), .Z(n940) );
  XOR U362 ( .A(a[19]), .B(b[19]), .Z(n272) );
  NANDN U363 ( .A(n984), .B(n272), .Z(n273) );
  NAND U364 ( .A(a[19]), .B(b[19]), .Z(n274) );
  AND U365 ( .A(n273), .B(n274), .Z(n1008) );
  XOR U366 ( .A(a[22]), .B(b[22]), .Z(n275) );
  NANDN U367 ( .A(n1052), .B(n275), .Z(n276) );
  NAND U368 ( .A(a[22]), .B(b[22]), .Z(n277) );
  AND U369 ( .A(n276), .B(n277), .Z(n1074) );
  XOR U370 ( .A(a[28]), .B(b[28]), .Z(n278) );
  NANDN U371 ( .A(n1115), .B(n278), .Z(n279) );
  NAND U372 ( .A(a[28]), .B(b[28]), .Z(n280) );
  AND U373 ( .A(n279), .B(n280), .Z(n1117) );
  XOR U374 ( .A(a[31]), .B(b[31]), .Z(n281) );
  NANDN U375 ( .A(n1123), .B(n281), .Z(n282) );
  NAND U376 ( .A(a[31]), .B(b[31]), .Z(n283) );
  AND U377 ( .A(n282), .B(n283), .Z(n1125) );
  XOR U378 ( .A(a[34]), .B(b[34]), .Z(n284) );
  NANDN U379 ( .A(n1129), .B(n284), .Z(n285) );
  NAND U380 ( .A(a[34]), .B(b[34]), .Z(n286) );
  AND U381 ( .A(n285), .B(n286), .Z(n1131) );
  XOR U382 ( .A(a[37]), .B(b[37]), .Z(n287) );
  NANDN U383 ( .A(n1135), .B(n287), .Z(n288) );
  NAND U384 ( .A(a[37]), .B(b[37]), .Z(n289) );
  AND U385 ( .A(n288), .B(n289), .Z(n1137) );
  XOR U386 ( .A(a[40]), .B(b[40]), .Z(n290) );
  NANDN U387 ( .A(n1143), .B(n290), .Z(n291) );
  NAND U388 ( .A(a[40]), .B(b[40]), .Z(n292) );
  AND U389 ( .A(n291), .B(n292), .Z(n1145) );
  XOR U390 ( .A(a[43]), .B(b[43]), .Z(n293) );
  NANDN U391 ( .A(n1149), .B(n293), .Z(n294) );
  NAND U392 ( .A(a[43]), .B(b[43]), .Z(n295) );
  AND U393 ( .A(n294), .B(n295), .Z(n1151) );
  XOR U394 ( .A(a[46]), .B(b[46]), .Z(n296) );
  NANDN U395 ( .A(n1155), .B(n296), .Z(n297) );
  NAND U396 ( .A(a[46]), .B(b[46]), .Z(n298) );
  AND U397 ( .A(n297), .B(n298), .Z(n1157) );
  XOR U398 ( .A(a[49]), .B(b[49]), .Z(n299) );
  NANDN U399 ( .A(n1161), .B(n299), .Z(n300) );
  NAND U400 ( .A(a[49]), .B(b[49]), .Z(n301) );
  AND U401 ( .A(n300), .B(n301), .Z(n1165) );
  XOR U402 ( .A(a[52]), .B(b[52]), .Z(n302) );
  NANDN U403 ( .A(n1169), .B(n302), .Z(n303) );
  NAND U404 ( .A(a[52]), .B(b[52]), .Z(n304) );
  AND U405 ( .A(n303), .B(n304), .Z(n1171) );
  XOR U406 ( .A(a[55]), .B(b[55]), .Z(n305) );
  NANDN U407 ( .A(n1175), .B(n305), .Z(n306) );
  NAND U408 ( .A(a[55]), .B(b[55]), .Z(n307) );
  AND U409 ( .A(n306), .B(n307), .Z(n1177) );
  XOR U410 ( .A(a[58]), .B(b[58]), .Z(n308) );
  NANDN U411 ( .A(n1181), .B(n308), .Z(n309) );
  NAND U412 ( .A(a[58]), .B(b[58]), .Z(n310) );
  AND U413 ( .A(n309), .B(n310), .Z(n1183) );
  XOR U414 ( .A(a[61]), .B(b[61]), .Z(n311) );
  NANDN U415 ( .A(n1189), .B(n311), .Z(n312) );
  NAND U416 ( .A(a[61]), .B(b[61]), .Z(n313) );
  AND U417 ( .A(n312), .B(n313), .Z(n1191) );
  XOR U418 ( .A(a[64]), .B(b[64]), .Z(n314) );
  NANDN U419 ( .A(n1195), .B(n314), .Z(n315) );
  NAND U420 ( .A(a[64]), .B(b[64]), .Z(n316) );
  AND U421 ( .A(n315), .B(n316), .Z(n1197) );
  XOR U422 ( .A(a[67]), .B(b[67]), .Z(n317) );
  NANDN U423 ( .A(n1201), .B(n317), .Z(n318) );
  NAND U424 ( .A(a[67]), .B(b[67]), .Z(n319) );
  AND U425 ( .A(n318), .B(n319), .Z(n1203) );
  XOR U426 ( .A(a[70]), .B(b[70]), .Z(n320) );
  NANDN U427 ( .A(n1209), .B(n320), .Z(n321) );
  NAND U428 ( .A(a[70]), .B(b[70]), .Z(n322) );
  AND U429 ( .A(n321), .B(n322), .Z(n1211) );
  XOR U430 ( .A(a[73]), .B(b[73]), .Z(n323) );
  NANDN U431 ( .A(n1215), .B(n323), .Z(n324) );
  NAND U432 ( .A(a[73]), .B(b[73]), .Z(n325) );
  AND U433 ( .A(n324), .B(n325), .Z(n1217) );
  XOR U434 ( .A(a[76]), .B(b[76]), .Z(n326) );
  NANDN U435 ( .A(n1221), .B(n326), .Z(n327) );
  NAND U436 ( .A(a[76]), .B(b[76]), .Z(n328) );
  AND U437 ( .A(n327), .B(n328), .Z(n1223) );
  XOR U438 ( .A(a[79]), .B(b[79]), .Z(n329) );
  NANDN U439 ( .A(n1227), .B(n329), .Z(n330) );
  NAND U440 ( .A(a[79]), .B(b[79]), .Z(n331) );
  AND U441 ( .A(n330), .B(n331), .Z(n1231) );
  XOR U442 ( .A(a[82]), .B(b[82]), .Z(n332) );
  NANDN U443 ( .A(n1235), .B(n332), .Z(n333) );
  NAND U444 ( .A(a[82]), .B(b[82]), .Z(n334) );
  AND U445 ( .A(n333), .B(n334), .Z(n1237) );
  XOR U446 ( .A(a[85]), .B(b[85]), .Z(n335) );
  NANDN U447 ( .A(n1241), .B(n335), .Z(n336) );
  NAND U448 ( .A(a[85]), .B(b[85]), .Z(n337) );
  AND U449 ( .A(n336), .B(n337), .Z(n1243) );
  XOR U450 ( .A(a[88]), .B(b[88]), .Z(n338) );
  NANDN U451 ( .A(n1247), .B(n338), .Z(n339) );
  NAND U452 ( .A(a[88]), .B(b[88]), .Z(n340) );
  AND U453 ( .A(n339), .B(n340), .Z(n1249) );
  XOR U454 ( .A(a[91]), .B(b[91]), .Z(n341) );
  NANDN U455 ( .A(n1255), .B(n341), .Z(n342) );
  NAND U456 ( .A(a[91]), .B(b[91]), .Z(n343) );
  AND U457 ( .A(n342), .B(n343), .Z(n1257) );
  XOR U458 ( .A(a[94]), .B(b[94]), .Z(n344) );
  NANDN U459 ( .A(n1261), .B(n344), .Z(n345) );
  NAND U460 ( .A(a[94]), .B(b[94]), .Z(n346) );
  AND U461 ( .A(n345), .B(n346), .Z(n1263) );
  XOR U462 ( .A(a[97]), .B(b[97]), .Z(n347) );
  NANDN U463 ( .A(n1267), .B(n347), .Z(n348) );
  NAND U464 ( .A(a[97]), .B(b[97]), .Z(n349) );
  AND U465 ( .A(n348), .B(n349), .Z(n1269) );
  XOR U466 ( .A(b[100]), .B(a[100]), .Z(n350) );
  NANDN U467 ( .A(n768), .B(n350), .Z(n351) );
  NAND U468 ( .A(b[100]), .B(a[100]), .Z(n352) );
  AND U469 ( .A(n351), .B(n352), .Z(n770) );
  XOR U470 ( .A(b[103]), .B(a[103]), .Z(n353) );
  NANDN U471 ( .A(n774), .B(n353), .Z(n354) );
  NAND U472 ( .A(b[103]), .B(a[103]), .Z(n355) );
  AND U473 ( .A(n354), .B(n355), .Z(n776) );
  XOR U474 ( .A(b[106]), .B(a[106]), .Z(n356) );
  NANDN U475 ( .A(n780), .B(n356), .Z(n357) );
  NAND U476 ( .A(b[106]), .B(a[106]), .Z(n358) );
  AND U477 ( .A(n357), .B(n358), .Z(n782) );
  XOR U478 ( .A(b[109]), .B(a[109]), .Z(n359) );
  NANDN U479 ( .A(n788), .B(n359), .Z(n360) );
  NAND U480 ( .A(b[109]), .B(a[109]), .Z(n361) );
  AND U481 ( .A(n360), .B(n361), .Z(n790) );
  XOR U482 ( .A(b[112]), .B(a[112]), .Z(n362) );
  NANDN U483 ( .A(n794), .B(n362), .Z(n363) );
  NAND U484 ( .A(b[112]), .B(a[112]), .Z(n364) );
  AND U485 ( .A(n363), .B(n364), .Z(n796) );
  XOR U486 ( .A(b[115]), .B(a[115]), .Z(n365) );
  NANDN U487 ( .A(n800), .B(n365), .Z(n366) );
  NAND U488 ( .A(b[115]), .B(a[115]), .Z(n367) );
  AND U489 ( .A(n366), .B(n367), .Z(n802) );
  XOR U490 ( .A(b[118]), .B(a[118]), .Z(n368) );
  NANDN U491 ( .A(n806), .B(n368), .Z(n369) );
  NAND U492 ( .A(b[118]), .B(a[118]), .Z(n370) );
  AND U493 ( .A(n369), .B(n370), .Z(n810) );
  XOR U494 ( .A(b[121]), .B(a[121]), .Z(n371) );
  NANDN U495 ( .A(n814), .B(n371), .Z(n372) );
  NAND U496 ( .A(b[121]), .B(a[121]), .Z(n373) );
  AND U497 ( .A(n372), .B(n373), .Z(n816) );
  XOR U498 ( .A(b[124]), .B(a[124]), .Z(n374) );
  NANDN U499 ( .A(n820), .B(n374), .Z(n375) );
  NAND U500 ( .A(b[124]), .B(a[124]), .Z(n376) );
  AND U501 ( .A(n375), .B(n376), .Z(n822) );
  XOR U502 ( .A(b[127]), .B(a[127]), .Z(n377) );
  NANDN U503 ( .A(n826), .B(n377), .Z(n378) );
  NAND U504 ( .A(b[127]), .B(a[127]), .Z(n379) );
  AND U505 ( .A(n378), .B(n379), .Z(n828) );
  XOR U506 ( .A(b[130]), .B(a[130]), .Z(n380) );
  NANDN U507 ( .A(n834), .B(n380), .Z(n381) );
  NAND U508 ( .A(b[130]), .B(a[130]), .Z(n382) );
  AND U509 ( .A(n381), .B(n382), .Z(n836) );
  XOR U510 ( .A(b[133]), .B(a[133]), .Z(n383) );
  NANDN U511 ( .A(n840), .B(n383), .Z(n384) );
  NAND U512 ( .A(b[133]), .B(a[133]), .Z(n385) );
  AND U513 ( .A(n384), .B(n385), .Z(n842) );
  XOR U514 ( .A(b[136]), .B(a[136]), .Z(n386) );
  NANDN U515 ( .A(n846), .B(n386), .Z(n387) );
  NAND U516 ( .A(b[136]), .B(a[136]), .Z(n388) );
  AND U517 ( .A(n387), .B(n388), .Z(n848) );
  XOR U518 ( .A(b[139]), .B(a[139]), .Z(n389) );
  NANDN U519 ( .A(n854), .B(n389), .Z(n390) );
  NAND U520 ( .A(b[139]), .B(a[139]), .Z(n391) );
  AND U521 ( .A(n390), .B(n391), .Z(n856) );
  XOR U522 ( .A(b[142]), .B(a[142]), .Z(n392) );
  NANDN U523 ( .A(n860), .B(n392), .Z(n393) );
  NAND U524 ( .A(b[142]), .B(a[142]), .Z(n394) );
  AND U525 ( .A(n393), .B(n394), .Z(n862) );
  XOR U526 ( .A(b[145]), .B(a[145]), .Z(n395) );
  NANDN U527 ( .A(n866), .B(n395), .Z(n396) );
  NAND U528 ( .A(b[145]), .B(a[145]), .Z(n397) );
  AND U529 ( .A(n396), .B(n397), .Z(n868) );
  XOR U530 ( .A(b[148]), .B(a[148]), .Z(n398) );
  NANDN U531 ( .A(n872), .B(n398), .Z(n399) );
  NAND U532 ( .A(b[148]), .B(a[148]), .Z(n400) );
  AND U533 ( .A(n399), .B(n400), .Z(n876) );
  XOR U534 ( .A(b[151]), .B(a[151]), .Z(n401) );
  NANDN U535 ( .A(n880), .B(n401), .Z(n402) );
  NAND U536 ( .A(b[151]), .B(a[151]), .Z(n403) );
  AND U537 ( .A(n402), .B(n403), .Z(n882) );
  XOR U538 ( .A(b[154]), .B(a[154]), .Z(n404) );
  NANDN U539 ( .A(n886), .B(n404), .Z(n405) );
  NAND U540 ( .A(b[154]), .B(a[154]), .Z(n406) );
  AND U541 ( .A(n405), .B(n406), .Z(n888) );
  XOR U542 ( .A(b[157]), .B(a[157]), .Z(n407) );
  NANDN U543 ( .A(n892), .B(n407), .Z(n408) );
  NAND U544 ( .A(b[157]), .B(a[157]), .Z(n409) );
  AND U545 ( .A(n408), .B(n409), .Z(n894) );
  XOR U546 ( .A(b[160]), .B(a[160]), .Z(n410) );
  NANDN U547 ( .A(n900), .B(n410), .Z(n411) );
  NAND U548 ( .A(b[160]), .B(a[160]), .Z(n412) );
  AND U549 ( .A(n411), .B(n412), .Z(n902) );
  XOR U550 ( .A(b[163]), .B(a[163]), .Z(n413) );
  NANDN U551 ( .A(n906), .B(n413), .Z(n414) );
  NAND U552 ( .A(b[163]), .B(a[163]), .Z(n415) );
  AND U553 ( .A(n414), .B(n415), .Z(n908) );
  XOR U554 ( .A(b[166]), .B(a[166]), .Z(n416) );
  NANDN U555 ( .A(n912), .B(n416), .Z(n417) );
  NAND U556 ( .A(b[166]), .B(a[166]), .Z(n418) );
  AND U557 ( .A(n417), .B(n418), .Z(n914) );
  XOR U558 ( .A(b[169]), .B(a[169]), .Z(n419) );
  NANDN U559 ( .A(n920), .B(n419), .Z(n420) );
  NAND U560 ( .A(b[169]), .B(a[169]), .Z(n421) );
  AND U561 ( .A(n420), .B(n421), .Z(n922) );
  XOR U562 ( .A(b[172]), .B(a[172]), .Z(n422) );
  NANDN U563 ( .A(n926), .B(n422), .Z(n423) );
  NAND U564 ( .A(b[172]), .B(a[172]), .Z(n424) );
  AND U565 ( .A(n423), .B(n424), .Z(n928) );
  XOR U566 ( .A(b[175]), .B(a[175]), .Z(n425) );
  NANDN U567 ( .A(n932), .B(n425), .Z(n426) );
  NAND U568 ( .A(b[175]), .B(a[175]), .Z(n427) );
  AND U569 ( .A(n426), .B(n427), .Z(n934) );
  XOR U570 ( .A(b[178]), .B(a[178]), .Z(n428) );
  NANDN U571 ( .A(n938), .B(n428), .Z(n429) );
  NAND U572 ( .A(b[178]), .B(a[178]), .Z(n430) );
  AND U573 ( .A(n429), .B(n430), .Z(n942) );
  XOR U574 ( .A(b[181]), .B(a[181]), .Z(n431) );
  NANDN U575 ( .A(n946), .B(n431), .Z(n432) );
  NAND U576 ( .A(b[181]), .B(a[181]), .Z(n433) );
  AND U577 ( .A(n432), .B(n433), .Z(n948) );
  XOR U578 ( .A(b[184]), .B(a[184]), .Z(n434) );
  NANDN U579 ( .A(n952), .B(n434), .Z(n435) );
  NAND U580 ( .A(b[184]), .B(a[184]), .Z(n436) );
  AND U581 ( .A(n435), .B(n436), .Z(n954) );
  XOR U582 ( .A(b[187]), .B(a[187]), .Z(n437) );
  NANDN U583 ( .A(n958), .B(n437), .Z(n438) );
  NAND U584 ( .A(b[187]), .B(a[187]), .Z(n439) );
  AND U585 ( .A(n438), .B(n439), .Z(n960) );
  XOR U586 ( .A(b[190]), .B(a[190]), .Z(n440) );
  NANDN U587 ( .A(n966), .B(n440), .Z(n441) );
  NAND U588 ( .A(b[190]), .B(a[190]), .Z(n442) );
  AND U589 ( .A(n441), .B(n442), .Z(n968) );
  XOR U590 ( .A(b[193]), .B(a[193]), .Z(n443) );
  NANDN U591 ( .A(n972), .B(n443), .Z(n444) );
  NAND U592 ( .A(b[193]), .B(a[193]), .Z(n445) );
  AND U593 ( .A(n444), .B(n445), .Z(n974) );
  XOR U594 ( .A(b[196]), .B(a[196]), .Z(n446) );
  NANDN U595 ( .A(n978), .B(n446), .Z(n447) );
  NAND U596 ( .A(b[196]), .B(a[196]), .Z(n448) );
  AND U597 ( .A(n447), .B(n448), .Z(n980) );
  XOR U598 ( .A(b[199]), .B(a[199]), .Z(n449) );
  NANDN U599 ( .A(n988), .B(n449), .Z(n450) );
  NAND U600 ( .A(b[199]), .B(a[199]), .Z(n451) );
  AND U601 ( .A(n450), .B(n451), .Z(n990) );
  XOR U602 ( .A(b[202]), .B(a[202]), .Z(n452) );
  NANDN U603 ( .A(n994), .B(n452), .Z(n453) );
  NAND U604 ( .A(b[202]), .B(a[202]), .Z(n454) );
  AND U605 ( .A(n453), .B(n454), .Z(n996) );
  XOR U606 ( .A(b[205]), .B(a[205]), .Z(n455) );
  NANDN U607 ( .A(n1000), .B(n455), .Z(n456) );
  NAND U608 ( .A(b[205]), .B(a[205]), .Z(n457) );
  AND U609 ( .A(n456), .B(n457), .Z(n1002) );
  XOR U610 ( .A(b[208]), .B(a[208]), .Z(n458) );
  NANDN U611 ( .A(n1006), .B(n458), .Z(n459) );
  NAND U612 ( .A(b[208]), .B(a[208]), .Z(n460) );
  AND U613 ( .A(n459), .B(n460), .Z(n1010) );
  XOR U614 ( .A(b[211]), .B(a[211]), .Z(n461) );
  NANDN U615 ( .A(n1014), .B(n461), .Z(n462) );
  NAND U616 ( .A(b[211]), .B(a[211]), .Z(n463) );
  AND U617 ( .A(n462), .B(n463), .Z(n1016) );
  XOR U618 ( .A(b[214]), .B(a[214]), .Z(n464) );
  NANDN U619 ( .A(n1020), .B(n464), .Z(n465) );
  NAND U620 ( .A(b[214]), .B(a[214]), .Z(n466) );
  AND U621 ( .A(n465), .B(n466), .Z(n1022) );
  XOR U622 ( .A(b[217]), .B(a[217]), .Z(n467) );
  NANDN U623 ( .A(n1026), .B(n467), .Z(n468) );
  NAND U624 ( .A(b[217]), .B(a[217]), .Z(n469) );
  AND U625 ( .A(n468), .B(n469), .Z(n1028) );
  XOR U626 ( .A(b[220]), .B(a[220]), .Z(n470) );
  NANDN U627 ( .A(n1034), .B(n470), .Z(n471) );
  NAND U628 ( .A(b[220]), .B(a[220]), .Z(n472) );
  AND U629 ( .A(n471), .B(n472), .Z(n1036) );
  XOR U630 ( .A(b[223]), .B(a[223]), .Z(n473) );
  NANDN U631 ( .A(n1040), .B(n473), .Z(n474) );
  NAND U632 ( .A(b[223]), .B(a[223]), .Z(n475) );
  AND U633 ( .A(n474), .B(n475), .Z(n1042) );
  XOR U634 ( .A(b[226]), .B(a[226]), .Z(n476) );
  NANDN U635 ( .A(n1046), .B(n476), .Z(n477) );
  NAND U636 ( .A(b[226]), .B(a[226]), .Z(n478) );
  AND U637 ( .A(n477), .B(n478), .Z(n1048) );
  XOR U638 ( .A(b[229]), .B(a[229]), .Z(n479) );
  NANDN U639 ( .A(n1054), .B(n479), .Z(n480) );
  NAND U640 ( .A(b[229]), .B(a[229]), .Z(n481) );
  AND U641 ( .A(n480), .B(n481), .Z(n1056) );
  XOR U642 ( .A(b[232]), .B(a[232]), .Z(n482) );
  NANDN U643 ( .A(n1060), .B(n482), .Z(n483) );
  NAND U644 ( .A(b[232]), .B(a[232]), .Z(n484) );
  AND U645 ( .A(n483), .B(n484), .Z(n1062) );
  XOR U646 ( .A(b[235]), .B(a[235]), .Z(n485) );
  NANDN U647 ( .A(n1066), .B(n485), .Z(n486) );
  NAND U648 ( .A(b[235]), .B(a[235]), .Z(n487) );
  AND U649 ( .A(n486), .B(n487), .Z(n1068) );
  XOR U650 ( .A(b[238]), .B(a[238]), .Z(n488) );
  NANDN U651 ( .A(n1072), .B(n488), .Z(n489) );
  NAND U652 ( .A(b[238]), .B(a[238]), .Z(n490) );
  AND U653 ( .A(n489), .B(n490), .Z(n1076) );
  XOR U654 ( .A(b[241]), .B(a[241]), .Z(n491) );
  NANDN U655 ( .A(n1080), .B(n491), .Z(n492) );
  NAND U656 ( .A(b[241]), .B(a[241]), .Z(n493) );
  AND U657 ( .A(n492), .B(n493), .Z(n1082) );
  XOR U658 ( .A(b[244]), .B(a[244]), .Z(n494) );
  NANDN U659 ( .A(n1086), .B(n494), .Z(n495) );
  NAND U660 ( .A(b[244]), .B(a[244]), .Z(n496) );
  AND U661 ( .A(n495), .B(n496), .Z(n1088) );
  XOR U662 ( .A(b[247]), .B(a[247]), .Z(n497) );
  NANDN U663 ( .A(n1092), .B(n497), .Z(n498) );
  NAND U664 ( .A(b[247]), .B(a[247]), .Z(n499) );
  AND U665 ( .A(n498), .B(n499), .Z(n1094) );
  XOR U666 ( .A(b[250]), .B(a[250]), .Z(n500) );
  NANDN U667 ( .A(n1100), .B(n500), .Z(n501) );
  NAND U668 ( .A(b[250]), .B(a[250]), .Z(n502) );
  AND U669 ( .A(n501), .B(n502), .Z(n1102) );
  XOR U670 ( .A(b[253]), .B(a[253]), .Z(n503) );
  NANDN U671 ( .A(n1106), .B(n503), .Z(n504) );
  NAND U672 ( .A(b[253]), .B(a[253]), .Z(n505) );
  AND U673 ( .A(n504), .B(n505), .Z(n1108) );
  XOR U674 ( .A(a[2]), .B(b[2]), .Z(n506) );
  NANDN U675 ( .A(n1119), .B(n506), .Z(n507) );
  NAND U676 ( .A(a[2]), .B(b[2]), .Z(n508) );
  AND U677 ( .A(n507), .B(n508), .Z(n1141) );
  XOR U678 ( .A(a[5]), .B(b[5]), .Z(n509) );
  NANDN U679 ( .A(n1185), .B(n509), .Z(n510) );
  NAND U680 ( .A(a[5]), .B(b[5]), .Z(n511) );
  AND U681 ( .A(n510), .B(n511), .Z(n1207) );
  XOR U682 ( .A(a[8]), .B(b[8]), .Z(n512) );
  NANDN U683 ( .A(n1251), .B(n512), .Z(n513) );
  NAND U684 ( .A(a[8]), .B(b[8]), .Z(n514) );
  AND U685 ( .A(n513), .B(n514), .Z(n1273) );
  XOR U686 ( .A(a[11]), .B(b[11]), .Z(n515) );
  NANDN U687 ( .A(n808), .B(n515), .Z(n516) );
  NAND U688 ( .A(a[11]), .B(b[11]), .Z(n517) );
  AND U689 ( .A(n516), .B(n517), .Z(n830) );
  XOR U690 ( .A(a[14]), .B(b[14]), .Z(n518) );
  NANDN U691 ( .A(n874), .B(n518), .Z(n519) );
  NAND U692 ( .A(a[14]), .B(b[14]), .Z(n520) );
  AND U693 ( .A(n519), .B(n520), .Z(n896) );
  XOR U694 ( .A(a[17]), .B(b[17]), .Z(n521) );
  NANDN U695 ( .A(n940), .B(n521), .Z(n522) );
  NAND U696 ( .A(a[17]), .B(b[17]), .Z(n523) );
  AND U697 ( .A(n522), .B(n523), .Z(n962) );
  XOR U698 ( .A(a[20]), .B(b[20]), .Z(n524) );
  NANDN U699 ( .A(n1008), .B(n524), .Z(n525) );
  NAND U700 ( .A(a[20]), .B(b[20]), .Z(n526) );
  AND U701 ( .A(n525), .B(n526), .Z(n1030) );
  XOR U702 ( .A(a[23]), .B(b[23]), .Z(n527) );
  NANDN U703 ( .A(n1074), .B(n527), .Z(n528) );
  NAND U704 ( .A(a[23]), .B(b[23]), .Z(n529) );
  AND U705 ( .A(n528), .B(n529), .Z(n1096) );
  XOR U706 ( .A(a[26]), .B(b[26]), .Z(n530) );
  NANDN U707 ( .A(n1111), .B(n530), .Z(n531) );
  NAND U708 ( .A(a[26]), .B(b[26]), .Z(n532) );
  AND U709 ( .A(n531), .B(n532), .Z(n1113) );
  XOR U710 ( .A(a[29]), .B(b[29]), .Z(n533) );
  NANDN U711 ( .A(n1117), .B(n533), .Z(n534) );
  NAND U712 ( .A(a[29]), .B(b[29]), .Z(n535) );
  AND U713 ( .A(n534), .B(n535), .Z(n1121) );
  XOR U714 ( .A(a[32]), .B(b[32]), .Z(n536) );
  NANDN U715 ( .A(n1125), .B(n536), .Z(n537) );
  NAND U716 ( .A(a[32]), .B(b[32]), .Z(n538) );
  AND U717 ( .A(n537), .B(n538), .Z(n1127) );
  XOR U718 ( .A(a[35]), .B(b[35]), .Z(n539) );
  NANDN U719 ( .A(n1131), .B(n539), .Z(n540) );
  NAND U720 ( .A(a[35]), .B(b[35]), .Z(n541) );
  AND U721 ( .A(n540), .B(n541), .Z(n1133) );
  XOR U722 ( .A(a[38]), .B(b[38]), .Z(n542) );
  NANDN U723 ( .A(n1137), .B(n542), .Z(n543) );
  NAND U724 ( .A(a[38]), .B(b[38]), .Z(n544) );
  AND U725 ( .A(n543), .B(n544), .Z(n1139) );
  XOR U726 ( .A(a[41]), .B(b[41]), .Z(n545) );
  NANDN U727 ( .A(n1145), .B(n545), .Z(n546) );
  NAND U728 ( .A(a[41]), .B(b[41]), .Z(n547) );
  AND U729 ( .A(n546), .B(n547), .Z(n1147) );
  XOR U730 ( .A(a[44]), .B(b[44]), .Z(n548) );
  NANDN U731 ( .A(n1151), .B(n548), .Z(n549) );
  NAND U732 ( .A(a[44]), .B(b[44]), .Z(n550) );
  AND U733 ( .A(n549), .B(n550), .Z(n1153) );
  XOR U734 ( .A(a[47]), .B(b[47]), .Z(n551) );
  NANDN U735 ( .A(n1157), .B(n551), .Z(n552) );
  NAND U736 ( .A(a[47]), .B(b[47]), .Z(n553) );
  AND U737 ( .A(n552), .B(n553), .Z(n1159) );
  XOR U738 ( .A(a[50]), .B(b[50]), .Z(n554) );
  NANDN U739 ( .A(n1165), .B(n554), .Z(n555) );
  NAND U740 ( .A(a[50]), .B(b[50]), .Z(n556) );
  AND U741 ( .A(n555), .B(n556), .Z(n1167) );
  XOR U742 ( .A(a[53]), .B(b[53]), .Z(n557) );
  NANDN U743 ( .A(n1171), .B(n557), .Z(n558) );
  NAND U744 ( .A(a[53]), .B(b[53]), .Z(n559) );
  AND U745 ( .A(n558), .B(n559), .Z(n1173) );
  XOR U746 ( .A(a[56]), .B(b[56]), .Z(n560) );
  NANDN U747 ( .A(n1177), .B(n560), .Z(n561) );
  NAND U748 ( .A(a[56]), .B(b[56]), .Z(n562) );
  AND U749 ( .A(n561), .B(n562), .Z(n1179) );
  XOR U750 ( .A(a[59]), .B(b[59]), .Z(n563) );
  NANDN U751 ( .A(n1183), .B(n563), .Z(n564) );
  NAND U752 ( .A(a[59]), .B(b[59]), .Z(n565) );
  AND U753 ( .A(n564), .B(n565), .Z(n1187) );
  XOR U754 ( .A(a[62]), .B(b[62]), .Z(n566) );
  NANDN U755 ( .A(n1191), .B(n566), .Z(n567) );
  NAND U756 ( .A(a[62]), .B(b[62]), .Z(n568) );
  AND U757 ( .A(n567), .B(n568), .Z(n1193) );
  XOR U758 ( .A(a[65]), .B(b[65]), .Z(n569) );
  NANDN U759 ( .A(n1197), .B(n569), .Z(n570) );
  NAND U760 ( .A(a[65]), .B(b[65]), .Z(n571) );
  AND U761 ( .A(n570), .B(n571), .Z(n1199) );
  XOR U762 ( .A(a[68]), .B(b[68]), .Z(n572) );
  NANDN U763 ( .A(n1203), .B(n572), .Z(n573) );
  NAND U764 ( .A(a[68]), .B(b[68]), .Z(n574) );
  AND U765 ( .A(n573), .B(n574), .Z(n1205) );
  XOR U766 ( .A(a[71]), .B(b[71]), .Z(n575) );
  NANDN U767 ( .A(n1211), .B(n575), .Z(n576) );
  NAND U768 ( .A(a[71]), .B(b[71]), .Z(n577) );
  AND U769 ( .A(n576), .B(n577), .Z(n1213) );
  XOR U770 ( .A(a[74]), .B(b[74]), .Z(n578) );
  NANDN U771 ( .A(n1217), .B(n578), .Z(n579) );
  NAND U772 ( .A(a[74]), .B(b[74]), .Z(n580) );
  AND U773 ( .A(n579), .B(n580), .Z(n1219) );
  XOR U774 ( .A(a[77]), .B(b[77]), .Z(n581) );
  NANDN U775 ( .A(n1223), .B(n581), .Z(n582) );
  NAND U776 ( .A(a[77]), .B(b[77]), .Z(n583) );
  AND U777 ( .A(n582), .B(n583), .Z(n1225) );
  XOR U778 ( .A(a[80]), .B(b[80]), .Z(n584) );
  NANDN U779 ( .A(n1231), .B(n584), .Z(n585) );
  NAND U780 ( .A(a[80]), .B(b[80]), .Z(n586) );
  AND U781 ( .A(n585), .B(n586), .Z(n1233) );
  XOR U782 ( .A(a[83]), .B(b[83]), .Z(n587) );
  NANDN U783 ( .A(n1237), .B(n587), .Z(n588) );
  NAND U784 ( .A(a[83]), .B(b[83]), .Z(n589) );
  AND U785 ( .A(n588), .B(n589), .Z(n1239) );
  XOR U786 ( .A(a[86]), .B(b[86]), .Z(n590) );
  NANDN U787 ( .A(n1243), .B(n590), .Z(n591) );
  NAND U788 ( .A(a[86]), .B(b[86]), .Z(n592) );
  AND U789 ( .A(n591), .B(n592), .Z(n1245) );
  XOR U790 ( .A(a[89]), .B(b[89]), .Z(n593) );
  NANDN U791 ( .A(n1249), .B(n593), .Z(n594) );
  NAND U792 ( .A(a[89]), .B(b[89]), .Z(n595) );
  AND U793 ( .A(n594), .B(n595), .Z(n1253) );
  XOR U794 ( .A(a[92]), .B(b[92]), .Z(n596) );
  NANDN U795 ( .A(n1257), .B(n596), .Z(n597) );
  NAND U796 ( .A(a[92]), .B(b[92]), .Z(n598) );
  AND U797 ( .A(n597), .B(n598), .Z(n1259) );
  XOR U798 ( .A(a[95]), .B(b[95]), .Z(n599) );
  NANDN U799 ( .A(n1263), .B(n599), .Z(n600) );
  NAND U800 ( .A(a[95]), .B(b[95]), .Z(n601) );
  AND U801 ( .A(n600), .B(n601), .Z(n1265) );
  XOR U802 ( .A(a[98]), .B(b[98]), .Z(n602) );
  NANDN U803 ( .A(n1269), .B(n602), .Z(n603) );
  NAND U804 ( .A(a[98]), .B(b[98]), .Z(n604) );
  AND U805 ( .A(n603), .B(n604), .Z(n1271) );
  XOR U806 ( .A(b[101]), .B(a[101]), .Z(n605) );
  NANDN U807 ( .A(n770), .B(n605), .Z(n606) );
  NAND U808 ( .A(b[101]), .B(a[101]), .Z(n607) );
  AND U809 ( .A(n606), .B(n607), .Z(n772) );
  XOR U810 ( .A(b[104]), .B(a[104]), .Z(n608) );
  NANDN U811 ( .A(n776), .B(n608), .Z(n609) );
  NAND U812 ( .A(b[104]), .B(a[104]), .Z(n610) );
  AND U813 ( .A(n609), .B(n610), .Z(n778) );
  XOR U814 ( .A(b[107]), .B(a[107]), .Z(n611) );
  NANDN U815 ( .A(n782), .B(n611), .Z(n612) );
  NAND U816 ( .A(b[107]), .B(a[107]), .Z(n613) );
  AND U817 ( .A(n612), .B(n613), .Z(n784) );
  XOR U818 ( .A(b[110]), .B(a[110]), .Z(n614) );
  NANDN U819 ( .A(n790), .B(n614), .Z(n615) );
  NAND U820 ( .A(b[110]), .B(a[110]), .Z(n616) );
  AND U821 ( .A(n615), .B(n616), .Z(n792) );
  XOR U822 ( .A(b[113]), .B(a[113]), .Z(n617) );
  NANDN U823 ( .A(n796), .B(n617), .Z(n618) );
  NAND U824 ( .A(b[113]), .B(a[113]), .Z(n619) );
  AND U825 ( .A(n618), .B(n619), .Z(n798) );
  XOR U826 ( .A(b[116]), .B(a[116]), .Z(n620) );
  NANDN U827 ( .A(n802), .B(n620), .Z(n621) );
  NAND U828 ( .A(b[116]), .B(a[116]), .Z(n622) );
  AND U829 ( .A(n621), .B(n622), .Z(n804) );
  XOR U830 ( .A(b[119]), .B(a[119]), .Z(n623) );
  NANDN U831 ( .A(n810), .B(n623), .Z(n624) );
  NAND U832 ( .A(b[119]), .B(a[119]), .Z(n625) );
  AND U833 ( .A(n624), .B(n625), .Z(n812) );
  XOR U834 ( .A(b[122]), .B(a[122]), .Z(n626) );
  NANDN U835 ( .A(n816), .B(n626), .Z(n627) );
  NAND U836 ( .A(b[122]), .B(a[122]), .Z(n628) );
  AND U837 ( .A(n627), .B(n628), .Z(n818) );
  XOR U838 ( .A(b[125]), .B(a[125]), .Z(n629) );
  NANDN U839 ( .A(n822), .B(n629), .Z(n630) );
  NAND U840 ( .A(b[125]), .B(a[125]), .Z(n631) );
  AND U841 ( .A(n630), .B(n631), .Z(n824) );
  XOR U842 ( .A(b[128]), .B(a[128]), .Z(n632) );
  NANDN U843 ( .A(n828), .B(n632), .Z(n633) );
  NAND U844 ( .A(b[128]), .B(a[128]), .Z(n634) );
  AND U845 ( .A(n633), .B(n634), .Z(n832) );
  XOR U846 ( .A(b[131]), .B(a[131]), .Z(n635) );
  NANDN U847 ( .A(n836), .B(n635), .Z(n636) );
  NAND U848 ( .A(b[131]), .B(a[131]), .Z(n637) );
  AND U849 ( .A(n636), .B(n637), .Z(n838) );
  XOR U850 ( .A(b[134]), .B(a[134]), .Z(n638) );
  NANDN U851 ( .A(n842), .B(n638), .Z(n639) );
  NAND U852 ( .A(b[134]), .B(a[134]), .Z(n640) );
  AND U853 ( .A(n639), .B(n640), .Z(n844) );
  XOR U854 ( .A(b[137]), .B(a[137]), .Z(n641) );
  NANDN U855 ( .A(n848), .B(n641), .Z(n642) );
  NAND U856 ( .A(b[137]), .B(a[137]), .Z(n643) );
  AND U857 ( .A(n642), .B(n643), .Z(n850) );
  XOR U858 ( .A(b[140]), .B(a[140]), .Z(n644) );
  NANDN U859 ( .A(n856), .B(n644), .Z(n645) );
  NAND U860 ( .A(b[140]), .B(a[140]), .Z(n646) );
  AND U861 ( .A(n645), .B(n646), .Z(n858) );
  XOR U862 ( .A(b[143]), .B(a[143]), .Z(n647) );
  NANDN U863 ( .A(n862), .B(n647), .Z(n648) );
  NAND U864 ( .A(b[143]), .B(a[143]), .Z(n649) );
  AND U865 ( .A(n648), .B(n649), .Z(n864) );
  XOR U866 ( .A(b[146]), .B(a[146]), .Z(n650) );
  NANDN U867 ( .A(n868), .B(n650), .Z(n651) );
  NAND U868 ( .A(b[146]), .B(a[146]), .Z(n652) );
  AND U869 ( .A(n651), .B(n652), .Z(n870) );
  XOR U870 ( .A(b[149]), .B(a[149]), .Z(n653) );
  NANDN U871 ( .A(n876), .B(n653), .Z(n654) );
  NAND U872 ( .A(b[149]), .B(a[149]), .Z(n655) );
  AND U873 ( .A(n654), .B(n655), .Z(n878) );
  XOR U874 ( .A(b[152]), .B(a[152]), .Z(n656) );
  NANDN U875 ( .A(n882), .B(n656), .Z(n657) );
  NAND U876 ( .A(b[152]), .B(a[152]), .Z(n658) );
  AND U877 ( .A(n657), .B(n658), .Z(n884) );
  XOR U878 ( .A(b[155]), .B(a[155]), .Z(n659) );
  NANDN U879 ( .A(n888), .B(n659), .Z(n660) );
  NAND U880 ( .A(b[155]), .B(a[155]), .Z(n661) );
  AND U881 ( .A(n660), .B(n661), .Z(n890) );
  XOR U882 ( .A(b[158]), .B(a[158]), .Z(n662) );
  NANDN U883 ( .A(n894), .B(n662), .Z(n663) );
  NAND U884 ( .A(b[158]), .B(a[158]), .Z(n664) );
  AND U885 ( .A(n663), .B(n664), .Z(n898) );
  XOR U886 ( .A(b[161]), .B(a[161]), .Z(n665) );
  NANDN U887 ( .A(n902), .B(n665), .Z(n666) );
  NAND U888 ( .A(b[161]), .B(a[161]), .Z(n667) );
  AND U889 ( .A(n666), .B(n667), .Z(n904) );
  XOR U890 ( .A(b[164]), .B(a[164]), .Z(n668) );
  NANDN U891 ( .A(n908), .B(n668), .Z(n669) );
  NAND U892 ( .A(b[164]), .B(a[164]), .Z(n670) );
  AND U893 ( .A(n669), .B(n670), .Z(n910) );
  XOR U894 ( .A(b[167]), .B(a[167]), .Z(n671) );
  NANDN U895 ( .A(n914), .B(n671), .Z(n672) );
  NAND U896 ( .A(b[167]), .B(a[167]), .Z(n673) );
  AND U897 ( .A(n672), .B(n673), .Z(n916) );
  XOR U898 ( .A(b[170]), .B(a[170]), .Z(n674) );
  NANDN U899 ( .A(n922), .B(n674), .Z(n675) );
  NAND U900 ( .A(b[170]), .B(a[170]), .Z(n676) );
  AND U901 ( .A(n675), .B(n676), .Z(n924) );
  XOR U902 ( .A(b[173]), .B(a[173]), .Z(n677) );
  NANDN U903 ( .A(n928), .B(n677), .Z(n678) );
  NAND U904 ( .A(b[173]), .B(a[173]), .Z(n679) );
  AND U905 ( .A(n678), .B(n679), .Z(n930) );
  XOR U906 ( .A(b[176]), .B(a[176]), .Z(n680) );
  NANDN U907 ( .A(n934), .B(n680), .Z(n681) );
  NAND U908 ( .A(b[176]), .B(a[176]), .Z(n682) );
  AND U909 ( .A(n681), .B(n682), .Z(n936) );
  XOR U910 ( .A(b[179]), .B(a[179]), .Z(n683) );
  NANDN U911 ( .A(n942), .B(n683), .Z(n684) );
  NAND U912 ( .A(b[179]), .B(a[179]), .Z(n685) );
  AND U913 ( .A(n684), .B(n685), .Z(n944) );
  XOR U914 ( .A(b[182]), .B(a[182]), .Z(n686) );
  NANDN U915 ( .A(n948), .B(n686), .Z(n687) );
  NAND U916 ( .A(b[182]), .B(a[182]), .Z(n688) );
  AND U917 ( .A(n687), .B(n688), .Z(n950) );
  XOR U918 ( .A(b[185]), .B(a[185]), .Z(n689) );
  NANDN U919 ( .A(n954), .B(n689), .Z(n690) );
  NAND U920 ( .A(b[185]), .B(a[185]), .Z(n691) );
  AND U921 ( .A(n690), .B(n691), .Z(n956) );
  XOR U922 ( .A(b[188]), .B(a[188]), .Z(n692) );
  NANDN U923 ( .A(n960), .B(n692), .Z(n693) );
  NAND U924 ( .A(b[188]), .B(a[188]), .Z(n694) );
  AND U925 ( .A(n693), .B(n694), .Z(n964) );
  XOR U926 ( .A(b[191]), .B(a[191]), .Z(n695) );
  NANDN U927 ( .A(n968), .B(n695), .Z(n696) );
  NAND U928 ( .A(b[191]), .B(a[191]), .Z(n697) );
  AND U929 ( .A(n696), .B(n697), .Z(n970) );
  XOR U930 ( .A(b[194]), .B(a[194]), .Z(n698) );
  NANDN U931 ( .A(n974), .B(n698), .Z(n699) );
  NAND U932 ( .A(b[194]), .B(a[194]), .Z(n700) );
  AND U933 ( .A(n699), .B(n700), .Z(n976) );
  XOR U934 ( .A(b[197]), .B(a[197]), .Z(n701) );
  NANDN U935 ( .A(n980), .B(n701), .Z(n702) );
  NAND U936 ( .A(b[197]), .B(a[197]), .Z(n703) );
  AND U937 ( .A(n702), .B(n703), .Z(n982) );
  XOR U938 ( .A(b[200]), .B(a[200]), .Z(n704) );
  NANDN U939 ( .A(n990), .B(n704), .Z(n705) );
  NAND U940 ( .A(b[200]), .B(a[200]), .Z(n706) );
  AND U941 ( .A(n705), .B(n706), .Z(n992) );
  XOR U942 ( .A(b[203]), .B(a[203]), .Z(n707) );
  NANDN U943 ( .A(n996), .B(n707), .Z(n708) );
  NAND U944 ( .A(b[203]), .B(a[203]), .Z(n709) );
  AND U945 ( .A(n708), .B(n709), .Z(n998) );
  XOR U946 ( .A(b[206]), .B(a[206]), .Z(n710) );
  NANDN U947 ( .A(n1002), .B(n710), .Z(n711) );
  NAND U948 ( .A(b[206]), .B(a[206]), .Z(n712) );
  AND U949 ( .A(n711), .B(n712), .Z(n1004) );
  XOR U950 ( .A(b[209]), .B(a[209]), .Z(n713) );
  NANDN U951 ( .A(n1010), .B(n713), .Z(n714) );
  NAND U952 ( .A(b[209]), .B(a[209]), .Z(n715) );
  AND U953 ( .A(n714), .B(n715), .Z(n1012) );
  XOR U954 ( .A(b[212]), .B(a[212]), .Z(n716) );
  NANDN U955 ( .A(n1016), .B(n716), .Z(n717) );
  NAND U956 ( .A(b[212]), .B(a[212]), .Z(n718) );
  AND U957 ( .A(n717), .B(n718), .Z(n1018) );
  XOR U958 ( .A(b[215]), .B(a[215]), .Z(n719) );
  NANDN U959 ( .A(n1022), .B(n719), .Z(n720) );
  NAND U960 ( .A(b[215]), .B(a[215]), .Z(n721) );
  AND U961 ( .A(n720), .B(n721), .Z(n1024) );
  XOR U962 ( .A(b[218]), .B(a[218]), .Z(n722) );
  NANDN U963 ( .A(n1028), .B(n722), .Z(n723) );
  NAND U964 ( .A(b[218]), .B(a[218]), .Z(n724) );
  AND U965 ( .A(n723), .B(n724), .Z(n1032) );
  XOR U966 ( .A(b[221]), .B(a[221]), .Z(n725) );
  NANDN U967 ( .A(n1036), .B(n725), .Z(n726) );
  NAND U968 ( .A(b[221]), .B(a[221]), .Z(n727) );
  AND U969 ( .A(n726), .B(n727), .Z(n1038) );
  XOR U970 ( .A(b[224]), .B(a[224]), .Z(n728) );
  NANDN U971 ( .A(n1042), .B(n728), .Z(n729) );
  NAND U972 ( .A(b[224]), .B(a[224]), .Z(n730) );
  AND U973 ( .A(n729), .B(n730), .Z(n1044) );
  XOR U974 ( .A(b[227]), .B(a[227]), .Z(n731) );
  NANDN U975 ( .A(n1048), .B(n731), .Z(n732) );
  NAND U976 ( .A(b[227]), .B(a[227]), .Z(n733) );
  AND U977 ( .A(n732), .B(n733), .Z(n1050) );
  XOR U978 ( .A(b[230]), .B(a[230]), .Z(n734) );
  NANDN U979 ( .A(n1056), .B(n734), .Z(n735) );
  NAND U980 ( .A(b[230]), .B(a[230]), .Z(n736) );
  AND U981 ( .A(n735), .B(n736), .Z(n1058) );
  XOR U982 ( .A(b[233]), .B(a[233]), .Z(n737) );
  NANDN U983 ( .A(n1062), .B(n737), .Z(n738) );
  NAND U984 ( .A(b[233]), .B(a[233]), .Z(n739) );
  AND U985 ( .A(n738), .B(n739), .Z(n1064) );
  XOR U986 ( .A(b[236]), .B(a[236]), .Z(n740) );
  NANDN U987 ( .A(n1068), .B(n740), .Z(n741) );
  NAND U988 ( .A(b[236]), .B(a[236]), .Z(n742) );
  AND U989 ( .A(n741), .B(n742), .Z(n1070) );
  XOR U990 ( .A(b[239]), .B(a[239]), .Z(n743) );
  NANDN U991 ( .A(n1076), .B(n743), .Z(n744) );
  NAND U992 ( .A(b[239]), .B(a[239]), .Z(n745) );
  AND U993 ( .A(n744), .B(n745), .Z(n1078) );
  XOR U994 ( .A(b[242]), .B(a[242]), .Z(n746) );
  NANDN U995 ( .A(n1082), .B(n746), .Z(n747) );
  NAND U996 ( .A(b[242]), .B(a[242]), .Z(n748) );
  AND U997 ( .A(n747), .B(n748), .Z(n1084) );
  XOR U998 ( .A(b[245]), .B(a[245]), .Z(n749) );
  NANDN U999 ( .A(n1088), .B(n749), .Z(n750) );
  NAND U1000 ( .A(b[245]), .B(a[245]), .Z(n751) );
  AND U1001 ( .A(n750), .B(n751), .Z(n1090) );
  XOR U1002 ( .A(b[248]), .B(a[248]), .Z(n752) );
  NANDN U1003 ( .A(n1094), .B(n752), .Z(n753) );
  NAND U1004 ( .A(b[248]), .B(a[248]), .Z(n754) );
  AND U1005 ( .A(n753), .B(n754), .Z(n1098) );
  XOR U1006 ( .A(b[251]), .B(a[251]), .Z(n755) );
  NANDN U1007 ( .A(n1102), .B(n755), .Z(n756) );
  NAND U1008 ( .A(b[251]), .B(a[251]), .Z(n757) );
  AND U1009 ( .A(n756), .B(n757), .Z(n1104) );
  NANDN U1010 ( .A(n1108), .B(b[254]), .Z(n758) );
  XNOR U1011 ( .A(n1108), .B(b[254]), .Z(n759) );
  NAND U1012 ( .A(a[254]), .B(n759), .Z(n760) );
  NAND U1013 ( .A(n758), .B(n760), .Z(n761) );
  XNOR U1014 ( .A(a[255]), .B(n761), .Z(n762) );
  XNOR U1015 ( .A(b[255]), .B(n762), .Z(c[255]) );
  XOR U1016 ( .A(a[0]), .B(b[0]), .Z(c[0]) );
  NAND U1017 ( .A(a[0]), .B(b[0]), .Z(n987) );
  IV U1018 ( .A(n763), .Z(n1110) );
  NAND U1019 ( .A(n1110), .B(b[25]), .Z(n766) );
  ANDN U1020 ( .B(n763), .A(b[25]), .Z(n764) );
  NANDN U1021 ( .A(n764), .B(a[25]), .Z(n765) );
  AND U1022 ( .A(n766), .B(n765), .Z(n1111) );
  XOR U1023 ( .A(a[100]), .B(n768), .Z(n767) );
  XNOR U1024 ( .A(b[100]), .B(n767), .Z(c[100]) );
  XOR U1025 ( .A(a[101]), .B(n770), .Z(n769) );
  XNOR U1026 ( .A(b[101]), .B(n769), .Z(c[101]) );
  XOR U1027 ( .A(a[102]), .B(n772), .Z(n771) );
  XNOR U1028 ( .A(b[102]), .B(n771), .Z(c[102]) );
  XOR U1029 ( .A(a[103]), .B(n774), .Z(n773) );
  XNOR U1030 ( .A(b[103]), .B(n773), .Z(c[103]) );
  XOR U1031 ( .A(a[104]), .B(n776), .Z(n775) );
  XNOR U1032 ( .A(b[104]), .B(n775), .Z(c[104]) );
  XOR U1033 ( .A(a[105]), .B(n778), .Z(n777) );
  XNOR U1034 ( .A(b[105]), .B(n777), .Z(c[105]) );
  XOR U1035 ( .A(a[106]), .B(n780), .Z(n779) );
  XNOR U1036 ( .A(b[106]), .B(n779), .Z(c[106]) );
  XOR U1037 ( .A(a[107]), .B(n782), .Z(n781) );
  XNOR U1038 ( .A(b[107]), .B(n781), .Z(c[107]) );
  XOR U1039 ( .A(a[108]), .B(n784), .Z(n783) );
  XNOR U1040 ( .A(b[108]), .B(n783), .Z(c[108]) );
  XOR U1041 ( .A(a[109]), .B(n788), .Z(n785) );
  XNOR U1042 ( .A(b[109]), .B(n785), .Z(c[109]) );
  XOR U1043 ( .A(b[10]), .B(n786), .Z(n787) );
  XNOR U1044 ( .A(a[10]), .B(n787), .Z(c[10]) );
  XOR U1045 ( .A(a[110]), .B(n790), .Z(n789) );
  XNOR U1046 ( .A(b[110]), .B(n789), .Z(c[110]) );
  XOR U1047 ( .A(a[111]), .B(n792), .Z(n791) );
  XNOR U1048 ( .A(b[111]), .B(n791), .Z(c[111]) );
  XOR U1049 ( .A(a[112]), .B(n794), .Z(n793) );
  XNOR U1050 ( .A(b[112]), .B(n793), .Z(c[112]) );
  XOR U1051 ( .A(a[113]), .B(n796), .Z(n795) );
  XNOR U1052 ( .A(b[113]), .B(n795), .Z(c[113]) );
  XOR U1053 ( .A(a[114]), .B(n798), .Z(n797) );
  XNOR U1054 ( .A(b[114]), .B(n797), .Z(c[114]) );
  XOR U1055 ( .A(a[115]), .B(n800), .Z(n799) );
  XNOR U1056 ( .A(b[115]), .B(n799), .Z(c[115]) );
  XOR U1057 ( .A(a[116]), .B(n802), .Z(n801) );
  XNOR U1058 ( .A(b[116]), .B(n801), .Z(c[116]) );
  XOR U1059 ( .A(a[117]), .B(n804), .Z(n803) );
  XNOR U1060 ( .A(b[117]), .B(n803), .Z(c[117]) );
  XOR U1061 ( .A(a[118]), .B(n806), .Z(n805) );
  XNOR U1062 ( .A(b[118]), .B(n805), .Z(c[118]) );
  XOR U1063 ( .A(a[119]), .B(n810), .Z(n807) );
  XNOR U1064 ( .A(b[119]), .B(n807), .Z(c[119]) );
  XOR U1065 ( .A(b[11]), .B(n808), .Z(n809) );
  XNOR U1066 ( .A(a[11]), .B(n809), .Z(c[11]) );
  XOR U1067 ( .A(a[120]), .B(n812), .Z(n811) );
  XNOR U1068 ( .A(b[120]), .B(n811), .Z(c[120]) );
  XOR U1069 ( .A(a[121]), .B(n814), .Z(n813) );
  XNOR U1070 ( .A(b[121]), .B(n813), .Z(c[121]) );
  XOR U1071 ( .A(a[122]), .B(n816), .Z(n815) );
  XNOR U1072 ( .A(b[122]), .B(n815), .Z(c[122]) );
  XOR U1073 ( .A(a[123]), .B(n818), .Z(n817) );
  XNOR U1074 ( .A(b[123]), .B(n817), .Z(c[123]) );
  XOR U1075 ( .A(a[124]), .B(n820), .Z(n819) );
  XNOR U1076 ( .A(b[124]), .B(n819), .Z(c[124]) );
  XOR U1077 ( .A(a[125]), .B(n822), .Z(n821) );
  XNOR U1078 ( .A(b[125]), .B(n821), .Z(c[125]) );
  XOR U1079 ( .A(a[126]), .B(n824), .Z(n823) );
  XNOR U1080 ( .A(b[126]), .B(n823), .Z(c[126]) );
  XOR U1081 ( .A(a[127]), .B(n826), .Z(n825) );
  XNOR U1082 ( .A(b[127]), .B(n825), .Z(c[127]) );
  XOR U1083 ( .A(a[128]), .B(n828), .Z(n827) );
  XNOR U1084 ( .A(b[128]), .B(n827), .Z(c[128]) );
  XOR U1085 ( .A(a[129]), .B(n832), .Z(n829) );
  XNOR U1086 ( .A(b[129]), .B(n829), .Z(c[129]) );
  XOR U1087 ( .A(b[12]), .B(n830), .Z(n831) );
  XNOR U1088 ( .A(a[12]), .B(n831), .Z(c[12]) );
  XOR U1089 ( .A(a[130]), .B(n834), .Z(n833) );
  XNOR U1090 ( .A(b[130]), .B(n833), .Z(c[130]) );
  XOR U1091 ( .A(a[131]), .B(n836), .Z(n835) );
  XNOR U1092 ( .A(b[131]), .B(n835), .Z(c[131]) );
  XOR U1093 ( .A(a[132]), .B(n838), .Z(n837) );
  XNOR U1094 ( .A(b[132]), .B(n837), .Z(c[132]) );
  XOR U1095 ( .A(a[133]), .B(n840), .Z(n839) );
  XNOR U1096 ( .A(b[133]), .B(n839), .Z(c[133]) );
  XOR U1097 ( .A(a[134]), .B(n842), .Z(n841) );
  XNOR U1098 ( .A(b[134]), .B(n841), .Z(c[134]) );
  XOR U1099 ( .A(a[135]), .B(n844), .Z(n843) );
  XNOR U1100 ( .A(b[135]), .B(n843), .Z(c[135]) );
  XOR U1101 ( .A(a[136]), .B(n846), .Z(n845) );
  XNOR U1102 ( .A(b[136]), .B(n845), .Z(c[136]) );
  XOR U1103 ( .A(a[137]), .B(n848), .Z(n847) );
  XNOR U1104 ( .A(b[137]), .B(n847), .Z(c[137]) );
  XOR U1105 ( .A(a[138]), .B(n850), .Z(n849) );
  XNOR U1106 ( .A(b[138]), .B(n849), .Z(c[138]) );
  XOR U1107 ( .A(a[139]), .B(n854), .Z(n851) );
  XNOR U1108 ( .A(b[139]), .B(n851), .Z(c[139]) );
  XOR U1109 ( .A(b[13]), .B(n852), .Z(n853) );
  XNOR U1110 ( .A(a[13]), .B(n853), .Z(c[13]) );
  XOR U1111 ( .A(a[140]), .B(n856), .Z(n855) );
  XNOR U1112 ( .A(b[140]), .B(n855), .Z(c[140]) );
  XOR U1113 ( .A(a[141]), .B(n858), .Z(n857) );
  XNOR U1114 ( .A(b[141]), .B(n857), .Z(c[141]) );
  XOR U1115 ( .A(a[142]), .B(n860), .Z(n859) );
  XNOR U1116 ( .A(b[142]), .B(n859), .Z(c[142]) );
  XOR U1117 ( .A(a[143]), .B(n862), .Z(n861) );
  XNOR U1118 ( .A(b[143]), .B(n861), .Z(c[143]) );
  XOR U1119 ( .A(a[144]), .B(n864), .Z(n863) );
  XNOR U1120 ( .A(b[144]), .B(n863), .Z(c[144]) );
  XOR U1121 ( .A(a[145]), .B(n866), .Z(n865) );
  XNOR U1122 ( .A(b[145]), .B(n865), .Z(c[145]) );
  XOR U1123 ( .A(a[146]), .B(n868), .Z(n867) );
  XNOR U1124 ( .A(b[146]), .B(n867), .Z(c[146]) );
  XOR U1125 ( .A(a[147]), .B(n870), .Z(n869) );
  XNOR U1126 ( .A(b[147]), .B(n869), .Z(c[147]) );
  XOR U1127 ( .A(a[148]), .B(n872), .Z(n871) );
  XNOR U1128 ( .A(b[148]), .B(n871), .Z(c[148]) );
  XOR U1129 ( .A(a[149]), .B(n876), .Z(n873) );
  XNOR U1130 ( .A(b[149]), .B(n873), .Z(c[149]) );
  XOR U1131 ( .A(b[14]), .B(n874), .Z(n875) );
  XNOR U1132 ( .A(a[14]), .B(n875), .Z(c[14]) );
  XOR U1133 ( .A(a[150]), .B(n878), .Z(n877) );
  XNOR U1134 ( .A(b[150]), .B(n877), .Z(c[150]) );
  XOR U1135 ( .A(a[151]), .B(n880), .Z(n879) );
  XNOR U1136 ( .A(b[151]), .B(n879), .Z(c[151]) );
  XOR U1137 ( .A(a[152]), .B(n882), .Z(n881) );
  XNOR U1138 ( .A(b[152]), .B(n881), .Z(c[152]) );
  XOR U1139 ( .A(a[153]), .B(n884), .Z(n883) );
  XNOR U1140 ( .A(b[153]), .B(n883), .Z(c[153]) );
  XOR U1141 ( .A(a[154]), .B(n886), .Z(n885) );
  XNOR U1142 ( .A(b[154]), .B(n885), .Z(c[154]) );
  XOR U1143 ( .A(a[155]), .B(n888), .Z(n887) );
  XNOR U1144 ( .A(b[155]), .B(n887), .Z(c[155]) );
  XOR U1145 ( .A(a[156]), .B(n890), .Z(n889) );
  XNOR U1146 ( .A(b[156]), .B(n889), .Z(c[156]) );
  XOR U1147 ( .A(a[157]), .B(n892), .Z(n891) );
  XNOR U1148 ( .A(b[157]), .B(n891), .Z(c[157]) );
  XOR U1149 ( .A(a[158]), .B(n894), .Z(n893) );
  XNOR U1150 ( .A(b[158]), .B(n893), .Z(c[158]) );
  XOR U1151 ( .A(a[159]), .B(n898), .Z(n895) );
  XNOR U1152 ( .A(b[159]), .B(n895), .Z(c[159]) );
  XOR U1153 ( .A(b[15]), .B(n896), .Z(n897) );
  XNOR U1154 ( .A(a[15]), .B(n897), .Z(c[15]) );
  XOR U1155 ( .A(a[160]), .B(n900), .Z(n899) );
  XNOR U1156 ( .A(b[160]), .B(n899), .Z(c[160]) );
  XOR U1157 ( .A(a[161]), .B(n902), .Z(n901) );
  XNOR U1158 ( .A(b[161]), .B(n901), .Z(c[161]) );
  XOR U1159 ( .A(a[162]), .B(n904), .Z(n903) );
  XNOR U1160 ( .A(b[162]), .B(n903), .Z(c[162]) );
  XOR U1161 ( .A(a[163]), .B(n906), .Z(n905) );
  XNOR U1162 ( .A(b[163]), .B(n905), .Z(c[163]) );
  XOR U1163 ( .A(a[164]), .B(n908), .Z(n907) );
  XNOR U1164 ( .A(b[164]), .B(n907), .Z(c[164]) );
  XOR U1165 ( .A(a[165]), .B(n910), .Z(n909) );
  XNOR U1166 ( .A(b[165]), .B(n909), .Z(c[165]) );
  XOR U1167 ( .A(a[166]), .B(n912), .Z(n911) );
  XNOR U1168 ( .A(b[166]), .B(n911), .Z(c[166]) );
  XOR U1169 ( .A(a[167]), .B(n914), .Z(n913) );
  XNOR U1170 ( .A(b[167]), .B(n913), .Z(c[167]) );
  XOR U1171 ( .A(a[168]), .B(n916), .Z(n915) );
  XNOR U1172 ( .A(b[168]), .B(n915), .Z(c[168]) );
  XOR U1173 ( .A(a[169]), .B(n920), .Z(n917) );
  XNOR U1174 ( .A(b[169]), .B(n917), .Z(c[169]) );
  XOR U1175 ( .A(b[16]), .B(n918), .Z(n919) );
  XNOR U1176 ( .A(a[16]), .B(n919), .Z(c[16]) );
  XOR U1177 ( .A(a[170]), .B(n922), .Z(n921) );
  XNOR U1178 ( .A(b[170]), .B(n921), .Z(c[170]) );
  XOR U1179 ( .A(a[171]), .B(n924), .Z(n923) );
  XNOR U1180 ( .A(b[171]), .B(n923), .Z(c[171]) );
  XOR U1181 ( .A(a[172]), .B(n926), .Z(n925) );
  XNOR U1182 ( .A(b[172]), .B(n925), .Z(c[172]) );
  XOR U1183 ( .A(a[173]), .B(n928), .Z(n927) );
  XNOR U1184 ( .A(b[173]), .B(n927), .Z(c[173]) );
  XOR U1185 ( .A(a[174]), .B(n930), .Z(n929) );
  XNOR U1186 ( .A(b[174]), .B(n929), .Z(c[174]) );
  XOR U1187 ( .A(a[175]), .B(n932), .Z(n931) );
  XNOR U1188 ( .A(b[175]), .B(n931), .Z(c[175]) );
  XOR U1189 ( .A(a[176]), .B(n934), .Z(n933) );
  XNOR U1190 ( .A(b[176]), .B(n933), .Z(c[176]) );
  XOR U1191 ( .A(a[177]), .B(n936), .Z(n935) );
  XNOR U1192 ( .A(b[177]), .B(n935), .Z(c[177]) );
  XOR U1193 ( .A(a[178]), .B(n938), .Z(n937) );
  XNOR U1194 ( .A(b[178]), .B(n937), .Z(c[178]) );
  XOR U1195 ( .A(a[179]), .B(n942), .Z(n939) );
  XNOR U1196 ( .A(b[179]), .B(n939), .Z(c[179]) );
  XOR U1197 ( .A(b[17]), .B(n940), .Z(n941) );
  XNOR U1198 ( .A(a[17]), .B(n941), .Z(c[17]) );
  XOR U1199 ( .A(a[180]), .B(n944), .Z(n943) );
  XNOR U1200 ( .A(b[180]), .B(n943), .Z(c[180]) );
  XOR U1201 ( .A(a[181]), .B(n946), .Z(n945) );
  XNOR U1202 ( .A(b[181]), .B(n945), .Z(c[181]) );
  XOR U1203 ( .A(a[182]), .B(n948), .Z(n947) );
  XNOR U1204 ( .A(b[182]), .B(n947), .Z(c[182]) );
  XOR U1205 ( .A(a[183]), .B(n950), .Z(n949) );
  XNOR U1206 ( .A(b[183]), .B(n949), .Z(c[183]) );
  XOR U1207 ( .A(a[184]), .B(n952), .Z(n951) );
  XNOR U1208 ( .A(b[184]), .B(n951), .Z(c[184]) );
  XOR U1209 ( .A(a[185]), .B(n954), .Z(n953) );
  XNOR U1210 ( .A(b[185]), .B(n953), .Z(c[185]) );
  XOR U1211 ( .A(a[186]), .B(n956), .Z(n955) );
  XNOR U1212 ( .A(b[186]), .B(n955), .Z(c[186]) );
  XOR U1213 ( .A(a[187]), .B(n958), .Z(n957) );
  XNOR U1214 ( .A(b[187]), .B(n957), .Z(c[187]) );
  XOR U1215 ( .A(a[188]), .B(n960), .Z(n959) );
  XNOR U1216 ( .A(b[188]), .B(n959), .Z(c[188]) );
  XOR U1217 ( .A(a[189]), .B(n964), .Z(n961) );
  XNOR U1218 ( .A(b[189]), .B(n961), .Z(c[189]) );
  XOR U1219 ( .A(b[18]), .B(n962), .Z(n963) );
  XNOR U1220 ( .A(a[18]), .B(n963), .Z(c[18]) );
  XOR U1221 ( .A(a[190]), .B(n966), .Z(n965) );
  XNOR U1222 ( .A(b[190]), .B(n965), .Z(c[190]) );
  XOR U1223 ( .A(a[191]), .B(n968), .Z(n967) );
  XNOR U1224 ( .A(b[191]), .B(n967), .Z(c[191]) );
  XOR U1225 ( .A(a[192]), .B(n970), .Z(n969) );
  XNOR U1226 ( .A(b[192]), .B(n969), .Z(c[192]) );
  XOR U1227 ( .A(a[193]), .B(n972), .Z(n971) );
  XNOR U1228 ( .A(b[193]), .B(n971), .Z(c[193]) );
  XOR U1229 ( .A(a[194]), .B(n974), .Z(n973) );
  XNOR U1230 ( .A(b[194]), .B(n973), .Z(c[194]) );
  XOR U1231 ( .A(a[195]), .B(n976), .Z(n975) );
  XNOR U1232 ( .A(b[195]), .B(n975), .Z(c[195]) );
  XOR U1233 ( .A(a[196]), .B(n978), .Z(n977) );
  XNOR U1234 ( .A(b[196]), .B(n977), .Z(c[196]) );
  XOR U1235 ( .A(a[197]), .B(n980), .Z(n979) );
  XNOR U1236 ( .A(b[197]), .B(n979), .Z(c[197]) );
  XOR U1237 ( .A(a[198]), .B(n982), .Z(n981) );
  XNOR U1238 ( .A(b[198]), .B(n981), .Z(c[198]) );
  XOR U1239 ( .A(a[199]), .B(n988), .Z(n983) );
  XNOR U1240 ( .A(b[199]), .B(n983), .Z(c[199]) );
  XOR U1241 ( .A(b[19]), .B(n984), .Z(n985) );
  XNOR U1242 ( .A(a[19]), .B(n985), .Z(c[19]) );
  XOR U1243 ( .A(a[1]), .B(b[1]), .Z(n986) );
  XNOR U1244 ( .A(n987), .B(n986), .Z(c[1]) );
  XOR U1245 ( .A(a[200]), .B(n990), .Z(n989) );
  XNOR U1246 ( .A(b[200]), .B(n989), .Z(c[200]) );
  XOR U1247 ( .A(a[201]), .B(n992), .Z(n991) );
  XNOR U1248 ( .A(b[201]), .B(n991), .Z(c[201]) );
  XOR U1249 ( .A(a[202]), .B(n994), .Z(n993) );
  XNOR U1250 ( .A(b[202]), .B(n993), .Z(c[202]) );
  XOR U1251 ( .A(a[203]), .B(n996), .Z(n995) );
  XNOR U1252 ( .A(b[203]), .B(n995), .Z(c[203]) );
  XOR U1253 ( .A(a[204]), .B(n998), .Z(n997) );
  XNOR U1254 ( .A(b[204]), .B(n997), .Z(c[204]) );
  XOR U1255 ( .A(a[205]), .B(n1000), .Z(n999) );
  XNOR U1256 ( .A(b[205]), .B(n999), .Z(c[205]) );
  XOR U1257 ( .A(a[206]), .B(n1002), .Z(n1001) );
  XNOR U1258 ( .A(b[206]), .B(n1001), .Z(c[206]) );
  XOR U1259 ( .A(a[207]), .B(n1004), .Z(n1003) );
  XNOR U1260 ( .A(b[207]), .B(n1003), .Z(c[207]) );
  XOR U1261 ( .A(a[208]), .B(n1006), .Z(n1005) );
  XNOR U1262 ( .A(b[208]), .B(n1005), .Z(c[208]) );
  XOR U1263 ( .A(a[209]), .B(n1010), .Z(n1007) );
  XNOR U1264 ( .A(b[209]), .B(n1007), .Z(c[209]) );
  XOR U1265 ( .A(b[20]), .B(n1008), .Z(n1009) );
  XNOR U1266 ( .A(a[20]), .B(n1009), .Z(c[20]) );
  XOR U1267 ( .A(a[210]), .B(n1012), .Z(n1011) );
  XNOR U1268 ( .A(b[210]), .B(n1011), .Z(c[210]) );
  XOR U1269 ( .A(a[211]), .B(n1014), .Z(n1013) );
  XNOR U1270 ( .A(b[211]), .B(n1013), .Z(c[211]) );
  XOR U1271 ( .A(a[212]), .B(n1016), .Z(n1015) );
  XNOR U1272 ( .A(b[212]), .B(n1015), .Z(c[212]) );
  XOR U1273 ( .A(a[213]), .B(n1018), .Z(n1017) );
  XNOR U1274 ( .A(b[213]), .B(n1017), .Z(c[213]) );
  XOR U1275 ( .A(a[214]), .B(n1020), .Z(n1019) );
  XNOR U1276 ( .A(b[214]), .B(n1019), .Z(c[214]) );
  XOR U1277 ( .A(a[215]), .B(n1022), .Z(n1021) );
  XNOR U1278 ( .A(b[215]), .B(n1021), .Z(c[215]) );
  XOR U1279 ( .A(a[216]), .B(n1024), .Z(n1023) );
  XNOR U1280 ( .A(b[216]), .B(n1023), .Z(c[216]) );
  XOR U1281 ( .A(a[217]), .B(n1026), .Z(n1025) );
  XNOR U1282 ( .A(b[217]), .B(n1025), .Z(c[217]) );
  XOR U1283 ( .A(a[218]), .B(n1028), .Z(n1027) );
  XNOR U1284 ( .A(b[218]), .B(n1027), .Z(c[218]) );
  XOR U1285 ( .A(a[219]), .B(n1032), .Z(n1029) );
  XNOR U1286 ( .A(b[219]), .B(n1029), .Z(c[219]) );
  XOR U1287 ( .A(b[21]), .B(n1030), .Z(n1031) );
  XNOR U1288 ( .A(a[21]), .B(n1031), .Z(c[21]) );
  XOR U1289 ( .A(a[220]), .B(n1034), .Z(n1033) );
  XNOR U1290 ( .A(b[220]), .B(n1033), .Z(c[220]) );
  XOR U1291 ( .A(a[221]), .B(n1036), .Z(n1035) );
  XNOR U1292 ( .A(b[221]), .B(n1035), .Z(c[221]) );
  XOR U1293 ( .A(a[222]), .B(n1038), .Z(n1037) );
  XNOR U1294 ( .A(b[222]), .B(n1037), .Z(c[222]) );
  XOR U1295 ( .A(a[223]), .B(n1040), .Z(n1039) );
  XNOR U1296 ( .A(b[223]), .B(n1039), .Z(c[223]) );
  XOR U1297 ( .A(a[224]), .B(n1042), .Z(n1041) );
  XNOR U1298 ( .A(b[224]), .B(n1041), .Z(c[224]) );
  XOR U1299 ( .A(a[225]), .B(n1044), .Z(n1043) );
  XNOR U1300 ( .A(b[225]), .B(n1043), .Z(c[225]) );
  XOR U1301 ( .A(a[226]), .B(n1046), .Z(n1045) );
  XNOR U1302 ( .A(b[226]), .B(n1045), .Z(c[226]) );
  XOR U1303 ( .A(a[227]), .B(n1048), .Z(n1047) );
  XNOR U1304 ( .A(b[227]), .B(n1047), .Z(c[227]) );
  XOR U1305 ( .A(a[228]), .B(n1050), .Z(n1049) );
  XNOR U1306 ( .A(b[228]), .B(n1049), .Z(c[228]) );
  XOR U1307 ( .A(a[229]), .B(n1054), .Z(n1051) );
  XNOR U1308 ( .A(b[229]), .B(n1051), .Z(c[229]) );
  XOR U1309 ( .A(b[22]), .B(n1052), .Z(n1053) );
  XNOR U1310 ( .A(a[22]), .B(n1053), .Z(c[22]) );
  XOR U1311 ( .A(a[230]), .B(n1056), .Z(n1055) );
  XNOR U1312 ( .A(b[230]), .B(n1055), .Z(c[230]) );
  XOR U1313 ( .A(a[231]), .B(n1058), .Z(n1057) );
  XNOR U1314 ( .A(b[231]), .B(n1057), .Z(c[231]) );
  XOR U1315 ( .A(a[232]), .B(n1060), .Z(n1059) );
  XNOR U1316 ( .A(b[232]), .B(n1059), .Z(c[232]) );
  XOR U1317 ( .A(a[233]), .B(n1062), .Z(n1061) );
  XNOR U1318 ( .A(b[233]), .B(n1061), .Z(c[233]) );
  XOR U1319 ( .A(a[234]), .B(n1064), .Z(n1063) );
  XNOR U1320 ( .A(b[234]), .B(n1063), .Z(c[234]) );
  XOR U1321 ( .A(a[235]), .B(n1066), .Z(n1065) );
  XNOR U1322 ( .A(b[235]), .B(n1065), .Z(c[235]) );
  XOR U1323 ( .A(a[236]), .B(n1068), .Z(n1067) );
  XNOR U1324 ( .A(b[236]), .B(n1067), .Z(c[236]) );
  XOR U1325 ( .A(a[237]), .B(n1070), .Z(n1069) );
  XNOR U1326 ( .A(b[237]), .B(n1069), .Z(c[237]) );
  XOR U1327 ( .A(a[238]), .B(n1072), .Z(n1071) );
  XNOR U1328 ( .A(b[238]), .B(n1071), .Z(c[238]) );
  XOR U1329 ( .A(a[239]), .B(n1076), .Z(n1073) );
  XNOR U1330 ( .A(b[239]), .B(n1073), .Z(c[239]) );
  XOR U1331 ( .A(b[23]), .B(n1074), .Z(n1075) );
  XNOR U1332 ( .A(a[23]), .B(n1075), .Z(c[23]) );
  XOR U1333 ( .A(a[240]), .B(n1078), .Z(n1077) );
  XNOR U1334 ( .A(b[240]), .B(n1077), .Z(c[240]) );
  XOR U1335 ( .A(a[241]), .B(n1080), .Z(n1079) );
  XNOR U1336 ( .A(b[241]), .B(n1079), .Z(c[241]) );
  XOR U1337 ( .A(a[242]), .B(n1082), .Z(n1081) );
  XNOR U1338 ( .A(b[242]), .B(n1081), .Z(c[242]) );
  XOR U1339 ( .A(a[243]), .B(n1084), .Z(n1083) );
  XNOR U1340 ( .A(b[243]), .B(n1083), .Z(c[243]) );
  XOR U1341 ( .A(a[244]), .B(n1086), .Z(n1085) );
  XNOR U1342 ( .A(b[244]), .B(n1085), .Z(c[244]) );
  XOR U1343 ( .A(a[245]), .B(n1088), .Z(n1087) );
  XNOR U1344 ( .A(b[245]), .B(n1087), .Z(c[245]) );
  XOR U1345 ( .A(a[246]), .B(n1090), .Z(n1089) );
  XNOR U1346 ( .A(b[246]), .B(n1089), .Z(c[246]) );
  XOR U1347 ( .A(a[247]), .B(n1092), .Z(n1091) );
  XNOR U1348 ( .A(b[247]), .B(n1091), .Z(c[247]) );
  XOR U1349 ( .A(a[248]), .B(n1094), .Z(n1093) );
  XNOR U1350 ( .A(b[248]), .B(n1093), .Z(c[248]) );
  XOR U1351 ( .A(a[249]), .B(n1098), .Z(n1095) );
  XNOR U1352 ( .A(b[249]), .B(n1095), .Z(c[249]) );
  XOR U1353 ( .A(b[24]), .B(n1096), .Z(n1097) );
  XNOR U1354 ( .A(a[24]), .B(n1097), .Z(c[24]) );
  XOR U1355 ( .A(a[250]), .B(n1100), .Z(n1099) );
  XNOR U1356 ( .A(b[250]), .B(n1099), .Z(c[250]) );
  XOR U1357 ( .A(a[251]), .B(n1102), .Z(n1101) );
  XNOR U1358 ( .A(b[251]), .B(n1101), .Z(c[251]) );
  XOR U1359 ( .A(a[252]), .B(n1104), .Z(n1103) );
  XNOR U1360 ( .A(b[252]), .B(n1103), .Z(c[252]) );
  XOR U1361 ( .A(a[253]), .B(n1106), .Z(n1105) );
  XNOR U1362 ( .A(b[253]), .B(n1105), .Z(c[253]) );
  XOR U1363 ( .A(a[254]), .B(n1108), .Z(n1107) );
  XNOR U1364 ( .A(b[254]), .B(n1107), .Z(c[254]) );
  XNOR U1365 ( .A(b[25]), .B(a[25]), .Z(n1109) );
  XNOR U1366 ( .A(n1110), .B(n1109), .Z(c[25]) );
  XOR U1367 ( .A(b[26]), .B(n1111), .Z(n1112) );
  XNOR U1368 ( .A(a[26]), .B(n1112), .Z(c[26]) );
  XOR U1369 ( .A(b[27]), .B(n1113), .Z(n1114) );
  XNOR U1370 ( .A(a[27]), .B(n1114), .Z(c[27]) );
  XOR U1371 ( .A(b[28]), .B(n1115), .Z(n1116) );
  XNOR U1372 ( .A(a[28]), .B(n1116), .Z(c[28]) );
  XOR U1373 ( .A(b[29]), .B(n1117), .Z(n1118) );
  XNOR U1374 ( .A(a[29]), .B(n1118), .Z(c[29]) );
  XOR U1375 ( .A(b[2]), .B(n1119), .Z(n1120) );
  XNOR U1376 ( .A(a[2]), .B(n1120), .Z(c[2]) );
  XOR U1377 ( .A(b[30]), .B(n1121), .Z(n1122) );
  XNOR U1378 ( .A(a[30]), .B(n1122), .Z(c[30]) );
  XOR U1379 ( .A(b[31]), .B(n1123), .Z(n1124) );
  XNOR U1380 ( .A(a[31]), .B(n1124), .Z(c[31]) );
  XOR U1381 ( .A(b[32]), .B(n1125), .Z(n1126) );
  XNOR U1382 ( .A(a[32]), .B(n1126), .Z(c[32]) );
  XOR U1383 ( .A(b[33]), .B(n1127), .Z(n1128) );
  XNOR U1384 ( .A(a[33]), .B(n1128), .Z(c[33]) );
  XOR U1385 ( .A(b[34]), .B(n1129), .Z(n1130) );
  XNOR U1386 ( .A(a[34]), .B(n1130), .Z(c[34]) );
  XOR U1387 ( .A(b[35]), .B(n1131), .Z(n1132) );
  XNOR U1388 ( .A(a[35]), .B(n1132), .Z(c[35]) );
  XOR U1389 ( .A(b[36]), .B(n1133), .Z(n1134) );
  XNOR U1390 ( .A(a[36]), .B(n1134), .Z(c[36]) );
  XOR U1391 ( .A(b[37]), .B(n1135), .Z(n1136) );
  XNOR U1392 ( .A(a[37]), .B(n1136), .Z(c[37]) );
  XOR U1393 ( .A(b[38]), .B(n1137), .Z(n1138) );
  XNOR U1394 ( .A(a[38]), .B(n1138), .Z(c[38]) );
  XOR U1395 ( .A(b[39]), .B(n1139), .Z(n1140) );
  XNOR U1396 ( .A(a[39]), .B(n1140), .Z(c[39]) );
  XOR U1397 ( .A(b[3]), .B(n1141), .Z(n1142) );
  XNOR U1398 ( .A(a[3]), .B(n1142), .Z(c[3]) );
  XOR U1399 ( .A(b[40]), .B(n1143), .Z(n1144) );
  XNOR U1400 ( .A(a[40]), .B(n1144), .Z(c[40]) );
  XOR U1401 ( .A(b[41]), .B(n1145), .Z(n1146) );
  XNOR U1402 ( .A(a[41]), .B(n1146), .Z(c[41]) );
  XOR U1403 ( .A(b[42]), .B(n1147), .Z(n1148) );
  XNOR U1404 ( .A(a[42]), .B(n1148), .Z(c[42]) );
  XOR U1405 ( .A(b[43]), .B(n1149), .Z(n1150) );
  XNOR U1406 ( .A(a[43]), .B(n1150), .Z(c[43]) );
  XOR U1407 ( .A(b[44]), .B(n1151), .Z(n1152) );
  XNOR U1408 ( .A(a[44]), .B(n1152), .Z(c[44]) );
  XOR U1409 ( .A(b[45]), .B(n1153), .Z(n1154) );
  XNOR U1410 ( .A(a[45]), .B(n1154), .Z(c[45]) );
  XOR U1411 ( .A(b[46]), .B(n1155), .Z(n1156) );
  XNOR U1412 ( .A(a[46]), .B(n1156), .Z(c[46]) );
  XOR U1413 ( .A(b[47]), .B(n1157), .Z(n1158) );
  XNOR U1414 ( .A(a[47]), .B(n1158), .Z(c[47]) );
  XOR U1415 ( .A(b[48]), .B(n1159), .Z(n1160) );
  XNOR U1416 ( .A(a[48]), .B(n1160), .Z(c[48]) );
  XOR U1417 ( .A(b[49]), .B(n1161), .Z(n1162) );
  XNOR U1418 ( .A(a[49]), .B(n1162), .Z(c[49]) );
  XOR U1419 ( .A(b[4]), .B(n1163), .Z(n1164) );
  XNOR U1420 ( .A(a[4]), .B(n1164), .Z(c[4]) );
  XOR U1421 ( .A(b[50]), .B(n1165), .Z(n1166) );
  XNOR U1422 ( .A(a[50]), .B(n1166), .Z(c[50]) );
  XOR U1423 ( .A(b[51]), .B(n1167), .Z(n1168) );
  XNOR U1424 ( .A(a[51]), .B(n1168), .Z(c[51]) );
  XOR U1425 ( .A(b[52]), .B(n1169), .Z(n1170) );
  XNOR U1426 ( .A(a[52]), .B(n1170), .Z(c[52]) );
  XOR U1427 ( .A(b[53]), .B(n1171), .Z(n1172) );
  XNOR U1428 ( .A(a[53]), .B(n1172), .Z(c[53]) );
  XOR U1429 ( .A(b[54]), .B(n1173), .Z(n1174) );
  XNOR U1430 ( .A(a[54]), .B(n1174), .Z(c[54]) );
  XOR U1431 ( .A(b[55]), .B(n1175), .Z(n1176) );
  XNOR U1432 ( .A(a[55]), .B(n1176), .Z(c[55]) );
  XOR U1433 ( .A(b[56]), .B(n1177), .Z(n1178) );
  XNOR U1434 ( .A(a[56]), .B(n1178), .Z(c[56]) );
  XOR U1435 ( .A(b[57]), .B(n1179), .Z(n1180) );
  XNOR U1436 ( .A(a[57]), .B(n1180), .Z(c[57]) );
  XOR U1437 ( .A(b[58]), .B(n1181), .Z(n1182) );
  XNOR U1438 ( .A(a[58]), .B(n1182), .Z(c[58]) );
  XOR U1439 ( .A(b[59]), .B(n1183), .Z(n1184) );
  XNOR U1440 ( .A(a[59]), .B(n1184), .Z(c[59]) );
  XOR U1441 ( .A(b[5]), .B(n1185), .Z(n1186) );
  XNOR U1442 ( .A(a[5]), .B(n1186), .Z(c[5]) );
  XOR U1443 ( .A(b[60]), .B(n1187), .Z(n1188) );
  XNOR U1444 ( .A(a[60]), .B(n1188), .Z(c[60]) );
  XOR U1445 ( .A(b[61]), .B(n1189), .Z(n1190) );
  XNOR U1446 ( .A(a[61]), .B(n1190), .Z(c[61]) );
  XOR U1447 ( .A(b[62]), .B(n1191), .Z(n1192) );
  XNOR U1448 ( .A(a[62]), .B(n1192), .Z(c[62]) );
  XOR U1449 ( .A(b[63]), .B(n1193), .Z(n1194) );
  XNOR U1450 ( .A(a[63]), .B(n1194), .Z(c[63]) );
  XOR U1451 ( .A(b[64]), .B(n1195), .Z(n1196) );
  XNOR U1452 ( .A(a[64]), .B(n1196), .Z(c[64]) );
  XOR U1453 ( .A(b[65]), .B(n1197), .Z(n1198) );
  XNOR U1454 ( .A(a[65]), .B(n1198), .Z(c[65]) );
  XOR U1455 ( .A(b[66]), .B(n1199), .Z(n1200) );
  XNOR U1456 ( .A(a[66]), .B(n1200), .Z(c[66]) );
  XOR U1457 ( .A(b[67]), .B(n1201), .Z(n1202) );
  XNOR U1458 ( .A(a[67]), .B(n1202), .Z(c[67]) );
  XOR U1459 ( .A(b[68]), .B(n1203), .Z(n1204) );
  XNOR U1460 ( .A(a[68]), .B(n1204), .Z(c[68]) );
  XOR U1461 ( .A(b[69]), .B(n1205), .Z(n1206) );
  XNOR U1462 ( .A(a[69]), .B(n1206), .Z(c[69]) );
  XOR U1463 ( .A(b[6]), .B(n1207), .Z(n1208) );
  XNOR U1464 ( .A(a[6]), .B(n1208), .Z(c[6]) );
  XOR U1465 ( .A(b[70]), .B(n1209), .Z(n1210) );
  XNOR U1466 ( .A(a[70]), .B(n1210), .Z(c[70]) );
  XOR U1467 ( .A(b[71]), .B(n1211), .Z(n1212) );
  XNOR U1468 ( .A(a[71]), .B(n1212), .Z(c[71]) );
  XOR U1469 ( .A(b[72]), .B(n1213), .Z(n1214) );
  XNOR U1470 ( .A(a[72]), .B(n1214), .Z(c[72]) );
  XOR U1471 ( .A(b[73]), .B(n1215), .Z(n1216) );
  XNOR U1472 ( .A(a[73]), .B(n1216), .Z(c[73]) );
  XOR U1473 ( .A(b[74]), .B(n1217), .Z(n1218) );
  XNOR U1474 ( .A(a[74]), .B(n1218), .Z(c[74]) );
  XOR U1475 ( .A(b[75]), .B(n1219), .Z(n1220) );
  XNOR U1476 ( .A(a[75]), .B(n1220), .Z(c[75]) );
  XOR U1477 ( .A(b[76]), .B(n1221), .Z(n1222) );
  XNOR U1478 ( .A(a[76]), .B(n1222), .Z(c[76]) );
  XOR U1479 ( .A(b[77]), .B(n1223), .Z(n1224) );
  XNOR U1480 ( .A(a[77]), .B(n1224), .Z(c[77]) );
  XOR U1481 ( .A(b[78]), .B(n1225), .Z(n1226) );
  XNOR U1482 ( .A(a[78]), .B(n1226), .Z(c[78]) );
  XOR U1483 ( .A(b[79]), .B(n1227), .Z(n1228) );
  XNOR U1484 ( .A(a[79]), .B(n1228), .Z(c[79]) );
  XOR U1485 ( .A(b[7]), .B(n1229), .Z(n1230) );
  XNOR U1486 ( .A(a[7]), .B(n1230), .Z(c[7]) );
  XOR U1487 ( .A(b[80]), .B(n1231), .Z(n1232) );
  XNOR U1488 ( .A(a[80]), .B(n1232), .Z(c[80]) );
  XOR U1489 ( .A(b[81]), .B(n1233), .Z(n1234) );
  XNOR U1490 ( .A(a[81]), .B(n1234), .Z(c[81]) );
  XOR U1491 ( .A(b[82]), .B(n1235), .Z(n1236) );
  XNOR U1492 ( .A(a[82]), .B(n1236), .Z(c[82]) );
  XOR U1493 ( .A(b[83]), .B(n1237), .Z(n1238) );
  XNOR U1494 ( .A(a[83]), .B(n1238), .Z(c[83]) );
  XOR U1495 ( .A(b[84]), .B(n1239), .Z(n1240) );
  XNOR U1496 ( .A(a[84]), .B(n1240), .Z(c[84]) );
  XOR U1497 ( .A(b[85]), .B(n1241), .Z(n1242) );
  XNOR U1498 ( .A(a[85]), .B(n1242), .Z(c[85]) );
  XOR U1499 ( .A(b[86]), .B(n1243), .Z(n1244) );
  XNOR U1500 ( .A(a[86]), .B(n1244), .Z(c[86]) );
  XOR U1501 ( .A(b[87]), .B(n1245), .Z(n1246) );
  XNOR U1502 ( .A(a[87]), .B(n1246), .Z(c[87]) );
  XOR U1503 ( .A(b[88]), .B(n1247), .Z(n1248) );
  XNOR U1504 ( .A(a[88]), .B(n1248), .Z(c[88]) );
  XOR U1505 ( .A(b[89]), .B(n1249), .Z(n1250) );
  XNOR U1506 ( .A(a[89]), .B(n1250), .Z(c[89]) );
  XOR U1507 ( .A(b[8]), .B(n1251), .Z(n1252) );
  XNOR U1508 ( .A(a[8]), .B(n1252), .Z(c[8]) );
  XOR U1509 ( .A(b[90]), .B(n1253), .Z(n1254) );
  XNOR U1510 ( .A(a[90]), .B(n1254), .Z(c[90]) );
  XOR U1511 ( .A(b[91]), .B(n1255), .Z(n1256) );
  XNOR U1512 ( .A(a[91]), .B(n1256), .Z(c[91]) );
  XOR U1513 ( .A(b[92]), .B(n1257), .Z(n1258) );
  XNOR U1514 ( .A(a[92]), .B(n1258), .Z(c[92]) );
  XOR U1515 ( .A(b[93]), .B(n1259), .Z(n1260) );
  XNOR U1516 ( .A(a[93]), .B(n1260), .Z(c[93]) );
  XOR U1517 ( .A(b[94]), .B(n1261), .Z(n1262) );
  XNOR U1518 ( .A(a[94]), .B(n1262), .Z(c[94]) );
  XOR U1519 ( .A(b[95]), .B(n1263), .Z(n1264) );
  XNOR U1520 ( .A(a[95]), .B(n1264), .Z(c[95]) );
  XOR U1521 ( .A(b[96]), .B(n1265), .Z(n1266) );
  XNOR U1522 ( .A(a[96]), .B(n1266), .Z(c[96]) );
  XOR U1523 ( .A(b[97]), .B(n1267), .Z(n1268) );
  XNOR U1524 ( .A(a[97]), .B(n1268), .Z(c[97]) );
  XOR U1525 ( .A(b[98]), .B(n1269), .Z(n1270) );
  XNOR U1526 ( .A(a[98]), .B(n1270), .Z(c[98]) );
  XOR U1527 ( .A(a[99]), .B(n1271), .Z(n1272) );
  XNOR U1528 ( .A(b[99]), .B(n1272), .Z(c[99]) );
  XOR U1529 ( .A(a[9]), .B(n1273), .Z(n1274) );
  XNOR U1530 ( .A(b[9]), .B(n1274), .Z(c[9]) );
endmodule

