
module mult_N256_CC256 ( clk, rst, a, b, c );
  input [255:0] a;
  input [0:0] b;
  output [511:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277;
  wire   [511:0] sreg;

  DFF \sreg_reg[510]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(sreg[510]) );
  DFF \sreg_reg[509]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(sreg[509]) );
  DFF \sreg_reg[508]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(sreg[508]) );
  DFF \sreg_reg[507]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(sreg[507]) );
  DFF \sreg_reg[506]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(sreg[506]) );
  DFF \sreg_reg[505]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(sreg[505]) );
  DFF \sreg_reg[504]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(sreg[504]) );
  DFF \sreg_reg[503]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(sreg[503]) );
  DFF \sreg_reg[502]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(sreg[502]) );
  DFF \sreg_reg[501]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(sreg[501]) );
  DFF \sreg_reg[500]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(sreg[500]) );
  DFF \sreg_reg[499]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(sreg[499]) );
  DFF \sreg_reg[498]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(sreg[498]) );
  DFF \sreg_reg[497]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(sreg[497]) );
  DFF \sreg_reg[496]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(sreg[496]) );
  DFF \sreg_reg[495]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(sreg[495]) );
  DFF \sreg_reg[494]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(sreg[494]) );
  DFF \sreg_reg[493]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(sreg[493]) );
  DFF \sreg_reg[492]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(sreg[492]) );
  DFF \sreg_reg[491]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(sreg[491]) );
  DFF \sreg_reg[490]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(sreg[490]) );
  DFF \sreg_reg[489]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(sreg[489]) );
  DFF \sreg_reg[488]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(sreg[488]) );
  DFF \sreg_reg[487]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(sreg[487]) );
  DFF \sreg_reg[486]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(sreg[486]) );
  DFF \sreg_reg[485]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(sreg[485]) );
  DFF \sreg_reg[484]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(sreg[484]) );
  DFF \sreg_reg[483]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(sreg[483]) );
  DFF \sreg_reg[482]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(sreg[482]) );
  DFF \sreg_reg[481]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(sreg[481]) );
  DFF \sreg_reg[480]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(sreg[480]) );
  DFF \sreg_reg[479]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[478]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[477]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[476]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[475]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[474]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[473]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[472]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[471]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[470]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[469]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[468]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[467]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[466]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[465]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[464]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[463]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[462]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[461]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[460]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[459]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[458]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[457]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[456]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[455]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[454]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[453]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[452]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[451]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[450]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[449]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[448]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[447]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[446]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[445]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[444]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[443]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[442]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[441]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[440]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[439]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[438]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[437]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[436]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[435]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[434]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[433]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[432]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[431]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[430]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[429]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[428]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[427]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[426]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[425]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[424]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[423]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[422]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[421]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[420]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[419]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[418]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[417]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[416]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[415]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[414]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[413]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[412]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[411]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[410]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[409]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[408]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[407]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[406]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[405]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[404]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[403]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[402]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[401]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[400]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[399]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[398]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[397]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[396]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[395]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[394]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[393]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[392]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[391]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[390]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[389]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[388]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[387]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[386]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[385]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[384]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[383]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[382]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[381]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[380]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[379]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[378]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[377]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[376]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[375]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[374]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[373]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[372]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[371]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[370]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[369]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[368]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[367]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[366]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[365]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[364]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[363]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[362]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[361]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[360]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[359]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[358]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[357]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[356]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[355]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[354]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[353]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[352]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[351]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[350]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[349]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[348]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[347]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[346]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[345]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[344]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[343]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[342]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[341]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[340]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[339]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[338]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[337]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[336]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[335]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[334]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[333]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[332]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[331]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[330]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[329]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[328]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[327]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[326]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[325]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[324]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[323]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[322]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[321]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[320]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[319]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[318]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[317]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[316]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[315]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[314]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[313]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[312]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[311]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[310]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[309]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[308]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[307]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[306]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[305]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[304]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[303]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[302]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[301]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[300]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[299]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[298]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[297]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[296]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[295]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[294]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[293]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[292]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[291]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[290]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[289]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[288]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[287]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[286]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[285]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[284]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[283]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[282]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[281]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[280]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[279]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[278]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[277]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[276]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[275]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[274]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[273]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[272]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[271]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[270]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[269]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[268]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[267]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[266]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[265]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[264]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[263]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[262]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[261]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[260]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[259]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[258]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[257]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[256]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[255]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(sreg[255]) );
  DFF \sreg_reg[254]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[254]) );
  DFF \sreg_reg[253]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[252]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[251]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[250]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[249]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[248]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[247]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[1]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U4 ( .A(b[0]), .B(a[0]), .Z(n1) );
  XNOR U5 ( .A(n1), .B(sreg[255]), .Z(c[255]) );
  NAND U6 ( .A(b[0]), .B(a[1]), .Z(n2) );
  XOR U7 ( .A(sreg[256]), .B(n2), .Z(n4) );
  NANDN U8 ( .A(n1), .B(sreg[255]), .Z(n3) );
  XOR U9 ( .A(n4), .B(n3), .Z(c[256]) );
  NAND U10 ( .A(b[0]), .B(a[2]), .Z(n7) );
  XOR U11 ( .A(sreg[257]), .B(n7), .Z(n9) );
  NANDN U12 ( .A(n2), .B(sreg[256]), .Z(n6) );
  OR U13 ( .A(n4), .B(n3), .Z(n5) );
  AND U14 ( .A(n6), .B(n5), .Z(n8) );
  XOR U15 ( .A(n9), .B(n8), .Z(c[257]) );
  NAND U16 ( .A(b[0]), .B(a[3]), .Z(n12) );
  XOR U17 ( .A(sreg[258]), .B(n12), .Z(n14) );
  NANDN U18 ( .A(n7), .B(sreg[257]), .Z(n11) );
  OR U19 ( .A(n9), .B(n8), .Z(n10) );
  AND U20 ( .A(n11), .B(n10), .Z(n13) );
  XOR U21 ( .A(n14), .B(n13), .Z(c[258]) );
  NAND U22 ( .A(b[0]), .B(a[4]), .Z(n17) );
  XOR U23 ( .A(sreg[259]), .B(n17), .Z(n19) );
  NANDN U24 ( .A(n12), .B(sreg[258]), .Z(n16) );
  OR U25 ( .A(n14), .B(n13), .Z(n15) );
  AND U26 ( .A(n16), .B(n15), .Z(n18) );
  XOR U27 ( .A(n19), .B(n18), .Z(c[259]) );
  NAND U28 ( .A(b[0]), .B(a[5]), .Z(n22) );
  XOR U29 ( .A(sreg[260]), .B(n22), .Z(n24) );
  NANDN U30 ( .A(n17), .B(sreg[259]), .Z(n21) );
  OR U31 ( .A(n19), .B(n18), .Z(n20) );
  AND U32 ( .A(n21), .B(n20), .Z(n23) );
  XOR U33 ( .A(n24), .B(n23), .Z(c[260]) );
  NAND U34 ( .A(b[0]), .B(a[6]), .Z(n27) );
  XOR U35 ( .A(sreg[261]), .B(n27), .Z(n29) );
  NANDN U36 ( .A(n22), .B(sreg[260]), .Z(n26) );
  OR U37 ( .A(n24), .B(n23), .Z(n25) );
  AND U38 ( .A(n26), .B(n25), .Z(n28) );
  XOR U39 ( .A(n29), .B(n28), .Z(c[261]) );
  NAND U40 ( .A(b[0]), .B(a[7]), .Z(n32) );
  XOR U41 ( .A(sreg[262]), .B(n32), .Z(n34) );
  NANDN U42 ( .A(n27), .B(sreg[261]), .Z(n31) );
  OR U43 ( .A(n29), .B(n28), .Z(n30) );
  AND U44 ( .A(n31), .B(n30), .Z(n33) );
  XOR U45 ( .A(n34), .B(n33), .Z(c[262]) );
  NAND U46 ( .A(b[0]), .B(a[8]), .Z(n37) );
  XOR U47 ( .A(sreg[263]), .B(n37), .Z(n39) );
  NANDN U48 ( .A(n32), .B(sreg[262]), .Z(n36) );
  OR U49 ( .A(n34), .B(n33), .Z(n35) );
  AND U50 ( .A(n36), .B(n35), .Z(n38) );
  XOR U51 ( .A(n39), .B(n38), .Z(c[263]) );
  NAND U52 ( .A(b[0]), .B(a[9]), .Z(n42) );
  XOR U53 ( .A(sreg[264]), .B(n42), .Z(n44) );
  NANDN U54 ( .A(n37), .B(sreg[263]), .Z(n41) );
  OR U55 ( .A(n39), .B(n38), .Z(n40) );
  AND U56 ( .A(n41), .B(n40), .Z(n43) );
  XOR U57 ( .A(n44), .B(n43), .Z(c[264]) );
  NAND U58 ( .A(b[0]), .B(a[10]), .Z(n47) );
  XOR U59 ( .A(sreg[265]), .B(n47), .Z(n49) );
  NANDN U60 ( .A(n42), .B(sreg[264]), .Z(n46) );
  OR U61 ( .A(n44), .B(n43), .Z(n45) );
  AND U62 ( .A(n46), .B(n45), .Z(n48) );
  XOR U63 ( .A(n49), .B(n48), .Z(c[265]) );
  NAND U64 ( .A(b[0]), .B(a[11]), .Z(n52) );
  XOR U65 ( .A(sreg[266]), .B(n52), .Z(n54) );
  NANDN U66 ( .A(n47), .B(sreg[265]), .Z(n51) );
  OR U67 ( .A(n49), .B(n48), .Z(n50) );
  AND U68 ( .A(n51), .B(n50), .Z(n53) );
  XOR U69 ( .A(n54), .B(n53), .Z(c[266]) );
  NAND U70 ( .A(b[0]), .B(a[12]), .Z(n57) );
  XOR U71 ( .A(sreg[267]), .B(n57), .Z(n59) );
  NANDN U72 ( .A(n52), .B(sreg[266]), .Z(n56) );
  OR U73 ( .A(n54), .B(n53), .Z(n55) );
  AND U74 ( .A(n56), .B(n55), .Z(n58) );
  XOR U75 ( .A(n59), .B(n58), .Z(c[267]) );
  NAND U76 ( .A(b[0]), .B(a[13]), .Z(n62) );
  XOR U77 ( .A(sreg[268]), .B(n62), .Z(n64) );
  NANDN U78 ( .A(n57), .B(sreg[267]), .Z(n61) );
  OR U79 ( .A(n59), .B(n58), .Z(n60) );
  AND U80 ( .A(n61), .B(n60), .Z(n63) );
  XOR U81 ( .A(n64), .B(n63), .Z(c[268]) );
  NAND U82 ( .A(b[0]), .B(a[14]), .Z(n67) );
  XOR U83 ( .A(sreg[269]), .B(n67), .Z(n69) );
  NANDN U84 ( .A(n62), .B(sreg[268]), .Z(n66) );
  OR U85 ( .A(n64), .B(n63), .Z(n65) );
  AND U86 ( .A(n66), .B(n65), .Z(n68) );
  XOR U87 ( .A(n69), .B(n68), .Z(c[269]) );
  NAND U88 ( .A(b[0]), .B(a[15]), .Z(n72) );
  XOR U89 ( .A(sreg[270]), .B(n72), .Z(n74) );
  NANDN U90 ( .A(n67), .B(sreg[269]), .Z(n71) );
  OR U91 ( .A(n69), .B(n68), .Z(n70) );
  AND U92 ( .A(n71), .B(n70), .Z(n73) );
  XOR U93 ( .A(n74), .B(n73), .Z(c[270]) );
  NAND U94 ( .A(b[0]), .B(a[16]), .Z(n77) );
  XOR U95 ( .A(sreg[271]), .B(n77), .Z(n79) );
  NANDN U96 ( .A(n72), .B(sreg[270]), .Z(n76) );
  OR U97 ( .A(n74), .B(n73), .Z(n75) );
  AND U98 ( .A(n76), .B(n75), .Z(n78) );
  XOR U99 ( .A(n79), .B(n78), .Z(c[271]) );
  NAND U100 ( .A(b[0]), .B(a[17]), .Z(n82) );
  XOR U101 ( .A(sreg[272]), .B(n82), .Z(n84) );
  NANDN U102 ( .A(n77), .B(sreg[271]), .Z(n81) );
  OR U103 ( .A(n79), .B(n78), .Z(n80) );
  AND U104 ( .A(n81), .B(n80), .Z(n83) );
  XOR U105 ( .A(n84), .B(n83), .Z(c[272]) );
  NAND U106 ( .A(b[0]), .B(a[18]), .Z(n87) );
  XOR U107 ( .A(sreg[273]), .B(n87), .Z(n89) );
  NANDN U108 ( .A(n82), .B(sreg[272]), .Z(n86) );
  OR U109 ( .A(n84), .B(n83), .Z(n85) );
  AND U110 ( .A(n86), .B(n85), .Z(n88) );
  XOR U111 ( .A(n89), .B(n88), .Z(c[273]) );
  NAND U112 ( .A(b[0]), .B(a[19]), .Z(n92) );
  XOR U113 ( .A(sreg[274]), .B(n92), .Z(n94) );
  NANDN U114 ( .A(n87), .B(sreg[273]), .Z(n91) );
  OR U115 ( .A(n89), .B(n88), .Z(n90) );
  AND U116 ( .A(n91), .B(n90), .Z(n93) );
  XOR U117 ( .A(n94), .B(n93), .Z(c[274]) );
  NAND U118 ( .A(b[0]), .B(a[20]), .Z(n97) );
  XOR U119 ( .A(sreg[275]), .B(n97), .Z(n99) );
  NANDN U120 ( .A(n92), .B(sreg[274]), .Z(n96) );
  OR U121 ( .A(n94), .B(n93), .Z(n95) );
  AND U122 ( .A(n96), .B(n95), .Z(n98) );
  XOR U123 ( .A(n99), .B(n98), .Z(c[275]) );
  NAND U124 ( .A(b[0]), .B(a[21]), .Z(n102) );
  XOR U125 ( .A(sreg[276]), .B(n102), .Z(n104) );
  NANDN U126 ( .A(n97), .B(sreg[275]), .Z(n101) );
  OR U127 ( .A(n99), .B(n98), .Z(n100) );
  AND U128 ( .A(n101), .B(n100), .Z(n103) );
  XOR U129 ( .A(n104), .B(n103), .Z(c[276]) );
  NAND U130 ( .A(b[0]), .B(a[22]), .Z(n107) );
  XOR U131 ( .A(sreg[277]), .B(n107), .Z(n109) );
  NANDN U132 ( .A(n102), .B(sreg[276]), .Z(n106) );
  OR U133 ( .A(n104), .B(n103), .Z(n105) );
  AND U134 ( .A(n106), .B(n105), .Z(n108) );
  XOR U135 ( .A(n109), .B(n108), .Z(c[277]) );
  NAND U136 ( .A(b[0]), .B(a[23]), .Z(n112) );
  XOR U137 ( .A(sreg[278]), .B(n112), .Z(n114) );
  NANDN U138 ( .A(n107), .B(sreg[277]), .Z(n111) );
  OR U139 ( .A(n109), .B(n108), .Z(n110) );
  AND U140 ( .A(n111), .B(n110), .Z(n113) );
  XOR U141 ( .A(n114), .B(n113), .Z(c[278]) );
  NAND U142 ( .A(b[0]), .B(a[24]), .Z(n117) );
  XOR U143 ( .A(sreg[279]), .B(n117), .Z(n119) );
  NANDN U144 ( .A(n112), .B(sreg[278]), .Z(n116) );
  OR U145 ( .A(n114), .B(n113), .Z(n115) );
  AND U146 ( .A(n116), .B(n115), .Z(n118) );
  XOR U147 ( .A(n119), .B(n118), .Z(c[279]) );
  NAND U148 ( .A(b[0]), .B(a[25]), .Z(n122) );
  XOR U149 ( .A(sreg[280]), .B(n122), .Z(n124) );
  NANDN U150 ( .A(n117), .B(sreg[279]), .Z(n121) );
  OR U151 ( .A(n119), .B(n118), .Z(n120) );
  AND U152 ( .A(n121), .B(n120), .Z(n123) );
  XOR U153 ( .A(n124), .B(n123), .Z(c[280]) );
  NAND U154 ( .A(b[0]), .B(a[26]), .Z(n127) );
  XOR U155 ( .A(sreg[281]), .B(n127), .Z(n129) );
  NANDN U156 ( .A(n122), .B(sreg[280]), .Z(n126) );
  OR U157 ( .A(n124), .B(n123), .Z(n125) );
  AND U158 ( .A(n126), .B(n125), .Z(n128) );
  XOR U159 ( .A(n129), .B(n128), .Z(c[281]) );
  NAND U160 ( .A(b[0]), .B(a[27]), .Z(n132) );
  XOR U161 ( .A(sreg[282]), .B(n132), .Z(n134) );
  NANDN U162 ( .A(n127), .B(sreg[281]), .Z(n131) );
  OR U163 ( .A(n129), .B(n128), .Z(n130) );
  AND U164 ( .A(n131), .B(n130), .Z(n133) );
  XOR U165 ( .A(n134), .B(n133), .Z(c[282]) );
  NAND U166 ( .A(b[0]), .B(a[28]), .Z(n137) );
  XOR U167 ( .A(sreg[283]), .B(n137), .Z(n139) );
  NANDN U168 ( .A(n132), .B(sreg[282]), .Z(n136) );
  OR U169 ( .A(n134), .B(n133), .Z(n135) );
  AND U170 ( .A(n136), .B(n135), .Z(n138) );
  XOR U171 ( .A(n139), .B(n138), .Z(c[283]) );
  NAND U172 ( .A(b[0]), .B(a[29]), .Z(n142) );
  XOR U173 ( .A(sreg[284]), .B(n142), .Z(n144) );
  NANDN U174 ( .A(n137), .B(sreg[283]), .Z(n141) );
  OR U175 ( .A(n139), .B(n138), .Z(n140) );
  AND U176 ( .A(n141), .B(n140), .Z(n143) );
  XOR U177 ( .A(n144), .B(n143), .Z(c[284]) );
  NAND U178 ( .A(b[0]), .B(a[30]), .Z(n147) );
  XOR U179 ( .A(sreg[285]), .B(n147), .Z(n149) );
  NANDN U180 ( .A(n142), .B(sreg[284]), .Z(n146) );
  OR U181 ( .A(n144), .B(n143), .Z(n145) );
  AND U182 ( .A(n146), .B(n145), .Z(n148) );
  XOR U183 ( .A(n149), .B(n148), .Z(c[285]) );
  NAND U184 ( .A(b[0]), .B(a[31]), .Z(n152) );
  XOR U185 ( .A(sreg[286]), .B(n152), .Z(n154) );
  NANDN U186 ( .A(n147), .B(sreg[285]), .Z(n151) );
  OR U187 ( .A(n149), .B(n148), .Z(n150) );
  AND U188 ( .A(n151), .B(n150), .Z(n153) );
  XOR U189 ( .A(n154), .B(n153), .Z(c[286]) );
  NAND U190 ( .A(b[0]), .B(a[32]), .Z(n157) );
  XOR U191 ( .A(sreg[287]), .B(n157), .Z(n159) );
  NANDN U192 ( .A(n152), .B(sreg[286]), .Z(n156) );
  OR U193 ( .A(n154), .B(n153), .Z(n155) );
  AND U194 ( .A(n156), .B(n155), .Z(n158) );
  XOR U195 ( .A(n159), .B(n158), .Z(c[287]) );
  NAND U196 ( .A(b[0]), .B(a[33]), .Z(n162) );
  XOR U197 ( .A(sreg[288]), .B(n162), .Z(n164) );
  NANDN U198 ( .A(n157), .B(sreg[287]), .Z(n161) );
  OR U199 ( .A(n159), .B(n158), .Z(n160) );
  AND U200 ( .A(n161), .B(n160), .Z(n163) );
  XOR U201 ( .A(n164), .B(n163), .Z(c[288]) );
  NAND U202 ( .A(b[0]), .B(a[34]), .Z(n167) );
  XOR U203 ( .A(sreg[289]), .B(n167), .Z(n169) );
  NANDN U204 ( .A(n162), .B(sreg[288]), .Z(n166) );
  OR U205 ( .A(n164), .B(n163), .Z(n165) );
  AND U206 ( .A(n166), .B(n165), .Z(n168) );
  XOR U207 ( .A(n169), .B(n168), .Z(c[289]) );
  NAND U208 ( .A(b[0]), .B(a[35]), .Z(n172) );
  XOR U209 ( .A(sreg[290]), .B(n172), .Z(n174) );
  NANDN U210 ( .A(n167), .B(sreg[289]), .Z(n171) );
  OR U211 ( .A(n169), .B(n168), .Z(n170) );
  AND U212 ( .A(n171), .B(n170), .Z(n173) );
  XOR U213 ( .A(n174), .B(n173), .Z(c[290]) );
  NAND U214 ( .A(b[0]), .B(a[36]), .Z(n177) );
  XOR U215 ( .A(sreg[291]), .B(n177), .Z(n179) );
  NANDN U216 ( .A(n172), .B(sreg[290]), .Z(n176) );
  OR U217 ( .A(n174), .B(n173), .Z(n175) );
  AND U218 ( .A(n176), .B(n175), .Z(n178) );
  XOR U219 ( .A(n179), .B(n178), .Z(c[291]) );
  NAND U220 ( .A(b[0]), .B(a[37]), .Z(n182) );
  XOR U221 ( .A(sreg[292]), .B(n182), .Z(n184) );
  NANDN U222 ( .A(n177), .B(sreg[291]), .Z(n181) );
  OR U223 ( .A(n179), .B(n178), .Z(n180) );
  AND U224 ( .A(n181), .B(n180), .Z(n183) );
  XOR U225 ( .A(n184), .B(n183), .Z(c[292]) );
  NAND U226 ( .A(b[0]), .B(a[38]), .Z(n187) );
  XOR U227 ( .A(sreg[293]), .B(n187), .Z(n189) );
  NANDN U228 ( .A(n182), .B(sreg[292]), .Z(n186) );
  OR U229 ( .A(n184), .B(n183), .Z(n185) );
  AND U230 ( .A(n186), .B(n185), .Z(n188) );
  XOR U231 ( .A(n189), .B(n188), .Z(c[293]) );
  NAND U232 ( .A(b[0]), .B(a[39]), .Z(n192) );
  XOR U233 ( .A(sreg[294]), .B(n192), .Z(n194) );
  NANDN U234 ( .A(n187), .B(sreg[293]), .Z(n191) );
  OR U235 ( .A(n189), .B(n188), .Z(n190) );
  AND U236 ( .A(n191), .B(n190), .Z(n193) );
  XOR U237 ( .A(n194), .B(n193), .Z(c[294]) );
  NAND U238 ( .A(b[0]), .B(a[40]), .Z(n197) );
  XOR U239 ( .A(sreg[295]), .B(n197), .Z(n199) );
  NANDN U240 ( .A(n192), .B(sreg[294]), .Z(n196) );
  OR U241 ( .A(n194), .B(n193), .Z(n195) );
  AND U242 ( .A(n196), .B(n195), .Z(n198) );
  XOR U243 ( .A(n199), .B(n198), .Z(c[295]) );
  NAND U244 ( .A(b[0]), .B(a[41]), .Z(n202) );
  XOR U245 ( .A(sreg[296]), .B(n202), .Z(n204) );
  NANDN U246 ( .A(n197), .B(sreg[295]), .Z(n201) );
  OR U247 ( .A(n199), .B(n198), .Z(n200) );
  AND U248 ( .A(n201), .B(n200), .Z(n203) );
  XOR U249 ( .A(n204), .B(n203), .Z(c[296]) );
  NAND U250 ( .A(b[0]), .B(a[42]), .Z(n207) );
  XOR U251 ( .A(sreg[297]), .B(n207), .Z(n209) );
  NANDN U252 ( .A(n202), .B(sreg[296]), .Z(n206) );
  OR U253 ( .A(n204), .B(n203), .Z(n205) );
  AND U254 ( .A(n206), .B(n205), .Z(n208) );
  XOR U255 ( .A(n209), .B(n208), .Z(c[297]) );
  NAND U256 ( .A(b[0]), .B(a[43]), .Z(n212) );
  XOR U257 ( .A(sreg[298]), .B(n212), .Z(n214) );
  NANDN U258 ( .A(n207), .B(sreg[297]), .Z(n211) );
  OR U259 ( .A(n209), .B(n208), .Z(n210) );
  AND U260 ( .A(n211), .B(n210), .Z(n213) );
  XOR U261 ( .A(n214), .B(n213), .Z(c[298]) );
  NAND U262 ( .A(b[0]), .B(a[44]), .Z(n217) );
  XOR U263 ( .A(sreg[299]), .B(n217), .Z(n219) );
  NANDN U264 ( .A(n212), .B(sreg[298]), .Z(n216) );
  OR U265 ( .A(n214), .B(n213), .Z(n215) );
  AND U266 ( .A(n216), .B(n215), .Z(n218) );
  XOR U267 ( .A(n219), .B(n218), .Z(c[299]) );
  NAND U268 ( .A(b[0]), .B(a[45]), .Z(n222) );
  XOR U269 ( .A(sreg[300]), .B(n222), .Z(n224) );
  NANDN U270 ( .A(n217), .B(sreg[299]), .Z(n221) );
  OR U271 ( .A(n219), .B(n218), .Z(n220) );
  AND U272 ( .A(n221), .B(n220), .Z(n223) );
  XOR U273 ( .A(n224), .B(n223), .Z(c[300]) );
  NAND U274 ( .A(b[0]), .B(a[46]), .Z(n227) );
  XOR U275 ( .A(sreg[301]), .B(n227), .Z(n229) );
  NANDN U276 ( .A(n222), .B(sreg[300]), .Z(n226) );
  OR U277 ( .A(n224), .B(n223), .Z(n225) );
  AND U278 ( .A(n226), .B(n225), .Z(n228) );
  XOR U279 ( .A(n229), .B(n228), .Z(c[301]) );
  NAND U280 ( .A(b[0]), .B(a[47]), .Z(n232) );
  XOR U281 ( .A(sreg[302]), .B(n232), .Z(n234) );
  NANDN U282 ( .A(n227), .B(sreg[301]), .Z(n231) );
  OR U283 ( .A(n229), .B(n228), .Z(n230) );
  AND U284 ( .A(n231), .B(n230), .Z(n233) );
  XOR U285 ( .A(n234), .B(n233), .Z(c[302]) );
  NAND U286 ( .A(b[0]), .B(a[48]), .Z(n237) );
  XOR U287 ( .A(sreg[303]), .B(n237), .Z(n239) );
  NANDN U288 ( .A(n232), .B(sreg[302]), .Z(n236) );
  OR U289 ( .A(n234), .B(n233), .Z(n235) );
  AND U290 ( .A(n236), .B(n235), .Z(n238) );
  XOR U291 ( .A(n239), .B(n238), .Z(c[303]) );
  NAND U292 ( .A(b[0]), .B(a[49]), .Z(n242) );
  XOR U293 ( .A(sreg[304]), .B(n242), .Z(n244) );
  NANDN U294 ( .A(n237), .B(sreg[303]), .Z(n241) );
  OR U295 ( .A(n239), .B(n238), .Z(n240) );
  AND U296 ( .A(n241), .B(n240), .Z(n243) );
  XOR U297 ( .A(n244), .B(n243), .Z(c[304]) );
  NAND U298 ( .A(b[0]), .B(a[50]), .Z(n247) );
  XOR U299 ( .A(sreg[305]), .B(n247), .Z(n249) );
  NANDN U300 ( .A(n242), .B(sreg[304]), .Z(n246) );
  OR U301 ( .A(n244), .B(n243), .Z(n245) );
  AND U302 ( .A(n246), .B(n245), .Z(n248) );
  XOR U303 ( .A(n249), .B(n248), .Z(c[305]) );
  NAND U304 ( .A(b[0]), .B(a[51]), .Z(n252) );
  XOR U305 ( .A(sreg[306]), .B(n252), .Z(n254) );
  NANDN U306 ( .A(n247), .B(sreg[305]), .Z(n251) );
  OR U307 ( .A(n249), .B(n248), .Z(n250) );
  AND U308 ( .A(n251), .B(n250), .Z(n253) );
  XOR U309 ( .A(n254), .B(n253), .Z(c[306]) );
  NAND U310 ( .A(b[0]), .B(a[52]), .Z(n257) );
  XOR U311 ( .A(sreg[307]), .B(n257), .Z(n259) );
  NANDN U312 ( .A(n252), .B(sreg[306]), .Z(n256) );
  OR U313 ( .A(n254), .B(n253), .Z(n255) );
  AND U314 ( .A(n256), .B(n255), .Z(n258) );
  XOR U315 ( .A(n259), .B(n258), .Z(c[307]) );
  NAND U316 ( .A(b[0]), .B(a[53]), .Z(n262) );
  XOR U317 ( .A(sreg[308]), .B(n262), .Z(n264) );
  NANDN U318 ( .A(n257), .B(sreg[307]), .Z(n261) );
  OR U319 ( .A(n259), .B(n258), .Z(n260) );
  AND U320 ( .A(n261), .B(n260), .Z(n263) );
  XOR U321 ( .A(n264), .B(n263), .Z(c[308]) );
  NAND U322 ( .A(b[0]), .B(a[54]), .Z(n267) );
  XOR U323 ( .A(sreg[309]), .B(n267), .Z(n269) );
  NANDN U324 ( .A(n262), .B(sreg[308]), .Z(n266) );
  OR U325 ( .A(n264), .B(n263), .Z(n265) );
  AND U326 ( .A(n266), .B(n265), .Z(n268) );
  XOR U327 ( .A(n269), .B(n268), .Z(c[309]) );
  NAND U328 ( .A(b[0]), .B(a[55]), .Z(n272) );
  XOR U329 ( .A(sreg[310]), .B(n272), .Z(n274) );
  NANDN U330 ( .A(n267), .B(sreg[309]), .Z(n271) );
  OR U331 ( .A(n269), .B(n268), .Z(n270) );
  AND U332 ( .A(n271), .B(n270), .Z(n273) );
  XOR U333 ( .A(n274), .B(n273), .Z(c[310]) );
  NAND U334 ( .A(b[0]), .B(a[56]), .Z(n277) );
  XOR U335 ( .A(sreg[311]), .B(n277), .Z(n279) );
  NANDN U336 ( .A(n272), .B(sreg[310]), .Z(n276) );
  OR U337 ( .A(n274), .B(n273), .Z(n275) );
  AND U338 ( .A(n276), .B(n275), .Z(n278) );
  XOR U339 ( .A(n279), .B(n278), .Z(c[311]) );
  NAND U340 ( .A(b[0]), .B(a[57]), .Z(n282) );
  XOR U341 ( .A(sreg[312]), .B(n282), .Z(n284) );
  NANDN U342 ( .A(n277), .B(sreg[311]), .Z(n281) );
  OR U343 ( .A(n279), .B(n278), .Z(n280) );
  AND U344 ( .A(n281), .B(n280), .Z(n283) );
  XOR U345 ( .A(n284), .B(n283), .Z(c[312]) );
  NAND U346 ( .A(b[0]), .B(a[58]), .Z(n287) );
  XOR U347 ( .A(sreg[313]), .B(n287), .Z(n289) );
  NANDN U348 ( .A(n282), .B(sreg[312]), .Z(n286) );
  OR U349 ( .A(n284), .B(n283), .Z(n285) );
  AND U350 ( .A(n286), .B(n285), .Z(n288) );
  XOR U351 ( .A(n289), .B(n288), .Z(c[313]) );
  NAND U352 ( .A(b[0]), .B(a[59]), .Z(n292) );
  XOR U353 ( .A(sreg[314]), .B(n292), .Z(n294) );
  NANDN U354 ( .A(n287), .B(sreg[313]), .Z(n291) );
  OR U355 ( .A(n289), .B(n288), .Z(n290) );
  AND U356 ( .A(n291), .B(n290), .Z(n293) );
  XOR U357 ( .A(n294), .B(n293), .Z(c[314]) );
  NAND U358 ( .A(b[0]), .B(a[60]), .Z(n297) );
  XOR U359 ( .A(sreg[315]), .B(n297), .Z(n299) );
  NANDN U360 ( .A(n292), .B(sreg[314]), .Z(n296) );
  OR U361 ( .A(n294), .B(n293), .Z(n295) );
  AND U362 ( .A(n296), .B(n295), .Z(n298) );
  XOR U363 ( .A(n299), .B(n298), .Z(c[315]) );
  NAND U364 ( .A(b[0]), .B(a[61]), .Z(n302) );
  XOR U365 ( .A(sreg[316]), .B(n302), .Z(n304) );
  NANDN U366 ( .A(n297), .B(sreg[315]), .Z(n301) );
  OR U367 ( .A(n299), .B(n298), .Z(n300) );
  AND U368 ( .A(n301), .B(n300), .Z(n303) );
  XOR U369 ( .A(n304), .B(n303), .Z(c[316]) );
  NAND U370 ( .A(b[0]), .B(a[62]), .Z(n307) );
  XOR U371 ( .A(sreg[317]), .B(n307), .Z(n309) );
  NANDN U372 ( .A(n302), .B(sreg[316]), .Z(n306) );
  OR U373 ( .A(n304), .B(n303), .Z(n305) );
  AND U374 ( .A(n306), .B(n305), .Z(n308) );
  XOR U375 ( .A(n309), .B(n308), .Z(c[317]) );
  NAND U376 ( .A(b[0]), .B(a[63]), .Z(n312) );
  XOR U377 ( .A(sreg[318]), .B(n312), .Z(n314) );
  NANDN U378 ( .A(n307), .B(sreg[317]), .Z(n311) );
  OR U379 ( .A(n309), .B(n308), .Z(n310) );
  AND U380 ( .A(n311), .B(n310), .Z(n313) );
  XOR U381 ( .A(n314), .B(n313), .Z(c[318]) );
  NAND U382 ( .A(b[0]), .B(a[64]), .Z(n317) );
  XOR U383 ( .A(sreg[319]), .B(n317), .Z(n319) );
  NANDN U384 ( .A(n312), .B(sreg[318]), .Z(n316) );
  OR U385 ( .A(n314), .B(n313), .Z(n315) );
  AND U386 ( .A(n316), .B(n315), .Z(n318) );
  XOR U387 ( .A(n319), .B(n318), .Z(c[319]) );
  NAND U388 ( .A(b[0]), .B(a[65]), .Z(n322) );
  XOR U389 ( .A(sreg[320]), .B(n322), .Z(n324) );
  NANDN U390 ( .A(n317), .B(sreg[319]), .Z(n321) );
  OR U391 ( .A(n319), .B(n318), .Z(n320) );
  AND U392 ( .A(n321), .B(n320), .Z(n323) );
  XOR U393 ( .A(n324), .B(n323), .Z(c[320]) );
  NAND U394 ( .A(b[0]), .B(a[66]), .Z(n327) );
  XOR U395 ( .A(sreg[321]), .B(n327), .Z(n329) );
  NANDN U396 ( .A(n322), .B(sreg[320]), .Z(n326) );
  OR U397 ( .A(n324), .B(n323), .Z(n325) );
  AND U398 ( .A(n326), .B(n325), .Z(n328) );
  XOR U399 ( .A(n329), .B(n328), .Z(c[321]) );
  NAND U400 ( .A(b[0]), .B(a[67]), .Z(n332) );
  XOR U401 ( .A(sreg[322]), .B(n332), .Z(n334) );
  NANDN U402 ( .A(n327), .B(sreg[321]), .Z(n331) );
  OR U403 ( .A(n329), .B(n328), .Z(n330) );
  AND U404 ( .A(n331), .B(n330), .Z(n333) );
  XOR U405 ( .A(n334), .B(n333), .Z(c[322]) );
  NAND U406 ( .A(b[0]), .B(a[68]), .Z(n337) );
  XOR U407 ( .A(sreg[323]), .B(n337), .Z(n339) );
  NANDN U408 ( .A(n332), .B(sreg[322]), .Z(n336) );
  OR U409 ( .A(n334), .B(n333), .Z(n335) );
  AND U410 ( .A(n336), .B(n335), .Z(n338) );
  XOR U411 ( .A(n339), .B(n338), .Z(c[323]) );
  NAND U412 ( .A(b[0]), .B(a[69]), .Z(n342) );
  XOR U413 ( .A(sreg[324]), .B(n342), .Z(n344) );
  NANDN U414 ( .A(n337), .B(sreg[323]), .Z(n341) );
  OR U415 ( .A(n339), .B(n338), .Z(n340) );
  AND U416 ( .A(n341), .B(n340), .Z(n343) );
  XOR U417 ( .A(n344), .B(n343), .Z(c[324]) );
  NAND U418 ( .A(b[0]), .B(a[70]), .Z(n347) );
  XOR U419 ( .A(sreg[325]), .B(n347), .Z(n349) );
  NANDN U420 ( .A(n342), .B(sreg[324]), .Z(n346) );
  OR U421 ( .A(n344), .B(n343), .Z(n345) );
  AND U422 ( .A(n346), .B(n345), .Z(n348) );
  XOR U423 ( .A(n349), .B(n348), .Z(c[325]) );
  NAND U424 ( .A(b[0]), .B(a[71]), .Z(n352) );
  XOR U425 ( .A(sreg[326]), .B(n352), .Z(n354) );
  NANDN U426 ( .A(n347), .B(sreg[325]), .Z(n351) );
  OR U427 ( .A(n349), .B(n348), .Z(n350) );
  AND U428 ( .A(n351), .B(n350), .Z(n353) );
  XOR U429 ( .A(n354), .B(n353), .Z(c[326]) );
  NAND U430 ( .A(b[0]), .B(a[72]), .Z(n357) );
  XOR U431 ( .A(sreg[327]), .B(n357), .Z(n359) );
  NANDN U432 ( .A(n352), .B(sreg[326]), .Z(n356) );
  OR U433 ( .A(n354), .B(n353), .Z(n355) );
  AND U434 ( .A(n356), .B(n355), .Z(n358) );
  XOR U435 ( .A(n359), .B(n358), .Z(c[327]) );
  NAND U436 ( .A(b[0]), .B(a[73]), .Z(n362) );
  XOR U437 ( .A(sreg[328]), .B(n362), .Z(n364) );
  NANDN U438 ( .A(n357), .B(sreg[327]), .Z(n361) );
  OR U439 ( .A(n359), .B(n358), .Z(n360) );
  AND U440 ( .A(n361), .B(n360), .Z(n363) );
  XOR U441 ( .A(n364), .B(n363), .Z(c[328]) );
  NAND U442 ( .A(b[0]), .B(a[74]), .Z(n367) );
  XOR U443 ( .A(sreg[329]), .B(n367), .Z(n369) );
  NANDN U444 ( .A(n362), .B(sreg[328]), .Z(n366) );
  OR U445 ( .A(n364), .B(n363), .Z(n365) );
  AND U446 ( .A(n366), .B(n365), .Z(n368) );
  XOR U447 ( .A(n369), .B(n368), .Z(c[329]) );
  NAND U448 ( .A(b[0]), .B(a[75]), .Z(n372) );
  XOR U449 ( .A(sreg[330]), .B(n372), .Z(n374) );
  NANDN U450 ( .A(n367), .B(sreg[329]), .Z(n371) );
  OR U451 ( .A(n369), .B(n368), .Z(n370) );
  AND U452 ( .A(n371), .B(n370), .Z(n373) );
  XOR U453 ( .A(n374), .B(n373), .Z(c[330]) );
  NAND U454 ( .A(b[0]), .B(a[76]), .Z(n377) );
  XOR U455 ( .A(sreg[331]), .B(n377), .Z(n379) );
  NANDN U456 ( .A(n372), .B(sreg[330]), .Z(n376) );
  OR U457 ( .A(n374), .B(n373), .Z(n375) );
  AND U458 ( .A(n376), .B(n375), .Z(n378) );
  XOR U459 ( .A(n379), .B(n378), .Z(c[331]) );
  NAND U460 ( .A(b[0]), .B(a[77]), .Z(n382) );
  XOR U461 ( .A(sreg[332]), .B(n382), .Z(n384) );
  NANDN U462 ( .A(n377), .B(sreg[331]), .Z(n381) );
  OR U463 ( .A(n379), .B(n378), .Z(n380) );
  AND U464 ( .A(n381), .B(n380), .Z(n383) );
  XOR U465 ( .A(n384), .B(n383), .Z(c[332]) );
  NAND U466 ( .A(b[0]), .B(a[78]), .Z(n387) );
  XOR U467 ( .A(sreg[333]), .B(n387), .Z(n389) );
  NANDN U468 ( .A(n382), .B(sreg[332]), .Z(n386) );
  OR U469 ( .A(n384), .B(n383), .Z(n385) );
  AND U470 ( .A(n386), .B(n385), .Z(n388) );
  XOR U471 ( .A(n389), .B(n388), .Z(c[333]) );
  NAND U472 ( .A(b[0]), .B(a[79]), .Z(n392) );
  XOR U473 ( .A(sreg[334]), .B(n392), .Z(n394) );
  NANDN U474 ( .A(n387), .B(sreg[333]), .Z(n391) );
  OR U475 ( .A(n389), .B(n388), .Z(n390) );
  AND U476 ( .A(n391), .B(n390), .Z(n393) );
  XOR U477 ( .A(n394), .B(n393), .Z(c[334]) );
  NAND U478 ( .A(b[0]), .B(a[80]), .Z(n397) );
  XOR U479 ( .A(sreg[335]), .B(n397), .Z(n399) );
  NANDN U480 ( .A(n392), .B(sreg[334]), .Z(n396) );
  OR U481 ( .A(n394), .B(n393), .Z(n395) );
  AND U482 ( .A(n396), .B(n395), .Z(n398) );
  XOR U483 ( .A(n399), .B(n398), .Z(c[335]) );
  NAND U484 ( .A(b[0]), .B(a[81]), .Z(n402) );
  XOR U485 ( .A(sreg[336]), .B(n402), .Z(n404) );
  NANDN U486 ( .A(n397), .B(sreg[335]), .Z(n401) );
  OR U487 ( .A(n399), .B(n398), .Z(n400) );
  AND U488 ( .A(n401), .B(n400), .Z(n403) );
  XOR U489 ( .A(n404), .B(n403), .Z(c[336]) );
  NAND U490 ( .A(b[0]), .B(a[82]), .Z(n407) );
  XOR U491 ( .A(sreg[337]), .B(n407), .Z(n409) );
  NANDN U492 ( .A(n402), .B(sreg[336]), .Z(n406) );
  OR U493 ( .A(n404), .B(n403), .Z(n405) );
  AND U494 ( .A(n406), .B(n405), .Z(n408) );
  XOR U495 ( .A(n409), .B(n408), .Z(c[337]) );
  NAND U496 ( .A(b[0]), .B(a[83]), .Z(n412) );
  XOR U497 ( .A(sreg[338]), .B(n412), .Z(n414) );
  NANDN U498 ( .A(n407), .B(sreg[337]), .Z(n411) );
  OR U499 ( .A(n409), .B(n408), .Z(n410) );
  AND U500 ( .A(n411), .B(n410), .Z(n413) );
  XOR U501 ( .A(n414), .B(n413), .Z(c[338]) );
  NAND U502 ( .A(b[0]), .B(a[84]), .Z(n417) );
  XOR U503 ( .A(sreg[339]), .B(n417), .Z(n419) );
  NANDN U504 ( .A(n412), .B(sreg[338]), .Z(n416) );
  OR U505 ( .A(n414), .B(n413), .Z(n415) );
  AND U506 ( .A(n416), .B(n415), .Z(n418) );
  XOR U507 ( .A(n419), .B(n418), .Z(c[339]) );
  NAND U508 ( .A(b[0]), .B(a[85]), .Z(n422) );
  XOR U509 ( .A(sreg[340]), .B(n422), .Z(n424) );
  NANDN U510 ( .A(n417), .B(sreg[339]), .Z(n421) );
  OR U511 ( .A(n419), .B(n418), .Z(n420) );
  AND U512 ( .A(n421), .B(n420), .Z(n423) );
  XOR U513 ( .A(n424), .B(n423), .Z(c[340]) );
  NAND U514 ( .A(b[0]), .B(a[86]), .Z(n427) );
  XOR U515 ( .A(sreg[341]), .B(n427), .Z(n429) );
  NANDN U516 ( .A(n422), .B(sreg[340]), .Z(n426) );
  OR U517 ( .A(n424), .B(n423), .Z(n425) );
  AND U518 ( .A(n426), .B(n425), .Z(n428) );
  XOR U519 ( .A(n429), .B(n428), .Z(c[341]) );
  NAND U520 ( .A(b[0]), .B(a[87]), .Z(n432) );
  XOR U521 ( .A(sreg[342]), .B(n432), .Z(n434) );
  NANDN U522 ( .A(n427), .B(sreg[341]), .Z(n431) );
  OR U523 ( .A(n429), .B(n428), .Z(n430) );
  AND U524 ( .A(n431), .B(n430), .Z(n433) );
  XOR U525 ( .A(n434), .B(n433), .Z(c[342]) );
  NAND U526 ( .A(b[0]), .B(a[88]), .Z(n437) );
  XOR U527 ( .A(sreg[343]), .B(n437), .Z(n439) );
  NANDN U528 ( .A(n432), .B(sreg[342]), .Z(n436) );
  OR U529 ( .A(n434), .B(n433), .Z(n435) );
  AND U530 ( .A(n436), .B(n435), .Z(n438) );
  XOR U531 ( .A(n439), .B(n438), .Z(c[343]) );
  NAND U532 ( .A(b[0]), .B(a[89]), .Z(n442) );
  XOR U533 ( .A(sreg[344]), .B(n442), .Z(n444) );
  NANDN U534 ( .A(n437), .B(sreg[343]), .Z(n441) );
  OR U535 ( .A(n439), .B(n438), .Z(n440) );
  AND U536 ( .A(n441), .B(n440), .Z(n443) );
  XOR U537 ( .A(n444), .B(n443), .Z(c[344]) );
  NAND U538 ( .A(b[0]), .B(a[90]), .Z(n447) );
  XOR U539 ( .A(sreg[345]), .B(n447), .Z(n449) );
  NANDN U540 ( .A(n442), .B(sreg[344]), .Z(n446) );
  OR U541 ( .A(n444), .B(n443), .Z(n445) );
  AND U542 ( .A(n446), .B(n445), .Z(n448) );
  XOR U543 ( .A(n449), .B(n448), .Z(c[345]) );
  NAND U544 ( .A(b[0]), .B(a[91]), .Z(n452) );
  XOR U545 ( .A(sreg[346]), .B(n452), .Z(n454) );
  NANDN U546 ( .A(n447), .B(sreg[345]), .Z(n451) );
  OR U547 ( .A(n449), .B(n448), .Z(n450) );
  AND U548 ( .A(n451), .B(n450), .Z(n453) );
  XOR U549 ( .A(n454), .B(n453), .Z(c[346]) );
  NAND U550 ( .A(b[0]), .B(a[92]), .Z(n457) );
  XOR U551 ( .A(sreg[347]), .B(n457), .Z(n459) );
  NANDN U552 ( .A(n452), .B(sreg[346]), .Z(n456) );
  OR U553 ( .A(n454), .B(n453), .Z(n455) );
  AND U554 ( .A(n456), .B(n455), .Z(n458) );
  XOR U555 ( .A(n459), .B(n458), .Z(c[347]) );
  NAND U556 ( .A(b[0]), .B(a[93]), .Z(n462) );
  XOR U557 ( .A(sreg[348]), .B(n462), .Z(n464) );
  NANDN U558 ( .A(n457), .B(sreg[347]), .Z(n461) );
  OR U559 ( .A(n459), .B(n458), .Z(n460) );
  AND U560 ( .A(n461), .B(n460), .Z(n463) );
  XOR U561 ( .A(n464), .B(n463), .Z(c[348]) );
  NAND U562 ( .A(b[0]), .B(a[94]), .Z(n467) );
  XOR U563 ( .A(sreg[349]), .B(n467), .Z(n469) );
  NANDN U564 ( .A(n462), .B(sreg[348]), .Z(n466) );
  OR U565 ( .A(n464), .B(n463), .Z(n465) );
  AND U566 ( .A(n466), .B(n465), .Z(n468) );
  XOR U567 ( .A(n469), .B(n468), .Z(c[349]) );
  NAND U568 ( .A(b[0]), .B(a[95]), .Z(n472) );
  XOR U569 ( .A(sreg[350]), .B(n472), .Z(n474) );
  NANDN U570 ( .A(n467), .B(sreg[349]), .Z(n471) );
  OR U571 ( .A(n469), .B(n468), .Z(n470) );
  AND U572 ( .A(n471), .B(n470), .Z(n473) );
  XOR U573 ( .A(n474), .B(n473), .Z(c[350]) );
  NAND U574 ( .A(b[0]), .B(a[96]), .Z(n477) );
  XOR U575 ( .A(sreg[351]), .B(n477), .Z(n479) );
  NANDN U576 ( .A(n472), .B(sreg[350]), .Z(n476) );
  OR U577 ( .A(n474), .B(n473), .Z(n475) );
  AND U578 ( .A(n476), .B(n475), .Z(n478) );
  XOR U579 ( .A(n479), .B(n478), .Z(c[351]) );
  NAND U580 ( .A(b[0]), .B(a[97]), .Z(n482) );
  XOR U581 ( .A(sreg[352]), .B(n482), .Z(n484) );
  NANDN U582 ( .A(n477), .B(sreg[351]), .Z(n481) );
  OR U583 ( .A(n479), .B(n478), .Z(n480) );
  AND U584 ( .A(n481), .B(n480), .Z(n483) );
  XOR U585 ( .A(n484), .B(n483), .Z(c[352]) );
  NAND U586 ( .A(b[0]), .B(a[98]), .Z(n487) );
  XOR U587 ( .A(sreg[353]), .B(n487), .Z(n489) );
  NANDN U588 ( .A(n482), .B(sreg[352]), .Z(n486) );
  OR U589 ( .A(n484), .B(n483), .Z(n485) );
  AND U590 ( .A(n486), .B(n485), .Z(n488) );
  XOR U591 ( .A(n489), .B(n488), .Z(c[353]) );
  NAND U592 ( .A(b[0]), .B(a[99]), .Z(n492) );
  XOR U593 ( .A(sreg[354]), .B(n492), .Z(n494) );
  NANDN U594 ( .A(n487), .B(sreg[353]), .Z(n491) );
  OR U595 ( .A(n489), .B(n488), .Z(n490) );
  AND U596 ( .A(n491), .B(n490), .Z(n493) );
  XOR U597 ( .A(n494), .B(n493), .Z(c[354]) );
  NAND U598 ( .A(b[0]), .B(a[100]), .Z(n497) );
  XOR U599 ( .A(sreg[355]), .B(n497), .Z(n499) );
  NANDN U600 ( .A(n492), .B(sreg[354]), .Z(n496) );
  OR U601 ( .A(n494), .B(n493), .Z(n495) );
  AND U602 ( .A(n496), .B(n495), .Z(n498) );
  XOR U603 ( .A(n499), .B(n498), .Z(c[355]) );
  NAND U604 ( .A(b[0]), .B(a[101]), .Z(n502) );
  XOR U605 ( .A(sreg[356]), .B(n502), .Z(n504) );
  NANDN U606 ( .A(n497), .B(sreg[355]), .Z(n501) );
  OR U607 ( .A(n499), .B(n498), .Z(n500) );
  AND U608 ( .A(n501), .B(n500), .Z(n503) );
  XOR U609 ( .A(n504), .B(n503), .Z(c[356]) );
  NAND U610 ( .A(b[0]), .B(a[102]), .Z(n507) );
  XOR U611 ( .A(sreg[357]), .B(n507), .Z(n509) );
  NANDN U612 ( .A(n502), .B(sreg[356]), .Z(n506) );
  OR U613 ( .A(n504), .B(n503), .Z(n505) );
  AND U614 ( .A(n506), .B(n505), .Z(n508) );
  XOR U615 ( .A(n509), .B(n508), .Z(c[357]) );
  NAND U616 ( .A(b[0]), .B(a[103]), .Z(n512) );
  XOR U617 ( .A(sreg[358]), .B(n512), .Z(n514) );
  NANDN U618 ( .A(n507), .B(sreg[357]), .Z(n511) );
  OR U619 ( .A(n509), .B(n508), .Z(n510) );
  AND U620 ( .A(n511), .B(n510), .Z(n513) );
  XOR U621 ( .A(n514), .B(n513), .Z(c[358]) );
  NAND U622 ( .A(b[0]), .B(a[104]), .Z(n517) );
  XOR U623 ( .A(sreg[359]), .B(n517), .Z(n519) );
  NANDN U624 ( .A(n512), .B(sreg[358]), .Z(n516) );
  OR U625 ( .A(n514), .B(n513), .Z(n515) );
  AND U626 ( .A(n516), .B(n515), .Z(n518) );
  XOR U627 ( .A(n519), .B(n518), .Z(c[359]) );
  NAND U628 ( .A(b[0]), .B(a[105]), .Z(n522) );
  XOR U629 ( .A(sreg[360]), .B(n522), .Z(n524) );
  NANDN U630 ( .A(n517), .B(sreg[359]), .Z(n521) );
  OR U631 ( .A(n519), .B(n518), .Z(n520) );
  AND U632 ( .A(n521), .B(n520), .Z(n523) );
  XOR U633 ( .A(n524), .B(n523), .Z(c[360]) );
  NAND U634 ( .A(b[0]), .B(a[106]), .Z(n527) );
  XOR U635 ( .A(sreg[361]), .B(n527), .Z(n529) );
  NANDN U636 ( .A(n522), .B(sreg[360]), .Z(n526) );
  OR U637 ( .A(n524), .B(n523), .Z(n525) );
  AND U638 ( .A(n526), .B(n525), .Z(n528) );
  XOR U639 ( .A(n529), .B(n528), .Z(c[361]) );
  NAND U640 ( .A(b[0]), .B(a[107]), .Z(n532) );
  XOR U641 ( .A(sreg[362]), .B(n532), .Z(n534) );
  NANDN U642 ( .A(n527), .B(sreg[361]), .Z(n531) );
  OR U643 ( .A(n529), .B(n528), .Z(n530) );
  AND U644 ( .A(n531), .B(n530), .Z(n533) );
  XOR U645 ( .A(n534), .B(n533), .Z(c[362]) );
  NAND U646 ( .A(b[0]), .B(a[108]), .Z(n537) );
  XOR U647 ( .A(sreg[363]), .B(n537), .Z(n539) );
  NANDN U648 ( .A(n532), .B(sreg[362]), .Z(n536) );
  OR U649 ( .A(n534), .B(n533), .Z(n535) );
  AND U650 ( .A(n536), .B(n535), .Z(n538) );
  XOR U651 ( .A(n539), .B(n538), .Z(c[363]) );
  NAND U652 ( .A(b[0]), .B(a[109]), .Z(n542) );
  XOR U653 ( .A(sreg[364]), .B(n542), .Z(n544) );
  NANDN U654 ( .A(n537), .B(sreg[363]), .Z(n541) );
  OR U655 ( .A(n539), .B(n538), .Z(n540) );
  AND U656 ( .A(n541), .B(n540), .Z(n543) );
  XOR U657 ( .A(n544), .B(n543), .Z(c[364]) );
  NAND U658 ( .A(b[0]), .B(a[110]), .Z(n547) );
  XOR U659 ( .A(sreg[365]), .B(n547), .Z(n549) );
  NANDN U660 ( .A(n542), .B(sreg[364]), .Z(n546) );
  OR U661 ( .A(n544), .B(n543), .Z(n545) );
  AND U662 ( .A(n546), .B(n545), .Z(n548) );
  XOR U663 ( .A(n549), .B(n548), .Z(c[365]) );
  NAND U664 ( .A(b[0]), .B(a[111]), .Z(n552) );
  XOR U665 ( .A(sreg[366]), .B(n552), .Z(n554) );
  NANDN U666 ( .A(n547), .B(sreg[365]), .Z(n551) );
  OR U667 ( .A(n549), .B(n548), .Z(n550) );
  AND U668 ( .A(n551), .B(n550), .Z(n553) );
  XOR U669 ( .A(n554), .B(n553), .Z(c[366]) );
  NAND U670 ( .A(b[0]), .B(a[112]), .Z(n557) );
  XOR U671 ( .A(sreg[367]), .B(n557), .Z(n559) );
  NANDN U672 ( .A(n552), .B(sreg[366]), .Z(n556) );
  OR U673 ( .A(n554), .B(n553), .Z(n555) );
  AND U674 ( .A(n556), .B(n555), .Z(n558) );
  XOR U675 ( .A(n559), .B(n558), .Z(c[367]) );
  NAND U676 ( .A(b[0]), .B(a[113]), .Z(n562) );
  XOR U677 ( .A(sreg[368]), .B(n562), .Z(n564) );
  NANDN U678 ( .A(n557), .B(sreg[367]), .Z(n561) );
  OR U679 ( .A(n559), .B(n558), .Z(n560) );
  AND U680 ( .A(n561), .B(n560), .Z(n563) );
  XOR U681 ( .A(n564), .B(n563), .Z(c[368]) );
  NAND U682 ( .A(b[0]), .B(a[114]), .Z(n567) );
  XOR U683 ( .A(sreg[369]), .B(n567), .Z(n569) );
  NANDN U684 ( .A(n562), .B(sreg[368]), .Z(n566) );
  OR U685 ( .A(n564), .B(n563), .Z(n565) );
  AND U686 ( .A(n566), .B(n565), .Z(n568) );
  XOR U687 ( .A(n569), .B(n568), .Z(c[369]) );
  NAND U688 ( .A(b[0]), .B(a[115]), .Z(n572) );
  XOR U689 ( .A(sreg[370]), .B(n572), .Z(n574) );
  NANDN U690 ( .A(n567), .B(sreg[369]), .Z(n571) );
  OR U691 ( .A(n569), .B(n568), .Z(n570) );
  AND U692 ( .A(n571), .B(n570), .Z(n573) );
  XOR U693 ( .A(n574), .B(n573), .Z(c[370]) );
  NAND U694 ( .A(b[0]), .B(a[116]), .Z(n577) );
  XOR U695 ( .A(sreg[371]), .B(n577), .Z(n579) );
  NANDN U696 ( .A(n572), .B(sreg[370]), .Z(n576) );
  OR U697 ( .A(n574), .B(n573), .Z(n575) );
  AND U698 ( .A(n576), .B(n575), .Z(n578) );
  XOR U699 ( .A(n579), .B(n578), .Z(c[371]) );
  NAND U700 ( .A(b[0]), .B(a[117]), .Z(n582) );
  XOR U701 ( .A(sreg[372]), .B(n582), .Z(n584) );
  NANDN U702 ( .A(n577), .B(sreg[371]), .Z(n581) );
  OR U703 ( .A(n579), .B(n578), .Z(n580) );
  AND U704 ( .A(n581), .B(n580), .Z(n583) );
  XOR U705 ( .A(n584), .B(n583), .Z(c[372]) );
  NAND U706 ( .A(b[0]), .B(a[118]), .Z(n587) );
  XOR U707 ( .A(sreg[373]), .B(n587), .Z(n589) );
  NANDN U708 ( .A(n582), .B(sreg[372]), .Z(n586) );
  OR U709 ( .A(n584), .B(n583), .Z(n585) );
  AND U710 ( .A(n586), .B(n585), .Z(n588) );
  XOR U711 ( .A(n589), .B(n588), .Z(c[373]) );
  NAND U712 ( .A(b[0]), .B(a[119]), .Z(n592) );
  XOR U713 ( .A(sreg[374]), .B(n592), .Z(n594) );
  NANDN U714 ( .A(n587), .B(sreg[373]), .Z(n591) );
  OR U715 ( .A(n589), .B(n588), .Z(n590) );
  AND U716 ( .A(n591), .B(n590), .Z(n593) );
  XOR U717 ( .A(n594), .B(n593), .Z(c[374]) );
  NAND U718 ( .A(b[0]), .B(a[120]), .Z(n597) );
  XOR U719 ( .A(sreg[375]), .B(n597), .Z(n599) );
  NANDN U720 ( .A(n592), .B(sreg[374]), .Z(n596) );
  OR U721 ( .A(n594), .B(n593), .Z(n595) );
  AND U722 ( .A(n596), .B(n595), .Z(n598) );
  XOR U723 ( .A(n599), .B(n598), .Z(c[375]) );
  NAND U724 ( .A(b[0]), .B(a[121]), .Z(n602) );
  XOR U725 ( .A(sreg[376]), .B(n602), .Z(n604) );
  NANDN U726 ( .A(n597), .B(sreg[375]), .Z(n601) );
  OR U727 ( .A(n599), .B(n598), .Z(n600) );
  AND U728 ( .A(n601), .B(n600), .Z(n603) );
  XOR U729 ( .A(n604), .B(n603), .Z(c[376]) );
  NAND U730 ( .A(b[0]), .B(a[122]), .Z(n607) );
  XOR U731 ( .A(sreg[377]), .B(n607), .Z(n609) );
  NANDN U732 ( .A(n602), .B(sreg[376]), .Z(n606) );
  OR U733 ( .A(n604), .B(n603), .Z(n605) );
  AND U734 ( .A(n606), .B(n605), .Z(n608) );
  XOR U735 ( .A(n609), .B(n608), .Z(c[377]) );
  NAND U736 ( .A(b[0]), .B(a[123]), .Z(n612) );
  XOR U737 ( .A(sreg[378]), .B(n612), .Z(n614) );
  NANDN U738 ( .A(n607), .B(sreg[377]), .Z(n611) );
  OR U739 ( .A(n609), .B(n608), .Z(n610) );
  AND U740 ( .A(n611), .B(n610), .Z(n613) );
  XOR U741 ( .A(n614), .B(n613), .Z(c[378]) );
  NAND U742 ( .A(b[0]), .B(a[124]), .Z(n617) );
  XOR U743 ( .A(sreg[379]), .B(n617), .Z(n619) );
  NANDN U744 ( .A(n612), .B(sreg[378]), .Z(n616) );
  OR U745 ( .A(n614), .B(n613), .Z(n615) );
  AND U746 ( .A(n616), .B(n615), .Z(n618) );
  XOR U747 ( .A(n619), .B(n618), .Z(c[379]) );
  NAND U748 ( .A(b[0]), .B(a[125]), .Z(n622) );
  XOR U749 ( .A(sreg[380]), .B(n622), .Z(n624) );
  NANDN U750 ( .A(n617), .B(sreg[379]), .Z(n621) );
  OR U751 ( .A(n619), .B(n618), .Z(n620) );
  AND U752 ( .A(n621), .B(n620), .Z(n623) );
  XOR U753 ( .A(n624), .B(n623), .Z(c[380]) );
  NAND U754 ( .A(b[0]), .B(a[126]), .Z(n627) );
  XOR U755 ( .A(sreg[381]), .B(n627), .Z(n629) );
  NANDN U756 ( .A(n622), .B(sreg[380]), .Z(n626) );
  OR U757 ( .A(n624), .B(n623), .Z(n625) );
  AND U758 ( .A(n626), .B(n625), .Z(n628) );
  XOR U759 ( .A(n629), .B(n628), .Z(c[381]) );
  NAND U760 ( .A(b[0]), .B(a[127]), .Z(n632) );
  XOR U761 ( .A(sreg[382]), .B(n632), .Z(n634) );
  NANDN U762 ( .A(n627), .B(sreg[381]), .Z(n631) );
  OR U763 ( .A(n629), .B(n628), .Z(n630) );
  AND U764 ( .A(n631), .B(n630), .Z(n633) );
  XOR U765 ( .A(n634), .B(n633), .Z(c[382]) );
  NAND U766 ( .A(b[0]), .B(a[128]), .Z(n637) );
  XOR U767 ( .A(sreg[383]), .B(n637), .Z(n639) );
  NANDN U768 ( .A(n632), .B(sreg[382]), .Z(n636) );
  OR U769 ( .A(n634), .B(n633), .Z(n635) );
  AND U770 ( .A(n636), .B(n635), .Z(n638) );
  XOR U771 ( .A(n639), .B(n638), .Z(c[383]) );
  NAND U772 ( .A(b[0]), .B(a[129]), .Z(n642) );
  XOR U773 ( .A(sreg[384]), .B(n642), .Z(n644) );
  NANDN U774 ( .A(n637), .B(sreg[383]), .Z(n641) );
  OR U775 ( .A(n639), .B(n638), .Z(n640) );
  AND U776 ( .A(n641), .B(n640), .Z(n643) );
  XOR U777 ( .A(n644), .B(n643), .Z(c[384]) );
  NAND U778 ( .A(b[0]), .B(a[130]), .Z(n647) );
  XOR U779 ( .A(sreg[385]), .B(n647), .Z(n649) );
  NANDN U780 ( .A(n642), .B(sreg[384]), .Z(n646) );
  OR U781 ( .A(n644), .B(n643), .Z(n645) );
  AND U782 ( .A(n646), .B(n645), .Z(n648) );
  XOR U783 ( .A(n649), .B(n648), .Z(c[385]) );
  NAND U784 ( .A(b[0]), .B(a[131]), .Z(n652) );
  XOR U785 ( .A(sreg[386]), .B(n652), .Z(n654) );
  NANDN U786 ( .A(n647), .B(sreg[385]), .Z(n651) );
  OR U787 ( .A(n649), .B(n648), .Z(n650) );
  AND U788 ( .A(n651), .B(n650), .Z(n653) );
  XOR U789 ( .A(n654), .B(n653), .Z(c[386]) );
  NAND U790 ( .A(b[0]), .B(a[132]), .Z(n657) );
  XOR U791 ( .A(sreg[387]), .B(n657), .Z(n659) );
  NANDN U792 ( .A(n652), .B(sreg[386]), .Z(n656) );
  OR U793 ( .A(n654), .B(n653), .Z(n655) );
  AND U794 ( .A(n656), .B(n655), .Z(n658) );
  XOR U795 ( .A(n659), .B(n658), .Z(c[387]) );
  NAND U796 ( .A(b[0]), .B(a[133]), .Z(n662) );
  XOR U797 ( .A(sreg[388]), .B(n662), .Z(n664) );
  NANDN U798 ( .A(n657), .B(sreg[387]), .Z(n661) );
  OR U799 ( .A(n659), .B(n658), .Z(n660) );
  AND U800 ( .A(n661), .B(n660), .Z(n663) );
  XOR U801 ( .A(n664), .B(n663), .Z(c[388]) );
  NAND U802 ( .A(b[0]), .B(a[134]), .Z(n667) );
  XOR U803 ( .A(sreg[389]), .B(n667), .Z(n669) );
  NANDN U804 ( .A(n662), .B(sreg[388]), .Z(n666) );
  OR U805 ( .A(n664), .B(n663), .Z(n665) );
  AND U806 ( .A(n666), .B(n665), .Z(n668) );
  XOR U807 ( .A(n669), .B(n668), .Z(c[389]) );
  NAND U808 ( .A(b[0]), .B(a[135]), .Z(n672) );
  XOR U809 ( .A(sreg[390]), .B(n672), .Z(n674) );
  NANDN U810 ( .A(n667), .B(sreg[389]), .Z(n671) );
  OR U811 ( .A(n669), .B(n668), .Z(n670) );
  AND U812 ( .A(n671), .B(n670), .Z(n673) );
  XOR U813 ( .A(n674), .B(n673), .Z(c[390]) );
  NAND U814 ( .A(b[0]), .B(a[136]), .Z(n677) );
  XOR U815 ( .A(sreg[391]), .B(n677), .Z(n679) );
  NANDN U816 ( .A(n672), .B(sreg[390]), .Z(n676) );
  OR U817 ( .A(n674), .B(n673), .Z(n675) );
  AND U818 ( .A(n676), .B(n675), .Z(n678) );
  XOR U819 ( .A(n679), .B(n678), .Z(c[391]) );
  NAND U820 ( .A(b[0]), .B(a[137]), .Z(n682) );
  XOR U821 ( .A(sreg[392]), .B(n682), .Z(n684) );
  NANDN U822 ( .A(n677), .B(sreg[391]), .Z(n681) );
  OR U823 ( .A(n679), .B(n678), .Z(n680) );
  AND U824 ( .A(n681), .B(n680), .Z(n683) );
  XOR U825 ( .A(n684), .B(n683), .Z(c[392]) );
  NAND U826 ( .A(b[0]), .B(a[138]), .Z(n687) );
  XOR U827 ( .A(sreg[393]), .B(n687), .Z(n689) );
  NANDN U828 ( .A(n682), .B(sreg[392]), .Z(n686) );
  OR U829 ( .A(n684), .B(n683), .Z(n685) );
  AND U830 ( .A(n686), .B(n685), .Z(n688) );
  XOR U831 ( .A(n689), .B(n688), .Z(c[393]) );
  NAND U832 ( .A(b[0]), .B(a[139]), .Z(n692) );
  XOR U833 ( .A(sreg[394]), .B(n692), .Z(n694) );
  NANDN U834 ( .A(n687), .B(sreg[393]), .Z(n691) );
  OR U835 ( .A(n689), .B(n688), .Z(n690) );
  AND U836 ( .A(n691), .B(n690), .Z(n693) );
  XOR U837 ( .A(n694), .B(n693), .Z(c[394]) );
  NAND U838 ( .A(b[0]), .B(a[140]), .Z(n697) );
  XOR U839 ( .A(sreg[395]), .B(n697), .Z(n699) );
  NANDN U840 ( .A(n692), .B(sreg[394]), .Z(n696) );
  OR U841 ( .A(n694), .B(n693), .Z(n695) );
  AND U842 ( .A(n696), .B(n695), .Z(n698) );
  XOR U843 ( .A(n699), .B(n698), .Z(c[395]) );
  NAND U844 ( .A(b[0]), .B(a[141]), .Z(n702) );
  XOR U845 ( .A(sreg[396]), .B(n702), .Z(n704) );
  NANDN U846 ( .A(n697), .B(sreg[395]), .Z(n701) );
  OR U847 ( .A(n699), .B(n698), .Z(n700) );
  AND U848 ( .A(n701), .B(n700), .Z(n703) );
  XOR U849 ( .A(n704), .B(n703), .Z(c[396]) );
  NAND U850 ( .A(b[0]), .B(a[142]), .Z(n707) );
  XOR U851 ( .A(sreg[397]), .B(n707), .Z(n709) );
  NANDN U852 ( .A(n702), .B(sreg[396]), .Z(n706) );
  OR U853 ( .A(n704), .B(n703), .Z(n705) );
  AND U854 ( .A(n706), .B(n705), .Z(n708) );
  XOR U855 ( .A(n709), .B(n708), .Z(c[397]) );
  NAND U856 ( .A(b[0]), .B(a[143]), .Z(n712) );
  XOR U857 ( .A(sreg[398]), .B(n712), .Z(n714) );
  NANDN U858 ( .A(n707), .B(sreg[397]), .Z(n711) );
  OR U859 ( .A(n709), .B(n708), .Z(n710) );
  AND U860 ( .A(n711), .B(n710), .Z(n713) );
  XOR U861 ( .A(n714), .B(n713), .Z(c[398]) );
  NAND U862 ( .A(b[0]), .B(a[144]), .Z(n717) );
  XOR U863 ( .A(sreg[399]), .B(n717), .Z(n719) );
  NANDN U864 ( .A(n712), .B(sreg[398]), .Z(n716) );
  OR U865 ( .A(n714), .B(n713), .Z(n715) );
  AND U866 ( .A(n716), .B(n715), .Z(n718) );
  XOR U867 ( .A(n719), .B(n718), .Z(c[399]) );
  NAND U868 ( .A(b[0]), .B(a[145]), .Z(n722) );
  XOR U869 ( .A(sreg[400]), .B(n722), .Z(n724) );
  NANDN U870 ( .A(n717), .B(sreg[399]), .Z(n721) );
  OR U871 ( .A(n719), .B(n718), .Z(n720) );
  AND U872 ( .A(n721), .B(n720), .Z(n723) );
  XOR U873 ( .A(n724), .B(n723), .Z(c[400]) );
  NAND U874 ( .A(b[0]), .B(a[146]), .Z(n727) );
  XOR U875 ( .A(sreg[401]), .B(n727), .Z(n729) );
  NANDN U876 ( .A(n722), .B(sreg[400]), .Z(n726) );
  OR U877 ( .A(n724), .B(n723), .Z(n725) );
  AND U878 ( .A(n726), .B(n725), .Z(n728) );
  XOR U879 ( .A(n729), .B(n728), .Z(c[401]) );
  NAND U880 ( .A(b[0]), .B(a[147]), .Z(n732) );
  XOR U881 ( .A(sreg[402]), .B(n732), .Z(n734) );
  NANDN U882 ( .A(n727), .B(sreg[401]), .Z(n731) );
  OR U883 ( .A(n729), .B(n728), .Z(n730) );
  AND U884 ( .A(n731), .B(n730), .Z(n733) );
  XOR U885 ( .A(n734), .B(n733), .Z(c[402]) );
  NAND U886 ( .A(b[0]), .B(a[148]), .Z(n737) );
  XOR U887 ( .A(sreg[403]), .B(n737), .Z(n739) );
  NANDN U888 ( .A(n732), .B(sreg[402]), .Z(n736) );
  OR U889 ( .A(n734), .B(n733), .Z(n735) );
  AND U890 ( .A(n736), .B(n735), .Z(n738) );
  XOR U891 ( .A(n739), .B(n738), .Z(c[403]) );
  NAND U892 ( .A(b[0]), .B(a[149]), .Z(n742) );
  XOR U893 ( .A(sreg[404]), .B(n742), .Z(n744) );
  NANDN U894 ( .A(n737), .B(sreg[403]), .Z(n741) );
  OR U895 ( .A(n739), .B(n738), .Z(n740) );
  AND U896 ( .A(n741), .B(n740), .Z(n743) );
  XOR U897 ( .A(n744), .B(n743), .Z(c[404]) );
  NAND U898 ( .A(b[0]), .B(a[150]), .Z(n747) );
  XOR U899 ( .A(sreg[405]), .B(n747), .Z(n749) );
  NANDN U900 ( .A(n742), .B(sreg[404]), .Z(n746) );
  OR U901 ( .A(n744), .B(n743), .Z(n745) );
  AND U902 ( .A(n746), .B(n745), .Z(n748) );
  XOR U903 ( .A(n749), .B(n748), .Z(c[405]) );
  NAND U904 ( .A(b[0]), .B(a[151]), .Z(n752) );
  XOR U905 ( .A(sreg[406]), .B(n752), .Z(n754) );
  NANDN U906 ( .A(n747), .B(sreg[405]), .Z(n751) );
  OR U907 ( .A(n749), .B(n748), .Z(n750) );
  AND U908 ( .A(n751), .B(n750), .Z(n753) );
  XOR U909 ( .A(n754), .B(n753), .Z(c[406]) );
  NAND U910 ( .A(b[0]), .B(a[152]), .Z(n757) );
  XOR U911 ( .A(sreg[407]), .B(n757), .Z(n759) );
  NANDN U912 ( .A(n752), .B(sreg[406]), .Z(n756) );
  OR U913 ( .A(n754), .B(n753), .Z(n755) );
  AND U914 ( .A(n756), .B(n755), .Z(n758) );
  XOR U915 ( .A(n759), .B(n758), .Z(c[407]) );
  NAND U916 ( .A(b[0]), .B(a[153]), .Z(n762) );
  XOR U917 ( .A(sreg[408]), .B(n762), .Z(n764) );
  NANDN U918 ( .A(n757), .B(sreg[407]), .Z(n761) );
  OR U919 ( .A(n759), .B(n758), .Z(n760) );
  AND U920 ( .A(n761), .B(n760), .Z(n763) );
  XOR U921 ( .A(n764), .B(n763), .Z(c[408]) );
  NAND U922 ( .A(b[0]), .B(a[154]), .Z(n767) );
  XOR U923 ( .A(sreg[409]), .B(n767), .Z(n769) );
  NANDN U924 ( .A(n762), .B(sreg[408]), .Z(n766) );
  OR U925 ( .A(n764), .B(n763), .Z(n765) );
  AND U926 ( .A(n766), .B(n765), .Z(n768) );
  XOR U927 ( .A(n769), .B(n768), .Z(c[409]) );
  NAND U928 ( .A(b[0]), .B(a[155]), .Z(n772) );
  XOR U929 ( .A(sreg[410]), .B(n772), .Z(n774) );
  NANDN U930 ( .A(n767), .B(sreg[409]), .Z(n771) );
  OR U931 ( .A(n769), .B(n768), .Z(n770) );
  AND U932 ( .A(n771), .B(n770), .Z(n773) );
  XOR U933 ( .A(n774), .B(n773), .Z(c[410]) );
  NAND U934 ( .A(b[0]), .B(a[156]), .Z(n777) );
  XOR U935 ( .A(sreg[411]), .B(n777), .Z(n779) );
  NANDN U936 ( .A(n772), .B(sreg[410]), .Z(n776) );
  OR U937 ( .A(n774), .B(n773), .Z(n775) );
  AND U938 ( .A(n776), .B(n775), .Z(n778) );
  XOR U939 ( .A(n779), .B(n778), .Z(c[411]) );
  NAND U940 ( .A(b[0]), .B(a[157]), .Z(n782) );
  XOR U941 ( .A(sreg[412]), .B(n782), .Z(n784) );
  NANDN U942 ( .A(n777), .B(sreg[411]), .Z(n781) );
  OR U943 ( .A(n779), .B(n778), .Z(n780) );
  AND U944 ( .A(n781), .B(n780), .Z(n783) );
  XOR U945 ( .A(n784), .B(n783), .Z(c[412]) );
  NAND U946 ( .A(b[0]), .B(a[158]), .Z(n787) );
  XOR U947 ( .A(sreg[413]), .B(n787), .Z(n789) );
  NANDN U948 ( .A(n782), .B(sreg[412]), .Z(n786) );
  OR U949 ( .A(n784), .B(n783), .Z(n785) );
  AND U950 ( .A(n786), .B(n785), .Z(n788) );
  XOR U951 ( .A(n789), .B(n788), .Z(c[413]) );
  NAND U952 ( .A(b[0]), .B(a[159]), .Z(n792) );
  XOR U953 ( .A(sreg[414]), .B(n792), .Z(n794) );
  NANDN U954 ( .A(n787), .B(sreg[413]), .Z(n791) );
  OR U955 ( .A(n789), .B(n788), .Z(n790) );
  AND U956 ( .A(n791), .B(n790), .Z(n793) );
  XOR U957 ( .A(n794), .B(n793), .Z(c[414]) );
  NAND U958 ( .A(b[0]), .B(a[160]), .Z(n797) );
  XOR U959 ( .A(sreg[415]), .B(n797), .Z(n799) );
  NANDN U960 ( .A(n792), .B(sreg[414]), .Z(n796) );
  OR U961 ( .A(n794), .B(n793), .Z(n795) );
  AND U962 ( .A(n796), .B(n795), .Z(n798) );
  XOR U963 ( .A(n799), .B(n798), .Z(c[415]) );
  NAND U964 ( .A(b[0]), .B(a[161]), .Z(n802) );
  XOR U965 ( .A(sreg[416]), .B(n802), .Z(n804) );
  NANDN U966 ( .A(n797), .B(sreg[415]), .Z(n801) );
  OR U967 ( .A(n799), .B(n798), .Z(n800) );
  AND U968 ( .A(n801), .B(n800), .Z(n803) );
  XOR U969 ( .A(n804), .B(n803), .Z(c[416]) );
  NAND U970 ( .A(b[0]), .B(a[162]), .Z(n807) );
  XOR U971 ( .A(sreg[417]), .B(n807), .Z(n809) );
  NANDN U972 ( .A(n802), .B(sreg[416]), .Z(n806) );
  OR U973 ( .A(n804), .B(n803), .Z(n805) );
  AND U974 ( .A(n806), .B(n805), .Z(n808) );
  XOR U975 ( .A(n809), .B(n808), .Z(c[417]) );
  NAND U976 ( .A(b[0]), .B(a[163]), .Z(n812) );
  XOR U977 ( .A(sreg[418]), .B(n812), .Z(n814) );
  NANDN U978 ( .A(n807), .B(sreg[417]), .Z(n811) );
  OR U979 ( .A(n809), .B(n808), .Z(n810) );
  AND U980 ( .A(n811), .B(n810), .Z(n813) );
  XOR U981 ( .A(n814), .B(n813), .Z(c[418]) );
  NAND U982 ( .A(b[0]), .B(a[164]), .Z(n817) );
  XOR U983 ( .A(sreg[419]), .B(n817), .Z(n819) );
  NANDN U984 ( .A(n812), .B(sreg[418]), .Z(n816) );
  OR U985 ( .A(n814), .B(n813), .Z(n815) );
  AND U986 ( .A(n816), .B(n815), .Z(n818) );
  XOR U987 ( .A(n819), .B(n818), .Z(c[419]) );
  NAND U988 ( .A(b[0]), .B(a[165]), .Z(n822) );
  XOR U989 ( .A(sreg[420]), .B(n822), .Z(n824) );
  NANDN U990 ( .A(n817), .B(sreg[419]), .Z(n821) );
  OR U991 ( .A(n819), .B(n818), .Z(n820) );
  AND U992 ( .A(n821), .B(n820), .Z(n823) );
  XOR U993 ( .A(n824), .B(n823), .Z(c[420]) );
  NAND U994 ( .A(b[0]), .B(a[166]), .Z(n827) );
  XOR U995 ( .A(sreg[421]), .B(n827), .Z(n829) );
  NANDN U996 ( .A(n822), .B(sreg[420]), .Z(n826) );
  OR U997 ( .A(n824), .B(n823), .Z(n825) );
  AND U998 ( .A(n826), .B(n825), .Z(n828) );
  XOR U999 ( .A(n829), .B(n828), .Z(c[421]) );
  NAND U1000 ( .A(b[0]), .B(a[167]), .Z(n832) );
  XOR U1001 ( .A(sreg[422]), .B(n832), .Z(n834) );
  NANDN U1002 ( .A(n827), .B(sreg[421]), .Z(n831) );
  OR U1003 ( .A(n829), .B(n828), .Z(n830) );
  AND U1004 ( .A(n831), .B(n830), .Z(n833) );
  XOR U1005 ( .A(n834), .B(n833), .Z(c[422]) );
  NAND U1006 ( .A(b[0]), .B(a[168]), .Z(n837) );
  XOR U1007 ( .A(sreg[423]), .B(n837), .Z(n839) );
  NANDN U1008 ( .A(n832), .B(sreg[422]), .Z(n836) );
  OR U1009 ( .A(n834), .B(n833), .Z(n835) );
  AND U1010 ( .A(n836), .B(n835), .Z(n838) );
  XOR U1011 ( .A(n839), .B(n838), .Z(c[423]) );
  NAND U1012 ( .A(b[0]), .B(a[169]), .Z(n842) );
  XOR U1013 ( .A(sreg[424]), .B(n842), .Z(n844) );
  NANDN U1014 ( .A(n837), .B(sreg[423]), .Z(n841) );
  OR U1015 ( .A(n839), .B(n838), .Z(n840) );
  AND U1016 ( .A(n841), .B(n840), .Z(n843) );
  XOR U1017 ( .A(n844), .B(n843), .Z(c[424]) );
  NAND U1018 ( .A(b[0]), .B(a[170]), .Z(n847) );
  XOR U1019 ( .A(sreg[425]), .B(n847), .Z(n849) );
  NANDN U1020 ( .A(n842), .B(sreg[424]), .Z(n846) );
  OR U1021 ( .A(n844), .B(n843), .Z(n845) );
  AND U1022 ( .A(n846), .B(n845), .Z(n848) );
  XOR U1023 ( .A(n849), .B(n848), .Z(c[425]) );
  NAND U1024 ( .A(b[0]), .B(a[171]), .Z(n852) );
  XOR U1025 ( .A(sreg[426]), .B(n852), .Z(n854) );
  NANDN U1026 ( .A(n847), .B(sreg[425]), .Z(n851) );
  OR U1027 ( .A(n849), .B(n848), .Z(n850) );
  AND U1028 ( .A(n851), .B(n850), .Z(n853) );
  XOR U1029 ( .A(n854), .B(n853), .Z(c[426]) );
  NAND U1030 ( .A(b[0]), .B(a[172]), .Z(n857) );
  XOR U1031 ( .A(sreg[427]), .B(n857), .Z(n859) );
  NANDN U1032 ( .A(n852), .B(sreg[426]), .Z(n856) );
  OR U1033 ( .A(n854), .B(n853), .Z(n855) );
  AND U1034 ( .A(n856), .B(n855), .Z(n858) );
  XOR U1035 ( .A(n859), .B(n858), .Z(c[427]) );
  NAND U1036 ( .A(b[0]), .B(a[173]), .Z(n862) );
  XOR U1037 ( .A(sreg[428]), .B(n862), .Z(n864) );
  NANDN U1038 ( .A(n857), .B(sreg[427]), .Z(n861) );
  OR U1039 ( .A(n859), .B(n858), .Z(n860) );
  AND U1040 ( .A(n861), .B(n860), .Z(n863) );
  XOR U1041 ( .A(n864), .B(n863), .Z(c[428]) );
  NAND U1042 ( .A(b[0]), .B(a[174]), .Z(n867) );
  XOR U1043 ( .A(sreg[429]), .B(n867), .Z(n869) );
  NANDN U1044 ( .A(n862), .B(sreg[428]), .Z(n866) );
  OR U1045 ( .A(n864), .B(n863), .Z(n865) );
  AND U1046 ( .A(n866), .B(n865), .Z(n868) );
  XOR U1047 ( .A(n869), .B(n868), .Z(c[429]) );
  NAND U1048 ( .A(b[0]), .B(a[175]), .Z(n872) );
  XOR U1049 ( .A(sreg[430]), .B(n872), .Z(n874) );
  NANDN U1050 ( .A(n867), .B(sreg[429]), .Z(n871) );
  OR U1051 ( .A(n869), .B(n868), .Z(n870) );
  AND U1052 ( .A(n871), .B(n870), .Z(n873) );
  XOR U1053 ( .A(n874), .B(n873), .Z(c[430]) );
  NAND U1054 ( .A(b[0]), .B(a[176]), .Z(n877) );
  XOR U1055 ( .A(sreg[431]), .B(n877), .Z(n879) );
  NANDN U1056 ( .A(n872), .B(sreg[430]), .Z(n876) );
  OR U1057 ( .A(n874), .B(n873), .Z(n875) );
  AND U1058 ( .A(n876), .B(n875), .Z(n878) );
  XOR U1059 ( .A(n879), .B(n878), .Z(c[431]) );
  NAND U1060 ( .A(b[0]), .B(a[177]), .Z(n882) );
  XOR U1061 ( .A(sreg[432]), .B(n882), .Z(n884) );
  NANDN U1062 ( .A(n877), .B(sreg[431]), .Z(n881) );
  OR U1063 ( .A(n879), .B(n878), .Z(n880) );
  AND U1064 ( .A(n881), .B(n880), .Z(n883) );
  XOR U1065 ( .A(n884), .B(n883), .Z(c[432]) );
  NAND U1066 ( .A(b[0]), .B(a[178]), .Z(n887) );
  XOR U1067 ( .A(sreg[433]), .B(n887), .Z(n889) );
  NANDN U1068 ( .A(n882), .B(sreg[432]), .Z(n886) );
  OR U1069 ( .A(n884), .B(n883), .Z(n885) );
  AND U1070 ( .A(n886), .B(n885), .Z(n888) );
  XOR U1071 ( .A(n889), .B(n888), .Z(c[433]) );
  NAND U1072 ( .A(b[0]), .B(a[179]), .Z(n892) );
  XOR U1073 ( .A(sreg[434]), .B(n892), .Z(n894) );
  NANDN U1074 ( .A(n887), .B(sreg[433]), .Z(n891) );
  OR U1075 ( .A(n889), .B(n888), .Z(n890) );
  AND U1076 ( .A(n891), .B(n890), .Z(n893) );
  XOR U1077 ( .A(n894), .B(n893), .Z(c[434]) );
  NAND U1078 ( .A(b[0]), .B(a[180]), .Z(n897) );
  XOR U1079 ( .A(sreg[435]), .B(n897), .Z(n899) );
  NANDN U1080 ( .A(n892), .B(sreg[434]), .Z(n896) );
  OR U1081 ( .A(n894), .B(n893), .Z(n895) );
  AND U1082 ( .A(n896), .B(n895), .Z(n898) );
  XOR U1083 ( .A(n899), .B(n898), .Z(c[435]) );
  NAND U1084 ( .A(b[0]), .B(a[181]), .Z(n902) );
  XOR U1085 ( .A(sreg[436]), .B(n902), .Z(n904) );
  NANDN U1086 ( .A(n897), .B(sreg[435]), .Z(n901) );
  OR U1087 ( .A(n899), .B(n898), .Z(n900) );
  AND U1088 ( .A(n901), .B(n900), .Z(n903) );
  XOR U1089 ( .A(n904), .B(n903), .Z(c[436]) );
  NAND U1090 ( .A(b[0]), .B(a[182]), .Z(n907) );
  XOR U1091 ( .A(sreg[437]), .B(n907), .Z(n909) );
  NANDN U1092 ( .A(n902), .B(sreg[436]), .Z(n906) );
  OR U1093 ( .A(n904), .B(n903), .Z(n905) );
  AND U1094 ( .A(n906), .B(n905), .Z(n908) );
  XOR U1095 ( .A(n909), .B(n908), .Z(c[437]) );
  NAND U1096 ( .A(b[0]), .B(a[183]), .Z(n912) );
  XOR U1097 ( .A(sreg[438]), .B(n912), .Z(n914) );
  NANDN U1098 ( .A(n907), .B(sreg[437]), .Z(n911) );
  OR U1099 ( .A(n909), .B(n908), .Z(n910) );
  AND U1100 ( .A(n911), .B(n910), .Z(n913) );
  XOR U1101 ( .A(n914), .B(n913), .Z(c[438]) );
  NAND U1102 ( .A(b[0]), .B(a[184]), .Z(n917) );
  XOR U1103 ( .A(sreg[439]), .B(n917), .Z(n919) );
  NANDN U1104 ( .A(n912), .B(sreg[438]), .Z(n916) );
  OR U1105 ( .A(n914), .B(n913), .Z(n915) );
  AND U1106 ( .A(n916), .B(n915), .Z(n918) );
  XOR U1107 ( .A(n919), .B(n918), .Z(c[439]) );
  NAND U1108 ( .A(b[0]), .B(a[185]), .Z(n922) );
  XOR U1109 ( .A(sreg[440]), .B(n922), .Z(n924) );
  NANDN U1110 ( .A(n917), .B(sreg[439]), .Z(n921) );
  OR U1111 ( .A(n919), .B(n918), .Z(n920) );
  AND U1112 ( .A(n921), .B(n920), .Z(n923) );
  XOR U1113 ( .A(n924), .B(n923), .Z(c[440]) );
  NAND U1114 ( .A(b[0]), .B(a[186]), .Z(n927) );
  XOR U1115 ( .A(sreg[441]), .B(n927), .Z(n929) );
  NANDN U1116 ( .A(n922), .B(sreg[440]), .Z(n926) );
  OR U1117 ( .A(n924), .B(n923), .Z(n925) );
  AND U1118 ( .A(n926), .B(n925), .Z(n928) );
  XOR U1119 ( .A(n929), .B(n928), .Z(c[441]) );
  NAND U1120 ( .A(b[0]), .B(a[187]), .Z(n932) );
  XOR U1121 ( .A(sreg[442]), .B(n932), .Z(n934) );
  NANDN U1122 ( .A(n927), .B(sreg[441]), .Z(n931) );
  OR U1123 ( .A(n929), .B(n928), .Z(n930) );
  AND U1124 ( .A(n931), .B(n930), .Z(n933) );
  XOR U1125 ( .A(n934), .B(n933), .Z(c[442]) );
  NAND U1126 ( .A(b[0]), .B(a[188]), .Z(n937) );
  XOR U1127 ( .A(sreg[443]), .B(n937), .Z(n939) );
  NANDN U1128 ( .A(n932), .B(sreg[442]), .Z(n936) );
  OR U1129 ( .A(n934), .B(n933), .Z(n935) );
  AND U1130 ( .A(n936), .B(n935), .Z(n938) );
  XOR U1131 ( .A(n939), .B(n938), .Z(c[443]) );
  NAND U1132 ( .A(b[0]), .B(a[189]), .Z(n942) );
  XOR U1133 ( .A(sreg[444]), .B(n942), .Z(n944) );
  NANDN U1134 ( .A(n937), .B(sreg[443]), .Z(n941) );
  OR U1135 ( .A(n939), .B(n938), .Z(n940) );
  AND U1136 ( .A(n941), .B(n940), .Z(n943) );
  XOR U1137 ( .A(n944), .B(n943), .Z(c[444]) );
  NAND U1138 ( .A(b[0]), .B(a[190]), .Z(n947) );
  XOR U1139 ( .A(sreg[445]), .B(n947), .Z(n949) );
  NANDN U1140 ( .A(n942), .B(sreg[444]), .Z(n946) );
  OR U1141 ( .A(n944), .B(n943), .Z(n945) );
  AND U1142 ( .A(n946), .B(n945), .Z(n948) );
  XOR U1143 ( .A(n949), .B(n948), .Z(c[445]) );
  NAND U1144 ( .A(b[0]), .B(a[191]), .Z(n952) );
  XOR U1145 ( .A(sreg[446]), .B(n952), .Z(n954) );
  NANDN U1146 ( .A(n947), .B(sreg[445]), .Z(n951) );
  OR U1147 ( .A(n949), .B(n948), .Z(n950) );
  AND U1148 ( .A(n951), .B(n950), .Z(n953) );
  XOR U1149 ( .A(n954), .B(n953), .Z(c[446]) );
  NAND U1150 ( .A(b[0]), .B(a[192]), .Z(n957) );
  XOR U1151 ( .A(sreg[447]), .B(n957), .Z(n959) );
  NANDN U1152 ( .A(n952), .B(sreg[446]), .Z(n956) );
  OR U1153 ( .A(n954), .B(n953), .Z(n955) );
  AND U1154 ( .A(n956), .B(n955), .Z(n958) );
  XOR U1155 ( .A(n959), .B(n958), .Z(c[447]) );
  NAND U1156 ( .A(b[0]), .B(a[193]), .Z(n962) );
  XOR U1157 ( .A(sreg[448]), .B(n962), .Z(n964) );
  NANDN U1158 ( .A(n957), .B(sreg[447]), .Z(n961) );
  OR U1159 ( .A(n959), .B(n958), .Z(n960) );
  AND U1160 ( .A(n961), .B(n960), .Z(n963) );
  XOR U1161 ( .A(n964), .B(n963), .Z(c[448]) );
  NAND U1162 ( .A(b[0]), .B(a[194]), .Z(n967) );
  XOR U1163 ( .A(sreg[449]), .B(n967), .Z(n969) );
  NANDN U1164 ( .A(n962), .B(sreg[448]), .Z(n966) );
  OR U1165 ( .A(n964), .B(n963), .Z(n965) );
  AND U1166 ( .A(n966), .B(n965), .Z(n968) );
  XOR U1167 ( .A(n969), .B(n968), .Z(c[449]) );
  NAND U1168 ( .A(b[0]), .B(a[195]), .Z(n972) );
  XOR U1169 ( .A(sreg[450]), .B(n972), .Z(n974) );
  NANDN U1170 ( .A(n967), .B(sreg[449]), .Z(n971) );
  OR U1171 ( .A(n969), .B(n968), .Z(n970) );
  AND U1172 ( .A(n971), .B(n970), .Z(n973) );
  XOR U1173 ( .A(n974), .B(n973), .Z(c[450]) );
  NAND U1174 ( .A(b[0]), .B(a[196]), .Z(n977) );
  XOR U1175 ( .A(sreg[451]), .B(n977), .Z(n979) );
  NANDN U1176 ( .A(n972), .B(sreg[450]), .Z(n976) );
  OR U1177 ( .A(n974), .B(n973), .Z(n975) );
  AND U1178 ( .A(n976), .B(n975), .Z(n978) );
  XOR U1179 ( .A(n979), .B(n978), .Z(c[451]) );
  NAND U1180 ( .A(b[0]), .B(a[197]), .Z(n982) );
  XOR U1181 ( .A(sreg[452]), .B(n982), .Z(n984) );
  NANDN U1182 ( .A(n977), .B(sreg[451]), .Z(n981) );
  OR U1183 ( .A(n979), .B(n978), .Z(n980) );
  AND U1184 ( .A(n981), .B(n980), .Z(n983) );
  XOR U1185 ( .A(n984), .B(n983), .Z(c[452]) );
  NAND U1186 ( .A(b[0]), .B(a[198]), .Z(n987) );
  XOR U1187 ( .A(sreg[453]), .B(n987), .Z(n989) );
  NANDN U1188 ( .A(n982), .B(sreg[452]), .Z(n986) );
  OR U1189 ( .A(n984), .B(n983), .Z(n985) );
  AND U1190 ( .A(n986), .B(n985), .Z(n988) );
  XOR U1191 ( .A(n989), .B(n988), .Z(c[453]) );
  NAND U1192 ( .A(b[0]), .B(a[199]), .Z(n992) );
  XOR U1193 ( .A(sreg[454]), .B(n992), .Z(n994) );
  NANDN U1194 ( .A(n987), .B(sreg[453]), .Z(n991) );
  OR U1195 ( .A(n989), .B(n988), .Z(n990) );
  AND U1196 ( .A(n991), .B(n990), .Z(n993) );
  XOR U1197 ( .A(n994), .B(n993), .Z(c[454]) );
  NAND U1198 ( .A(b[0]), .B(a[200]), .Z(n997) );
  XOR U1199 ( .A(sreg[455]), .B(n997), .Z(n999) );
  NANDN U1200 ( .A(n992), .B(sreg[454]), .Z(n996) );
  OR U1201 ( .A(n994), .B(n993), .Z(n995) );
  AND U1202 ( .A(n996), .B(n995), .Z(n998) );
  XOR U1203 ( .A(n999), .B(n998), .Z(c[455]) );
  NAND U1204 ( .A(b[0]), .B(a[201]), .Z(n1002) );
  XOR U1205 ( .A(sreg[456]), .B(n1002), .Z(n1004) );
  NANDN U1206 ( .A(n997), .B(sreg[455]), .Z(n1001) );
  OR U1207 ( .A(n999), .B(n998), .Z(n1000) );
  AND U1208 ( .A(n1001), .B(n1000), .Z(n1003) );
  XOR U1209 ( .A(n1004), .B(n1003), .Z(c[456]) );
  NAND U1210 ( .A(b[0]), .B(a[202]), .Z(n1007) );
  XOR U1211 ( .A(sreg[457]), .B(n1007), .Z(n1009) );
  NANDN U1212 ( .A(n1002), .B(sreg[456]), .Z(n1006) );
  OR U1213 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U1214 ( .A(n1006), .B(n1005), .Z(n1008) );
  XOR U1215 ( .A(n1009), .B(n1008), .Z(c[457]) );
  NAND U1216 ( .A(b[0]), .B(a[203]), .Z(n1012) );
  XOR U1217 ( .A(sreg[458]), .B(n1012), .Z(n1014) );
  NANDN U1218 ( .A(n1007), .B(sreg[457]), .Z(n1011) );
  OR U1219 ( .A(n1009), .B(n1008), .Z(n1010) );
  AND U1220 ( .A(n1011), .B(n1010), .Z(n1013) );
  XOR U1221 ( .A(n1014), .B(n1013), .Z(c[458]) );
  NAND U1222 ( .A(b[0]), .B(a[204]), .Z(n1017) );
  XOR U1223 ( .A(sreg[459]), .B(n1017), .Z(n1019) );
  NANDN U1224 ( .A(n1012), .B(sreg[458]), .Z(n1016) );
  OR U1225 ( .A(n1014), .B(n1013), .Z(n1015) );
  AND U1226 ( .A(n1016), .B(n1015), .Z(n1018) );
  XOR U1227 ( .A(n1019), .B(n1018), .Z(c[459]) );
  NAND U1228 ( .A(b[0]), .B(a[205]), .Z(n1022) );
  XOR U1229 ( .A(sreg[460]), .B(n1022), .Z(n1024) );
  NANDN U1230 ( .A(n1017), .B(sreg[459]), .Z(n1021) );
  OR U1231 ( .A(n1019), .B(n1018), .Z(n1020) );
  AND U1232 ( .A(n1021), .B(n1020), .Z(n1023) );
  XOR U1233 ( .A(n1024), .B(n1023), .Z(c[460]) );
  NAND U1234 ( .A(b[0]), .B(a[206]), .Z(n1027) );
  XOR U1235 ( .A(sreg[461]), .B(n1027), .Z(n1029) );
  NANDN U1236 ( .A(n1022), .B(sreg[460]), .Z(n1026) );
  OR U1237 ( .A(n1024), .B(n1023), .Z(n1025) );
  AND U1238 ( .A(n1026), .B(n1025), .Z(n1028) );
  XOR U1239 ( .A(n1029), .B(n1028), .Z(c[461]) );
  NAND U1240 ( .A(b[0]), .B(a[207]), .Z(n1032) );
  XOR U1241 ( .A(sreg[462]), .B(n1032), .Z(n1034) );
  NANDN U1242 ( .A(n1027), .B(sreg[461]), .Z(n1031) );
  OR U1243 ( .A(n1029), .B(n1028), .Z(n1030) );
  AND U1244 ( .A(n1031), .B(n1030), .Z(n1033) );
  XOR U1245 ( .A(n1034), .B(n1033), .Z(c[462]) );
  NAND U1246 ( .A(b[0]), .B(a[208]), .Z(n1037) );
  XOR U1247 ( .A(sreg[463]), .B(n1037), .Z(n1039) );
  NANDN U1248 ( .A(n1032), .B(sreg[462]), .Z(n1036) );
  OR U1249 ( .A(n1034), .B(n1033), .Z(n1035) );
  AND U1250 ( .A(n1036), .B(n1035), .Z(n1038) );
  XOR U1251 ( .A(n1039), .B(n1038), .Z(c[463]) );
  NAND U1252 ( .A(b[0]), .B(a[209]), .Z(n1042) );
  XOR U1253 ( .A(sreg[464]), .B(n1042), .Z(n1044) );
  NANDN U1254 ( .A(n1037), .B(sreg[463]), .Z(n1041) );
  OR U1255 ( .A(n1039), .B(n1038), .Z(n1040) );
  AND U1256 ( .A(n1041), .B(n1040), .Z(n1043) );
  XOR U1257 ( .A(n1044), .B(n1043), .Z(c[464]) );
  NAND U1258 ( .A(b[0]), .B(a[210]), .Z(n1047) );
  XOR U1259 ( .A(sreg[465]), .B(n1047), .Z(n1049) );
  NANDN U1260 ( .A(n1042), .B(sreg[464]), .Z(n1046) );
  OR U1261 ( .A(n1044), .B(n1043), .Z(n1045) );
  AND U1262 ( .A(n1046), .B(n1045), .Z(n1048) );
  XOR U1263 ( .A(n1049), .B(n1048), .Z(c[465]) );
  NAND U1264 ( .A(b[0]), .B(a[211]), .Z(n1052) );
  XOR U1265 ( .A(sreg[466]), .B(n1052), .Z(n1054) );
  NANDN U1266 ( .A(n1047), .B(sreg[465]), .Z(n1051) );
  OR U1267 ( .A(n1049), .B(n1048), .Z(n1050) );
  AND U1268 ( .A(n1051), .B(n1050), .Z(n1053) );
  XOR U1269 ( .A(n1054), .B(n1053), .Z(c[466]) );
  NAND U1270 ( .A(b[0]), .B(a[212]), .Z(n1057) );
  XOR U1271 ( .A(sreg[467]), .B(n1057), .Z(n1059) );
  NANDN U1272 ( .A(n1052), .B(sreg[466]), .Z(n1056) );
  OR U1273 ( .A(n1054), .B(n1053), .Z(n1055) );
  AND U1274 ( .A(n1056), .B(n1055), .Z(n1058) );
  XOR U1275 ( .A(n1059), .B(n1058), .Z(c[467]) );
  NAND U1276 ( .A(b[0]), .B(a[213]), .Z(n1062) );
  XOR U1277 ( .A(sreg[468]), .B(n1062), .Z(n1064) );
  NANDN U1278 ( .A(n1057), .B(sreg[467]), .Z(n1061) );
  OR U1279 ( .A(n1059), .B(n1058), .Z(n1060) );
  AND U1280 ( .A(n1061), .B(n1060), .Z(n1063) );
  XOR U1281 ( .A(n1064), .B(n1063), .Z(c[468]) );
  NAND U1282 ( .A(b[0]), .B(a[214]), .Z(n1067) );
  XOR U1283 ( .A(sreg[469]), .B(n1067), .Z(n1069) );
  NANDN U1284 ( .A(n1062), .B(sreg[468]), .Z(n1066) );
  OR U1285 ( .A(n1064), .B(n1063), .Z(n1065) );
  AND U1286 ( .A(n1066), .B(n1065), .Z(n1068) );
  XOR U1287 ( .A(n1069), .B(n1068), .Z(c[469]) );
  NAND U1288 ( .A(b[0]), .B(a[215]), .Z(n1072) );
  XOR U1289 ( .A(sreg[470]), .B(n1072), .Z(n1074) );
  NANDN U1290 ( .A(n1067), .B(sreg[469]), .Z(n1071) );
  OR U1291 ( .A(n1069), .B(n1068), .Z(n1070) );
  AND U1292 ( .A(n1071), .B(n1070), .Z(n1073) );
  XOR U1293 ( .A(n1074), .B(n1073), .Z(c[470]) );
  NAND U1294 ( .A(b[0]), .B(a[216]), .Z(n1077) );
  XOR U1295 ( .A(sreg[471]), .B(n1077), .Z(n1079) );
  NANDN U1296 ( .A(n1072), .B(sreg[470]), .Z(n1076) );
  OR U1297 ( .A(n1074), .B(n1073), .Z(n1075) );
  AND U1298 ( .A(n1076), .B(n1075), .Z(n1078) );
  XOR U1299 ( .A(n1079), .B(n1078), .Z(c[471]) );
  NAND U1300 ( .A(b[0]), .B(a[217]), .Z(n1082) );
  XOR U1301 ( .A(sreg[472]), .B(n1082), .Z(n1084) );
  NANDN U1302 ( .A(n1077), .B(sreg[471]), .Z(n1081) );
  OR U1303 ( .A(n1079), .B(n1078), .Z(n1080) );
  AND U1304 ( .A(n1081), .B(n1080), .Z(n1083) );
  XOR U1305 ( .A(n1084), .B(n1083), .Z(c[472]) );
  NAND U1306 ( .A(b[0]), .B(a[218]), .Z(n1087) );
  XOR U1307 ( .A(sreg[473]), .B(n1087), .Z(n1089) );
  NANDN U1308 ( .A(n1082), .B(sreg[472]), .Z(n1086) );
  OR U1309 ( .A(n1084), .B(n1083), .Z(n1085) );
  AND U1310 ( .A(n1086), .B(n1085), .Z(n1088) );
  XOR U1311 ( .A(n1089), .B(n1088), .Z(c[473]) );
  NAND U1312 ( .A(b[0]), .B(a[219]), .Z(n1092) );
  XOR U1313 ( .A(sreg[474]), .B(n1092), .Z(n1094) );
  NANDN U1314 ( .A(n1087), .B(sreg[473]), .Z(n1091) );
  OR U1315 ( .A(n1089), .B(n1088), .Z(n1090) );
  AND U1316 ( .A(n1091), .B(n1090), .Z(n1093) );
  XOR U1317 ( .A(n1094), .B(n1093), .Z(c[474]) );
  NAND U1318 ( .A(b[0]), .B(a[220]), .Z(n1097) );
  XOR U1319 ( .A(sreg[475]), .B(n1097), .Z(n1099) );
  NANDN U1320 ( .A(n1092), .B(sreg[474]), .Z(n1096) );
  OR U1321 ( .A(n1094), .B(n1093), .Z(n1095) );
  AND U1322 ( .A(n1096), .B(n1095), .Z(n1098) );
  XOR U1323 ( .A(n1099), .B(n1098), .Z(c[475]) );
  NAND U1324 ( .A(b[0]), .B(a[221]), .Z(n1102) );
  XOR U1325 ( .A(sreg[476]), .B(n1102), .Z(n1104) );
  NANDN U1326 ( .A(n1097), .B(sreg[475]), .Z(n1101) );
  OR U1327 ( .A(n1099), .B(n1098), .Z(n1100) );
  AND U1328 ( .A(n1101), .B(n1100), .Z(n1103) );
  XOR U1329 ( .A(n1104), .B(n1103), .Z(c[476]) );
  NAND U1330 ( .A(b[0]), .B(a[222]), .Z(n1107) );
  XOR U1331 ( .A(sreg[477]), .B(n1107), .Z(n1109) );
  NANDN U1332 ( .A(n1102), .B(sreg[476]), .Z(n1106) );
  OR U1333 ( .A(n1104), .B(n1103), .Z(n1105) );
  AND U1334 ( .A(n1106), .B(n1105), .Z(n1108) );
  XOR U1335 ( .A(n1109), .B(n1108), .Z(c[477]) );
  NAND U1336 ( .A(b[0]), .B(a[223]), .Z(n1112) );
  XOR U1337 ( .A(sreg[478]), .B(n1112), .Z(n1114) );
  NANDN U1338 ( .A(n1107), .B(sreg[477]), .Z(n1111) );
  OR U1339 ( .A(n1109), .B(n1108), .Z(n1110) );
  AND U1340 ( .A(n1111), .B(n1110), .Z(n1113) );
  XOR U1341 ( .A(n1114), .B(n1113), .Z(c[478]) );
  NAND U1342 ( .A(b[0]), .B(a[224]), .Z(n1117) );
  XOR U1343 ( .A(sreg[479]), .B(n1117), .Z(n1119) );
  NANDN U1344 ( .A(n1112), .B(sreg[478]), .Z(n1116) );
  OR U1345 ( .A(n1114), .B(n1113), .Z(n1115) );
  AND U1346 ( .A(n1116), .B(n1115), .Z(n1118) );
  XOR U1347 ( .A(n1119), .B(n1118), .Z(c[479]) );
  NAND U1348 ( .A(b[0]), .B(a[225]), .Z(n1122) );
  XOR U1349 ( .A(sreg[480]), .B(n1122), .Z(n1124) );
  NANDN U1350 ( .A(n1117), .B(sreg[479]), .Z(n1121) );
  OR U1351 ( .A(n1119), .B(n1118), .Z(n1120) );
  AND U1352 ( .A(n1121), .B(n1120), .Z(n1123) );
  XOR U1353 ( .A(n1124), .B(n1123), .Z(c[480]) );
  NAND U1354 ( .A(b[0]), .B(a[226]), .Z(n1127) );
  XOR U1355 ( .A(sreg[481]), .B(n1127), .Z(n1129) );
  NANDN U1356 ( .A(n1122), .B(sreg[480]), .Z(n1126) );
  OR U1357 ( .A(n1124), .B(n1123), .Z(n1125) );
  AND U1358 ( .A(n1126), .B(n1125), .Z(n1128) );
  XOR U1359 ( .A(n1129), .B(n1128), .Z(c[481]) );
  NAND U1360 ( .A(b[0]), .B(a[227]), .Z(n1132) );
  XOR U1361 ( .A(sreg[482]), .B(n1132), .Z(n1134) );
  NANDN U1362 ( .A(n1127), .B(sreg[481]), .Z(n1131) );
  OR U1363 ( .A(n1129), .B(n1128), .Z(n1130) );
  AND U1364 ( .A(n1131), .B(n1130), .Z(n1133) );
  XOR U1365 ( .A(n1134), .B(n1133), .Z(c[482]) );
  NAND U1366 ( .A(b[0]), .B(a[228]), .Z(n1137) );
  XOR U1367 ( .A(sreg[483]), .B(n1137), .Z(n1139) );
  NANDN U1368 ( .A(n1132), .B(sreg[482]), .Z(n1136) );
  OR U1369 ( .A(n1134), .B(n1133), .Z(n1135) );
  AND U1370 ( .A(n1136), .B(n1135), .Z(n1138) );
  XOR U1371 ( .A(n1139), .B(n1138), .Z(c[483]) );
  NAND U1372 ( .A(b[0]), .B(a[229]), .Z(n1142) );
  XOR U1373 ( .A(sreg[484]), .B(n1142), .Z(n1144) );
  NANDN U1374 ( .A(n1137), .B(sreg[483]), .Z(n1141) );
  OR U1375 ( .A(n1139), .B(n1138), .Z(n1140) );
  AND U1376 ( .A(n1141), .B(n1140), .Z(n1143) );
  XOR U1377 ( .A(n1144), .B(n1143), .Z(c[484]) );
  NAND U1378 ( .A(b[0]), .B(a[230]), .Z(n1147) );
  XOR U1379 ( .A(sreg[485]), .B(n1147), .Z(n1149) );
  NANDN U1380 ( .A(n1142), .B(sreg[484]), .Z(n1146) );
  OR U1381 ( .A(n1144), .B(n1143), .Z(n1145) );
  AND U1382 ( .A(n1146), .B(n1145), .Z(n1148) );
  XOR U1383 ( .A(n1149), .B(n1148), .Z(c[485]) );
  NAND U1384 ( .A(b[0]), .B(a[231]), .Z(n1152) );
  XOR U1385 ( .A(sreg[486]), .B(n1152), .Z(n1154) );
  NANDN U1386 ( .A(n1147), .B(sreg[485]), .Z(n1151) );
  OR U1387 ( .A(n1149), .B(n1148), .Z(n1150) );
  AND U1388 ( .A(n1151), .B(n1150), .Z(n1153) );
  XOR U1389 ( .A(n1154), .B(n1153), .Z(c[486]) );
  NAND U1390 ( .A(b[0]), .B(a[232]), .Z(n1157) );
  XOR U1391 ( .A(sreg[487]), .B(n1157), .Z(n1159) );
  NANDN U1392 ( .A(n1152), .B(sreg[486]), .Z(n1156) );
  OR U1393 ( .A(n1154), .B(n1153), .Z(n1155) );
  AND U1394 ( .A(n1156), .B(n1155), .Z(n1158) );
  XOR U1395 ( .A(n1159), .B(n1158), .Z(c[487]) );
  NAND U1396 ( .A(b[0]), .B(a[233]), .Z(n1162) );
  XOR U1397 ( .A(sreg[488]), .B(n1162), .Z(n1164) );
  NANDN U1398 ( .A(n1157), .B(sreg[487]), .Z(n1161) );
  OR U1399 ( .A(n1159), .B(n1158), .Z(n1160) );
  AND U1400 ( .A(n1161), .B(n1160), .Z(n1163) );
  XOR U1401 ( .A(n1164), .B(n1163), .Z(c[488]) );
  NAND U1402 ( .A(b[0]), .B(a[234]), .Z(n1167) );
  XOR U1403 ( .A(sreg[489]), .B(n1167), .Z(n1169) );
  NANDN U1404 ( .A(n1162), .B(sreg[488]), .Z(n1166) );
  OR U1405 ( .A(n1164), .B(n1163), .Z(n1165) );
  AND U1406 ( .A(n1166), .B(n1165), .Z(n1168) );
  XOR U1407 ( .A(n1169), .B(n1168), .Z(c[489]) );
  NAND U1408 ( .A(b[0]), .B(a[235]), .Z(n1172) );
  XOR U1409 ( .A(sreg[490]), .B(n1172), .Z(n1174) );
  NANDN U1410 ( .A(n1167), .B(sreg[489]), .Z(n1171) );
  OR U1411 ( .A(n1169), .B(n1168), .Z(n1170) );
  AND U1412 ( .A(n1171), .B(n1170), .Z(n1173) );
  XOR U1413 ( .A(n1174), .B(n1173), .Z(c[490]) );
  NAND U1414 ( .A(b[0]), .B(a[236]), .Z(n1177) );
  XOR U1415 ( .A(sreg[491]), .B(n1177), .Z(n1179) );
  NANDN U1416 ( .A(n1172), .B(sreg[490]), .Z(n1176) );
  OR U1417 ( .A(n1174), .B(n1173), .Z(n1175) );
  AND U1418 ( .A(n1176), .B(n1175), .Z(n1178) );
  XOR U1419 ( .A(n1179), .B(n1178), .Z(c[491]) );
  NAND U1420 ( .A(b[0]), .B(a[237]), .Z(n1182) );
  XOR U1421 ( .A(sreg[492]), .B(n1182), .Z(n1184) );
  NANDN U1422 ( .A(n1177), .B(sreg[491]), .Z(n1181) );
  OR U1423 ( .A(n1179), .B(n1178), .Z(n1180) );
  AND U1424 ( .A(n1181), .B(n1180), .Z(n1183) );
  XOR U1425 ( .A(n1184), .B(n1183), .Z(c[492]) );
  NAND U1426 ( .A(b[0]), .B(a[238]), .Z(n1187) );
  XOR U1427 ( .A(sreg[493]), .B(n1187), .Z(n1189) );
  NANDN U1428 ( .A(n1182), .B(sreg[492]), .Z(n1186) );
  OR U1429 ( .A(n1184), .B(n1183), .Z(n1185) );
  AND U1430 ( .A(n1186), .B(n1185), .Z(n1188) );
  XOR U1431 ( .A(n1189), .B(n1188), .Z(c[493]) );
  NAND U1432 ( .A(b[0]), .B(a[239]), .Z(n1192) );
  XOR U1433 ( .A(sreg[494]), .B(n1192), .Z(n1194) );
  NANDN U1434 ( .A(n1187), .B(sreg[493]), .Z(n1191) );
  OR U1435 ( .A(n1189), .B(n1188), .Z(n1190) );
  AND U1436 ( .A(n1191), .B(n1190), .Z(n1193) );
  XOR U1437 ( .A(n1194), .B(n1193), .Z(c[494]) );
  NAND U1438 ( .A(b[0]), .B(a[240]), .Z(n1197) );
  XOR U1439 ( .A(sreg[495]), .B(n1197), .Z(n1199) );
  NANDN U1440 ( .A(n1192), .B(sreg[494]), .Z(n1196) );
  OR U1441 ( .A(n1194), .B(n1193), .Z(n1195) );
  AND U1442 ( .A(n1196), .B(n1195), .Z(n1198) );
  XOR U1443 ( .A(n1199), .B(n1198), .Z(c[495]) );
  NAND U1444 ( .A(b[0]), .B(a[241]), .Z(n1202) );
  XOR U1445 ( .A(sreg[496]), .B(n1202), .Z(n1204) );
  NANDN U1446 ( .A(n1197), .B(sreg[495]), .Z(n1201) );
  OR U1447 ( .A(n1199), .B(n1198), .Z(n1200) );
  AND U1448 ( .A(n1201), .B(n1200), .Z(n1203) );
  XOR U1449 ( .A(n1204), .B(n1203), .Z(c[496]) );
  NAND U1450 ( .A(b[0]), .B(a[242]), .Z(n1207) );
  XOR U1451 ( .A(sreg[497]), .B(n1207), .Z(n1209) );
  NANDN U1452 ( .A(n1202), .B(sreg[496]), .Z(n1206) );
  OR U1453 ( .A(n1204), .B(n1203), .Z(n1205) );
  AND U1454 ( .A(n1206), .B(n1205), .Z(n1208) );
  XOR U1455 ( .A(n1209), .B(n1208), .Z(c[497]) );
  NAND U1456 ( .A(b[0]), .B(a[243]), .Z(n1212) );
  XOR U1457 ( .A(sreg[498]), .B(n1212), .Z(n1214) );
  NANDN U1458 ( .A(n1207), .B(sreg[497]), .Z(n1211) );
  OR U1459 ( .A(n1209), .B(n1208), .Z(n1210) );
  AND U1460 ( .A(n1211), .B(n1210), .Z(n1213) );
  XOR U1461 ( .A(n1214), .B(n1213), .Z(c[498]) );
  NAND U1462 ( .A(b[0]), .B(a[244]), .Z(n1217) );
  XOR U1463 ( .A(sreg[499]), .B(n1217), .Z(n1219) );
  NANDN U1464 ( .A(n1212), .B(sreg[498]), .Z(n1216) );
  OR U1465 ( .A(n1214), .B(n1213), .Z(n1215) );
  AND U1466 ( .A(n1216), .B(n1215), .Z(n1218) );
  XOR U1467 ( .A(n1219), .B(n1218), .Z(c[499]) );
  NAND U1468 ( .A(b[0]), .B(a[245]), .Z(n1222) );
  XOR U1469 ( .A(sreg[500]), .B(n1222), .Z(n1224) );
  NANDN U1470 ( .A(n1217), .B(sreg[499]), .Z(n1221) );
  OR U1471 ( .A(n1219), .B(n1218), .Z(n1220) );
  AND U1472 ( .A(n1221), .B(n1220), .Z(n1223) );
  XOR U1473 ( .A(n1224), .B(n1223), .Z(c[500]) );
  NAND U1474 ( .A(b[0]), .B(a[246]), .Z(n1227) );
  XOR U1475 ( .A(sreg[501]), .B(n1227), .Z(n1229) );
  NANDN U1476 ( .A(n1222), .B(sreg[500]), .Z(n1226) );
  OR U1477 ( .A(n1224), .B(n1223), .Z(n1225) );
  AND U1478 ( .A(n1226), .B(n1225), .Z(n1228) );
  XOR U1479 ( .A(n1229), .B(n1228), .Z(c[501]) );
  NAND U1480 ( .A(b[0]), .B(a[247]), .Z(n1232) );
  XOR U1481 ( .A(sreg[502]), .B(n1232), .Z(n1234) );
  NANDN U1482 ( .A(n1227), .B(sreg[501]), .Z(n1231) );
  OR U1483 ( .A(n1229), .B(n1228), .Z(n1230) );
  AND U1484 ( .A(n1231), .B(n1230), .Z(n1233) );
  XOR U1485 ( .A(n1234), .B(n1233), .Z(c[502]) );
  NAND U1486 ( .A(b[0]), .B(a[248]), .Z(n1237) );
  XOR U1487 ( .A(sreg[503]), .B(n1237), .Z(n1239) );
  NANDN U1488 ( .A(n1232), .B(sreg[502]), .Z(n1236) );
  OR U1489 ( .A(n1234), .B(n1233), .Z(n1235) );
  AND U1490 ( .A(n1236), .B(n1235), .Z(n1238) );
  XOR U1491 ( .A(n1239), .B(n1238), .Z(c[503]) );
  NAND U1492 ( .A(b[0]), .B(a[249]), .Z(n1242) );
  XOR U1493 ( .A(sreg[504]), .B(n1242), .Z(n1244) );
  NANDN U1494 ( .A(n1237), .B(sreg[503]), .Z(n1241) );
  OR U1495 ( .A(n1239), .B(n1238), .Z(n1240) );
  AND U1496 ( .A(n1241), .B(n1240), .Z(n1243) );
  XOR U1497 ( .A(n1244), .B(n1243), .Z(c[504]) );
  NAND U1498 ( .A(b[0]), .B(a[250]), .Z(n1247) );
  XOR U1499 ( .A(sreg[505]), .B(n1247), .Z(n1249) );
  NANDN U1500 ( .A(n1242), .B(sreg[504]), .Z(n1246) );
  OR U1501 ( .A(n1244), .B(n1243), .Z(n1245) );
  AND U1502 ( .A(n1246), .B(n1245), .Z(n1248) );
  XOR U1503 ( .A(n1249), .B(n1248), .Z(c[505]) );
  NAND U1504 ( .A(b[0]), .B(a[251]), .Z(n1252) );
  XOR U1505 ( .A(sreg[506]), .B(n1252), .Z(n1254) );
  NANDN U1506 ( .A(n1247), .B(sreg[505]), .Z(n1251) );
  OR U1507 ( .A(n1249), .B(n1248), .Z(n1250) );
  AND U1508 ( .A(n1251), .B(n1250), .Z(n1253) );
  XOR U1509 ( .A(n1254), .B(n1253), .Z(c[506]) );
  NAND U1510 ( .A(b[0]), .B(a[252]), .Z(n1257) );
  XOR U1511 ( .A(sreg[507]), .B(n1257), .Z(n1259) );
  NANDN U1512 ( .A(n1252), .B(sreg[506]), .Z(n1256) );
  OR U1513 ( .A(n1254), .B(n1253), .Z(n1255) );
  AND U1514 ( .A(n1256), .B(n1255), .Z(n1258) );
  XOR U1515 ( .A(n1259), .B(n1258), .Z(c[507]) );
  NAND U1516 ( .A(b[0]), .B(a[253]), .Z(n1262) );
  XOR U1517 ( .A(sreg[508]), .B(n1262), .Z(n1264) );
  NANDN U1518 ( .A(n1257), .B(sreg[507]), .Z(n1261) );
  OR U1519 ( .A(n1259), .B(n1258), .Z(n1260) );
  AND U1520 ( .A(n1261), .B(n1260), .Z(n1263) );
  XOR U1521 ( .A(n1264), .B(n1263), .Z(c[508]) );
  NAND U1522 ( .A(b[0]), .B(a[254]), .Z(n1267) );
  XOR U1523 ( .A(sreg[509]), .B(n1267), .Z(n1269) );
  NANDN U1524 ( .A(n1262), .B(sreg[508]), .Z(n1266) );
  OR U1525 ( .A(n1264), .B(n1263), .Z(n1265) );
  AND U1526 ( .A(n1266), .B(n1265), .Z(n1268) );
  XOR U1527 ( .A(n1269), .B(n1268), .Z(c[509]) );
  NANDN U1528 ( .A(n1267), .B(sreg[509]), .Z(n1271) );
  OR U1529 ( .A(n1269), .B(n1268), .Z(n1270) );
  AND U1530 ( .A(n1271), .B(n1270), .Z(n1275) );
  AND U1531 ( .A(a[255]), .B(b[0]), .Z(n1273) );
  XNOR U1532 ( .A(sreg[510]), .B(n1273), .Z(n1272) );
  XOR U1533 ( .A(n1275), .B(n1272), .Z(c[510]) );
  NAND U1534 ( .A(sreg[510]), .B(n1273), .Z(n1277) );
  XOR U1535 ( .A(n1273), .B(sreg[510]), .Z(n1274) );
  NANDN U1536 ( .A(n1275), .B(n1274), .Z(n1276) );
  NAND U1537 ( .A(n1277), .B(n1276), .Z(c[511]) );
endmodule

