
module hamming_N160_CC2 ( clk, rst, x, y, o );
  input [79:0] x;
  input [79:0] y;
  output [7:0] o;
  input clk, rst;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457;
  wire   [7:0] oglobal;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[7]) );
  XOR U92 ( .A(n361), .B(n360), .Z(n358) );
  XOR U93 ( .A(n317), .B(n316), .Z(n314) );
  XOR U94 ( .A(n449), .B(n448), .Z(n446) );
  XOR U95 ( .A(n375), .B(n374), .Z(n385) );
  XNOR U96 ( .A(n212), .B(n326), .Z(n185) );
  XOR U97 ( .A(n159), .B(n161), .Z(n180) );
  XOR U98 ( .A(n337), .B(n336), .Z(n357) );
  XOR U99 ( .A(n427), .B(n426), .Z(n445) );
  XOR U100 ( .A(n406), .B(n405), .Z(n384) );
  XOR U101 ( .A(n91), .B(n93), .Z(n112) );
  XOR U102 ( .A(n241), .B(n243), .Z(n277) );
  XOR U103 ( .A(n314), .B(n313), .Z(n346) );
  XNOR U104 ( .A(n74), .B(n113), .Z(n75) );
  XOR U105 ( .A(oglobal[7]), .B(n10), .Z(o[7]) );
  NAND U106 ( .A(n11), .B(n12), .Z(n10) );
  NANDN U107 ( .A(n13), .B(oglobal[6]), .Z(n12) );
  NANDN U108 ( .A(n14), .B(oglobal[6]), .Z(n11) );
  XNOR U109 ( .A(n13), .B(n15), .Z(o[6]) );
  XNOR U110 ( .A(oglobal[6]), .B(n14), .Z(n15) );
  AND U111 ( .A(n16), .B(n17), .Z(n14) );
  NANDN U112 ( .A(n18), .B(oglobal[5]), .Z(n17) );
  NAND U113 ( .A(n19), .B(n20), .Z(n16) );
  NAND U114 ( .A(n21), .B(n18), .Z(n19) );
  OR U115 ( .A(n22), .B(n23), .Z(n13) );
  XNOR U116 ( .A(n20), .B(n24), .Z(o[5]) );
  XNOR U117 ( .A(n21), .B(n18), .Z(n24) );
  AND U118 ( .A(n25), .B(n26), .Z(n18) );
  NANDN U119 ( .A(n27), .B(oglobal[4]), .Z(n26) );
  NAND U120 ( .A(n28), .B(n29), .Z(n25) );
  NANDN U121 ( .A(oglobal[4]), .B(n27), .Z(n28) );
  IV U122 ( .A(oglobal[5]), .Z(n21) );
  XOR U123 ( .A(n22), .B(n23), .Z(n20) );
  AND U124 ( .A(n30), .B(n31), .Z(n23) );
  OR U125 ( .A(n32), .B(n33), .Z(n31) );
  XOR U126 ( .A(n34), .B(n35), .Z(n30) );
  ANDN U127 ( .B(n36), .A(n37), .Z(n34) );
  XOR U128 ( .A(n38), .B(n39), .Z(n36) );
  OR U129 ( .A(n40), .B(n41), .Z(n22) );
  XOR U130 ( .A(n29), .B(n42), .Z(o[4]) );
  XNOR U131 ( .A(oglobal[4]), .B(n27), .Z(n42) );
  AND U132 ( .A(n43), .B(n44), .Z(n27) );
  NANDN U133 ( .A(n45), .B(oglobal[3]), .Z(n44) );
  NANDN U134 ( .A(n46), .B(n47), .Z(n43) );
  NANDN U135 ( .A(oglobal[3]), .B(n45), .Z(n47) );
  XNOR U136 ( .A(n37), .B(n39), .Z(n29) );
  XOR U137 ( .A(n40), .B(n41), .Z(n39) );
  AND U138 ( .A(n48), .B(n49), .Z(n41) );
  OR U139 ( .A(n50), .B(n51), .Z(n49) );
  XOR U140 ( .A(n52), .B(n53), .Z(n48) );
  ANDN U141 ( .B(n54), .A(n55), .Z(n52) );
  XOR U142 ( .A(n56), .B(n57), .Z(n54) );
  OR U143 ( .A(n58), .B(n59), .Z(n40) );
  XOR U144 ( .A(n35), .B(n60), .Z(n37) );
  XOR U145 ( .A(n32), .B(n33), .Z(n60) );
  AND U146 ( .A(n61), .B(n62), .Z(n33) );
  OR U147 ( .A(n63), .B(n64), .Z(n62) );
  XOR U148 ( .A(n65), .B(n66), .Z(n61) );
  ANDN U149 ( .B(n67), .A(n68), .Z(n65) );
  XNOR U150 ( .A(n69), .B(n70), .Z(n67) );
  OR U151 ( .A(n71), .B(n72), .Z(n32) );
  IV U152 ( .A(n38), .Z(n35) );
  XOR U153 ( .A(n73), .B(n74), .Z(n38) );
  AND U154 ( .A(n75), .B(n76), .Z(n73) );
  XOR U155 ( .A(n74), .B(n77), .Z(n76) );
  XNOR U156 ( .A(n46), .B(n78), .Z(o[3]) );
  XNOR U157 ( .A(oglobal[3]), .B(n45), .Z(n78) );
  AND U158 ( .A(n79), .B(n80), .Z(n45) );
  NANDN U159 ( .A(n81), .B(oglobal[2]), .Z(n80) );
  NANDN U160 ( .A(n82), .B(n83), .Z(n79) );
  NANDN U161 ( .A(oglobal[2]), .B(n81), .Z(n83) );
  XNOR U162 ( .A(n75), .B(n77), .Z(n46) );
  XNOR U163 ( .A(n55), .B(n57), .Z(n77) );
  XOR U164 ( .A(n58), .B(n59), .Z(n57) );
  AND U165 ( .A(n84), .B(n85), .Z(n59) );
  OR U166 ( .A(n86), .B(n87), .Z(n85) );
  XOR U167 ( .A(n88), .B(n89), .Z(n84) );
  AND U168 ( .A(n90), .B(n91), .Z(n88) );
  XOR U169 ( .A(n92), .B(n93), .Z(n90) );
  OR U170 ( .A(n94), .B(n95), .Z(n58) );
  XOR U171 ( .A(n53), .B(n96), .Z(n55) );
  XOR U172 ( .A(n50), .B(n51), .Z(n96) );
  AND U173 ( .A(n97), .B(n98), .Z(n51) );
  OR U174 ( .A(n99), .B(n100), .Z(n98) );
  XOR U175 ( .A(n101), .B(n102), .Z(n97) );
  AND U176 ( .A(n103), .B(n104), .Z(n101) );
  XNOR U177 ( .A(n105), .B(n102), .Z(n104) );
  OR U178 ( .A(n106), .B(n107), .Z(n50) );
  IV U179 ( .A(n56), .Z(n53) );
  XNOR U180 ( .A(n108), .B(n109), .Z(n56) );
  AND U181 ( .A(n110), .B(n111), .Z(n108) );
  XNOR U182 ( .A(n109), .B(n112), .Z(n111) );
  XNOR U183 ( .A(n68), .B(n70), .Z(n113) );
  XNOR U184 ( .A(n71), .B(n72), .Z(n70) );
  AND U185 ( .A(n114), .B(n115), .Z(n72) );
  OR U186 ( .A(n116), .B(n117), .Z(n115) );
  XOR U187 ( .A(n118), .B(n119), .Z(n114) );
  AND U188 ( .A(n120), .B(n121), .Z(n118) );
  XOR U189 ( .A(n119), .B(n122), .Z(n121) );
  OR U190 ( .A(n123), .B(n124), .Z(n71) );
  XOR U191 ( .A(n66), .B(n125), .Z(n68) );
  XOR U192 ( .A(n63), .B(n64), .Z(n125) );
  AND U193 ( .A(n126), .B(n127), .Z(n64) );
  OR U194 ( .A(n128), .B(n129), .Z(n127) );
  XOR U195 ( .A(n130), .B(n131), .Z(n126) );
  ANDN U196 ( .B(n132), .A(n133), .Z(n130) );
  XOR U197 ( .A(n131), .B(n134), .Z(n132) );
  OR U198 ( .A(n135), .B(n136), .Z(n63) );
  IV U199 ( .A(n69), .Z(n66) );
  XNOR U200 ( .A(n137), .B(n138), .Z(n69) );
  AND U201 ( .A(n139), .B(n140), .Z(n137) );
  XOR U202 ( .A(n138), .B(n141), .Z(n140) );
  XNOR U203 ( .A(n142), .B(n143), .Z(n74) );
  ANDN U204 ( .B(n144), .A(n145), .Z(n142) );
  XNOR U205 ( .A(n143), .B(n146), .Z(n144) );
  XNOR U206 ( .A(n82), .B(n147), .Z(o[2]) );
  XNOR U207 ( .A(oglobal[2]), .B(n81), .Z(n147) );
  AND U208 ( .A(n148), .B(n149), .Z(n81) );
  NANDN U209 ( .A(n150), .B(oglobal[1]), .Z(n149) );
  NANDN U210 ( .A(n151), .B(n152), .Z(n148) );
  NANDN U211 ( .A(oglobal[1]), .B(n150), .Z(n152) );
  XOR U212 ( .A(n145), .B(n146), .Z(n82) );
  XOR U213 ( .A(n110), .B(n112), .Z(n146) );
  XOR U214 ( .A(n94), .B(n95), .Z(n93) );
  AND U215 ( .A(n153), .B(n154), .Z(n95) );
  OR U216 ( .A(n155), .B(n156), .Z(n154) );
  XOR U217 ( .A(n157), .B(n158), .Z(n153) );
  NAND U218 ( .A(n159), .B(n160), .Z(n158) );
  XOR U219 ( .A(n157), .B(n161), .Z(n160) );
  OR U220 ( .A(n162), .B(n163), .Z(n94) );
  XOR U221 ( .A(n92), .B(n164), .Z(n91) );
  XOR U222 ( .A(n86), .B(n87), .Z(n164) );
  AND U223 ( .A(n165), .B(n166), .Z(n87) );
  OR U224 ( .A(n167), .B(n168), .Z(n166) );
  XOR U225 ( .A(n169), .B(n170), .Z(n165) );
  NAND U226 ( .A(n171), .B(n172), .Z(n170) );
  XNOR U227 ( .A(n169), .B(n173), .Z(n171) );
  OR U228 ( .A(n174), .B(n175), .Z(n86) );
  IV U229 ( .A(n89), .Z(n92) );
  XOR U230 ( .A(n176), .B(n177), .Z(n89) );
  NAND U231 ( .A(n178), .B(n179), .Z(n177) );
  XOR U232 ( .A(n176), .B(n180), .Z(n178) );
  XOR U233 ( .A(n103), .B(n181), .Z(n110) );
  XNOR U234 ( .A(n105), .B(n109), .Z(n181) );
  XNOR U235 ( .A(n182), .B(n183), .Z(n109) );
  NAND U236 ( .A(n184), .B(n185), .Z(n183) );
  XNOR U237 ( .A(n182), .B(n186), .Z(n184) );
  XOR U238 ( .A(n106), .B(n107), .Z(n105) );
  AND U239 ( .A(n187), .B(n188), .Z(n107) );
  OR U240 ( .A(n189), .B(n190), .Z(n188) );
  XOR U241 ( .A(n191), .B(n192), .Z(n187) );
  NAND U242 ( .A(n193), .B(n194), .Z(n192) );
  XNOR U243 ( .A(n191), .B(n195), .Z(n193) );
  OR U244 ( .A(n196), .B(n197), .Z(n106) );
  XNOR U245 ( .A(n102), .B(n198), .Z(n103) );
  XOR U246 ( .A(n99), .B(n100), .Z(n198) );
  AND U247 ( .A(n199), .B(n200), .Z(n100) );
  OR U248 ( .A(n201), .B(n202), .Z(n200) );
  XOR U249 ( .A(n203), .B(n204), .Z(n199) );
  NAND U250 ( .A(n205), .B(n206), .Z(n204) );
  XNOR U251 ( .A(n203), .B(n207), .Z(n205) );
  OR U252 ( .A(n208), .B(n209), .Z(n99) );
  XNOR U253 ( .A(n210), .B(n211), .Z(n102) );
  NAND U254 ( .A(n212), .B(n213), .Z(n211) );
  XOR U255 ( .A(n210), .B(n214), .Z(n213) );
  XNOR U256 ( .A(n143), .B(n215), .Z(n145) );
  XOR U257 ( .A(n139), .B(n141), .Z(n215) );
  XOR U258 ( .A(n120), .B(n122), .Z(n141) );
  XNOR U259 ( .A(n123), .B(n124), .Z(n122) );
  AND U260 ( .A(n216), .B(n217), .Z(n124) );
  OR U261 ( .A(n218), .B(n219), .Z(n217) );
  XOR U262 ( .A(n220), .B(n221), .Z(n216) );
  NAND U263 ( .A(n222), .B(n223), .Z(n221) );
  XNOR U264 ( .A(n220), .B(n224), .Z(n222) );
  OR U265 ( .A(n225), .B(n226), .Z(n123) );
  XNOR U266 ( .A(n119), .B(n227), .Z(n120) );
  XOR U267 ( .A(n116), .B(n117), .Z(n227) );
  AND U268 ( .A(n228), .B(n229), .Z(n117) );
  OR U269 ( .A(n230), .B(n231), .Z(n229) );
  XOR U270 ( .A(n232), .B(n233), .Z(n228) );
  NAND U271 ( .A(n234), .B(n235), .Z(n233) );
  XNOR U272 ( .A(n232), .B(n236), .Z(n234) );
  OR U273 ( .A(n237), .B(n238), .Z(n116) );
  XNOR U274 ( .A(n239), .B(n240), .Z(n119) );
  NAND U275 ( .A(n241), .B(n242), .Z(n240) );
  XOR U276 ( .A(n239), .B(n243), .Z(n242) );
  XOR U277 ( .A(n138), .B(n244), .Z(n139) );
  XNOR U278 ( .A(n133), .B(n134), .Z(n244) );
  XNOR U279 ( .A(n135), .B(n136), .Z(n134) );
  AND U280 ( .A(n245), .B(n246), .Z(n136) );
  OR U281 ( .A(n247), .B(n248), .Z(n246) );
  XOR U282 ( .A(n249), .B(n250), .Z(n245) );
  NANDN U283 ( .A(n251), .B(n252), .Z(n250) );
  XNOR U284 ( .A(n249), .B(n253), .Z(n252) );
  OR U285 ( .A(n254), .B(n255), .Z(n135) );
  XOR U286 ( .A(n131), .B(n256), .Z(n133) );
  XOR U287 ( .A(n128), .B(n129), .Z(n256) );
  AND U288 ( .A(n257), .B(n258), .Z(n129) );
  OR U289 ( .A(n259), .B(n260), .Z(n258) );
  XOR U290 ( .A(n261), .B(n262), .Z(n257) );
  NANDN U291 ( .A(n263), .B(n264), .Z(n262) );
  XOR U292 ( .A(n261), .B(n265), .Z(n264) );
  OR U293 ( .A(n266), .B(n267), .Z(n128) );
  XNOR U294 ( .A(n268), .B(n269), .Z(n131) );
  NAND U295 ( .A(n270), .B(n271), .Z(n269) );
  XOR U296 ( .A(n268), .B(n272), .Z(n270) );
  XNOR U297 ( .A(n273), .B(n274), .Z(n138) );
  NANDN U298 ( .A(n275), .B(n276), .Z(n274) );
  XOR U299 ( .A(n273), .B(n277), .Z(n276) );
  XNOR U300 ( .A(n278), .B(n279), .Z(n143) );
  NAND U301 ( .A(n280), .B(n281), .Z(n279) );
  XNOR U302 ( .A(n278), .B(n282), .Z(n280) );
  XNOR U303 ( .A(n151), .B(n283), .Z(o[1]) );
  XNOR U304 ( .A(oglobal[1]), .B(n150), .Z(n283) );
  NANDN U305 ( .A(n284), .B(oglobal[0]), .Z(n150) );
  XNOR U306 ( .A(n281), .B(n282), .Z(n151) );
  XOR U307 ( .A(n185), .B(n186), .Z(n282) );
  XOR U308 ( .A(n179), .B(n180), .Z(n186) );
  XOR U309 ( .A(n162), .B(n163), .Z(n161) );
  AND U310 ( .A(n285), .B(n286), .Z(n163) );
  OR U311 ( .A(n287), .B(n288), .Z(n286) );
  NANDN U312 ( .A(n289), .B(n290), .Z(n285) );
  OR U313 ( .A(n291), .B(n292), .Z(n162) );
  XOR U314 ( .A(n156), .B(n293), .Z(n159) );
  XOR U315 ( .A(n155), .B(n157), .Z(n293) );
  ANDN U316 ( .B(n294), .A(n295), .Z(n157) );
  OR U317 ( .A(n296), .B(n297), .Z(n155) );
  AND U318 ( .A(n298), .B(n299), .Z(n156) );
  OR U319 ( .A(n300), .B(n301), .Z(n299) );
  OR U320 ( .A(n302), .B(n303), .Z(n298) );
  XOR U321 ( .A(n172), .B(n304), .Z(n179) );
  XNOR U322 ( .A(n176), .B(n173), .Z(n304) );
  XNOR U323 ( .A(n174), .B(n175), .Z(n173) );
  AND U324 ( .A(n305), .B(n306), .Z(n175) );
  OR U325 ( .A(n307), .B(n308), .Z(n306) );
  OR U326 ( .A(n309), .B(n310), .Z(n305) );
  OR U327 ( .A(n311), .B(n312), .Z(n174) );
  ANDN U328 ( .B(n313), .A(n314), .Z(n176) );
  XOR U329 ( .A(n168), .B(n315), .Z(n172) );
  XOR U330 ( .A(n167), .B(n169), .Z(n315) );
  ANDN U331 ( .B(n316), .A(n317), .Z(n169) );
  OR U332 ( .A(n318), .B(n319), .Z(n167) );
  AND U333 ( .A(n320), .B(n321), .Z(n168) );
  OR U334 ( .A(n322), .B(n323), .Z(n321) );
  OR U335 ( .A(n324), .B(n325), .Z(n320) );
  XNOR U336 ( .A(n182), .B(n214), .Z(n326) );
  XOR U337 ( .A(n194), .B(n195), .Z(n214) );
  XNOR U338 ( .A(n196), .B(n197), .Z(n195) );
  AND U339 ( .A(n327), .B(n328), .Z(n197) );
  OR U340 ( .A(n329), .B(n330), .Z(n328) );
  OR U341 ( .A(n331), .B(n332), .Z(n327) );
  OR U342 ( .A(n333), .B(n334), .Z(n196) );
  XOR U343 ( .A(n190), .B(n335), .Z(n194) );
  XOR U344 ( .A(n189), .B(n191), .Z(n335) );
  ANDN U345 ( .B(n336), .A(n337), .Z(n191) );
  OR U346 ( .A(n338), .B(n339), .Z(n189) );
  AND U347 ( .A(n340), .B(n341), .Z(n190) );
  OR U348 ( .A(n342), .B(n343), .Z(n341) );
  OR U349 ( .A(n344), .B(n345), .Z(n340) );
  OR U350 ( .A(n346), .B(n347), .Z(n182) );
  XOR U351 ( .A(n206), .B(n348), .Z(n212) );
  XOR U352 ( .A(n210), .B(n207), .Z(n348) );
  XNOR U353 ( .A(n208), .B(n209), .Z(n207) );
  AND U354 ( .A(n349), .B(n350), .Z(n209) );
  OR U355 ( .A(n351), .B(n352), .Z(n350) );
  OR U356 ( .A(n353), .B(n354), .Z(n349) );
  OR U357 ( .A(n355), .B(n356), .Z(n208) );
  OR U358 ( .A(n357), .B(n358), .Z(n210) );
  XOR U359 ( .A(n202), .B(n359), .Z(n206) );
  XOR U360 ( .A(n201), .B(n203), .Z(n359) );
  ANDN U361 ( .B(n360), .A(n361), .Z(n203) );
  OR U362 ( .A(n362), .B(n363), .Z(n201) );
  AND U363 ( .A(n364), .B(n365), .Z(n202) );
  OR U364 ( .A(n366), .B(n367), .Z(n365) );
  OR U365 ( .A(n368), .B(n369), .Z(n364) );
  XOR U366 ( .A(n277), .B(n370), .Z(n281) );
  XNOR U367 ( .A(n278), .B(n275), .Z(n370) );
  XNOR U368 ( .A(n272), .B(n371), .Z(n275) );
  XOR U369 ( .A(n273), .B(n271), .Z(n371) );
  XOR U370 ( .A(n265), .B(n372), .Z(n271) );
  XOR U371 ( .A(n268), .B(n263), .Z(n372) );
  XNOR U372 ( .A(n260), .B(n373), .Z(n263) );
  XOR U373 ( .A(n259), .B(n261), .Z(n373) );
  ANDN U374 ( .B(n374), .A(n375), .Z(n261) );
  OR U375 ( .A(n376), .B(n377), .Z(n259) );
  AND U376 ( .A(n378), .B(n379), .Z(n260) );
  OR U377 ( .A(n380), .B(n381), .Z(n379) );
  OR U378 ( .A(n382), .B(n383), .Z(n378) );
  OR U379 ( .A(n384), .B(n385), .Z(n268) );
  XOR U380 ( .A(n266), .B(n267), .Z(n265) );
  AND U381 ( .A(n386), .B(n387), .Z(n267) );
  OR U382 ( .A(n388), .B(n389), .Z(n387) );
  OR U383 ( .A(n390), .B(n391), .Z(n386) );
  OR U384 ( .A(n392), .B(n393), .Z(n266) );
  OR U385 ( .A(n394), .B(n395), .Z(n273) );
  XNOR U386 ( .A(n251), .B(n253), .Z(n272) );
  XNOR U387 ( .A(n254), .B(n255), .Z(n253) );
  AND U388 ( .A(n396), .B(n397), .Z(n255) );
  OR U389 ( .A(n398), .B(n399), .Z(n397) );
  OR U390 ( .A(n400), .B(n401), .Z(n396) );
  OR U391 ( .A(n402), .B(n403), .Z(n254) );
  XNOR U392 ( .A(n248), .B(n404), .Z(n251) );
  XOR U393 ( .A(n247), .B(n249), .Z(n404) );
  ANDN U394 ( .B(n405), .A(n406), .Z(n249) );
  OR U395 ( .A(n407), .B(n408), .Z(n247) );
  AND U396 ( .A(n409), .B(n410), .Z(n248) );
  OR U397 ( .A(n411), .B(n412), .Z(n410) );
  OR U398 ( .A(n413), .B(n414), .Z(n409) );
  OR U399 ( .A(n415), .B(n416), .Z(n278) );
  XOR U400 ( .A(n223), .B(n224), .Z(n243) );
  XNOR U401 ( .A(n225), .B(n226), .Z(n224) );
  AND U402 ( .A(n417), .B(n418), .Z(n226) );
  OR U403 ( .A(n419), .B(n420), .Z(n418) );
  OR U404 ( .A(n421), .B(n422), .Z(n417) );
  OR U405 ( .A(n423), .B(n424), .Z(n225) );
  XOR U406 ( .A(n219), .B(n425), .Z(n223) );
  XOR U407 ( .A(n218), .B(n220), .Z(n425) );
  ANDN U408 ( .B(n426), .A(n427), .Z(n220) );
  OR U409 ( .A(n428), .B(n429), .Z(n218) );
  AND U410 ( .A(n430), .B(n431), .Z(n219) );
  OR U411 ( .A(n432), .B(n433), .Z(n431) );
  OR U412 ( .A(n434), .B(n435), .Z(n430) );
  XOR U413 ( .A(n235), .B(n436), .Z(n241) );
  XOR U414 ( .A(n239), .B(n236), .Z(n436) );
  XNOR U415 ( .A(n237), .B(n238), .Z(n236) );
  AND U416 ( .A(n437), .B(n438), .Z(n238) );
  OR U417 ( .A(n439), .B(n440), .Z(n438) );
  OR U418 ( .A(n441), .B(n442), .Z(n437) );
  OR U419 ( .A(n443), .B(n444), .Z(n237) );
  OR U420 ( .A(n445), .B(n446), .Z(n239) );
  XOR U421 ( .A(n231), .B(n447), .Z(n235) );
  XOR U422 ( .A(n230), .B(n232), .Z(n447) );
  ANDN U423 ( .B(n448), .A(n449), .Z(n232) );
  OR U424 ( .A(n450), .B(n451), .Z(n230) );
  AND U425 ( .A(n452), .B(n453), .Z(n231) );
  OR U426 ( .A(n454), .B(n455), .Z(n453) );
  OR U427 ( .A(n456), .B(n457), .Z(n452) );
  XNOR U428 ( .A(oglobal[0]), .B(n284), .Z(o[0]) );
  XNOR U429 ( .A(n416), .B(n415), .Z(n284) );
  XNOR U430 ( .A(n395), .B(n394), .Z(n415) );
  XNOR U431 ( .A(n446), .B(n445), .Z(n394) );
  XOR U432 ( .A(n421), .B(n422), .Z(n426) );
  XNOR U433 ( .A(n424), .B(n423), .Z(n422) );
  XNOR U434 ( .A(y[31]), .B(x[31]), .Z(n423) );
  XNOR U435 ( .A(y[30]), .B(x[30]), .Z(n424) );
  XNOR U436 ( .A(n419), .B(n420), .Z(n421) );
  XNOR U437 ( .A(y[29]), .B(x[29]), .Z(n420) );
  XNOR U438 ( .A(y[28]), .B(x[28]), .Z(n419) );
  XNOR U439 ( .A(n434), .B(n435), .Z(n427) );
  XNOR U440 ( .A(n429), .B(n428), .Z(n435) );
  XNOR U441 ( .A(y[27]), .B(x[27]), .Z(n428) );
  XNOR U442 ( .A(y[26]), .B(x[26]), .Z(n429) );
  XNOR U443 ( .A(n432), .B(n433), .Z(n434) );
  XNOR U444 ( .A(y[25]), .B(x[25]), .Z(n433) );
  XNOR U445 ( .A(y[24]), .B(x[24]), .Z(n432) );
  XOR U446 ( .A(n441), .B(n442), .Z(n448) );
  XNOR U447 ( .A(n444), .B(n443), .Z(n442) );
  XNOR U448 ( .A(y[23]), .B(x[23]), .Z(n443) );
  XNOR U449 ( .A(y[22]), .B(x[22]), .Z(n444) );
  XNOR U450 ( .A(n439), .B(n440), .Z(n441) );
  XNOR U451 ( .A(y[21]), .B(x[21]), .Z(n440) );
  XNOR U452 ( .A(y[20]), .B(x[20]), .Z(n439) );
  XNOR U453 ( .A(n456), .B(n457), .Z(n449) );
  XNOR U454 ( .A(n451), .B(n450), .Z(n457) );
  XNOR U455 ( .A(y[19]), .B(x[19]), .Z(n450) );
  XNOR U456 ( .A(y[18]), .B(x[18]), .Z(n451) );
  XNOR U457 ( .A(n454), .B(n455), .Z(n456) );
  XNOR U458 ( .A(y[17]), .B(x[17]), .Z(n455) );
  XNOR U459 ( .A(y[16]), .B(x[16]), .Z(n454) );
  XNOR U460 ( .A(n385), .B(n384), .Z(n395) );
  XOR U461 ( .A(n400), .B(n401), .Z(n405) );
  XNOR U462 ( .A(n403), .B(n402), .Z(n401) );
  XNOR U463 ( .A(y[15]), .B(x[15]), .Z(n402) );
  XNOR U464 ( .A(y[14]), .B(x[14]), .Z(n403) );
  XNOR U465 ( .A(n398), .B(n399), .Z(n400) );
  XNOR U466 ( .A(y[13]), .B(x[13]), .Z(n399) );
  XNOR U467 ( .A(y[12]), .B(x[12]), .Z(n398) );
  XNOR U468 ( .A(n413), .B(n414), .Z(n406) );
  XNOR U469 ( .A(n408), .B(n407), .Z(n414) );
  XNOR U470 ( .A(y[11]), .B(x[11]), .Z(n407) );
  XNOR U471 ( .A(y[10]), .B(x[10]), .Z(n408) );
  XNOR U472 ( .A(n411), .B(n412), .Z(n413) );
  XNOR U473 ( .A(y[9]), .B(x[9]), .Z(n412) );
  XNOR U474 ( .A(y[8]), .B(x[8]), .Z(n411) );
  XOR U475 ( .A(n390), .B(n391), .Z(n374) );
  XNOR U476 ( .A(n393), .B(n392), .Z(n391) );
  XNOR U477 ( .A(y[7]), .B(x[7]), .Z(n392) );
  XNOR U478 ( .A(y[6]), .B(x[6]), .Z(n393) );
  XNOR U479 ( .A(n388), .B(n389), .Z(n390) );
  XNOR U480 ( .A(y[5]), .B(x[5]), .Z(n389) );
  XNOR U481 ( .A(y[4]), .B(x[4]), .Z(n388) );
  XNOR U482 ( .A(n382), .B(n383), .Z(n375) );
  XNOR U483 ( .A(n377), .B(n376), .Z(n383) );
  XNOR U484 ( .A(y[3]), .B(x[3]), .Z(n376) );
  XNOR U485 ( .A(y[2]), .B(x[2]), .Z(n377) );
  XNOR U486 ( .A(n380), .B(n381), .Z(n382) );
  XNOR U487 ( .A(y[1]), .B(x[1]), .Z(n381) );
  XNOR U488 ( .A(y[0]), .B(x[0]), .Z(n380) );
  XNOR U489 ( .A(n347), .B(n346), .Z(n416) );
  XNOR U490 ( .A(n294), .B(n295), .Z(n313) );
  XOR U491 ( .A(n289), .B(n290), .Z(n295) );
  XOR U492 ( .A(n291), .B(n292), .Z(n290) );
  XNOR U493 ( .A(y[63]), .B(x[63]), .Z(n292) );
  XNOR U494 ( .A(y[62]), .B(x[62]), .Z(n291) );
  XNOR U495 ( .A(n287), .B(n288), .Z(n289) );
  XNOR U496 ( .A(y[61]), .B(x[61]), .Z(n288) );
  XNOR U497 ( .A(y[60]), .B(x[60]), .Z(n287) );
  XOR U498 ( .A(n302), .B(n303), .Z(n294) );
  XNOR U499 ( .A(n297), .B(n296), .Z(n303) );
  XNOR U500 ( .A(y[59]), .B(x[59]), .Z(n296) );
  XNOR U501 ( .A(y[58]), .B(x[58]), .Z(n297) );
  XNOR U502 ( .A(n300), .B(n301), .Z(n302) );
  XNOR U503 ( .A(y[57]), .B(x[57]), .Z(n301) );
  XNOR U504 ( .A(y[56]), .B(x[56]), .Z(n300) );
  XOR U505 ( .A(n309), .B(n310), .Z(n316) );
  XNOR U506 ( .A(n312), .B(n311), .Z(n310) );
  XNOR U507 ( .A(y[55]), .B(x[55]), .Z(n311) );
  XNOR U508 ( .A(y[54]), .B(x[54]), .Z(n312) );
  XNOR U509 ( .A(n307), .B(n308), .Z(n309) );
  XNOR U510 ( .A(y[53]), .B(x[53]), .Z(n308) );
  XNOR U511 ( .A(y[52]), .B(x[52]), .Z(n307) );
  XNOR U512 ( .A(n324), .B(n325), .Z(n317) );
  XNOR U513 ( .A(n319), .B(n318), .Z(n325) );
  XNOR U514 ( .A(y[51]), .B(x[51]), .Z(n318) );
  XNOR U515 ( .A(y[50]), .B(x[50]), .Z(n319) );
  XNOR U516 ( .A(n322), .B(n323), .Z(n324) );
  XNOR U517 ( .A(y[49]), .B(x[49]), .Z(n323) );
  XNOR U518 ( .A(y[48]), .B(x[48]), .Z(n322) );
  XNOR U519 ( .A(n358), .B(n357), .Z(n347) );
  XOR U520 ( .A(n331), .B(n332), .Z(n336) );
  XNOR U521 ( .A(n334), .B(n333), .Z(n332) );
  XNOR U522 ( .A(y[47]), .B(x[47]), .Z(n333) );
  XNOR U523 ( .A(y[46]), .B(x[46]), .Z(n334) );
  XNOR U524 ( .A(n329), .B(n330), .Z(n331) );
  XNOR U525 ( .A(y[45]), .B(x[45]), .Z(n330) );
  XNOR U526 ( .A(y[44]), .B(x[44]), .Z(n329) );
  XNOR U527 ( .A(n344), .B(n345), .Z(n337) );
  XNOR U528 ( .A(n339), .B(n338), .Z(n345) );
  XNOR U529 ( .A(y[43]), .B(x[43]), .Z(n338) );
  XNOR U530 ( .A(y[42]), .B(x[42]), .Z(n339) );
  XNOR U531 ( .A(n342), .B(n343), .Z(n344) );
  XNOR U532 ( .A(y[41]), .B(x[41]), .Z(n343) );
  XNOR U533 ( .A(y[40]), .B(x[40]), .Z(n342) );
  XOR U534 ( .A(n353), .B(n354), .Z(n360) );
  XNOR U535 ( .A(n356), .B(n355), .Z(n354) );
  XNOR U536 ( .A(y[39]), .B(x[39]), .Z(n355) );
  XNOR U537 ( .A(y[38]), .B(x[38]), .Z(n356) );
  XNOR U538 ( .A(n351), .B(n352), .Z(n353) );
  XNOR U539 ( .A(y[37]), .B(x[37]), .Z(n352) );
  XNOR U540 ( .A(y[36]), .B(x[36]), .Z(n351) );
  XNOR U541 ( .A(n368), .B(n369), .Z(n361) );
  XNOR U542 ( .A(n363), .B(n362), .Z(n369) );
  XNOR U543 ( .A(y[35]), .B(x[35]), .Z(n362) );
  XNOR U544 ( .A(y[34]), .B(x[34]), .Z(n363) );
  XNOR U545 ( .A(n366), .B(n367), .Z(n368) );
  XNOR U546 ( .A(y[33]), .B(x[33]), .Z(n367) );
  XNOR U547 ( .A(y[32]), .B(x[32]), .Z(n366) );
endmodule

