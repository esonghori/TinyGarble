
module hamming ( x, y, o );
  input [1023:0] x;
  input [1023:0] y;
  output [10:0] o;
  wire   n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442,
         n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450,
         n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458,
         n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466,
         n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474,
         n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482,
         n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490,
         n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498,
         n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506,
         n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514,
         n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522,
         n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530,
         n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538,
         n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546,
         n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554,
         n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562,
         n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570,
         n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578,
         n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586,
         n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594,
         n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602,
         n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610,
         n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618,
         n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626,
         n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634,
         n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642,
         n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650,
         n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658,
         n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666,
         n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674,
         n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682,
         n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690,
         n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698,
         n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706,
         n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714,
         n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722,
         n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730,
         n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738,
         n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746,
         n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754,
         n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762,
         n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770,
         n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778,
         n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786,
         n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794,
         n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802,
         n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810,
         n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818,
         n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826,
         n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834,
         n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842,
         n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850,
         n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858,
         n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866,
         n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874,
         n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882,
         n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890,
         n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898,
         n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906,
         n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914,
         n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
         n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930,
         n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938,
         n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946,
         n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954,
         n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962,
         n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970,
         n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978,
         n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986,
         n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994,
         n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002,
         n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010,
         n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018,
         n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026,
         n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034,
         n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042,
         n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050,
         n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058,
         n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066,
         n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074,
         n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082,
         n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090,
         n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098,
         n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106,
         n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
         n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122,
         n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130,
         n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
         n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146,
         n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154,
         n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
         n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170,
         n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178,
         n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186,
         n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194,
         n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202,
         n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
         n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218,
         n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
         n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
         n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242,
         n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
         n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
         n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
         n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
         n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
         n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
         n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
         n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
         n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
         n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
         n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
         n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
         n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
         n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
         n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362,
         n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
         n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378,
         n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386,
         n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394,
         n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
         n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410,
         n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418,
         n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426,
         n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434,
         n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
         n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450,
         n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458,
         n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466,
         n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
         n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482,
         n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490,
         n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498,
         n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506,
         n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514,
         n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522,
         n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530,
         n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538,
         n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
         n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554,
         n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562,
         n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
         n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578,
         n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586,
         n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594,
         n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602,
         n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610,
         n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618,
         n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626,
         n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634,
         n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642,
         n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650,
         n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658,
         n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666,
         n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674,
         n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682,
         n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690,
         n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698,
         n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706,
         n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714,
         n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722,
         n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730,
         n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738,
         n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746,
         n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754,
         n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762,
         n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770,
         n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778,
         n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786,
         n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794,
         n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802,
         n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810,
         n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818,
         n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826,
         n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834,
         n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842,
         n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850,
         n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858,
         n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866,
         n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874,
         n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882,
         n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890,
         n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898,
         n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906,
         n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914,
         n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922,
         n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930,
         n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938,
         n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946,
         n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954,
         n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962,
         n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970,
         n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978,
         n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986,
         n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994,
         n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002,
         n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010,
         n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018,
         n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026,
         n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034,
         n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042,
         n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050,
         n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058,
         n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066,
         n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074,
         n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082,
         n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090,
         n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098,
         n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106,
         n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114,
         n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122,
         n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130,
         n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138,
         n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146,
         n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154,
         n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162,
         n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170,
         n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178,
         n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186,
         n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194,
         n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202,
         n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210,
         n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218,
         n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226,
         n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234,
         n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242,
         n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250,
         n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258,
         n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266,
         n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274,
         n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282,
         n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290,
         n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298,
         n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306,
         n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314,
         n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322,
         n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330,
         n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338,
         n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346,
         n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354,
         n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362,
         n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370,
         n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
         n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386,
         n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394,
         n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402,
         n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410,
         n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418,
         n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426,
         n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434,
         n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442,
         n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
         n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458,
         n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466,
         n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474,
         n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482,
         n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
         n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498,
         n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506,
         n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514,
         n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
         n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530,
         n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538,
         n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546,
         n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554,
         n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562,
         n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570,
         n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578,
         n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586,
         n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
         n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
         n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610,
         n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618,
         n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
         n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634,
         n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642,
         n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650,
         n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658,
         n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
         n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674,
         n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682,
         n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690,
         n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698,
         n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706,
         n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714,
         n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722,
         n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730,
         n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
         n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746,
         n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754,
         n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762,
         n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
         n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778,
         n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786,
         n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794,
         n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802,
         n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
         n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818,
         n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826,
         n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834,
         n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
         n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850,
         n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858,
         n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866,
         n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874,
         n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882,
         n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890,
         n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898,
         n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906,
         n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
         n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922,
         n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930,
         n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938,
         n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946,
         n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954,
         n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962,
         n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970,
         n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
         n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986,
         n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994,
         n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002,
         n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
         n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018,
         n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026,
         n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034,
         n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042,
         n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050,
         n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058,
         n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066,
         n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074,
         n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
         n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090,
         n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098,
         n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106,
         n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114,
         n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122,
         n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130,
         n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138,
         n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146,
         n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154,
         n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162,
         n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170,
         n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178,
         n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186,
         n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194,
         n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202,
         n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210,
         n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218,
         n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226,
         n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234,
         n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242,
         n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250,
         n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258,
         n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266,
         n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274,
         n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282,
         n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290,
         n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298,
         n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306,
         n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314,
         n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322,
         n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330,
         n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338,
         n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346,
         n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354,
         n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362,
         n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370,
         n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378,
         n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386,
         n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394,
         n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402,
         n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410,
         n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418,
         n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426,
         n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434,
         n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442,
         n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450,
         n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458,
         n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466,
         n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474,
         n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482,
         n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490,
         n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498,
         n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506,
         n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514,
         n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522,
         n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530,
         n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538,
         n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546,
         n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554,
         n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562,
         n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570,
         n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578,
         n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586,
         n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594,
         n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602,
         n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610,
         n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618,
         n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626,
         n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634,
         n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642,
         n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650,
         n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658,
         n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666,
         n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674,
         n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682,
         n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690,
         n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698,
         n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706,
         n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714,
         n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722,
         n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730,
         n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738,
         n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746,
         n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754,
         n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762,
         n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770,
         n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778,
         n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786,
         n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794,
         n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802,
         n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810,
         n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818,
         n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826,
         n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834,
         n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842,
         n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850,
         n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858,
         n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866,
         n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874,
         n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882,
         n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890,
         n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898,
         n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906,
         n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914,
         n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922,
         n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930,
         n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938,
         n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946,
         n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954,
         n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962,
         n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970,
         n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978,
         n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986,
         n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994,
         n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002,
         n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010,
         n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018,
         n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026,
         n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034,
         n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042,
         n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050,
         n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058,
         n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066,
         n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074,
         n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082,
         n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090,
         n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098,
         n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106,
         n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114,
         n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122,
         n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130,
         n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138,
         n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146,
         n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154,
         n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162,
         n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170,
         n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178,
         n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186,
         n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194,
         n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202,
         n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210,
         n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218,
         n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226,
         n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234,
         n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242,
         n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250,
         n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258,
         n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266,
         n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274,
         n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282,
         n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290,
         n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298,
         n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306,
         n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314,
         n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322,
         n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330,
         n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338,
         n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346,
         n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354,
         n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362,
         n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370,
         n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378,
         n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386,
         n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394,
         n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402,
         n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410,
         n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418,
         n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426,
         n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434,
         n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442,
         n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450,
         n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458,
         n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466,
         n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474,
         n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482,
         n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490,
         n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498,
         n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506,
         n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514,
         n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522,
         n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530,
         n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538,
         n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546,
         n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554,
         n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562,
         n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570,
         n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578,
         n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586,
         n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594,
         n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602,
         n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610,
         n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618,
         n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626,
         n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634,
         n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642,
         n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650,
         n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658,
         n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666,
         n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674,
         n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682,
         n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690,
         n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698,
         n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706,
         n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714,
         n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722,
         n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730,
         n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738,
         n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746,
         n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754,
         n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762,
         n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770,
         n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778,
         n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786,
         n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794,
         n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802,
         n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810,
         n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818,
         n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826,
         n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834,
         n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842,
         n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850,
         n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858,
         n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866,
         n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874,
         n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882,
         n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890,
         n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898,
         n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906,
         n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914,
         n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922,
         n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930,
         n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938,
         n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946,
         n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954,
         n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962,
         n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970,
         n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978,
         n28979, n28980, n28981, n28982, n28983, n28984, n28985, n28986,
         n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994,
         n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002,
         n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010,
         n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018,
         n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026,
         n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034,
         n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042,
         n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050,
         n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058,
         n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066,
         n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074,
         n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082,
         n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090,
         n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098,
         n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106,
         n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114,
         n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122,
         n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130,
         n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138,
         n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146,
         n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154,
         n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162,
         n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170,
         n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178,
         n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186,
         n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194,
         n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202,
         n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210,
         n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218,
         n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226,
         n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234,
         n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242,
         n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250,
         n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258,
         n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266,
         n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274,
         n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282,
         n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290,
         n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298,
         n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306,
         n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314,
         n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322,
         n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330,
         n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338,
         n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346,
         n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354,
         n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362,
         n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370,
         n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378,
         n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386,
         n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394,
         n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402,
         n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410,
         n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418,
         n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426,
         n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434,
         n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442,
         n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450,
         n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458,
         n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466,
         n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474,
         n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482,
         n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490,
         n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498,
         n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506,
         n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514,
         n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522,
         n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
         n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538,
         n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546,
         n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554,
         n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562,
         n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570,
         n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578,
         n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586,
         n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594,
         n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602,
         n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610,
         n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618,
         n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626,
         n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634,
         n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642,
         n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650,
         n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658,
         n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666,
         n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674,
         n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682,
         n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690,
         n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698,
         n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706,
         n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714,
         n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722,
         n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730,
         n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738,
         n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746,
         n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754,
         n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762,
         n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770,
         n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778,
         n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786,
         n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794,
         n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802,
         n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810,
         n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818,
         n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826,
         n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834,
         n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842,
         n29843, n29844, n29845, n29846, n29847, n29848, n29849, n29850,
         n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858,
         n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866,
         n29867, n29868, n29869, n29870, n29871, n29872, n29873, n29874,
         n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882,
         n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890,
         n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898,
         n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906,
         n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914,
         n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922,
         n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29930,
         n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938,
         n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946,
         n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954,
         n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962,
         n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970,
         n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978,
         n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986,
         n29987, n29988, n29989, n29990, n29991, n29992, n29993, n29994,
         n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002,
         n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010,
         n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30018,
         n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026,
         n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034,
         n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042,
         n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050,
         n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058,
         n30059, n30060, n30061, n30062, n30063, n30064, n30065, n30066,
         n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074,
         n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082,
         n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090,
         n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098,
         n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106,
         n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114,
         n30115, n30116, n30117, n30118, n30119, n30120, n30121, n30122,
         n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130,
         n30131, n30132, n30133, n30134, n30135, n30136, n30137, n30138,
         n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146,
         n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154,
         n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162,
         n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170,
         n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178,
         n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186,
         n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194,
         n30195, n30196, n30197, n30198, n30199, n30200, n30201, n30202,
         n30203, n30204, n30205, n30206, n30207, n30208, n30209, n30210,
         n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218,
         n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226,
         n30227, n30228, n30229, n30230, n30231, n30232, n30233, n30234,
         n30235, n30236, n30237, n30238, n30239, n30240, n30241, n30242,
         n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250,
         n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258,
         n30259, n30260, n30261, n30262, n30263, n30264, n30265, n30266,
         n30267, n30268, n30269, n30270, n30271, n30272, n30273, n30274,
         n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282,
         n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290,
         n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298,
         n30299, n30300, n30301, n30302, n30303, n30304, n30305, n30306,
         n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314,
         n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322,
         n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330,
         n30331, n30332, n30333, n30334, n30335, n30336, n30337, n30338,
         n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346,
         n30347, n30348, n30349, n30350, n30351, n30352, n30353, n30354,
         n30355, n30356, n30357, n30358, n30359, n30360, n30361, n30362,
         n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370,
         n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378,
         n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386,
         n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394,
         n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402,
         n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410,
         n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418,
         n30419, n30420, n30421, n30422, n30423, n30424, n30425, n30426,
         n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434,
         n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442,
         n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450,
         n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458,
         n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466,
         n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474,
         n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482,
         n30483, n30484, n30485, n30486, n30487, n30488, n30489, n30490,
         n30491, n30492, n30493, n30494, n30495, n30496, n30497, n30498,
         n30499, n30500, n30501, n30502, n30503, n30504, n30505, n30506,
         n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514,
         n30515, n30516, n30517, n30518, n30519, n30520, n30521, n30522,
         n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530,
         n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538,
         n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546,
         n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554,
         n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562,
         n30563, n30564, n30565, n30566, n30567, n30568, n30569, n30570,
         n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578,
         n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586,
         n30587, n30588, n30589, n30590, n30591, n30592, n30593, n30594,
         n30595, n30596, n30597, n30598, n30599, n30600, n30601, n30602,
         n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610,
         n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618,
         n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626,
         n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634,
         n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30642,
         n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650,
         n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658,
         n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666,
         n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674,
         n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682,
         n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690,
         n30691, n30692, n30693, n30694, n30695, n30696, n30697, n30698,
         n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706,
         n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30714,
         n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722,
         n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730,
         n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738,
         n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746,
         n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754,
         n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762,
         n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770,
         n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778,
         n30779, n30780, n30781, n30782, n30783, n30784, n30785, n30786,
         n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794,
         n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802,
         n30803, n30804, n30805, n30806, n30807, n30808, n30809, n30810,
         n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818,
         n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826,
         n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834,
         n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842,
         n30843, n30844, n30845, n30846, n30847, n30848, n30849, n30850,
         n30851, n30852, n30853, n30854, n30855, n30856, n30857, n30858,
         n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866,
         n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874,
         n30875, n30876, n30877, n30878, n30879, n30880, n30881, n30882,
         n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890,
         n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898,
         n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906,
         n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914,
         n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922,
         n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930,
         n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938,
         n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946,
         n30947, n30948, n30949, n30950, n30951, n30952, n30953, n30954,
         n30955, n30956, n30957, n30958, n30959, n30960, n30961, n30962,
         n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970,
         n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978,
         n30979, n30980, n30981, n30982, n30983, n30984, n30985, n30986,
         n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994,
         n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002,
         n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010,
         n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018,
         n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026,
         n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034,
         n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042,
         n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050,
         n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058,
         n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066,
         n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31074,
         n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31082,
         n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090,
         n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098,
         n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106,
         n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114,
         n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122,
         n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130,
         n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138,
         n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146,
         n31147, n31148, n31149, n31150, n31151, n31152, n31153, n31154,
         n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162,
         n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170,
         n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178,
         n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186,
         n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194,
         n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202,
         n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210,
         n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218,
         n31219, n31220, n31221, n31222, n31223, n31224, n31225, n31226,
         n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234,
         n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242,
         n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250,
         n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258,
         n31259, n31260, n31261, n31262, n31263, n31264, n31265, n31266,
         n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274,
         n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282,
         n31283, n31284, n31285, n31286, n31287, n31288, n31289, n31290,
         n31291, n31292, n31293, n31294, n31295, n31296, n31297, n31298,
         n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306,
         n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314,
         n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322,
         n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330,
         n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338,
         n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346,
         n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354,
         n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362,
         n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370,
         n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378,
         n31379, n31380, n31381, n31382, n31383, n31384, n31385, n31386,
         n31387, n31388, n31389, n31390, n31391, n31392, n31393, n31394,
         n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402,
         n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410,
         n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418,
         n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426,
         n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434,
         n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442,
         n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450,
         n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458,
         n31459, n31460, n31461, n31462, n31463, n31464, n31465, n31466,
         n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474,
         n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482,
         n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490,
         n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498,
         n31499, n31500, n31501, n31502, n31503, n31504, n31505, n31506,
         n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514,
         n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522,
         n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530,
         n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538,
         n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546,
         n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554,
         n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562,
         n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570,
         n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578,
         n31579, n31580, n31581, n31582, n31583, n31584, n31585, n31586,
         n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594,
         n31595, n31596, n31597, n31598, n31599, n31600, n31601, n31602,
         n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610,
         n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618,
         n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626,
         n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634,
         n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642,
         n31643, n31644, n31645, n31646, n31647, n31648, n31649, n31650,
         n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658,
         n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666,
         n31667, n31668, n31669, n31670, n31671, n31672, n31673, n31674,
         n31675, n31676, n31677, n31678, n31679, n31680, n31681, n31682,
         n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690,
         n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698,
         n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706,
         n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714,
         n31715, n31716, n31717, n31718, n31719, n31720, n31721, n31722,
         n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730,
         n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738,
         n31739, n31740, n31741, n31742, n31743, n31744, n31745, n31746,
         n31747, n31748, n31749, n31750, n31751, n31752, n31753, n31754,
         n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762,
         n31763, n31764, n31765, n31766, n31767, n31768, n31769, n31770,
         n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778,
         n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786,
         n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794,
         n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802,
         n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810,
         n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818,
         n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826,
         n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834,
         n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842,
         n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850,
         n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858,
         n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866,
         n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874,
         n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882,
         n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890,
         n31891, n31892, n31893, n31894, n31895, n31896, n31897, n31898,
         n31899, n31900, n31901, n31902, n31903, n31904, n31905, n31906,
         n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914,
         n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922,
         n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930,
         n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938,
         n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946,
         n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954,
         n31955, n31956, n31957, n31958, n31959, n31960, n31961, n31962,
         n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970,
         n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978,
         n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986,
         n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994,
         n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002,
         n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010,
         n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018,
         n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026,
         n32027, n32028, n32029, n32030, n32031, n32032, n32033, n32034,
         n32035, n32036, n32037, n32038, n32039, n32040, n32041, n32042,
         n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050,
         n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058,
         n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066,
         n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074,
         n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082,
         n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090,
         n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098,
         n32099, n32100, n32101, n32102, n32103, n32104, n32105, n32106,
         n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114,
         n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122,
         n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130,
         n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138,
         n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146,
         n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154,
         n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162,
         n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170,
         n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178,
         n32179, n32180, n32181, n32182, n32183, n32184, n32185, n32186,
         n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194,
         n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202,
         n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210,
         n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218,
         n32219, n32220, n32221, n32222, n32223, n32224, n32225, n32226,
         n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234,
         n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242,
         n32243, n32244, n32245, n32246, n32247, n32248, n32249, n32250,
         n32251, n32252, n32253, n32254, n32255, n32256, n32257, n32258,
         n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266,
         n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274,
         n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282,
         n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290,
         n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298,
         n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306,
         n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314,
         n32315, n32316, n32317, n32318, n32319, n32320, n32321, n32322,
         n32323, n32324, n32325, n32326, n32327, n32328, n32329, n32330,
         n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338,
         n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346,
         n32347, n32348, n32349, n32350, n32351, n32352, n32353, n32354,
         n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362,
         n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370,
         n32371, n32372, n32373, n32374, n32375, n32376, n32377, n32378,
         n32379, n32380, n32381, n32382, n32383, n32384, n32385, n32386,
         n32387, n32388, n32389, n32390, n32391, n32392, n32393, n32394,
         n32395, n32396, n32397, n32398, n32399, n32400, n32401, n32402,
         n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410,
         n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418,
         n32419, n32420, n32421, n32422, n32423, n32424, n32425, n32426,
         n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434,
         n32435, n32436, n32437, n32438, n32439, n32440, n32441, n32442,
         n32443, n32444, n32445, n32446, n32447, n32448, n32449, n32450,
         n32451, n32452, n32453, n32454, n32455, n32456, n32457, n32458,
         n32459, n32460, n32461, n32462, n32463, n32464, n32465, n32466,
         n32467, n32468, n32469, n32470, n32471, n32472, n32473, n32474,
         n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482,
         n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490,
         n32491, n32492, n32493, n32494, n32495, n32496, n32497, n32498,
         n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506,
         n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514,
         n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522,
         n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530,
         n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32538,
         n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546,
         n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554,
         n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562,
         n32563, n32564, n32565, n32566, n32567, n32568, n32569, n32570,
         n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578,
         n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586,
         n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594,
         n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602,
         n32603, n32604, n32605, n32606, n32607, n32608, n32609, n32610,
         n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618,
         n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626,
         n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634,
         n32635, n32636, n32637, n32638, n32639, n32640, n32641, n32642,
         n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650,
         n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658,
         n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666,
         n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674,
         n32675, n32676, n32677, n32678, n32679, n32680, n32681, n32682,
         n32683, n32684, n32685, n32686, n32687, n32688, n32689, n32690,
         n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698,
         n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706,
         n32707, n32708, n32709, n32710, n32711, n32712, n32713, n32714,
         n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722,
         n32723, n32724, n32725, n32726, n32727, n32728, n32729, n32730,
         n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738,
         n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746,
         n32747, n32748, n32749, n32750, n32751, n32752, n32753, n32754,
         n32755, n32756, n32757, n32758, n32759, n32760, n32761, n32762,
         n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770,
         n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778,
         n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786,
         n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794,
         n32795, n32796, n32797, n32798, n32799, n32800, n32801, n32802,
         n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810,
         n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818,
         n32819, n32820, n32821, n32822, n32823, n32824, n32825, n32826,
         n32827, n32828, n32829, n32830, n32831, n32832, n32833, n32834,
         n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842,
         n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850,
         n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858,
         n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866,
         n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874,
         n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882,
         n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890,
         n32891, n32892, n32893, n32894, n32895, n32896, n32897, n32898,
         n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906,
         n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914,
         n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922,
         n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930,
         n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938,
         n32939, n32940, n32941, n32942, n32943, n32944, n32945, n32946,
         n32947, n32948, n32949, n32950, n32951, n32952, n32953, n32954,
         n32955, n32956, n32957, n32958, n32959, n32960, n32961, n32962,
         n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32970,
         n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978,
         n32979, n32980, n32981, n32982, n32983, n32984, n32985, n32986,
         n32987, n32988, n32989, n32990, n32991, n32992, n32993, n32994,
         n32995, n32996, n32997, n32998, n32999, n33000, n33001, n33002,
         n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010,
         n33011, n33012, n33013, n33014, n33015, n33016, n33017, n33018,
         n33019, n33020, n33021, n33022, n33023, n33024, n33025, n33026,
         n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034,
         n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042,
         n33043, n33044, n33045, n33046, n33047, n33048, n33049, n33050,
         n33051, n33052, n33053, n33054, n33055, n33056, n33057, n33058,
         n33059, n33060, n33061, n33062, n33063, n33064, n33065, n33066,
         n33067, n33068, n33069, n33070, n33071, n33072, n33073, n33074,
         n33075, n33076, n33077, n33078, n33079, n33080, n33081, n33082,
         n33083, n33084, n33085, n33086, n33087, n33088, n33089, n33090,
         n33091, n33092, n33093, n33094, n33095, n33096, n33097, n33098,
         n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106,
         n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114,
         n33115, n33116, n33117, n33118, n33119, n33120, n33121, n33122,
         n33123, n33124, n33125, n33126, n33127, n33128, n33129, n33130,
         n33131, n33132, n33133, n33134, n33135, n33136, n33137, n33138,
         n33139, n33140, n33141, n33142, n33143, n33144, n33145, n33146,
         n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154,
         n33155, n33156, n33157, n33158, n33159, n33160, n33161, n33162,
         n33163, n33164, n33165, n33166, n33167, n33168, n33169, n33170,
         n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178,
         n33179, n33180, n33181, n33182, n33183, n33184, n33185, n33186,
         n33187, n33188, n33189, n33190, n33191, n33192, n33193, n33194,
         n33195, n33196, n33197, n33198, n33199, n33200, n33201, n33202,
         n33203, n33204, n33205, n33206, n33207, n33208, n33209, n33210,
         n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218,
         n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226,
         n33227, n33228, n33229, n33230, n33231, n33232, n33233, n33234,
         n33235, n33236, n33237, n33238, n33239, n33240, n33241, n33242,
         n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250,
         n33251, n33252, n33253, n33254, n33255, n33256, n33257, n33258,
         n33259, n33260, n33261, n33262, n33263, n33264, n33265, n33266,
         n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274,
         n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282,
         n33283, n33284, n33285, n33286, n33287, n33288, n33289, n33290,
         n33291, n33292, n33293, n33294, n33295, n33296, n33297, n33298,
         n33299, n33300, n33301, n33302, n33303, n33304, n33305, n33306,
         n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33314,
         n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322,
         n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330,
         n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338,
         n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346,
         n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354,
         n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362,
         n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370,
         n33371, n33372, n33373, n33374, n33375, n33376, n33377, n33378,
         n33379, n33380, n33381, n33382, n33383, n33384, n33385, n33386,
         n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394,
         n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402,
         n33403, n33404, n33405, n33406, n33407, n33408, n33409, n33410,
         n33411, n33412, n33413, n33414, n33415, n33416, n33417, n33418,
         n33419, n33420, n33421, n33422, n33423, n33424, n33425, n33426,
         n33427, n33428, n33429, n33430, n33431, n33432, n33433, n33434,
         n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442,
         n33443, n33444, n33445, n33446, n33447, n33448, n33449, n33450,
         n33451, n33452, n33453, n33454, n33455, n33456, n33457, n33458,
         n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466,
         n33467, n33468, n33469, n33470, n33471, n33472, n33473, n33474,
         n33475, n33476, n33477, n33478, n33479, n33480, n33481, n33482,
         n33483, n33484, n33485, n33486, n33487, n33488, n33489, n33490,
         n33491, n33492, n33493, n33494, n33495, n33496, n33497, n33498,
         n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506,
         n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514,
         n33515, n33516, n33517, n33518, n33519, n33520, n33521, n33522,
         n33523, n33524, n33525, n33526, n33527, n33528, n33529, n33530,
         n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538,
         n33539, n33540, n33541, n33542, n33543, n33544, n33545, n33546,
         n33547, n33548, n33549, n33550, n33551, n33552, n33553, n33554,
         n33555, n33556, n33557, n33558, n33559, n33560, n33561, n33562,
         n33563, n33564, n33565, n33566, n33567, n33568, n33569, n33570,
         n33571, n33572, n33573, n33574, n33575, n33576, n33577, n33578,
         n33579, n33580, n33581, n33582, n33583, n33584, n33585, n33586,
         n33587, n33588, n33589, n33590, n33591, n33592, n33593, n33594,
         n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602,
         n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610,
         n33611, n33612, n33613, n33614, n33615, n33616, n33617, n33618,
         n33619, n33620, n33621, n33622, n33623, n33624, n33625, n33626,
         n33627, n33628, n33629, n33630, n33631, n33632, n33633, n33634,
         n33635, n33636, n33637, n33638, n33639, n33640, n33641, n33642,
         n33643, n33644, n33645, n33646, n33647, n33648, n33649, n33650,
         n33651, n33652, n33653, n33654, n33655, n33656, n33657, n33658,
         n33659, n33660, n33661, n33662, n33663, n33664, n33665, n33666,
         n33667, n33668, n33669, n33670, n33671, n33672, n33673, n33674,
         n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682,
         n33683, n33684, n33685, n33686, n33687, n33688, n33689, n33690,
         n33691, n33692, n33693, n33694, n33695, n33696, n33697, n33698,
         n33699, n33700, n33701, n33702, n33703, n33704, n33705, n33706,
         n33707, n33708, n33709, n33710, n33711, n33712, n33713, n33714,
         n33715, n33716, n33717, n33718, n33719, n33720, n33721, n33722,
         n33723, n33724, n33725, n33726, n33727, n33728, n33729, n33730,
         n33731, n33732, n33733, n33734, n33735, n33736, n33737, n33738,
         n33739, n33740, n33741, n33742, n33743, n33744, n33745, n33746,
         n33747, n33748, n33749, n33750, n33751, n33752, n33753, n33754,
         n33755, n33756, n33757, n33758, n33759, n33760, n33761, n33762,
         n33763, n33764, n33765, n33766, n33767, n33768, n33769, n33770,
         n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778,
         n33779, n33780, n33781, n33782, n33783, n33784, n33785, n33786,
         n33787, n33788, n33789, n33790, n33791, n33792, n33793, n33794,
         n33795, n33796, n33797, n33798, n33799, n33800, n33801, n33802,
         n33803, n33804, n33805, n33806, n33807, n33808, n33809, n33810,
         n33811, n33812, n33813, n33814, n33815, n33816, n33817, n33818,
         n33819, n33820, n33821, n33822, n33823, n33824, n33825, n33826,
         n33827, n33828, n33829, n33830, n33831, n33832, n33833, n33834,
         n33835, n33836, n33837, n33838, n33839, n33840, n33841, n33842,
         n33843, n33844, n33845, n33846, n33847, n33848, n33849, n33850,
         n33851, n33852, n33853, n33854, n33855, n33856, n33857, n33858,
         n33859, n33860, n33861, n33862, n33863, n33864, n33865, n33866,
         n33867, n33868, n33869, n33870, n33871, n33872, n33873, n33874,
         n33875, n33876, n33877, n33878, n33879, n33880, n33881, n33882,
         n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890,
         n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33898,
         n33899, n33900, n33901, n33902, n33903, n33904, n33905, n33906,
         n33907, n33908, n33909, n33910, n33911, n33912, n33913, n33914,
         n33915, n33916, n33917, n33918, n33919, n33920, n33921, n33922,
         n33923, n33924, n33925, n33926, n33927, n33928, n33929, n33930,
         n33931, n33932, n33933, n33934, n33935, n33936, n33937, n33938,
         n33939, n33940, n33941, n33942, n33943, n33944, n33945, n33946,
         n33947, n33948, n33949, n33950, n33951, n33952, n33953, n33954,
         n33955, n33956, n33957, n33958, n33959, n33960, n33961, n33962,
         n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970,
         n33971, n33972, n33973, n33974, n33975, n33976, n33977, n33978,
         n33979, n33980, n33981, n33982, n33983, n33984, n33985, n33986,
         n33987, n33988, n33989, n33990, n33991, n33992, n33993, n33994,
         n33995, n33996, n33997, n33998, n33999, n34000, n34001, n34002,
         n34003, n34004, n34005, n34006, n34007, n34008, n34009, n34010,
         n34011, n34012, n34013, n34014, n34015, n34016, n34017, n34018,
         n34019, n34020, n34021, n34022, n34023, n34024, n34025, n34026,
         n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034,
         n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042,
         n34043, n34044, n34045, n34046, n34047, n34048, n34049, n34050,
         n34051, n34052, n34053, n34054, n34055, n34056, n34057, n34058,
         n34059, n34060, n34061, n34062, n34063, n34064, n34065, n34066,
         n34067, n34068, n34069, n34070, n34071, n34072, n34073, n34074,
         n34075, n34076, n34077, n34078, n34079, n34080, n34081, n34082,
         n34083, n34084, n34085, n34086, n34087, n34088, n34089, n34090,
         n34091, n34092, n34093, n34094, n34095, n34096, n34097, n34098,
         n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106,
         n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114,
         n34115, n34116, n34117, n34118, n34119, n34120, n34121, n34122,
         n34123, n34124, n34125, n34126, n34127, n34128, n34129, n34130,
         n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138,
         n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34146,
         n34147, n34148, n34149, n34150, n34151, n34152, n34153, n34154,
         n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162,
         n34163, n34164, n34165, n34166, n34167, n34168, n34169, n34170,
         n34171, n34172, n34173, n34174, n34175, n34176, n34177, n34178,
         n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186,
         n34187, n34188, n34189, n34190, n34191, n34192, n34193, n34194,
         n34195, n34196, n34197, n34198, n34199, n34200, n34201, n34202,
         n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210,
         n34211, n34212, n34213, n34214, n34215, n34216, n34217, n34218,
         n34219, n34220, n34221, n34222, n34223, n34224, n34225, n34226,
         n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234,
         n34235, n34236, n34237, n34238, n34239, n34240, n34241, n34242,
         n34243, n34244, n34245, n34246, n34247, n34248, n34249, n34250,
         n34251, n34252, n34253, n34254, n34255, n34256, n34257, n34258,
         n34259, n34260, n34261, n34262, n34263, n34264, n34265, n34266,
         n34267, n34268, n34269, n34270, n34271, n34272, n34273, n34274,
         n34275, n34276, n34277, n34278, n34279, n34280, n34281, n34282,
         n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290,
         n34291, n34292, n34293, n34294, n34295, n34296, n34297, n34298,
         n34299, n34300, n34301, n34302, n34303, n34304, n34305, n34306,
         n34307, n34308, n34309, n34310, n34311, n34312, n34313, n34314,
         n34315, n34316, n34317, n34318, n34319, n34320, n34321, n34322,
         n34323, n34324, n34325, n34326, n34327, n34328, n34329, n34330,
         n34331, n34332, n34333, n34334, n34335, n34336, n34337, n34338,
         n34339, n34340, n34341, n34342, n34343, n34344, n34345, n34346,
         n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354,
         n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362,
         n34363, n34364, n34365, n34366, n34367, n34368, n34369, n34370,
         n34371, n34372, n34373, n34374, n34375, n34376, n34377, n34378,
         n34379, n34380, n34381, n34382, n34383, n34384, n34385, n34386,
         n34387, n34388, n34389, n34390, n34391, n34392, n34393, n34394,
         n34395, n34396, n34397, n34398, n34399, n34400, n34401, n34402,
         n34403, n34404, n34405, n34406, n34407, n34408, n34409, n34410,
         n34411, n34412, n34413, n34414, n34415, n34416, n34417, n34418,
         n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426,
         n34427, n34428, n34429, n34430, n34431, n34432, n34433, n34434,
         n34435, n34436, n34437, n34438, n34439, n34440, n34441, n34442,
         n34443, n34444, n34445, n34446, n34447, n34448, n34449, n34450,
         n34451, n34452, n34453, n34454, n34455, n34456, n34457, n34458,
         n34459, n34460, n34461, n34462, n34463, n34464, n34465, n34466,
         n34467, n34468, n34469, n34470, n34471, n34472, n34473, n34474,
         n34475, n34476, n34477, n34478, n34479, n34480, n34481, n34482,
         n34483, n34484, n34485, n34486, n34487, n34488, n34489, n34490,
         n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498,
         n34499, n34500, n34501, n34502, n34503, n34504, n34505, n34506,
         n34507, n34508, n34509, n34510, n34511, n34512, n34513, n34514,
         n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522,
         n34523, n34524, n34525, n34526, n34527, n34528, n34529, n34530,
         n34531, n34532, n34533, n34534, n34535, n34536, n34537, n34538,
         n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546,
         n34547, n34548, n34549, n34550, n34551, n34552, n34553, n34554,
         n34555, n34556, n34557, n34558, n34559, n34560, n34561, n34562,
         n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570,
         n34571, n34572, n34573, n34574, n34575, n34576, n34577, n34578,
         n34579, n34580, n34581, n34582, n34583, n34584, n34585, n34586,
         n34587, n34588, n34589, n34590, n34591, n34592, n34593, n34594,
         n34595, n34596, n34597, n34598, n34599, n34600, n34601, n34602,
         n34603, n34604, n34605, n34606, n34607, n34608, n34609, n34610,
         n34611, n34612, n34613, n34614, n34615, n34616, n34617, n34618,
         n34619, n34620, n34621, n34622, n34623, n34624, n34625, n34626,
         n34627, n34628, n34629, n34630, n34631, n34632, n34633, n34634,
         n34635, n34636, n34637, n34638, n34639, n34640, n34641, n34642,
         n34643, n34644, n34645, n34646, n34647, n34648, n34649, n34650,
         n34651, n34652, n34653, n34654, n34655, n34656, n34657, n34658,
         n34659, n34660, n34661, n34662, n34663, n34664, n34665, n34666,
         n34667, n34668, n34669, n34670, n34671, n34672, n34673, n34674,
         n34675, n34676, n34677, n34678, n34679, n34680, n34681, n34682,
         n34683, n34684, n34685, n34686, n34687, n34688, n34689, n34690,
         n34691, n34692, n34693, n34694, n34695, n34696, n34697, n34698,
         n34699, n34700, n34701, n34702, n34703, n34704, n34705, n34706,
         n34707, n34708, n34709, n34710, n34711, n34712, n34713, n34714,
         n34715, n34716, n34717, n34718, n34719, n34720, n34721, n34722,
         n34723, n34724, n34725, n34726, n34727, n34728, n34729, n34730,
         n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738,
         n34739, n34740, n34741, n34742, n34743, n34744, n34745, n34746,
         n34747, n34748, n34749, n34750, n34751, n34752, n34753, n34754,
         n34755, n34756, n34757, n34758, n34759, n34760, n34761, n34762,
         n34763, n34764, n34765, n34766, n34767, n34768, n34769, n34770,
         n34771, n34772, n34773, n34774, n34775, n34776, n34777, n34778,
         n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786,
         n34787, n34788, n34789, n34790, n34791, n34792, n34793, n34794,
         n34795, n34796, n34797, n34798, n34799, n34800, n34801, n34802,
         n34803, n34804, n34805, n34806, n34807, n34808, n34809, n34810,
         n34811, n34812, n34813, n34814, n34815, n34816, n34817, n34818,
         n34819, n34820, n34821, n34822, n34823, n34824, n34825, n34826,
         n34827, n34828, n34829, n34830, n34831, n34832, n34833, n34834,
         n34835, n34836, n34837, n34838, n34839, n34840, n34841, n34842,
         n34843, n34844, n34845, n34846, n34847, n34848, n34849, n34850,
         n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858,
         n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866,
         n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874,
         n34875, n34876, n34877, n34878, n34879, n34880, n34881, n34882,
         n34883, n34884, n34885, n34886, n34887, n34888, n34889, n34890,
         n34891, n34892, n34893, n34894, n34895, n34896, n34897, n34898,
         n34899, n34900, n34901, n34902, n34903, n34904, n34905, n34906,
         n34907, n34908, n34909, n34910, n34911, n34912, n34913, n34914,
         n34915, n34916, n34917, n34918, n34919, n34920, n34921, n34922,
         n34923, n34924, n34925, n34926, n34927, n34928, n34929, n34930,
         n34931, n34932, n34933, n34934, n34935, n34936, n34937, n34938,
         n34939, n34940, n34941, n34942, n34943, n34944, n34945, n34946,
         n34947, n34948, n34949, n34950, n34951, n34952, n34953, n34954,
         n34955, n34956, n34957, n34958, n34959, n34960, n34961, n34962,
         n34963, n34964, n34965, n34966, n34967, n34968, n34969, n34970,
         n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978,
         n34979, n34980, n34981, n34982, n34983, n34984, n34985, n34986,
         n34987, n34988, n34989, n34990, n34991, n34992, n34993, n34994,
         n34995, n34996, n34997, n34998, n34999, n35000, n35001, n35002,
         n35003, n35004, n35005, n35006, n35007, n35008, n35009, n35010,
         n35011, n35012, n35013, n35014, n35015, n35016, n35017, n35018,
         n35019, n35020, n35021, n35022, n35023, n35024, n35025, n35026,
         n35027, n35028, n35029, n35030, n35031, n35032, n35033, n35034,
         n35035, n35036, n35037, n35038, n35039, n35040, n35041, n35042,
         n35043, n35044, n35045, n35046, n35047, n35048, n35049, n35050,
         n35051, n35052, n35053, n35054, n35055, n35056, n35057, n35058,
         n35059, n35060, n35061, n35062, n35063, n35064, n35065, n35066,
         n35067, n35068, n35069, n35070, n35071, n35072, n35073, n35074,
         n35075, n35076, n35077, n35078, n35079, n35080, n35081, n35082,
         n35083, n35084, n35085, n35086, n35087, n35088, n35089, n35090,
         n35091, n35092, n35093, n35094, n35095, n35096, n35097, n35098,
         n35099, n35100, n35101, n35102, n35103, n35104, n35105, n35106,
         n35107, n35108, n35109, n35110, n35111, n35112, n35113, n35114,
         n35115, n35116, n35117, n35118, n35119, n35120, n35121, n35122,
         n35123, n35124, n35125, n35126, n35127, n35128, n35129, n35130,
         n35131, n35132, n35133, n35134, n35135, n35136, n35137, n35138,
         n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146,
         n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154,
         n35155, n35156, n35157, n35158, n35159, n35160, n35161, n35162,
         n35163, n35164, n35165, n35166, n35167, n35168, n35169, n35170,
         n35171, n35172, n35173, n35174, n35175, n35176, n35177, n35178,
         n35179, n35180, n35181, n35182, n35183, n35184, n35185, n35186,
         n35187, n35188, n35189, n35190, n35191, n35192, n35193, n35194,
         n35195, n35196, n35197, n35198, n35199, n35200, n35201, n35202,
         n35203, n35204, n35205, n35206, n35207, n35208, n35209, n35210,
         n35211, n35212, n35213, n35214, n35215, n35216, n35217, n35218,
         n35219, n35220, n35221, n35222, n35223, n35224, n35225, n35226,
         n35227, n35228, n35229, n35230, n35231, n35232, n35233, n35234,
         n35235, n35236, n35237, n35238, n35239, n35240, n35241, n35242,
         n35243, n35244, n35245, n35246, n35247, n35248, n35249, n35250,
         n35251, n35252, n35253, n35254, n35255, n35256, n35257, n35258,
         n35259, n35260, n35261, n35262, n35263, n35264, n35265, n35266,
         n35267, n35268, n35269, n35270, n35271, n35272, n35273, n35274,
         n35275, n35276, n35277, n35278, n35279, n35280, n35281, n35282,
         n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290,
         n35291, n35292, n35293, n35294, n35295, n35296, n35297, n35298,
         n35299, n35300, n35301, n35302, n35303, n35304, n35305, n35306,
         n35307, n35308, n35309, n35310, n35311, n35312, n35313, n35314,
         n35315, n35316, n35317, n35318, n35319, n35320, n35321, n35322,
         n35323, n35324, n35325, n35326, n35327, n35328, n35329, n35330,
         n35331, n35332, n35333, n35334, n35335, n35336, n35337, n35338,
         n35339, n35340, n35341, n35342, n35343, n35344, n35345, n35346,
         n35347, n35348, n35349, n35350, n35351, n35352, n35353, n35354,
         n35355, n35356, n35357, n35358, n35359, n35360, n35361, n35362,
         n35363, n35364, n35365, n35366, n35367, n35368, n35369, n35370,
         n35371, n35372, n35373, n35374, n35375, n35376, n35377, n35378,
         n35379, n35380, n35381, n35382, n35383, n35384, n35385, n35386,
         n35387, n35388, n35389, n35390, n35391, n35392, n35393, n35394,
         n35395, n35396, n35397, n35398, n35399, n35400, n35401, n35402,
         n35403, n35404, n35405, n35406, n35407, n35408, n35409, n35410,
         n35411, n35412, n35413, n35414, n35415, n35416, n35417, n35418,
         n35419, n35420, n35421, n35422, n35423, n35424, n35425, n35426,
         n35427, n35428, n35429, n35430, n35431, n35432, n35433, n35434,
         n35435, n35436, n35437, n35438, n35439, n35440, n35441, n35442,
         n35443, n35444, n35445, n35446, n35447, n35448, n35449, n35450,
         n35451, n35452, n35453, n35454, n35455, n35456, n35457, n35458,
         n35459, n35460, n35461, n35462, n35463, n35464, n35465, n35466,
         n35467, n35468, n35469, n35470, n35471, n35472, n35473, n35474,
         n35475, n35476, n35477, n35478, n35479, n35480, n35481, n35482,
         n35483, n35484, n35485, n35486, n35487, n35488, n35489, n35490,
         n35491, n35492, n35493, n35494, n35495, n35496, n35497, n35498,
         n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506,
         n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514,
         n35515, n35516, n35517, n35518, n35519, n35520, n35521, n35522,
         n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530,
         n35531, n35532, n35533, n35534, n35535, n35536, n35537, n35538,
         n35539, n35540, n35541, n35542, n35543, n35544, n35545, n35546,
         n35547, n35548, n35549, n35550, n35551, n35552, n35553, n35554,
         n35555, n35556, n35557, n35558, n35559, n35560, n35561, n35562,
         n35563, n35564, n35565, n35566, n35567, n35568, n35569, n35570,
         n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578,
         n35579, n35580, n35581, n35582, n35583, n35584, n35585, n35586,
         n35587, n35588, n35589, n35590, n35591, n35592, n35593, n35594,
         n35595, n35596, n35597, n35598, n35599, n35600, n35601, n35602,
         n35603, n35604, n35605, n35606, n35607, n35608, n35609, n35610,
         n35611, n35612, n35613, n35614, n35615, n35616, n35617, n35618,
         n35619, n35620, n35621, n35622, n35623, n35624, n35625, n35626,
         n35627, n35628, n35629, n35630, n35631, n35632, n35633, n35634,
         n35635, n35636, n35637, n35638, n35639, n35640, n35641, n35642,
         n35643, n35644, n35645, n35646, n35647, n35648, n35649, n35650,
         n35651, n35652, n35653, n35654, n35655, n35656, n35657, n35658,
         n35659, n35660, n35661, n35662, n35663, n35664, n35665, n35666,
         n35667, n35668, n35669, n35670, n35671, n35672, n35673, n35674,
         n35675, n35676, n35677, n35678, n35679, n35680, n35681, n35682,
         n35683, n35684, n35685, n35686, n35687, n35688, n35689, n35690,
         n35691, n35692, n35693, n35694, n35695, n35696, n35697, n35698,
         n35699, n35700, n35701, n35702, n35703, n35704, n35705, n35706,
         n35707, n35708, n35709, n35710, n35711, n35712, n35713, n35714,
         n35715, n35716, n35717, n35718, n35719, n35720, n35721, n35722,
         n35723, n35724, n35725, n35726, n35727, n35728, n35729, n35730,
         n35731, n35732, n35733, n35734, n35735, n35736, n35737, n35738,
         n35739, n35740, n35741, n35742, n35743, n35744, n35745, n35746,
         n35747, n35748, n35749, n35750, n35751, n35752, n35753, n35754,
         n35755, n35756, n35757, n35758, n35759, n35760, n35761, n35762,
         n35763, n35764, n35765, n35766, n35767, n35768, n35769, n35770,
         n35771, n35772, n35773, n35774, n35775, n35776, n35777, n35778,
         n35779, n35780, n35781, n35782, n35783, n35784, n35785, n35786,
         n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794,
         n35795, n35796, n35797, n35798, n35799, n35800, n35801, n35802,
         n35803, n35804, n35805, n35806, n35807, n35808, n35809, n35810,
         n35811, n35812, n35813, n35814, n35815, n35816, n35817, n35818,
         n35819, n35820, n35821, n35822, n35823, n35824, n35825, n35826,
         n35827, n35828, n35829, n35830, n35831, n35832, n35833, n35834,
         n35835, n35836, n35837, n35838, n35839, n35840, n35841, n35842,
         n35843, n35844, n35845, n35846, n35847, n35848, n35849, n35850,
         n35851, n35852, n35853, n35854, n35855, n35856, n35857, n35858,
         n35859, n35860, n35861, n35862, n35863, n35864, n35865, n35866,
         n35867, n35868, n35869, n35870, n35871, n35872, n35873, n35874,
         n35875, n35876, n35877, n35878, n35879, n35880, n35881, n35882,
         n35883, n35884, n35885, n35886, n35887, n35888, n35889, n35890,
         n35891, n35892, n35893, n35894, n35895, n35896, n35897, n35898,
         n35899, n35900, n35901, n35902, n35903, n35904, n35905, n35906,
         n35907, n35908, n35909, n35910, n35911, n35912, n35913, n35914,
         n35915, n35916, n35917, n35918, n35919, n35920, n35921, n35922,
         n35923, n35924, n35925, n35926, n35927, n35928, n35929, n35930,
         n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938,
         n35939, n35940, n35941, n35942, n35943, n35944, n35945, n35946,
         n35947, n35948, n35949, n35950, n35951, n35952, n35953, n35954,
         n35955, n35956, n35957, n35958, n35959, n35960, n35961, n35962,
         n35963, n35964, n35965, n35966, n35967, n35968, n35969, n35970,
         n35971, n35972, n35973, n35974, n35975, n35976, n35977, n35978,
         n35979, n35980, n35981, n35982, n35983, n35984, n35985, n35986,
         n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994,
         n35995, n35996, n35997, n35998, n35999, n36000, n36001, n36002,
         n36003, n36004, n36005, n36006, n36007, n36008, n36009, n36010,
         n36011, n36012, n36013, n36014, n36015, n36016, n36017, n36018,
         n36019, n36020, n36021, n36022, n36023, n36024, n36025, n36026,
         n36027, n36028, n36029, n36030, n36031, n36032, n36033, n36034,
         n36035, n36036, n36037, n36038, n36039, n36040, n36041, n36042,
         n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050,
         n36051, n36052, n36053, n36054, n36055, n36056, n36057, n36058,
         n36059, n36060, n36061, n36062, n36063, n36064, n36065, n36066,
         n36067, n36068, n36069, n36070, n36071, n36072, n36073, n36074,
         n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082,
         n36083, n36084, n36085, n36086, n36087, n36088, n36089, n36090,
         n36091, n36092, n36093, n36094, n36095, n36096, n36097, n36098,
         n36099, n36100, n36101, n36102, n36103, n36104, n36105, n36106,
         n36107, n36108, n36109, n36110, n36111, n36112, n36113, n36114,
         n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122,
         n36123, n36124, n36125, n36126, n36127, n36128, n36129, n36130,
         n36131, n36132, n36133, n36134, n36135, n36136, n36137, n36138,
         n36139, n36140, n36141, n36142, n36143, n36144, n36145, n36146,
         n36147, n36148, n36149, n36150, n36151, n36152, n36153, n36154,
         n36155, n36156, n36157, n36158, n36159, n36160, n36161, n36162,
         n36163, n36164, n36165, n36166, n36167, n36168, n36169, n36170,
         n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178,
         n36179, n36180, n36181, n36182, n36183, n36184, n36185, n36186,
         n36187, n36188, n36189, n36190, n36191, n36192, n36193, n36194,
         n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202,
         n36203, n36204, n36205, n36206, n36207, n36208, n36209, n36210,
         n36211, n36212, n36213, n36214, n36215, n36216, n36217, n36218,
         n36219, n36220, n36221, n36222, n36223, n36224, n36225, n36226,
         n36227, n36228, n36229, n36230, n36231, n36232, n36233, n36234,
         n36235, n36236, n36237, n36238, n36239, n36240, n36241, n36242,
         n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250,
         n36251, n36252, n36253, n36254, n36255, n36256, n36257, n36258,
         n36259, n36260, n36261, n36262, n36263, n36264, n36265, n36266,
         n36267, n36268, n36269, n36270, n36271, n36272, n36273, n36274,
         n36275, n36276, n36277, n36278, n36279, n36280, n36281, n36282,
         n36283, n36284, n36285, n36286, n36287, n36288, n36289, n36290,
         n36291, n36292, n36293, n36294, n36295, n36296, n36297, n36298,
         n36299, n36300, n36301, n36302, n36303, n36304, n36305, n36306,
         n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314,
         n36315, n36316, n36317, n36318, n36319, n36320, n36321, n36322,
         n36323, n36324, n36325, n36326, n36327, n36328, n36329, n36330,
         n36331, n36332, n36333, n36334, n36335, n36336, n36337, n36338,
         n36339, n36340, n36341, n36342, n36343, n36344, n36345, n36346,
         n36347, n36348, n36349, n36350, n36351, n36352, n36353, n36354,
         n36355, n36356, n36357, n36358, n36359, n36360, n36361, n36362,
         n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370,
         n36371, n36372, n36373, n36374, n36375, n36376, n36377, n36378,
         n36379, n36380, n36381, n36382, n36383, n36384, n36385, n36386,
         n36387, n36388, n36389, n36390, n36391, n36392, n36393, n36394,
         n36395, n36396, n36397, n36398, n36399, n36400, n36401, n36402,
         n36403, n36404, n36405, n36406, n36407, n36408, n36409, n36410,
         n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418,
         n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36426,
         n36427, n36428, n36429, n36430, n36431, n36432, n36433, n36434,
         n36435, n36436, n36437, n36438, n36439, n36440, n36441, n36442,
         n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450,
         n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458,
         n36459, n36460, n36461, n36462, n36463, n36464, n36465, n36466,
         n36467, n36468, n36469, n36470, n36471, n36472, n36473, n36474,
         n36475, n36476, n36477, n36478, n36479, n36480, n36481, n36482,
         n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490,
         n36491, n36492, n36493, n36494, n36495, n36496, n36497, n36498,
         n36499, n36500, n36501, n36502, n36503, n36504, n36505, n36506,
         n36507, n36508, n36509, n36510, n36511, n36512, n36513, n36514,
         n36515, n36516, n36517, n36518, n36519, n36520, n36521, n36522,
         n36523, n36524, n36525, n36526, n36527, n36528, n36529, n36530,
         n36531, n36532, n36533, n36534, n36535, n36536, n36537, n36538,
         n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546,
         n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554,
         n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562,
         n36563, n36564, n36565, n36566, n36567, n36568, n36569, n36570,
         n36571, n36572, n36573, n36574, n36575, n36576, n36577, n36578,
         n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586,
         n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594,
         n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602,
         n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610,
         n36611, n36612, n36613, n36614, n36615, n36616, n36617, n36618,
         n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626,
         n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634,
         n36635, n36636, n36637, n36638, n36639, n36640, n36641, n36642,
         n36643, n36644, n36645, n36646, n36647, n36648, n36649, n36650,
         n36651, n36652, n36653, n36654, n36655, n36656, n36657, n36658,
         n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666,
         n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674,
         n36675, n36676, n36677, n36678, n36679, n36680, n36681, n36682,
         n36683, n36684, n36685, n36686, n36687, n36688, n36689, n36690,
         n36691, n36692, n36693, n36694, n36695, n36696, n36697, n36698,
         n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706,
         n36707, n36708, n36709, n36710, n36711, n36712, n36713, n36714,
         n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722,
         n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730,
         n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738,
         n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746,
         n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754,
         n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762,
         n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770,
         n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778,
         n36779, n36780, n36781, n36782, n36783, n36784, n36785, n36786,
         n36787, n36788, n36789, n36790, n36791, n36792, n36793, n36794,
         n36795, n36796, n36797, n36798, n36799, n36800, n36801, n36802,
         n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810,
         n36811, n36812, n36813, n36814, n36815, n36816, n36817, n36818,
         n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826,
         n36827, n36828, n36829, n36830, n36831, n36832, n36833, n36834,
         n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842,
         n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850,
         n36851, n36852, n36853, n36854, n36855, n36856, n36857, n36858,
         n36859, n36860, n36861, n36862, n36863, n36864, n36865, n36866,
         n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874,
         n36875, n36876, n36877, n36878, n36879, n36880, n36881, n36882,
         n36883, n36884, n36885, n36886, n36887, n36888, n36889, n36890,
         n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898,
         n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906,
         n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914,
         n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922,
         n36923, n36924, n36925, n36926, n36927, n36928, n36929, n36930,
         n36931, n36932, n36933, n36934, n36935, n36936, n36937, n36938,
         n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946,
         n36947, n36948, n36949, n36950, n36951, n36952, n36953, n36954,
         n36955, n36956, n36957, n36958, n36959, n36960, n36961, n36962,
         n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970,
         n36971, n36972, n36973, n36974, n36975, n36976, n36977, n36978,
         n36979, n36980, n36981, n36982, n36983, n36984, n36985, n36986,
         n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994,
         n36995, n36996, n36997, n36998, n36999, n37000, n37001, n37002,
         n37003, n37004, n37005, n37006, n37007, n37008, n37009, n37010,
         n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018,
         n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026,
         n37027, n37028, n37029, n37030, n37031, n37032, n37033, n37034,
         n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042,
         n37043, n37044, n37045, n37046, n37047, n37048, n37049, n37050,
         n37051, n37052, n37053, n37054, n37055, n37056, n37057, n37058,
         n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066,
         n37067, n37068, n37069, n37070, n37071, n37072, n37073, n37074,
         n37075, n37076, n37077, n37078, n37079, n37080, n37081, n37082,
         n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090,
         n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098,
         n37099, n37100, n37101, n37102, n37103, n37104, n37105, n37106,
         n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114,
         n37115, n37116, n37117, n37118, n37119, n37120, n37121, n37122,
         n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130,
         n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138,
         n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146,
         n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154,
         n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162,
         n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170,
         n37171, n37172, n37173, n37174, n37175, n37176, n37177, n37178,
         n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186,
         n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194,
         n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202,
         n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210,
         n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218,
         n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226,
         n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234,
         n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242,
         n37243, n37244, n37245, n37246, n37247, n37248, n37249, n37250,
         n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258,
         n37259, n37260, n37261, n37262, n37263, n37264, n37265, n37266,
         n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274,
         n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282,
         n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290,
         n37291, n37292, n37293, n37294, n37295, n37296, n37297, n37298,
         n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306,
         n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314,
         n37315, n37316, n37317, n37318, n37319, n37320, n37321, n37322,
         n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330,
         n37331, n37332, n37333, n37334, n37335, n37336, n37337, n37338,
         n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346,
         n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354,
         n37355, n37356, n37357, n37358, n37359, n37360, n37361, n37362,
         n37363, n37364, n37365, n37366, n37367, n37368, n37369, n37370,
         n37371, n37372, n37373, n37374, n37375, n37376, n37377, n37378,
         n37379, n37380, n37381, n37382, n37383, n37384, n37385, n37386,
         n37387, n37388, n37389, n37390, n37391, n37392, n37393, n37394,
         n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402,
         n37403, n37404, n37405, n37406, n37407, n37408, n37409, n37410,
         n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418,
         n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426,
         n37427, n37428, n37429, n37430, n37431, n37432, n37433, n37434,
         n37435, n37436, n37437, n37438, n37439, n37440, n37441, n37442,
         n37443, n37444, n37445, n37446, n37447, n37448, n37449, n37450,
         n37451, n37452, n37453, n37454, n37455, n37456, n37457, n37458,
         n37459, n37460, n37461, n37462, n37463, n37464, n37465, n37466,
         n37467, n37468, n37469, n37470, n37471, n37472, n37473, n37474,
         n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482,
         n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490,
         n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498,
         n37499, n37500, n37501, n37502, n37503, n37504, n37505, n37506,
         n37507, n37508, n37509, n37510, n37511, n37512, n37513, n37514,
         n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522,
         n37523, n37524, n37525, n37526, n37527, n37528, n37529, n37530,
         n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538,
         n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546,
         n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554,
         n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562,
         n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570,
         n37571, n37572, n37573, n37574, n37575, n37576, n37577, n37578,
         n37579, n37580, n37581, n37582, n37583, n37584, n37585, n37586,
         n37587, n37588, n37589, n37590, n37591, n37592, n37593, n37594,
         n37595, n37596, n37597, n37598, n37599, n37600, n37601, n37602,
         n37603, n37604, n37605, n37606, n37607, n37608, n37609, n37610,
         n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618,
         n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626,
         n37627, n37628, n37629, n37630, n37631, n37632, n37633, n37634,
         n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642,
         n37643, n37644, n37645, n37646, n37647, n37648, n37649, n37650,
         n37651, n37652, n37653, n37654, n37655, n37656, n37657, n37658,
         n37659, n37660, n37661, n37662, n37663, n37664, n37665, n37666,
         n37667, n37668, n37669, n37670, n37671, n37672, n37673, n37674,
         n37675, n37676, n37677, n37678, n37679, n37680, n37681, n37682,
         n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690,
         n37691, n37692, n37693, n37694, n37695, n37696, n37697, n37698,
         n37699, n37700, n37701, n37702, n37703, n37704, n37705, n37706,
         n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714,
         n37715, n37716, n37717, n37718, n37719, n37720, n37721, n37722,
         n37723, n37724, n37725, n37726, n37727, n37728, n37729, n37730,
         n37731, n37732, n37733, n37734, n37735, n37736, n37737, n37738,
         n37739, n37740, n37741, n37742, n37743, n37744, n37745, n37746,
         n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754,
         n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762,
         n37763, n37764, n37765, n37766, n37767, n37768, n37769, n37770,
         n37771, n37772, n37773, n37774, n37775, n37776, n37777, n37778,
         n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786,
         n37787, n37788, n37789, n37790, n37791, n37792, n37793, n37794,
         n37795, n37796, n37797, n37798, n37799, n37800, n37801, n37802,
         n37803, n37804, n37805, n37806, n37807, n37808, n37809, n37810,
         n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818,
         n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37826,
         n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834,
         n37835, n37836, n37837, n37838, n37839, n37840, n37841, n37842,
         n37843, n37844, n37845, n37846, n37847, n37848, n37849, n37850,
         n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858,
         n37859, n37860, n37861, n37862, n37863, n37864, n37865, n37866,
         n37867, n37868, n37869, n37870, n37871, n37872, n37873, n37874,
         n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882,
         n37883, n37884, n37885, n37886, n37887, n37888, n37889, n37890,
         n37891, n37892, n37893, n37894, n37895, n37896, n37897, n37898,
         n37899, n37900, n37901, n37902, n37903, n37904, n37905, n37906,
         n37907, n37908, n37909, n37910, n37911, n37912, n37913, n37914,
         n37915, n37916, n37917, n37918, n37919, n37920, n37921, n37922,
         n37923, n37924, n37925, n37926, n37927, n37928, n37929, n37930,
         n37931, n37932, n37933, n37934, n37935, n37936, n37937, n37938,
         n37939, n37940, n37941, n37942, n37943, n37944, n37945, n37946,
         n37947, n37948, n37949, n37950, n37951, n37952, n37953, n37954,
         n37955, n37956, n37957, n37958, n37959, n37960, n37961, n37962,
         n37963, n37964, n37965, n37966, n37967, n37968, n37969, n37970,
         n37971, n37972, n37973, n37974, n37975, n37976, n37977, n37978,
         n37979, n37980, n37981, n37982, n37983, n37984, n37985, n37986,
         n37987, n37988, n37989, n37990, n37991, n37992, n37993, n37994,
         n37995, n37996, n37997, n37998, n37999, n38000, n38001, n38002,
         n38003, n38004, n38005, n38006, n38007, n38008, n38009, n38010,
         n38011, n38012, n38013, n38014, n38015, n38016, n38017, n38018,
         n38019, n38020, n38021, n38022, n38023, n38024, n38025, n38026,
         n38027, n38028, n38029, n38030, n38031, n38032, n38033, n38034,
         n38035, n38036, n38037, n38038, n38039, n38040, n38041, n38042,
         n38043, n38044, n38045, n38046, n38047, n38048, n38049, n38050,
         n38051, n38052, n38053, n38054, n38055, n38056, n38057, n38058,
         n38059, n38060, n38061, n38062, n38063, n38064, n38065, n38066,
         n38067, n38068, n38069, n38070, n38071, n38072, n38073, n38074,
         n38075, n38076, n38077, n38078, n38079, n38080, n38081, n38082,
         n38083, n38084, n38085, n38086, n38087, n38088, n38089, n38090,
         n38091, n38092, n38093, n38094, n38095, n38096, n38097, n38098,
         n38099, n38100, n38101, n38102, n38103, n38104, n38105, n38106,
         n38107, n38108, n38109, n38110, n38111, n38112, n38113, n38114,
         n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122,
         n38123, n38124, n38125, n38126, n38127, n38128, n38129, n38130,
         n38131, n38132, n38133, n38134, n38135, n38136, n38137, n38138,
         n38139, n38140, n38141, n38142, n38143, n38144, n38145, n38146,
         n38147, n38148, n38149, n38150, n38151, n38152, n38153, n38154,
         n38155, n38156, n38157, n38158, n38159, n38160, n38161, n38162,
         n38163, n38164, n38165, n38166, n38167, n38168, n38169, n38170,
         n38171, n38172, n38173, n38174, n38175, n38176, n38177, n38178,
         n38179, n38180, n38181, n38182, n38183, n38184, n38185, n38186,
         n38187, n38188, n38189, n38190, n38191, n38192, n38193, n38194,
         n38195, n38196, n38197, n38198, n38199, n38200, n38201, n38202,
         n38203, n38204, n38205, n38206, n38207, n38208, n38209, n38210,
         n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218,
         n38219, n38220, n38221, n38222, n38223, n38224, n38225, n38226,
         n38227, n38228, n38229, n38230, n38231, n38232, n38233, n38234,
         n38235, n38236, n38237, n38238, n38239, n38240, n38241, n38242,
         n38243, n38244, n38245, n38246, n38247, n38248, n38249, n38250,
         n38251, n38252, n38253, n38254, n38255, n38256, n38257, n38258,
         n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38266,
         n38267, n38268, n38269, n38270, n38271, n38272, n38273, n38274,
         n38275, n38276, n38277, n38278, n38279, n38280, n38281, n38282,
         n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290,
         n38291, n38292, n38293, n38294, n38295, n38296, n38297, n38298,
         n38299, n38300, n38301, n38302, n38303, n38304, n38305, n38306,
         n38307, n38308, n38309, n38310, n38311, n38312, n38313, n38314,
         n38315, n38316, n38317, n38318, n38319, n38320, n38321, n38322,
         n38323, n38324, n38325, n38326, n38327, n38328, n38329, n38330,
         n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338,
         n38339, n38340, n38341, n38342, n38343, n38344, n38345, n38346,
         n38347, n38348, n38349, n38350, n38351, n38352, n38353, n38354,
         n38355, n38356, n38357, n38358, n38359, n38360, n38361, n38362,
         n38363, n38364, n38365, n38366, n38367, n38368, n38369, n38370,
         n38371, n38372, n38373, n38374, n38375, n38376, n38377, n38378,
         n38379, n38380, n38381, n38382, n38383, n38384, n38385, n38386,
         n38387, n38388, n38389, n38390, n38391, n38392, n38393, n38394,
         n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402,
         n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410,
         n38411, n38412, n38413, n38414, n38415, n38416, n38417, n38418,
         n38419, n38420, n38421, n38422, n38423, n38424, n38425, n38426,
         n38427, n38428, n38429, n38430, n38431, n38432, n38433, n38434,
         n38435, n38436, n38437, n38438, n38439, n38440, n38441, n38442,
         n38443, n38444, n38445, n38446, n38447, n38448, n38449, n38450,
         n38451, n38452, n38453, n38454, n38455, n38456, n38457, n38458,
         n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466,
         n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474,
         n38475, n38476, n38477, n38478, n38479, n38480, n38481, n38482,
         n38483, n38484, n38485, n38486, n38487, n38488, n38489, n38490,
         n38491, n38492, n38493, n38494, n38495, n38496, n38497, n38498,
         n38499, n38500, n38501, n38502, n38503, n38504, n38505, n38506,
         n38507, n38508, n38509, n38510, n38511, n38512, n38513, n38514,
         n38515, n38516, n38517, n38518, n38519, n38520, n38521, n38522,
         n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530,
         n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538,
         n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546,
         n38547, n38548, n38549, n38550, n38551, n38552, n38553, n38554,
         n38555, n38556, n38557, n38558, n38559, n38560, n38561, n38562,
         n38563, n38564, n38565, n38566, n38567, n38568, n38569, n38570,
         n38571, n38572, n38573, n38574, n38575, n38576, n38577, n38578,
         n38579, n38580, n38581, n38582, n38583, n38584, n38585, n38586,
         n38587, n38588, n38589, n38590, n38591, n38592, n38593, n38594,
         n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602,
         n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610,
         n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618,
         n38619, n38620, n38621, n38622, n38623, n38624, n38625, n38626,
         n38627, n38628, n38629, n38630, n38631, n38632, n38633, n38634,
         n38635, n38636, n38637, n38638, n38639, n38640, n38641, n38642,
         n38643, n38644, n38645, n38646, n38647, n38648, n38649, n38650,
         n38651, n38652, n38653, n38654, n38655, n38656, n38657, n38658,
         n38659, n38660, n38661, n38662, n38663, n38664, n38665, n38666,
         n38667, n38668, n38669, n38670, n38671, n38672, n38673, n38674,
         n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682,
         n38683, n38684, n38685, n38686, n38687, n38688, n38689, n38690,
         n38691, n38692, n38693, n38694, n38695, n38696, n38697, n38698,
         n38699, n38700, n38701, n38702, n38703, n38704, n38705, n38706,
         n38707, n38708, n38709, n38710, n38711, n38712, n38713, n38714,
         n38715, n38716, n38717, n38718, n38719, n38720, n38721, n38722,
         n38723, n38724, n38725, n38726, n38727, n38728, n38729, n38730,
         n38731, n38732, n38733, n38734, n38735, n38736, n38737, n38738,
         n38739, n38740, n38741, n38742, n38743, n38744, n38745, n38746,
         n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754,
         n38755, n38756, n38757, n38758, n38759, n38760, n38761, n38762,
         n38763, n38764, n38765, n38766, n38767, n38768, n38769, n38770,
         n38771, n38772, n38773, n38774, n38775, n38776, n38777, n38778,
         n38779, n38780, n38781, n38782, n38783, n38784, n38785, n38786,
         n38787, n38788, n38789, n38790, n38791, n38792, n38793, n38794,
         n38795, n38796, n38797, n38798, n38799, n38800, n38801, n38802,
         n38803, n38804, n38805, n38806, n38807, n38808, n38809, n38810,
         n38811, n38812, n38813, n38814, n38815, n38816, n38817, n38818,
         n38819, n38820, n38821, n38822, n38823, n38824, n38825, n38826,
         n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834,
         n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842,
         n38843, n38844, n38845, n38846, n38847, n38848, n38849, n38850,
         n38851, n38852, n38853, n38854, n38855, n38856, n38857, n38858,
         n38859, n38860, n38861, n38862, n38863, n38864, n38865, n38866,
         n38867, n38868, n38869, n38870, n38871, n38872, n38873, n38874,
         n38875, n38876, n38877, n38878, n38879, n38880, n38881, n38882,
         n38883, n38884, n38885, n38886, n38887, n38888, n38889, n38890,
         n38891, n38892, n38893, n38894, n38895, n38896, n38897, n38898,
         n38899, n38900, n38901, n38902, n38903, n38904, n38905, n38906,
         n38907, n38908, n38909, n38910, n38911, n38912, n38913, n38914,
         n38915, n38916, n38917, n38918, n38919, n38920, n38921, n38922,
         n38923, n38924, n38925, n38926, n38927, n38928, n38929, n38930,
         n38931, n38932, n38933, n38934, n38935, n38936, n38937, n38938,
         n38939, n38940, n38941, n38942, n38943, n38944, n38945, n38946,
         n38947, n38948, n38949, n38950, n38951, n38952, n38953, n38954,
         n38955, n38956, n38957, n38958, n38959, n38960, n38961, n38962,
         n38963, n38964, n38965, n38966, n38967, n38968, n38969, n38970,
         n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38978,
         n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986,
         n38987, n38988, n38989, n38990, n38991, n38992, n38993, n38994,
         n38995, n38996, n38997, n38998, n38999, n39000, n39001, n39002,
         n39003, n39004, n39005, n39006, n39007, n39008, n39009, n39010,
         n39011, n39012, n39013, n39014, n39015, n39016, n39017, n39018,
         n39019, n39020, n39021, n39022, n39023, n39024, n39025, n39026,
         n39027, n39028, n39029, n39030, n39031, n39032, n39033, n39034,
         n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042,
         n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050,
         n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058,
         n39059, n39060, n39061, n39062, n39063, n39064, n39065, n39066,
         n39067, n39068, n39069, n39070, n39071, n39072, n39073, n39074,
         n39075, n39076, n39077, n39078, n39079, n39080, n39081, n39082,
         n39083, n39084, n39085, n39086, n39087, n39088, n39089, n39090,
         n39091, n39092, n39093, n39094, n39095, n39096, n39097, n39098,
         n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106,
         n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114,
         n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122,
         n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130,
         n39131, n39132, n39133, n39134, n39135, n39136, n39137, n39138,
         n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146,
         n39147, n39148, n39149, n39150, n39151, n39152, n39153, n39154,
         n39155, n39156, n39157, n39158, n39159, n39160, n39161, n39162,
         n39163, n39164, n39165, n39166, n39167, n39168, n39169, n39170,
         n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178,
         n39179, n39180, n39181, n39182, n39183, n39184, n39185, n39186,
         n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39194,
         n39195, n39196, n39197, n39198, n39199, n39200, n39201, n39202,
         n39203, n39204, n39205, n39206, n39207, n39208, n39209, n39210,
         n39211, n39212, n39213, n39214, n39215, n39216, n39217, n39218,
         n39219, n39220, n39221, n39222, n39223, n39224, n39225, n39226,
         n39227, n39228, n39229, n39230, n39231, n39232, n39233, n39234,
         n39235, n39236, n39237, n39238, n39239, n39240, n39241, n39242,
         n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250,
         n39251, n39252, n39253, n39254, n39255, n39256, n39257, n39258,
         n39259, n39260, n39261, n39262, n39263, n39264, n39265, n39266,
         n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39274,
         n39275, n39276, n39277, n39278, n39279, n39280, n39281, n39282,
         n39283, n39284, n39285, n39286, n39287, n39288, n39289, n39290,
         n39291, n39292, n39293, n39294, n39295, n39296, n39297, n39298,
         n39299, n39300, n39301, n39302, n39303, n39304, n39305, n39306,
         n39307, n39308, n39309, n39310, n39311, n39312, n39313, n39314,
         n39315, n39316, n39317, n39318, n39319, n39320, n39321, n39322,
         n39323, n39324, n39325, n39326, n39327, n39328, n39329, n39330,
         n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338,
         n39339, n39340, n39341, n39342, n39343, n39344, n39345, n39346,
         n39347, n39348, n39349, n39350, n39351, n39352, n39353, n39354,
         n39355, n39356, n39357, n39358, n39359, n39360, n39361, n39362,
         n39363, n39364, n39365, n39366, n39367, n39368, n39369, n39370,
         n39371, n39372, n39373, n39374, n39375, n39376, n39377, n39378,
         n39379, n39380, n39381, n39382, n39383, n39384, n39385, n39386,
         n39387, n39388, n39389, n39390, n39391, n39392, n39393, n39394,
         n39395, n39396, n39397, n39398, n39399, n39400, n39401, n39402,
         n39403, n39404, n39405, n39406, n39407, n39408, n39409, n39410,
         n39411, n39412, n39413, n39414, n39415, n39416, n39417, n39418,
         n39419, n39420, n39421, n39422, n39423, n39424, n39425, n39426,
         n39427, n39428, n39429, n39430, n39431, n39432, n39433, n39434,
         n39435, n39436, n39437, n39438, n39439, n39440, n39441, n39442,
         n39443, n39444, n39445, n39446, n39447, n39448, n39449, n39450,
         n39451, n39452, n39453, n39454, n39455, n39456, n39457, n39458,
         n39459, n39460, n39461, n39462, n39463, n39464, n39465, n39466,
         n39467, n39468, n39469, n39470, n39471, n39472, n39473, n39474,
         n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482,
         n39483, n39484, n39485, n39486, n39487, n39488, n39489, n39490,
         n39491, n39492, n39493, n39494, n39495, n39496, n39497, n39498,
         n39499, n39500, n39501, n39502, n39503, n39504, n39505, n39506,
         n39507, n39508, n39509, n39510, n39511, n39512, n39513, n39514,
         n39515, n39516, n39517, n39518, n39519, n39520, n39521, n39522,
         n39523, n39524, n39525, n39526, n39527, n39528, n39529, n39530,
         n39531, n39532, n39533, n39534, n39535, n39536, n39537, n39538,
         n39539, n39540, n39541, n39542, n39543, n39544, n39545, n39546,
         n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554,
         n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562,
         n39563, n39564, n39565, n39566, n39567, n39568, n39569, n39570,
         n39571, n39572, n39573, n39574, n39575, n39576, n39577, n39578,
         n39579, n39580, n39581, n39582, n39583, n39584, n39585, n39586,
         n39587, n39588, n39589, n39590, n39591, n39592, n39593, n39594,
         n39595, n39596, n39597, n39598, n39599, n39600, n39601, n39602,
         n39603, n39604, n39605, n39606, n39607, n39608, n39609, n39610,
         n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39618,
         n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626,
         n39627, n39628, n39629, n39630, n39631, n39632, n39633, n39634,
         n39635, n39636, n39637, n39638, n39639, n39640, n39641, n39642,
         n39643, n39644, n39645, n39646, n39647, n39648, n39649, n39650,
         n39651, n39652, n39653, n39654, n39655, n39656, n39657, n39658,
         n39659, n39660, n39661, n39662, n39663, n39664, n39665, n39666,
         n39667, n39668, n39669, n39670, n39671, n39672, n39673, n39674,
         n39675, n39676, n39677, n39678, n39679, n39680, n39681, n39682,
         n39683, n39684, n39685, n39686, n39687, n39688, n39689, n39690,
         n39691, n39692, n39693, n39694, n39695, n39696, n39697, n39698,
         n39699, n39700, n39701, n39702, n39703, n39704, n39705, n39706,
         n39707, n39708, n39709, n39710, n39711, n39712, n39713, n39714,
         n39715, n39716, n39717, n39718, n39719, n39720, n39721, n39722,
         n39723, n39724, n39725, n39726, n39727, n39728, n39729, n39730,
         n39731, n39732, n39733, n39734, n39735, n39736, n39737, n39738,
         n39739, n39740, n39741, n39742, n39743, n39744, n39745, n39746,
         n39747, n39748, n39749, n39750, n39751, n39752, n39753, n39754,
         n39755, n39756, n39757, n39758, n39759, n39760, n39761, n39762,
         n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770,
         n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778,
         n39779, n39780, n39781, n39782, n39783, n39784, n39785, n39786,
         n39787, n39788, n39789, n39790, n39791, n39792, n39793, n39794,
         n39795, n39796, n39797, n39798, n39799, n39800, n39801, n39802,
         n39803, n39804, n39805, n39806, n39807, n39808, n39809, n39810,
         n39811, n39812, n39813, n39814, n39815, n39816, n39817, n39818,
         n39819, n39820, n39821, n39822, n39823, n39824, n39825, n39826,
         n39827, n39828, n39829, n39830, n39831, n39832, n39833, n39834,
         n39835, n39836, n39837, n39838, n39839, n39840, n39841, n39842,
         n39843, n39844, n39845, n39846, n39847, n39848, n39849, n39850,
         n39851, n39852, n39853, n39854, n39855, n39856, n39857, n39858,
         n39859, n39860, n39861, n39862, n39863, n39864, n39865, n39866,
         n39867, n39868, n39869, n39870, n39871, n39872, n39873, n39874,
         n39875, n39876, n39877, n39878, n39879, n39880, n39881, n39882,
         n39883, n39884, n39885, n39886, n39887, n39888, n39889, n39890,
         n39891, n39892, n39893, n39894, n39895, n39896, n39897, n39898,
         n39899, n39900, n39901, n39902, n39903, n39904, n39905, n39906,
         n39907, n39908, n39909, n39910, n39911, n39912, n39913, n39914,
         n39915, n39916, n39917, n39918, n39919, n39920, n39921, n39922,
         n39923, n39924, n39925, n39926, n39927, n39928, n39929, n39930,
         n39931, n39932, n39933, n39934, n39935, n39936, n39937, n39938,
         n39939, n39940, n39941, n39942, n39943, n39944, n39945, n39946,
         n39947, n39948, n39949, n39950, n39951, n39952, n39953, n39954,
         n39955, n39956, n39957, n39958, n39959, n39960, n39961, n39962,
         n39963, n39964, n39965, n39966, n39967, n39968, n39969, n39970,
         n39971, n39972, n39973, n39974, n39975, n39976, n39977, n39978,
         n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39986,
         n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994,
         n39995, n39996, n39997, n39998, n39999, n40000, n40001, n40002,
         n40003, n40004, n40005, n40006, n40007, n40008, n40009, n40010,
         n40011, n40012, n40013, n40014, n40015, n40016, n40017, n40018,
         n40019, n40020, n40021, n40022, n40023, n40024, n40025, n40026,
         n40027, n40028, n40029, n40030, n40031, n40032, n40033, n40034,
         n40035, n40036, n40037, n40038, n40039, n40040, n40041, n40042,
         n40043, n40044, n40045, n40046, n40047, n40048, n40049, n40050,
         n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058,
         n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066,
         n40067, n40068, n40069, n40070, n40071, n40072, n40073, n40074,
         n40075, n40076, n40077, n40078, n40079, n40080, n40081, n40082,
         n40083, n40084, n40085, n40086, n40087, n40088, n40089, n40090,
         n40091, n40092, n40093, n40094, n40095, n40096, n40097, n40098,
         n40099, n40100, n40101, n40102, n40103, n40104, n40105, n40106,
         n40107, n40108, n40109, n40110, n40111, n40112, n40113, n40114,
         n40115, n40116, n40117, n40118, n40119, n40120, n40121, n40122,
         n40123, n40124, n40125, n40126, n40127, n40128, n40129, n40130,
         n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138,
         n40139, n40140, n40141, n40142, n40143, n40144, n40145, n40146,
         n40147, n40148, n40149, n40150, n40151, n40152, n40153, n40154,
         n40155, n40156, n40157, n40158, n40159, n40160, n40161, n40162,
         n40163, n40164, n40165, n40166, n40167, n40168, n40169, n40170,
         n40171, n40172, n40173, n40174, n40175, n40176, n40177, n40178,
         n40179, n40180, n40181, n40182, n40183, n40184, n40185, n40186,
         n40187, n40188, n40189, n40190, n40191, n40192, n40193, n40194,
         n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202,
         n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210,
         n40211, n40212, n40213, n40214, n40215, n40216, n40217, n40218,
         n40219, n40220, n40221, n40222, n40223, n40224, n40225, n40226,
         n40227, n40228, n40229, n40230, n40231, n40232, n40233, n40234,
         n40235, n40236, n40237, n40238, n40239, n40240, n40241, n40242,
         n40243, n40244, n40245, n40246, n40247, n40248, n40249, n40250,
         n40251, n40252, n40253, n40254, n40255, n40256, n40257, n40258,
         n40259, n40260, n40261, n40262, n40263, n40264, n40265, n40266,
         n40267, n40268, n40269, n40270, n40271, n40272, n40273, n40274,
         n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282,
         n40283, n40284, n40285, n40286, n40287, n40288, n40289, n40290,
         n40291, n40292, n40293, n40294, n40295, n40296, n40297, n40298,
         n40299, n40300, n40301, n40302, n40303, n40304, n40305, n40306,
         n40307, n40308, n40309, n40310, n40311, n40312, n40313, n40314,
         n40315, n40316, n40317, n40318, n40319, n40320, n40321, n40322,
         n40323, n40324, n40325, n40326, n40327, n40328, n40329, n40330,
         n40331, n40332, n40333, n40334, n40335, n40336, n40337, n40338,
         n40339, n40340, n40341, n40342, n40343, n40344, n40345, n40346,
         n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354,
         n40355, n40356, n40357, n40358, n40359, n40360, n40361, n40362,
         n40363, n40364, n40365, n40366, n40367, n40368, n40369, n40370,
         n40371, n40372, n40373, n40374, n40375, n40376, n40377, n40378,
         n40379, n40380, n40381, n40382, n40383, n40384, n40385, n40386,
         n40387, n40388, n40389, n40390, n40391, n40392, n40393, n40394,
         n40395, n40396, n40397, n40398, n40399, n40400, n40401, n40402,
         n40403, n40404, n40405, n40406, n40407, n40408, n40409, n40410,
         n40411, n40412, n40413, n40414, n40415, n40416, n40417, n40418,
         n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426,
         n40427, n40428, n40429, n40430, n40431, n40432, n40433, n40434,
         n40435, n40436, n40437, n40438, n40439, n40440, n40441, n40442,
         n40443, n40444, n40445, n40446, n40447, n40448, n40449, n40450,
         n40451, n40452, n40453, n40454, n40455, n40456, n40457, n40458,
         n40459, n40460, n40461, n40462, n40463, n40464, n40465, n40466,
         n40467, n40468, n40469, n40470, n40471, n40472, n40473, n40474,
         n40475, n40476, n40477, n40478, n40479, n40480, n40481, n40482,
         n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490,
         n40491, n40492, n40493, n40494, n40495, n40496, n40497, n40498,
         n40499, n40500, n40501, n40502, n40503, n40504, n40505, n40506,
         n40507, n40508, n40509, n40510, n40511, n40512, n40513, n40514,
         n40515, n40516, n40517, n40518, n40519, n40520, n40521, n40522,
         n40523, n40524, n40525, n40526, n40527, n40528, n40529, n40530,
         n40531, n40532, n40533, n40534, n40535, n40536, n40537, n40538,
         n40539, n40540, n40541, n40542, n40543, n40544, n40545, n40546,
         n40547, n40548, n40549, n40550, n40551, n40552, n40553, n40554,
         n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562,
         n40563, n40564, n40565, n40566, n40567, n40568, n40569, n40570,
         n40571, n40572, n40573, n40574, n40575, n40576, n40577, n40578,
         n40579, n40580, n40581, n40582, n40583, n40584, n40585, n40586,
         n40587, n40588, n40589, n40590, n40591, n40592, n40593, n40594,
         n40595, n40596, n40597, n40598, n40599, n40600, n40601, n40602,
         n40603, n40604, n40605, n40606, n40607, n40608, n40609, n40610,
         n40611, n40612, n40613, n40614, n40615, n40616, n40617, n40618,
         n40619, n40620, n40621, n40622, n40623, n40624, n40625, n40626,
         n40627, n40628, n40629, n40630, n40631, n40632, n40633, n40634,
         n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642,
         n40643, n40644, n40645, n40646, n40647, n40648, n40649, n40650,
         n40651, n40652, n40653, n40654, n40655, n40656, n40657, n40658,
         n40659, n40660, n40661, n40662, n40663, n40664, n40665, n40666,
         n40667, n40668, n40669, n40670, n40671, n40672, n40673, n40674,
         n40675, n40676, n40677, n40678, n40679, n40680, n40681, n40682,
         n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690,
         n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698,
         n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706,
         n40707, n40708, n40709, n40710, n40711, n40712, n40713, n40714,
         n40715, n40716, n40717, n40718, n40719, n40720, n40721, n40722,
         n40723, n40724, n40725, n40726, n40727, n40728, n40729, n40730,
         n40731, n40732, n40733, n40734, n40735, n40736, n40737, n40738,
         n40739, n40740, n40741, n40742, n40743, n40744, n40745, n40746,
         n40747, n40748, n40749, n40750, n40751, n40752, n40753, n40754,
         n40755, n40756, n40757, n40758, n40759, n40760, n40761, n40762,
         n40763, n40764, n40765, n40766, n40767, n40768, n40769, n40770,
         n40771, n40772, n40773, n40774, n40775, n40776, n40777, n40778,
         n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786,
         n40787, n40788, n40789, n40790, n40791, n40792, n40793, n40794,
         n40795, n40796, n40797, n40798, n40799, n40800, n40801, n40802,
         n40803, n40804, n40805, n40806, n40807, n40808, n40809, n40810,
         n40811, n40812, n40813, n40814, n40815, n40816, n40817, n40818,
         n40819, n40820, n40821, n40822, n40823, n40824, n40825, n40826,
         n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834,
         n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842,
         n40843, n40844, n40845, n40846, n40847, n40848, n40849, n40850,
         n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40858,
         n40859, n40860, n40861, n40862, n40863, n40864, n40865, n40866,
         n40867, n40868, n40869, n40870, n40871, n40872, n40873, n40874,
         n40875, n40876, n40877, n40878, n40879, n40880, n40881, n40882,
         n40883, n40884, n40885, n40886, n40887, n40888, n40889, n40890,
         n40891, n40892, n40893, n40894, n40895, n40896, n40897, n40898,
         n40899, n40900, n40901, n40902, n40903, n40904, n40905, n40906,
         n40907, n40908, n40909, n40910, n40911, n40912, n40913, n40914,
         n40915, n40916, n40917, n40918, n40919, n40920, n40921, n40922,
         n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930,
         n40931, n40932, n40933, n40934, n40935, n40936, n40937, n40938,
         n40939, n40940, n40941, n40942, n40943, n40944, n40945, n40946,
         n40947, n40948, n40949, n40950, n40951, n40952, n40953, n40954,
         n40955, n40956, n40957, n40958, n40959, n40960, n40961, n40962,
         n40963, n40964, n40965, n40966, n40967, n40968, n40969, n40970,
         n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40978,
         n40979, n40980, n40981, n40982, n40983, n40984, n40985, n40986,
         n40987, n40988, n40989, n40990, n40991, n40992, n40993, n40994,
         n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002,
         n41003, n41004, n41005, n41006, n41007, n41008, n41009, n41010,
         n41011, n41012, n41013, n41014, n41015, n41016, n41017, n41018,
         n41019, n41020, n41021, n41022, n41023, n41024, n41025, n41026,
         n41027, n41028, n41029, n41030, n41031, n41032, n41033, n41034,
         n41035, n41036, n41037, n41038, n41039, n41040, n41041, n41042,
         n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050,
         n41051, n41052, n41053, n41054, n41055, n41056, n41057, n41058,
         n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066,
         n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074,
         n41075, n41076, n41077, n41078, n41079, n41080, n41081, n41082,
         n41083, n41084, n41085, n41086, n41087, n41088, n41089, n41090,
         n41091, n41092, n41093, n41094, n41095, n41096, n41097, n41098,
         n41099, n41100, n41101, n41102, n41103, n41104, n41105, n41106,
         n41107, n41108, n41109, n41110, n41111, n41112, n41113, n41114,
         n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122,
         n41123, n41124, n41125, n41126, n41127, n41128, n41129, n41130,
         n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138,
         n41139, n41140, n41141, n41142, n41143, n41144, n41145, n41146,
         n41147, n41148, n41149, n41150, n41151, n41152, n41153, n41154,
         n41155, n41156, n41157, n41158, n41159, n41160, n41161, n41162,
         n41163, n41164, n41165, n41166, n41167, n41168, n41169, n41170,
         n41171, n41172, n41173, n41174, n41175, n41176, n41177, n41178,
         n41179, n41180, n41181, n41182, n41183, n41184, n41185, n41186,
         n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194,
         n41195, n41196, n41197, n41198, n41199, n41200, n41201, n41202,
         n41203, n41204, n41205, n41206, n41207, n41208, n41209, n41210,
         n41211, n41212, n41213, n41214, n41215, n41216, n41217, n41218,
         n41219, n41220, n41221, n41222, n41223, n41224, n41225, n41226,
         n41227, n41228, n41229, n41230, n41231, n41232, n41233, n41234,
         n41235, n41236, n41237, n41238, n41239, n41240, n41241, n41242,
         n41243, n41244, n41245, n41246, n41247, n41248, n41249, n41250,
         n41251, n41252, n41253, n41254, n41255, n41256, n41257, n41258,
         n41259, n41260, n41261, n41262, n41263, n41264, n41265, n41266,
         n41267, n41268, n41269, n41270, n41271, n41272, n41273, n41274,
         n41275, n41276, n41277, n41278, n41279, n41280, n41281, n41282,
         n41283, n41284, n41285, n41286, n41287, n41288, n41289, n41290,
         n41291, n41292, n41293, n41294, n41295, n41296, n41297, n41298,
         n41299, n41300, n41301, n41302, n41303, n41304, n41305, n41306,
         n41307, n41308, n41309, n41310, n41311, n41312, n41313, n41314,
         n41315, n41316, n41317, n41318, n41319, n41320, n41321, n41322,
         n41323, n41324, n41325, n41326, n41327, n41328, n41329, n41330,
         n41331, n41332, n41333, n41334, n41335, n41336, n41337, n41338,
         n41339, n41340, n41341, n41342, n41343, n41344, n41345, n41346,
         n41347, n41348, n41349, n41350, n41351, n41352, n41353, n41354,
         n41355, n41356, n41357, n41358, n41359, n41360, n41361, n41362,
         n41363, n41364, n41365, n41366, n41367, n41368, n41369, n41370,
         n41371, n41372, n41373, n41374, n41375, n41376, n41377, n41378,
         n41379, n41380, n41381, n41382, n41383, n41384, n41385, n41386,
         n41387, n41388, n41389, n41390, n41391, n41392, n41393, n41394,
         n41395, n41396, n41397, n41398, n41399, n41400, n41401, n41402,
         n41403, n41404, n41405, n41406, n41407, n41408, n41409, n41410,
         n41411, n41412, n41413, n41414, n41415, n41416, n41417, n41418,
         n41419, n41420, n41421, n41422, n41423, n41424, n41425, n41426,
         n41427, n41428, n41429, n41430, n41431, n41432, n41433, n41434,
         n41435, n41436, n41437, n41438, n41439, n41440, n41441, n41442,
         n41443, n41444, n41445, n41446, n41447, n41448, n41449, n41450,
         n41451, n41452, n41453, n41454, n41455, n41456, n41457, n41458,
         n41459, n41460, n41461, n41462, n41463, n41464, n41465, n41466,
         n41467, n41468, n41469, n41470, n41471, n41472, n41473, n41474,
         n41475, n41476, n41477, n41478, n41479, n41480, n41481, n41482,
         n41483, n41484, n41485, n41486, n41487, n41488, n41489, n41490,
         n41491, n41492, n41493, n41494, n41495, n41496, n41497, n41498,
         n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506,
         n41507, n41508, n41509, n41510, n41511, n41512, n41513, n41514,
         n41515, n41516, n41517, n41518, n41519, n41520, n41521, n41522,
         n41523, n41524, n41525, n41526, n41527, n41528, n41529, n41530,
         n41531, n41532, n41533, n41534, n41535, n41536, n41537, n41538,
         n41539, n41540, n41541, n41542, n41543, n41544, n41545, n41546,
         n41547, n41548, n41549, n41550, n41551, n41552, n41553, n41554,
         n41555, n41556, n41557, n41558, n41559, n41560, n41561, n41562,
         n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570,
         n41571, n41572, n41573, n41574, n41575, n41576, n41577, n41578,
         n41579, n41580, n41581, n41582, n41583, n41584, n41585, n41586,
         n41587, n41588, n41589, n41590, n41591, n41592, n41593, n41594,
         n41595, n41596, n41597, n41598, n41599, n41600, n41601, n41602,
         n41603, n41604, n41605, n41606, n41607, n41608, n41609, n41610,
         n41611, n41612, n41613, n41614, n41615, n41616, n41617, n41618,
         n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626,
         n41627, n41628, n41629, n41630, n41631, n41632, n41633, n41634,
         n41635, n41636, n41637, n41638, n41639, n41640, n41641, n41642,
         n41643, n41644, n41645, n41646, n41647, n41648, n41649, n41650,
         n41651, n41652, n41653, n41654, n41655, n41656, n41657, n41658,
         n41659, n41660, n41661, n41662, n41663, n41664, n41665, n41666,
         n41667, n41668, n41669, n41670, n41671, n41672, n41673, n41674,
         n41675, n41676, n41677, n41678, n41679, n41680, n41681, n41682,
         n41683, n41684, n41685, n41686, n41687, n41688, n41689, n41690,
         n41691, n41692, n41693, n41694, n41695, n41696, n41697, n41698,
         n41699, n41700, n41701, n41702, n41703, n41704, n41705, n41706,
         n41707, n41708, n41709, n41710, n41711, n41712, n41713, n41714,
         n41715, n41716, n41717, n41718, n41719, n41720, n41721, n41722,
         n41723, n41724, n41725, n41726, n41727, n41728, n41729, n41730,
         n41731, n41732, n41733, n41734, n41735, n41736, n41737, n41738,
         n41739, n41740, n41741, n41742, n41743, n41744, n41745, n41746,
         n41747, n41748, n41749, n41750, n41751, n41752, n41753, n41754,
         n41755, n41756, n41757, n41758, n41759, n41760, n41761, n41762,
         n41763, n41764, n41765, n41766, n41767, n41768, n41769, n41770,
         n41771, n41772, n41773, n41774, n41775, n41776, n41777, n41778,
         n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786,
         n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794,
         n41795, n41796, n41797, n41798, n41799, n41800, n41801, n41802,
         n41803, n41804, n41805, n41806, n41807, n41808, n41809, n41810,
         n41811, n41812, n41813, n41814, n41815, n41816, n41817, n41818,
         n41819, n41820, n41821, n41822, n41823, n41824, n41825, n41826,
         n41827, n41828, n41829, n41830, n41831, n41832, n41833, n41834,
         n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842,
         n41843, n41844, n41845, n41846, n41847, n41848, n41849, n41850,
         n41851, n41852, n41853, n41854, n41855, n41856, n41857, n41858,
         n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866,
         n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874,
         n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882,
         n41883, n41884, n41885, n41886, n41887, n41888, n41889, n41890,
         n41891, n41892, n41893, n41894, n41895, n41896, n41897, n41898,
         n41899, n41900, n41901, n41902, n41903, n41904, n41905, n41906,
         n41907, n41908, n41909, n41910, n41911, n41912, n41913, n41914,
         n41915, n41916, n41917, n41918, n41919, n41920, n41921, n41922,
         n41923, n41924, n41925, n41926, n41927, n41928, n41929, n41930,
         n41931, n41932, n41933, n41934, n41935, n41936, n41937, n41938,
         n41939, n41940, n41941, n41942, n41943, n41944, n41945, n41946,
         n41947, n41948, n41949, n41950, n41951, n41952, n41953, n41954,
         n41955, n41956, n41957, n41958, n41959, n41960, n41961, n41962,
         n41963, n41964, n41965, n41966, n41967, n41968, n41969, n41970,
         n41971, n41972, n41973, n41974, n41975, n41976, n41977, n41978,
         n41979, n41980, n41981, n41982, n41983, n41984, n41985, n41986,
         n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41994,
         n41995, n41996, n41997, n41998, n41999, n42000, n42001, n42002,
         n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010,
         n42011, n42012, n42013, n42014, n42015, n42016, n42017, n42018,
         n42019, n42020, n42021, n42022, n42023, n42024, n42025, n42026,
         n42027, n42028, n42029, n42030, n42031, n42032, n42033, n42034,
         n42035, n42036, n42037, n42038, n42039, n42040, n42041, n42042,
         n42043, n42044, n42045, n42046, n42047, n42048, n42049, n42050,
         n42051, n42052, n42053, n42054, n42055, n42056, n42057, n42058,
         n42059, n42060, n42061, n42062, n42063, n42064, n42065, n42066,
         n42067, n42068, n42069, n42070, n42071, n42072, n42073, n42074,
         n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082,
         n42083, n42084, n42085, n42086, n42087, n42088, n42089, n42090,
         n42091, n42092, n42093, n42094, n42095, n42096, n42097, n42098,
         n42099, n42100, n42101, n42102, n42103, n42104, n42105, n42106,
         n42107, n42108, n42109, n42110, n42111, n42112, n42113, n42114,
         n42115, n42116, n42117, n42118, n42119, n42120, n42121, n42122,
         n42123, n42124, n42125, n42126, n42127, n42128, n42129, n42130,
         n42131, n42132, n42133, n42134, n42135, n42136, n42137, n42138,
         n42139, n42140, n42141, n42142, n42143, n42144, n42145, n42146,
         n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154,
         n42155, n42156, n42157, n42158, n42159, n42160, n42161, n42162,
         n42163, n42164, n42165, n42166, n42167, n42168, n42169, n42170,
         n42171, n42172, n42173, n42174, n42175, n42176, n42177, n42178,
         n42179, n42180, n42181, n42182, n42183, n42184, n42185, n42186,
         n42187, n42188, n42189, n42190, n42191, n42192, n42193, n42194,
         n42195, n42196, n42197, n42198, n42199, n42200, n42201, n42202,
         n42203, n42204, n42205, n42206, n42207, n42208, n42209, n42210,
         n42211, n42212, n42213, n42214, n42215, n42216, n42217, n42218,
         n42219, n42220, n42221, n42222, n42223, n42224, n42225, n42226,
         n42227, n42228, n42229, n42230, n42231, n42232, n42233, n42234,
         n42235, n42236, n42237, n42238, n42239, n42240, n42241, n42242,
         n42243, n42244, n42245, n42246, n42247, n42248, n42249, n42250,
         n42251, n42252, n42253, n42254, n42255, n42256, n42257, n42258,
         n42259, n42260, n42261, n42262, n42263, n42264, n42265, n42266,
         n42267, n42268, n42269, n42270, n42271, n42272, n42273, n42274,
         n42275, n42276, n42277, n42278, n42279, n42280, n42281, n42282,
         n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290,
         n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298,
         n42299, n42300, n42301, n42302, n42303, n42304, n42305, n42306,
         n42307, n42308, n42309, n42310, n42311, n42312, n42313, n42314,
         n42315, n42316, n42317, n42318, n42319, n42320, n42321, n42322,
         n42323, n42324, n42325, n42326, n42327, n42328, n42329, n42330,
         n42331, n42332, n42333, n42334, n42335, n42336, n42337, n42338,
         n42339, n42340, n42341, n42342, n42343, n42344, n42345, n42346,
         n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354,
         n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362,
         n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370,
         n42371, n42372, n42373, n42374, n42375, n42376, n42377, n42378,
         n42379, n42380, n42381, n42382, n42383, n42384, n42385, n42386,
         n42387, n42388, n42389, n42390, n42391, n42392, n42393, n42394,
         n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402,
         n42403, n42404, n42405, n42406, n42407, n42408, n42409, n42410,
         n42411, n42412, n42413, n42414, n42415, n42416, n42417, n42418,
         n42419, n42420, n42421, n42422, n42423, n42424, n42425, n42426,
         n42427, n42428, n42429, n42430, n42431, n42432, n42433, n42434,
         n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442,
         n42443, n42444, n42445, n42446, n42447, n42448, n42449, n42450,
         n42451, n42452, n42453, n42454, n42455, n42456, n42457, n42458,
         n42459, n42460, n42461, n42462, n42463, n42464, n42465, n42466,
         n42467, n42468, n42469, n42470, n42471, n42472, n42473, n42474,
         n42475, n42476, n42477, n42478, n42479, n42480, n42481, n42482,
         n42483, n42484, n42485, n42486, n42487, n42488, n42489, n42490,
         n42491, n42492, n42493, n42494, n42495, n42496, n42497, n42498,
         n42499, n42500, n42501, n42502, n42503, n42504, n42505, n42506,
         n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514,
         n42515, n42516, n42517, n42518, n42519, n42520, n42521, n42522,
         n42523, n42524, n42525, n42526, n42527, n42528, n42529, n42530,
         n42531, n42532, n42533, n42534, n42535, n42536, n42537, n42538,
         n42539, n42540, n42541, n42542, n42543, n42544, n42545, n42546,
         n42547, n42548, n42549, n42550, n42551, n42552, n42553, n42554,
         n42555, n42556, n42557, n42558, n42559, n42560, n42561, n42562,
         n42563, n42564, n42565, n42566, n42567, n42568, n42569, n42570,
         n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42578,
         n42579, n42580, n42581, n42582, n42583, n42584, n42585, n42586,
         n42587, n42588, n42589, n42590, n42591, n42592, n42593, n42594,
         n42595, n42596, n42597, n42598, n42599, n42600, n42601, n42602,
         n42603, n42604, n42605, n42606, n42607, n42608, n42609, n42610,
         n42611, n42612, n42613, n42614, n42615, n42616, n42617, n42618,
         n42619, n42620, n42621, n42622, n42623, n42624, n42625, n42626,
         n42627, n42628, n42629, n42630, n42631, n42632, n42633, n42634,
         n42635, n42636, n42637, n42638, n42639, n42640, n42641, n42642,
         n42643, n42644, n42645, n42646, n42647, n42648, n42649, n42650,
         n42651, n42652, n42653, n42654, n42655, n42656, n42657, n42658,
         n42659, n42660, n42661, n42662, n42663, n42664, n42665, n42666,
         n42667, n42668, n42669, n42670, n42671, n42672, n42673, n42674,
         n42675, n42676, n42677, n42678, n42679, n42680, n42681, n42682,
         n42683, n42684, n42685, n42686, n42687, n42688, n42689, n42690,
         n42691, n42692, n42693, n42694, n42695, n42696, n42697, n42698,
         n42699, n42700, n42701, n42702, n42703, n42704, n42705, n42706,
         n42707, n42708, n42709, n42710, n42711, n42712, n42713, n42714,
         n42715, n42716, n42717, n42718, n42719, n42720, n42721, n42722,
         n42723, n42724, n42725, n42726, n42727, n42728, n42729, n42730,
         n42731, n42732, n42733, n42734, n42735, n42736, n42737, n42738,
         n42739, n42740, n42741, n42742, n42743, n42744, n42745, n42746,
         n42747, n42748, n42749, n42750, n42751, n42752, n42753, n42754,
         n42755, n42756, n42757, n42758, n42759, n42760, n42761, n42762,
         n42763, n42764, n42765, n42766, n42767, n42768, n42769, n42770,
         n42771, n42772, n42773, n42774, n42775, n42776, n42777, n42778,
         n42779, n42780, n42781, n42782, n42783, n42784, n42785, n42786,
         n42787, n42788, n42789, n42790, n42791, n42792, n42793, n42794,
         n42795, n42796, n42797, n42798, n42799, n42800, n42801, n42802,
         n42803, n42804, n42805, n42806, n42807, n42808, n42809, n42810,
         n42811, n42812, n42813, n42814, n42815, n42816, n42817, n42818,
         n42819, n42820, n42821, n42822, n42823, n42824, n42825, n42826,
         n42827, n42828, n42829, n42830, n42831, n42832, n42833, n42834,
         n42835, n42836, n42837, n42838, n42839, n42840, n42841, n42842,
         n42843, n42844, n42845, n42846, n42847, n42848, n42849, n42850,
         n42851, n42852, n42853, n42854, n42855, n42856, n42857, n42858,
         n42859, n42860, n42861, n42862, n42863, n42864, n42865, n42866,
         n42867, n42868, n42869, n42870, n42871, n42872, n42873, n42874,
         n42875, n42876, n42877, n42878, n42879, n42880, n42881, n42882,
         n42883, n42884, n42885, n42886, n42887, n42888, n42889, n42890,
         n42891, n42892, n42893, n42894, n42895, n42896, n42897, n42898,
         n42899, n42900, n42901, n42902, n42903, n42904, n42905, n42906,
         n42907, n42908, n42909, n42910, n42911, n42912, n42913, n42914,
         n42915, n42916, n42917, n42918, n42919, n42920, n42921, n42922,
         n42923, n42924, n42925, n42926, n42927, n42928, n42929, n42930,
         n42931, n42932, n42933, n42934, n42935, n42936, n42937, n42938,
         n42939, n42940, n42941, n42942, n42943, n42944, n42945, n42946,
         n42947, n42948, n42949, n42950, n42951, n42952, n42953, n42954,
         n42955, n42956, n42957, n42958, n42959, n42960, n42961, n42962,
         n42963, n42964, n42965, n42966, n42967, n42968, n42969, n42970,
         n42971, n42972, n42973, n42974, n42975, n42976, n42977, n42978,
         n42979, n42980, n42981, n42982, n42983, n42984, n42985, n42986,
         n42987, n42988, n42989, n42990, n42991, n42992, n42993, n42994,
         n42995, n42996, n42997, n42998, n42999, n43000, n43001, n43002,
         n43003, n43004, n43005, n43006, n43007, n43008, n43009, n43010,
         n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018,
         n43019, n43020, n43021, n43022, n43023, n43024, n43025, n43026,
         n43027, n43028, n43029, n43030, n43031, n43032, n43033, n43034,
         n43035, n43036, n43037, n43038, n43039, n43040, n43041, n43042,
         n43043, n43044, n43045, n43046, n43047, n43048, n43049, n43050,
         n43051, n43052, n43053, n43054, n43055, n43056, n43057, n43058,
         n43059, n43060, n43061, n43062, n43063, n43064, n43065, n43066,
         n43067, n43068, n43069, n43070, n43071, n43072, n43073, n43074,
         n43075, n43076, n43077, n43078, n43079, n43080, n43081, n43082,
         n43083, n43084, n43085, n43086, n43087, n43088, n43089, n43090,
         n43091, n43092, n43093, n43094, n43095, n43096, n43097, n43098,
         n43099, n43100, n43101, n43102, n43103, n43104, n43105, n43106,
         n43107, n43108, n43109, n43110, n43111, n43112, n43113, n43114,
         n43115, n43116, n43117, n43118, n43119, n43120, n43121, n43122,
         n43123, n43124, n43125, n43126, n43127, n43128, n43129, n43130,
         n43131, n43132, n43133, n43134, n43135, n43136, n43137, n43138,
         n43139, n43140, n43141, n43142, n43143, n43144, n43145, n43146,
         n43147, n43148, n43149, n43150, n43151, n43152, n43153, n43154,
         n43155, n43156, n43157, n43158, n43159, n43160, n43161, n43162,
         n43163, n43164, n43165, n43166, n43167, n43168, n43169, n43170,
         n43171, n43172, n43173, n43174, n43175, n43176, n43177, n43178,
         n43179, n43180, n43181, n43182, n43183, n43184, n43185, n43186,
         n43187, n43188, n43189, n43190, n43191, n43192, n43193, n43194,
         n43195, n43196, n43197, n43198, n43199, n43200, n43201, n43202,
         n43203, n43204, n43205, n43206, n43207, n43208, n43209, n43210,
         n43211, n43212, n43213, n43214, n43215, n43216, n43217, n43218,
         n43219, n43220, n43221, n43222, n43223, n43224, n43225, n43226,
         n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234,
         n43235, n43236, n43237, n43238, n43239, n43240, n43241, n43242,
         n43243, n43244, n43245, n43246, n43247, n43248, n43249, n43250,
         n43251, n43252, n43253, n43254, n43255, n43256, n43257, n43258,
         n43259, n43260, n43261, n43262, n43263, n43264, n43265, n43266,
         n43267, n43268, n43269, n43270, n43271, n43272, n43273, n43274,
         n43275, n43276, n43277, n43278, n43279, n43280, n43281, n43282,
         n43283, n43284, n43285, n43286, n43287, n43288, n43289, n43290,
         n43291, n43292, n43293, n43294, n43295, n43296, n43297, n43298,
         n43299, n43300, n43301, n43302, n43303, n43304, n43305, n43306,
         n43307, n43308, n43309, n43310, n43311, n43312, n43313, n43314,
         n43315, n43316, n43317, n43318, n43319, n43320, n43321, n43322,
         n43323, n43324, n43325, n43326, n43327, n43328, n43329, n43330,
         n43331, n43332, n43333, n43334, n43335, n43336, n43337, n43338,
         n43339, n43340, n43341, n43342, n43343, n43344, n43345, n43346,
         n43347, n43348, n43349, n43350, n43351, n43352, n43353, n43354,
         n43355, n43356, n43357, n43358, n43359, n43360, n43361, n43362,
         n43363, n43364, n43365, n43366, n43367, n43368, n43369, n43370,
         n43371, n43372, n43373, n43374, n43375, n43376, n43377, n43378,
         n43379, n43380, n43381, n43382, n43383, n43384, n43385, n43386,
         n43387, n43388, n43389, n43390, n43391, n43392, n43393, n43394,
         n43395, n43396, n43397, n43398, n43399, n43400, n43401, n43402,
         n43403, n43404, n43405, n43406, n43407, n43408, n43409, n43410,
         n43411, n43412, n43413, n43414, n43415, n43416, n43417, n43418,
         n43419, n43420, n43421, n43422, n43423, n43424, n43425, n43426,
         n43427, n43428, n43429, n43430, n43431, n43432, n43433, n43434,
         n43435, n43436, n43437, n43438, n43439, n43440, n43441, n43442,
         n43443, n43444, n43445, n43446, n43447, n43448, n43449, n43450,
         n43451, n43452, n43453, n43454, n43455, n43456, n43457, n43458,
         n43459, n43460, n43461, n43462, n43463, n43464, n43465, n43466,
         n43467, n43468, n43469, n43470, n43471, n43472, n43473, n43474,
         n43475, n43476, n43477, n43478, n43479, n43480, n43481, n43482,
         n43483, n43484, n43485, n43486, n43487, n43488, n43489, n43490,
         n43491, n43492, n43493, n43494, n43495, n43496, n43497, n43498,
         n43499, n43500, n43501, n43502, n43503, n43504, n43505, n43506,
         n43507, n43508, n43509, n43510, n43511, n43512, n43513, n43514,
         n43515, n43516, n43517, n43518, n43519, n43520, n43521, n43522,
         n43523, n43524, n43525, n43526, n43527, n43528, n43529, n43530,
         n43531, n43532, n43533, n43534, n43535, n43536, n43537, n43538,
         n43539, n43540, n43541, n43542, n43543, n43544, n43545, n43546,
         n43547, n43548, n43549, n43550, n43551, n43552, n43553, n43554,
         n43555, n43556, n43557, n43558, n43559, n43560, n43561, n43562,
         n43563, n43564, n43565, n43566, n43567, n43568, n43569, n43570,
         n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578,
         n43579, n43580, n43581, n43582, n43583, n43584, n43585, n43586,
         n43587, n43588, n43589, n43590, n43591, n43592, n43593, n43594,
         n43595, n43596, n43597, n43598, n43599, n43600, n43601, n43602,
         n43603, n43604, n43605, n43606, n43607, n43608, n43609, n43610,
         n43611, n43612, n43613, n43614, n43615, n43616, n43617, n43618,
         n43619, n43620, n43621, n43622, n43623, n43624, n43625, n43626,
         n43627, n43628, n43629, n43630, n43631, n43632, n43633, n43634,
         n43635, n43636, n43637, n43638, n43639, n43640, n43641, n43642,
         n43643, n43644, n43645, n43646, n43647, n43648, n43649, n43650,
         n43651, n43652, n43653, n43654, n43655, n43656, n43657, n43658,
         n43659, n43660, n43661, n43662, n43663, n43664, n43665, n43666,
         n43667, n43668, n43669, n43670, n43671, n43672, n43673, n43674,
         n43675, n43676, n43677, n43678, n43679, n43680, n43681, n43682,
         n43683, n43684, n43685, n43686, n43687, n43688, n43689, n43690,
         n43691, n43692, n43693, n43694, n43695, n43696, n43697, n43698,
         n43699, n43700, n43701, n43702, n43703, n43704, n43705, n43706,
         n43707, n43708, n43709, n43710, n43711, n43712, n43713, n43714,
         n43715, n43716, n43717, n43718, n43719, n43720, n43721, n43722,
         n43723, n43724, n43725, n43726, n43727, n43728, n43729, n43730,
         n43731, n43732, n43733, n43734, n43735, n43736, n43737, n43738,
         n43739, n43740, n43741, n43742, n43743, n43744, n43745, n43746,
         n43747, n43748, n43749, n43750, n43751, n43752, n43753, n43754,
         n43755, n43756, n43757, n43758, n43759, n43760, n43761, n43762,
         n43763, n43764, n43765, n43766, n43767, n43768, n43769, n43770,
         n43771, n43772, n43773, n43774, n43775, n43776, n43777, n43778,
         n43779, n43780, n43781, n43782, n43783, n43784, n43785, n43786,
         n43787, n43788, n43789, n43790, n43791, n43792, n43793, n43794,
         n43795, n43796, n43797, n43798, n43799, n43800, n43801, n43802,
         n43803, n43804, n43805, n43806, n43807, n43808, n43809, n43810,
         n43811, n43812, n43813, n43814, n43815, n43816, n43817, n43818,
         n43819, n43820, n43821, n43822, n43823, n43824, n43825, n43826,
         n43827, n43828, n43829, n43830, n43831, n43832, n43833, n43834,
         n43835, n43836, n43837, n43838, n43839, n43840, n43841, n43842,
         n43843, n43844, n43845, n43846, n43847, n43848, n43849, n43850,
         n43851, n43852, n43853, n43854, n43855, n43856, n43857, n43858,
         n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866,
         n43867, n43868, n43869, n43870, n43871, n43872, n43873, n43874,
         n43875, n43876, n43877, n43878, n43879, n43880, n43881, n43882,
         n43883, n43884, n43885, n43886, n43887, n43888, n43889, n43890,
         n43891, n43892, n43893, n43894, n43895, n43896, n43897, n43898,
         n43899, n43900, n43901, n43902, n43903, n43904, n43905, n43906,
         n43907, n43908, n43909, n43910, n43911, n43912, n43913, n43914,
         n43915, n43916, n43917, n43918, n43919, n43920, n43921, n43922,
         n43923, n43924, n43925, n43926, n43927, n43928, n43929, n43930,
         n43931, n43932, n43933, n43934, n43935, n43936, n43937, n43938,
         n43939, n43940, n43941, n43942, n43943, n43944, n43945, n43946,
         n43947, n43948, n43949, n43950, n43951, n43952, n43953, n43954,
         n43955, n43956, n43957, n43958, n43959, n43960, n43961, n43962,
         n43963, n43964, n43965, n43966, n43967, n43968, n43969, n43970,
         n43971, n43972, n43973, n43974, n43975, n43976, n43977, n43978,
         n43979, n43980, n43981, n43982, n43983, n43984, n43985, n43986,
         n43987, n43988, n43989, n43990, n43991, n43992, n43993, n43994,
         n43995, n43996, n43997, n43998, n43999, n44000, n44001, n44002,
         n44003, n44004, n44005, n44006, n44007, n44008, n44009, n44010,
         n44011, n44012, n44013, n44014, n44015, n44016, n44017, n44018,
         n44019, n44020, n44021, n44022, n44023, n44024, n44025, n44026,
         n44027, n44028, n44029, n44030, n44031, n44032, n44033, n44034,
         n44035, n44036, n44037, n44038, n44039, n44040, n44041, n44042,
         n44043, n44044, n44045, n44046, n44047, n44048, n44049, n44050,
         n44051, n44052, n44053, n44054, n44055, n44056, n44057, n44058,
         n44059, n44060, n44061, n44062, n44063, n44064, n44065, n44066,
         n44067, n44068, n44069, n44070, n44071, n44072, n44073, n44074,
         n44075, n44076, n44077, n44078, n44079, n44080, n44081, n44082,
         n44083, n44084, n44085, n44086, n44087, n44088, n44089, n44090,
         n44091, n44092, n44093, n44094, n44095, n44096, n44097, n44098,
         n44099, n44100, n44101, n44102, n44103, n44104, n44105, n44106,
         n44107, n44108, n44109, n44110, n44111, n44112, n44113, n44114,
         n44115, n44116, n44117, n44118, n44119, n44120, n44121, n44122,
         n44123, n44124, n44125, n44126, n44127, n44128, n44129, n44130,
         n44131, n44132, n44133, n44134, n44135, n44136, n44137, n44138,
         n44139, n44140, n44141, n44142, n44143, n44144, n44145, n44146,
         n44147, n44148, n44149, n44150, n44151, n44152, n44153, n44154,
         n44155, n44156, n44157, n44158, n44159, n44160, n44161, n44162,
         n44163, n44164, n44165, n44166, n44167, n44168, n44169, n44170,
         n44171, n44172, n44173, n44174, n44175, n44176, n44177, n44178,
         n44179, n44180, n44181, n44182, n44183, n44184, n44185, n44186,
         n44187, n44188, n44189, n44190, n44191, n44192, n44193, n44194,
         n44195, n44196, n44197, n44198, n44199, n44200, n44201, n44202,
         n44203, n44204, n44205, n44206, n44207, n44208, n44209, n44210,
         n44211, n44212, n44213, n44214, n44215, n44216, n44217, n44218,
         n44219, n44220, n44221, n44222, n44223, n44224, n44225, n44226,
         n44227, n44228, n44229, n44230, n44231, n44232, n44233, n44234,
         n44235, n44236, n44237, n44238, n44239, n44240, n44241, n44242,
         n44243, n44244, n44245, n44246, n44247, n44248, n44249, n44250,
         n44251, n44252, n44253, n44254, n44255, n44256, n44257, n44258,
         n44259, n44260, n44261, n44262, n44263, n44264, n44265, n44266,
         n44267, n44268, n44269, n44270, n44271, n44272, n44273, n44274,
         n44275, n44276, n44277, n44278, n44279, n44280, n44281, n44282,
         n44283, n44284, n44285, n44286, n44287, n44288, n44289, n44290,
         n44291, n44292, n44293, n44294, n44295, n44296, n44297, n44298,
         n44299, n44300, n44301, n44302, n44303, n44304, n44305, n44306,
         n44307, n44308, n44309, n44310, n44311, n44312, n44313, n44314,
         n44315, n44316, n44317, n44318, n44319, n44320, n44321, n44322,
         n44323, n44324, n44325, n44326, n44327, n44328, n44329, n44330,
         n44331, n44332, n44333, n44334, n44335, n44336, n44337, n44338,
         n44339, n44340, n44341, n44342, n44343, n44344, n44345, n44346,
         n44347, n44348, n44349, n44350, n44351, n44352, n44353, n44354,
         n44355, n44356, n44357, n44358, n44359, n44360, n44361, n44362,
         n44363, n44364, n44365, n44366, n44367, n44368, n44369, n44370,
         n44371, n44372, n44373, n44374, n44375, n44376, n44377, n44378,
         n44379, n44380, n44381, n44382, n44383, n44384, n44385, n44386,
         n44387, n44388, n44389, n44390, n44391, n44392, n44393, n44394,
         n44395, n44396, n44397, n44398, n44399, n44400, n44401, n44402,
         n44403, n44404, n44405, n44406, n44407, n44408, n44409, n44410,
         n44411, n44412, n44413, n44414, n44415, n44416, n44417, n44418,
         n44419, n44420, n44421, n44422, n44423, n44424, n44425, n44426,
         n44427, n44428, n44429, n44430, n44431, n44432, n44433, n44434,
         n44435, n44436, n44437, n44438, n44439, n44440, n44441, n44442,
         n44443, n44444, n44445, n44446, n44447, n44448, n44449, n44450,
         n44451, n44452, n44453, n44454, n44455, n44456, n44457, n44458,
         n44459, n44460, n44461, n44462, n44463, n44464, n44465, n44466,
         n44467, n44468, n44469, n44470, n44471, n44472, n44473, n44474,
         n44475, n44476, n44477, n44478, n44479, n44480, n44481, n44482,
         n44483, n44484, n44485, n44486, n44487, n44488, n44489, n44490,
         n44491, n44492, n44493, n44494, n44495, n44496, n44497, n44498,
         n44499, n44500, n44501, n44502, n44503, n44504, n44505, n44506,
         n44507, n44508, n44509, n44510, n44511, n44512, n44513, n44514,
         n44515, n44516, n44517, n44518, n44519, n44520, n44521, n44522,
         n44523, n44524, n44525, n44526, n44527, n44528, n44529, n44530,
         n44531, n44532, n44533, n44534, n44535, n44536, n44537, n44538,
         n44539, n44540, n44541, n44542, n44543, n44544, n44545, n44546,
         n44547, n44548, n44549, n44550, n44551, n44552, n44553, n44554,
         n44555, n44556, n44557, n44558, n44559, n44560, n44561, n44562,
         n44563, n44564, n44565, n44566, n44567, n44568, n44569, n44570,
         n44571, n44572, n44573, n44574, n44575, n44576, n44577, n44578,
         n44579, n44580, n44581, n44582, n44583, n44584, n44585, n44586,
         n44587, n44588, n44589, n44590, n44591, n44592, n44593, n44594,
         n44595, n44596, n44597, n44598, n44599, n44600, n44601, n44602,
         n44603, n44604, n44605, n44606, n44607, n44608, n44609, n44610,
         n44611, n44612, n44613, n44614, n44615, n44616, n44617, n44618,
         n44619, n44620, n44621, n44622, n44623, n44624, n44625, n44626,
         n44627, n44628, n44629, n44630, n44631, n44632, n44633, n44634,
         n44635, n44636, n44637, n44638, n44639, n44640, n44641, n44642,
         n44643, n44644, n44645, n44646, n44647, n44648, n44649, n44650,
         n44651, n44652, n44653, n44654, n44655, n44656, n44657, n44658,
         n44659, n44660, n44661, n44662, n44663, n44664, n44665, n44666,
         n44667, n44668, n44669, n44670, n44671, n44672, n44673, n44674,
         n44675, n44676, n44677, n44678, n44679, n44680, n44681, n44682,
         n44683, n44684, n44685, n44686, n44687, n44688, n44689, n44690,
         n44691, n44692, n44693, n44694, n44695, n44696, n44697, n44698,
         n44699, n44700, n44701, n44702, n44703, n44704, n44705, n44706,
         n44707, n44708, n44709, n44710, n44711, n44712, n44713, n44714,
         n44715, n44716, n44717, n44718, n44719, n44720, n44721, n44722,
         n44723, n44724, n44725, n44726, n44727, n44728, n44729, n44730,
         n44731, n44732, n44733, n44734, n44735, n44736, n44737, n44738,
         n44739, n44740, n44741, n44742, n44743, n44744, n44745, n44746,
         n44747, n44748, n44749, n44750, n44751, n44752, n44753, n44754,
         n44755, n44756, n44757, n44758, n44759, n44760, n44761, n44762,
         n44763, n44764, n44765, n44766, n44767, n44768, n44769, n44770,
         n44771, n44772, n44773, n44774, n44775, n44776, n44777, n44778,
         n44779, n44780, n44781, n44782, n44783, n44784, n44785, n44786,
         n44787, n44788, n44789, n44790, n44791, n44792, n44793, n44794,
         n44795, n44796, n44797, n44798, n44799, n44800, n44801, n44802,
         n44803, n44804, n44805, n44806, n44807, n44808, n44809, n44810,
         n44811, n44812, n44813, n44814, n44815, n44816, n44817, n44818,
         n44819, n44820, n44821, n44822, n44823, n44824, n44825, n44826,
         n44827, n44828, n44829, n44830, n44831, n44832, n44833, n44834,
         n44835, n44836, n44837, n44838, n44839, n44840, n44841, n44842,
         n44843, n44844, n44845, n44846, n44847, n44848, n44849, n44850,
         n44851, n44852, n44853, n44854, n44855, n44856, n44857, n44858,
         n44859, n44860, n44861, n44862, n44863, n44864, n44865, n44866,
         n44867, n44868, n44869, n44870, n44871, n44872, n44873, n44874,
         n44875, n44876, n44877, n44878, n44879, n44880, n44881, n44882,
         n44883, n44884, n44885, n44886, n44887, n44888, n44889, n44890,
         n44891, n44892, n44893, n44894, n44895, n44896, n44897, n44898,
         n44899, n44900, n44901, n44902, n44903, n44904, n44905, n44906,
         n44907, n44908, n44909, n44910, n44911, n44912, n44913, n44914,
         n44915, n44916, n44917, n44918, n44919, n44920, n44921, n44922,
         n44923, n44924, n44925, n44926, n44927, n44928, n44929, n44930,
         n44931, n44932, n44933, n44934, n44935, n44936, n44937, n44938,
         n44939, n44940, n44941, n44942, n44943, n44944, n44945, n44946,
         n44947, n44948, n44949, n44950, n44951, n44952, n44953, n44954,
         n44955, n44956, n44957, n44958, n44959, n44960, n44961, n44962,
         n44963, n44964, n44965, n44966, n44967, n44968, n44969, n44970,
         n44971, n44972, n44973, n44974, n44975, n44976, n44977, n44978,
         n44979, n44980, n44981, n44982, n44983, n44984, n44985, n44986,
         n44987, n44988, n44989, n44990, n44991, n44992, n44993, n44994,
         n44995, n44996, n44997, n44998, n44999, n45000, n45001, n45002,
         n45003, n45004, n45005, n45006, n45007, n45008, n45009, n45010,
         n45011, n45012, n45013, n45014, n45015, n45016, n45017, n45018,
         n45019, n45020, n45021, n45022, n45023, n45024, n45025, n45026,
         n45027, n45028, n45029, n45030, n45031, n45032, n45033, n45034,
         n45035, n45036, n45037, n45038, n45039, n45040, n45041, n45042,
         n45043, n45044, n45045, n45046, n45047, n45048, n45049, n45050,
         n45051, n45052, n45053, n45054, n45055, n45056, n45057, n45058,
         n45059, n45060, n45061, n45062, n45063, n45064, n45065, n45066,
         n45067, n45068, n45069, n45070, n45071, n45072, n45073, n45074,
         n45075, n45076, n45077, n45078, n45079, n45080, n45081, n45082,
         n45083, n45084, n45085, n45086, n45087, n45088, n45089, n45090,
         n45091, n45092, n45093, n45094, n45095, n45096, n45097, n45098,
         n45099, n45100, n45101, n45102, n45103, n45104, n45105, n45106,
         n45107, n45108, n45109, n45110, n45111, n45112, n45113, n45114,
         n45115, n45116, n45117, n45118, n45119, n45120, n45121, n45122,
         n45123, n45124, n45125, n45126, n45127, n45128, n45129, n45130,
         n45131, n45132, n45133, n45134, n45135, n45136, n45137, n45138,
         n45139, n45140, n45141, n45142, n45143, n45144, n45145, n45146,
         n45147, n45148, n45149, n45150, n45151, n45152, n45153, n45154,
         n45155, n45156, n45157, n45158, n45159, n45160, n45161, n45162,
         n45163, n45164, n45165, n45166, n45167, n45168, n45169, n45170,
         n45171, n45172, n45173, n45174, n45175, n45176, n45177, n45178,
         n45179, n45180, n45181, n45182, n45183, n45184, n45185, n45186,
         n45187, n45188, n45189, n45190, n45191, n45192, n45193, n45194,
         n45195, n45196, n45197, n45198, n45199, n45200, n45201, n45202,
         n45203, n45204, n45205, n45206, n45207, n45208, n45209, n45210,
         n45211, n45212, n45213, n45214, n45215, n45216, n45217, n45218,
         n45219, n45220, n45221, n45222, n45223, n45224, n45225, n45226,
         n45227, n45228, n45229, n45230, n45231, n45232, n45233, n45234,
         n45235, n45236, n45237, n45238, n45239, n45240, n45241, n45242,
         n45243, n45244, n45245, n45246, n45247, n45248, n45249, n45250,
         n45251, n45252, n45253, n45254, n45255, n45256, n45257, n45258,
         n45259, n45260, n45261, n45262, n45263, n45264, n45265, n45266,
         n45267, n45268, n45269, n45270, n45271, n45272, n45273, n45274,
         n45275, n45276, n45277, n45278, n45279, n45280, n45281, n45282,
         n45283, n45284, n45285, n45286, n45287, n45288, n45289, n45290,
         n45291, n45292, n45293, n45294, n45295, n45296, n45297, n45298,
         n45299, n45300, n45301, n45302, n45303, n45304, n45305, n45306,
         n45307, n45308, n45309, n45310, n45311, n45312, n45313, n45314,
         n45315, n45316, n45317, n45318, n45319, n45320, n45321, n45322,
         n45323, n45324, n45325, n45326, n45327, n45328, n45329, n45330,
         n45331, n45332, n45333, n45334, n45335, n45336, n45337, n45338,
         n45339, n45340, n45341, n45342, n45343, n45344, n45345, n45346,
         n45347, n45348, n45349, n45350, n45351, n45352, n45353, n45354,
         n45355, n45356, n45357, n45358, n45359, n45360, n45361, n45362,
         n45363, n45364, n45365, n45366, n45367, n45368, n45369, n45370,
         n45371, n45372, n45373, n45374, n45375, n45376, n45377, n45378,
         n45379, n45380, n45381, n45382, n45383, n45384, n45385, n45386,
         n45387, n45388, n45389, n45390, n45391, n45392, n45393, n45394,
         n45395, n45396, n45397, n45398, n45399, n45400, n45401, n45402,
         n45403, n45404, n45405, n45406, n45407, n45408, n45409, n45410,
         n45411, n45412, n45413, n45414, n45415, n45416, n45417, n45418,
         n45419, n45420, n45421, n45422, n45423, n45424, n45425, n45426,
         n45427, n45428, n45429, n45430, n45431, n45432, n45433, n45434,
         n45435, n45436, n45437, n45438, n45439, n45440, n45441, n45442,
         n45443, n45444, n45445, n45446, n45447, n45448, n45449, n45450,
         n45451, n45452, n45453, n45454, n45455, n45456, n45457, n45458,
         n45459, n45460, n45461, n45462, n45463, n45464, n45465, n45466,
         n45467, n45468, n45469, n45470, n45471, n45472, n45473, n45474,
         n45475, n45476, n45477, n45478, n45479, n45480, n45481, n45482,
         n45483, n45484, n45485, n45486, n45487, n45488, n45489, n45490,
         n45491, n45492, n45493, n45494, n45495, n45496, n45497, n45498,
         n45499, n45500, n45501, n45502, n45503, n45504, n45505, n45506,
         n45507, n45508, n45509, n45510, n45511, n45512, n45513, n45514,
         n45515, n45516, n45517, n45518, n45519, n45520, n45521, n45522,
         n45523, n45524, n45525, n45526, n45527, n45528, n45529, n45530,
         n45531, n45532, n45533, n45534, n45535, n45536, n45537, n45538,
         n45539, n45540, n45541, n45542, n45543, n45544, n45545, n45546,
         n45547, n45548, n45549, n45550, n45551, n45552, n45553, n45554,
         n45555, n45556, n45557, n45558, n45559, n45560, n45561, n45562,
         n45563, n45564, n45565, n45566, n45567, n45568, n45569, n45570,
         n45571, n45572, n45573, n45574, n45575, n45576, n45577, n45578,
         n45579, n45580, n45581, n45582, n45583, n45584, n45585, n45586,
         n45587, n45588, n45589, n45590, n45591, n45592, n45593, n45594,
         n45595, n45596, n45597, n45598, n45599, n45600, n45601, n45602,
         n45603, n45604, n45605, n45606, n45607, n45608, n45609, n45610,
         n45611, n45612, n45613, n45614, n45615, n45616, n45617, n45618,
         n45619, n45620, n45621, n45622, n45623, n45624, n45625, n45626,
         n45627, n45628, n45629, n45630, n45631, n45632, n45633, n45634,
         n45635, n45636, n45637, n45638, n45639, n45640, n45641, n45642,
         n45643, n45644, n45645, n45646, n45647, n45648, n45649, n45650,
         n45651, n45652, n45653, n45654, n45655, n45656, n45657, n45658,
         n45659, n45660, n45661, n45662, n45663, n45664, n45665, n45666,
         n45667, n45668, n45669, n45670, n45671, n45672, n45673, n45674,
         n45675, n45676, n45677, n45678, n45679, n45680, n45681, n45682,
         n45683, n45684, n45685, n45686, n45687, n45688, n45689, n45690,
         n45691, n45692, n45693, n45694, n45695, n45696, n45697, n45698,
         n45699, n45700, n45701, n45702, n45703, n45704, n45705, n45706,
         n45707, n45708, n45709, n45710, n45711, n45712, n45713, n45714,
         n45715, n45716, n45717, n45718, n45719, n45720, n45721, n45722,
         n45723, n45724, n45725, n45726, n45727, n45728, n45729, n45730,
         n45731, n45732, n45733, n45734, n45735, n45736, n45737, n45738,
         n45739, n45740, n45741, n45742, n45743, n45744, n45745, n45746,
         n45747, n45748, n45749, n45750, n45751, n45752, n45753, n45754,
         n45755, n45756, n45757, n45758, n45759, n45760, n45761, n45762,
         n45763, n45764, n45765, n45766, n45767, n45768, n45769, n45770,
         n45771, n45772, n45773, n45774, n45775, n45776, n45777, n45778,
         n45779, n45780, n45781, n45782, n45783, n45784, n45785, n45786,
         n45787, n45788, n45789, n45790, n45791, n45792, n45793, n45794,
         n45795, n45796, n45797, n45798, n45799, n45800, n45801, n45802,
         n45803, n45804, n45805, n45806, n45807, n45808, n45809, n45810,
         n45811, n45812, n45813, n45814, n45815, n45816, n45817, n45818,
         n45819, n45820, n45821, n45822, n45823, n45824, n45825, n45826,
         n45827, n45828, n45829, n45830, n45831, n45832, n45833, n45834,
         n45835, n45836, n45837, n45838, n45839, n45840, n45841, n45842,
         n45843, n45844, n45845, n45846, n45847, n45848, n45849, n45850,
         n45851, n45852, n45853, n45854, n45855, n45856, n45857, n45858,
         n45859, n45860, n45861, n45862, n45863, n45864, n45865, n45866,
         n45867, n45868, n45869, n45870, n45871, n45872, n45873, n45874,
         n45875, n45876, n45877, n45878, n45879, n45880, n45881, n45882,
         n45883, n45884, n45885, n45886, n45887, n45888, n45889, n45890,
         n45891, n45892, n45893, n45894, n45895, n45896, n45897, n45898,
         n45899, n45900, n45901, n45902, n45903, n45904, n45905, n45906,
         n45907, n45908, n45909, n45910, n45911, n45912, n45913, n45914,
         n45915, n45916, n45917, n45918, n45919, n45920, n45921, n45922,
         n45923, n45924, n45925, n45926, n45927, n45928, n45929, n45930,
         n45931, n45932, n45933, n45934, n45935, n45936, n45937, n45938,
         n45939, n45940, n45941, n45942, n45943, n45944, n45945, n45946,
         n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45954,
         n45955, n45956, n45957, n45958, n45959, n45960, n45961, n45962,
         n45963, n45964, n45965, n45966, n45967, n45968, n45969, n45970,
         n45971, n45972, n45973, n45974, n45975, n45976, n45977, n45978,
         n45979, n45980, n45981, n45982, n45983, n45984, n45985, n45986,
         n45987, n45988, n45989, n45990, n45991, n45992, n45993, n45994,
         n45995, n45996, n45997, n45998, n45999, n46000, n46001, n46002,
         n46003, n46004, n46005, n46006, n46007, n46008, n46009, n46010,
         n46011, n46012, n46013, n46014, n46015, n46016, n46017, n46018,
         n46019, n46020, n46021, n46022, n46023, n46024, n46025, n46026,
         n46027, n46028, n46029, n46030, n46031, n46032, n46033, n46034,
         n46035, n46036, n46037, n46038, n46039, n46040, n46041, n46042,
         n46043, n46044, n46045, n46046, n46047, n46048, n46049, n46050,
         n46051, n46052, n46053, n46054, n46055, n46056, n46057, n46058,
         n46059, n46060, n46061, n46062, n46063, n46064, n46065, n46066,
         n46067, n46068, n46069, n46070, n46071, n46072, n46073, n46074,
         n46075, n46076, n46077, n46078, n46079, n46080, n46081, n46082,
         n46083, n46084, n46085, n46086, n46087, n46088, n46089, n46090,
         n46091, n46092, n46093, n46094, n46095, n46096, n46097, n46098,
         n46099, n46100, n46101, n46102, n46103, n46104, n46105, n46106,
         n46107, n46108, n46109, n46110, n46111, n46112, n46113, n46114,
         n46115, n46116, n46117, n46118, n46119, n46120, n46121, n46122,
         n46123, n46124, n46125, n46126, n46127, n46128, n46129, n46130,
         n46131, n46132, n46133, n46134, n46135, n46136, n46137, n46138,
         n46139, n46140, n46141, n46142, n46143, n46144, n46145, n46146,
         n46147, n46148, n46149, n46150, n46151, n46152, n46153, n46154,
         n46155, n46156, n46157, n46158, n46159, n46160, n46161, n46162,
         n46163, n46164, n46165, n46166, n46167, n46168, n46169, n46170,
         n46171, n46172, n46173, n46174, n46175, n46176, n46177, n46178,
         n46179, n46180, n46181, n46182, n46183, n46184, n46185, n46186,
         n46187, n46188, n46189, n46190, n46191, n46192, n46193, n46194,
         n46195, n46196, n46197, n46198, n46199, n46200, n46201, n46202,
         n46203, n46204, n46205, n46206, n46207, n46208, n46209, n46210,
         n46211, n46212, n46213, n46214, n46215, n46216, n46217, n46218,
         n46219, n46220, n46221, n46222, n46223, n46224, n46225, n46226,
         n46227, n46228, n46229, n46230, n46231, n46232, n46233, n46234,
         n46235, n46236, n46237, n46238, n46239, n46240, n46241, n46242,
         n46243, n46244, n46245, n46246, n46247, n46248, n46249, n46250,
         n46251, n46252, n46253, n46254, n46255, n46256, n46257, n46258,
         n46259, n46260, n46261, n46262, n46263, n46264, n46265, n46266,
         n46267, n46268, n46269, n46270, n46271, n46272, n46273, n46274,
         n46275, n46276, n46277, n46278, n46279, n46280, n46281, n46282,
         n46283, n46284, n46285, n46286, n46287, n46288, n46289, n46290,
         n46291, n46292, n46293, n46294, n46295, n46296, n46297, n46298,
         n46299, n46300, n46301, n46302, n46303, n46304, n46305, n46306,
         n46307, n46308, n46309, n46310, n46311, n46312, n46313, n46314,
         n46315, n46316, n46317, n46318, n46319, n46320, n46321, n46322,
         n46323, n46324, n46325, n46326, n46327, n46328, n46329, n46330,
         n46331, n46332, n46333, n46334, n46335, n46336, n46337, n46338,
         n46339, n46340, n46341, n46342, n46343, n46344, n46345, n46346,
         n46347, n46348, n46349, n46350, n46351, n46352, n46353, n46354,
         n46355, n46356, n46357, n46358, n46359, n46360, n46361, n46362,
         n46363, n46364, n46365, n46366, n46367, n46368, n46369, n46370,
         n46371, n46372, n46373, n46374, n46375, n46376, n46377, n46378,
         n46379, n46380, n46381, n46382, n46383, n46384, n46385, n46386,
         n46387, n46388, n46389, n46390, n46391, n46392, n46393, n46394,
         n46395, n46396, n46397, n46398, n46399, n46400, n46401, n46402,
         n46403, n46404, n46405, n46406, n46407, n46408, n46409, n46410,
         n46411, n46412, n46413, n46414, n46415, n46416, n46417, n46418,
         n46419, n46420, n46421, n46422, n46423, n46424, n46425, n46426,
         n46427, n46428, n46429, n46430, n46431, n46432, n46433, n46434,
         n46435, n46436, n46437, n46438, n46439, n46440, n46441, n46442,
         n46443, n46444, n46445, n46446, n46447, n46448, n46449, n46450,
         n46451, n46452, n46453, n46454, n46455, n46456, n46457, n46458,
         n46459, n46460, n46461, n46462, n46463, n46464, n46465, n46466,
         n46467, n46468, n46469, n46470, n46471, n46472, n46473, n46474,
         n46475, n46476, n46477, n46478, n46479, n46480, n46481, n46482,
         n46483, n46484, n46485, n46486, n46487, n46488, n46489, n46490,
         n46491, n46492, n46493, n46494, n46495, n46496, n46497, n46498,
         n46499, n46500, n46501, n46502, n46503, n46504, n46505, n46506,
         n46507, n46508, n46509, n46510, n46511, n46512, n46513, n46514,
         n46515, n46516, n46517, n46518, n46519, n46520, n46521, n46522,
         n46523, n46524, n46525, n46526, n46527, n46528, n46529, n46530,
         n46531, n46532, n46533, n46534, n46535, n46536, n46537, n46538,
         n46539, n46540, n46541, n46542, n46543, n46544, n46545, n46546,
         n46547, n46548, n46549, n46550, n46551, n46552, n46553, n46554,
         n46555, n46556, n46557, n46558, n46559, n46560, n46561, n46562,
         n46563, n46564, n46565, n46566, n46567, n46568, n46569, n46570,
         n46571, n46572, n46573, n46574, n46575, n46576, n46577, n46578,
         n46579, n46580, n46581, n46582, n46583, n46584, n46585, n46586,
         n46587, n46588, n46589, n46590, n46591, n46592, n46593, n46594,
         n46595, n46596, n46597, n46598, n46599, n46600, n46601, n46602,
         n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610,
         n46611, n46612, n46613, n46614, n46615, n46616, n46617, n46618,
         n46619, n46620, n46621, n46622, n46623, n46624, n46625, n46626,
         n46627, n46628, n46629, n46630, n46631, n46632, n46633, n46634,
         n46635, n46636, n46637, n46638, n46639, n46640, n46641, n46642,
         n46643, n46644, n46645, n46646, n46647, n46648, n46649, n46650,
         n46651, n46652, n46653, n46654, n46655, n46656, n46657, n46658,
         n46659, n46660, n46661, n46662, n46663, n46664, n46665, n46666,
         n46667, n46668, n46669, n46670, n46671, n46672, n46673, n46674,
         n46675, n46676, n46677, n46678, n46679, n46680, n46681, n46682,
         n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690,
         n46691, n46692, n46693, n46694, n46695, n46696, n46697, n46698,
         n46699, n46700, n46701, n46702, n46703, n46704, n46705, n46706,
         n46707, n46708, n46709, n46710, n46711, n46712, n46713, n46714,
         n46715, n46716, n46717, n46718, n46719, n46720, n46721, n46722,
         n46723, n46724, n46725, n46726, n46727, n46728, n46729, n46730,
         n46731, n46732, n46733, n46734, n46735, n46736, n46737, n46738,
         n46739, n46740, n46741, n46742, n46743, n46744, n46745, n46746,
         n46747, n46748, n46749, n46750, n46751, n46752, n46753, n46754,
         n46755, n46756, n46757, n46758, n46759, n46760, n46761, n46762,
         n46763, n46764, n46765, n46766, n46767, n46768, n46769, n46770,
         n46771, n46772, n46773, n46774, n46775, n46776, n46777, n46778,
         n46779, n46780, n46781, n46782, n46783, n46784, n46785, n46786,
         n46787, n46788, n46789, n46790, n46791, n46792, n46793, n46794,
         n46795, n46796, n46797, n46798, n46799, n46800, n46801, n46802,
         n46803, n46804, n46805, n46806, n46807, n46808, n46809, n46810,
         n46811, n46812, n46813, n46814, n46815, n46816, n46817, n46818,
         n46819, n46820, n46821, n46822, n46823, n46824, n46825, n46826,
         n46827, n46828, n46829, n46830, n46831, n46832, n46833, n46834,
         n46835, n46836, n46837, n46838, n46839, n46840, n46841, n46842,
         n46843, n46844, n46845, n46846, n46847, n46848, n46849, n46850,
         n46851, n46852, n46853, n46854, n46855, n46856, n46857, n46858,
         n46859, n46860, n46861, n46862, n46863, n46864, n46865, n46866,
         n46867, n46868, n46869, n46870, n46871, n46872, n46873, n46874,
         n46875, n46876, n46877, n46878, n46879, n46880, n46881, n46882,
         n46883, n46884, n46885, n46886, n46887, n46888, n46889, n46890,
         n46891, n46892, n46893, n46894, n46895, n46896, n46897, n46898,
         n46899, n46900, n46901, n46902, n46903, n46904, n46905, n46906,
         n46907, n46908, n46909, n46910, n46911, n46912, n46913, n46914,
         n46915, n46916, n46917, n46918, n46919, n46920, n46921, n46922,
         n46923, n46924, n46925, n46926, n46927, n46928, n46929, n46930,
         n46931, n46932, n46933, n46934, n46935, n46936, n46937, n46938,
         n46939, n46940, n46941, n46942, n46943, n46944, n46945, n46946,
         n46947, n46948, n46949, n46950, n46951, n46952, n46953, n46954,
         n46955, n46956, n46957, n46958, n46959, n46960, n46961, n46962,
         n46963, n46964, n46965, n46966, n46967, n46968, n46969, n46970,
         n46971, n46972, n46973, n46974, n46975, n46976, n46977, n46978,
         n46979, n46980, n46981, n46982, n46983, n46984, n46985, n46986,
         n46987, n46988, n46989, n46990, n46991, n46992, n46993, n46994,
         n46995, n46996, n46997, n46998, n46999, n47000, n47001, n47002,
         n47003, n47004, n47005, n47006, n47007, n47008, n47009, n47010,
         n47011, n47012, n47013, n47014, n47015, n47016, n47017, n47018,
         n47019, n47020, n47021, n47022, n47023, n47024, n47025, n47026,
         n47027, n47028, n47029, n47030, n47031, n47032, n47033, n47034,
         n47035, n47036, n47037, n47038, n47039, n47040, n47041, n47042,
         n47043, n47044, n47045, n47046, n47047, n47048, n47049, n47050,
         n47051, n47052, n47053, n47054, n47055, n47056, n47057, n47058,
         n47059, n47060, n47061, n47062, n47063, n47064, n47065, n47066,
         n47067, n47068, n47069, n47070, n47071, n47072, n47073, n47074,
         n47075, n47076, n47077, n47078, n47079, n47080, n47081, n47082,
         n47083, n47084, n47085, n47086, n47087, n47088, n47089, n47090,
         n47091, n47092, n47093, n47094, n47095, n47096, n47097, n47098,
         n47099, n47100, n47101, n47102, n47103, n47104, n47105, n47106,
         n47107, n47108, n47109, n47110, n47111, n47112, n47113, n47114,
         n47115, n47116, n47117, n47118, n47119, n47120, n47121, n47122,
         n47123, n47124, n47125, n47126, n47127, n47128, n47129, n47130,
         n47131, n47132, n47133, n47134, n47135, n47136, n47137, n47138,
         n47139, n47140, n47141, n47142, n47143, n47144, n47145, n47146,
         n47147, n47148, n47149, n47150, n47151, n47152, n47153, n47154,
         n47155, n47156, n47157, n47158, n47159, n47160, n47161, n47162,
         n47163, n47164, n47165, n47166, n47167, n47168, n47169, n47170,
         n47171, n47172, n47173, n47174, n47175, n47176, n47177, n47178,
         n47179, n47180, n47181, n47182, n47183, n47184, n47185, n47186,
         n47187, n47188, n47189, n47190, n47191, n47192, n47193, n47194,
         n47195, n47196, n47197, n47198, n47199, n47200, n47201, n47202,
         n47203, n47204, n47205, n47206, n47207, n47208, n47209, n47210,
         n47211, n47212, n47213, n47214, n47215, n47216, n47217, n47218,
         n47219, n47220, n47221, n47222, n47223, n47224, n47225, n47226,
         n47227, n47228, n47229, n47230, n47231, n47232, n47233, n47234,
         n47235, n47236, n47237, n47238, n47239, n47240, n47241, n47242,
         n47243, n47244, n47245, n47246, n47247, n47248, n47249, n47250,
         n47251, n47252, n47253, n47254, n47255, n47256, n47257, n47258,
         n47259, n47260, n47261, n47262, n47263, n47264, n47265, n47266,
         n47267, n47268, n47269, n47270, n47271, n47272, n47273, n47274,
         n47275, n47276, n47277, n47278, n47279, n47280, n47281, n47282,
         n47283, n47284, n47285, n47286, n47287, n47288, n47289, n47290,
         n47291, n47292, n47293, n47294, n47295, n47296, n47297, n47298,
         n47299, n47300, n47301, n47302, n47303, n47304, n47305, n47306,
         n47307, n47308, n47309, n47310, n47311, n47312, n47313, n47314,
         n47315, n47316, n47317, n47318, n47319, n47320, n47321, n47322,
         n47323, n47324, n47325, n47326, n47327, n47328, n47329, n47330,
         n47331, n47332, n47333, n47334, n47335, n47336, n47337, n47338,
         n47339, n47340, n47341, n47342, n47343, n47344, n47345, n47346,
         n47347, n47348, n47349, n47350, n47351, n47352, n47353, n47354,
         n47355, n47356, n47357, n47358, n47359, n47360, n47361, n47362,
         n47363, n47364, n47365, n47366, n47367, n47368, n47369, n47370,
         n47371, n47372, n47373, n47374, n47375, n47376, n47377, n47378,
         n47379, n47380, n47381, n47382, n47383, n47384, n47385, n47386,
         n47387, n47388, n47389, n47390, n47391, n47392, n47393, n47394,
         n47395, n47396, n47397, n47398, n47399, n47400, n47401, n47402,
         n47403, n47404, n47405, n47406, n47407, n47408, n47409, n47410,
         n47411, n47412, n47413, n47414, n47415, n47416, n47417, n47418,
         n47419, n47420, n47421, n47422, n47423, n47424, n47425, n47426,
         n47427, n47428, n47429, n47430, n47431, n47432, n47433, n47434,
         n47435, n47436, n47437, n47438, n47439, n47440, n47441, n47442,
         n47443, n47444, n47445, n47446, n47447, n47448, n47449, n47450,
         n47451, n47452, n47453, n47454, n47455, n47456, n47457, n47458,
         n47459, n47460, n47461, n47462, n47463, n47464, n47465, n47466,
         n47467, n47468, n47469, n47470, n47471, n47472, n47473, n47474,
         n47475, n47476, n47477, n47478, n47479, n47480, n47481, n47482,
         n47483, n47484, n47485, n47486, n47487, n47488, n47489, n47490,
         n47491, n47492, n47493, n47494, n47495, n47496, n47497, n47498,
         n47499, n47500, n47501, n47502, n47503, n47504, n47505, n47506,
         n47507, n47508, n47509, n47510, n47511, n47512, n47513, n47514,
         n47515, n47516, n47517, n47518, n47519, n47520, n47521, n47522,
         n47523, n47524, n47525, n47526, n47527, n47528, n47529, n47530,
         n47531, n47532, n47533, n47534, n47535, n47536, n47537, n47538,
         n47539, n47540, n47541, n47542, n47543, n47544, n47545, n47546,
         n47547, n47548, n47549, n47550, n47551, n47552, n47553, n47554,
         n47555, n47556, n47557, n47558, n47559, n47560, n47561, n47562,
         n47563, n47564, n47565, n47566, n47567, n47568, n47569, n47570,
         n47571, n47572, n47573, n47574, n47575, n47576, n47577, n47578,
         n47579, n47580, n47581, n47582, n47583, n47584, n47585, n47586,
         n47587, n47588, n47589, n47590, n47591, n47592, n47593, n47594,
         n47595, n47596, n47597, n47598, n47599, n47600, n47601, n47602,
         n47603, n47604, n47605, n47606, n47607, n47608, n47609, n47610,
         n47611, n47612, n47613, n47614, n47615, n47616, n47617, n47618,
         n47619, n47620, n47621, n47622, n47623, n47624, n47625, n47626,
         n47627, n47628, n47629, n47630, n47631, n47632, n47633, n47634,
         n47635, n47636, n47637, n47638, n47639, n47640, n47641, n47642,
         n47643, n47644, n47645, n47646, n47647, n47648, n47649, n47650,
         n47651, n47652, n47653, n47654, n47655, n47656, n47657, n47658,
         n47659, n47660, n47661, n47662, n47663, n47664, n47665, n47666,
         n47667, n47668, n47669, n47670, n47671, n47672, n47673, n47674,
         n47675, n47676, n47677, n47678, n47679, n47680, n47681, n47682,
         n47683, n47684, n47685, n47686, n47687, n47688, n47689, n47690,
         n47691, n47692, n47693, n47694, n47695, n47696, n47697, n47698,
         n47699, n47700, n47701, n47702, n47703, n47704, n47705, n47706,
         n47707, n47708, n47709, n47710, n47711, n47712, n47713, n47714,
         n47715, n47716, n47717, n47718, n47719, n47720, n47721, n47722,
         n47723, n47724, n47725, n47726, n47727, n47728, n47729, n47730,
         n47731, n47732, n47733, n47734, n47735, n47736, n47737, n47738,
         n47739, n47740, n47741, n47742, n47743, n47744, n47745, n47746,
         n47747, n47748, n47749, n47750, n47751, n47752, n47753, n47754,
         n47755, n47756, n47757, n47758, n47759, n47760, n47761, n47762,
         n47763, n47764, n47765, n47766, n47767, n47768, n47769, n47770,
         n47771, n47772, n47773, n47774, n47775, n47776, n47777, n47778,
         n47779, n47780, n47781, n47782, n47783, n47784, n47785, n47786,
         n47787, n47788, n47789, n47790, n47791, n47792, n47793, n47794,
         n47795, n47796, n47797, n47798, n47799, n47800, n47801, n47802,
         n47803, n47804, n47805, n47806, n47807, n47808, n47809, n47810,
         n47811, n47812, n47813, n47814, n47815, n47816, n47817, n47818,
         n47819, n47820, n47821, n47822, n47823, n47824, n47825, n47826,
         n47827, n47828, n47829, n47830, n47831, n47832, n47833, n47834,
         n47835, n47836, n47837, n47838, n47839, n47840, n47841, n47842,
         n47843, n47844, n47845, n47846, n47847, n47848, n47849, n47850,
         n47851, n47852, n47853, n47854, n47855, n47856, n47857, n47858,
         n47859, n47860, n47861, n47862, n47863, n47864, n47865, n47866,
         n47867, n47868, n47869, n47870, n47871, n47872, n47873, n47874,
         n47875, n47876, n47877, n47878, n47879, n47880, n47881, n47882,
         n47883, n47884, n47885, n47886, n47887, n47888, n47889, n47890,
         n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898,
         n47899, n47900, n47901, n47902, n47903, n47904, n47905, n47906,
         n47907, n47908, n47909, n47910, n47911, n47912, n47913, n47914,
         n47915, n47916, n47917, n47918, n47919, n47920, n47921, n47922,
         n47923, n47924, n47925, n47926, n47927, n47928, n47929, n47930,
         n47931, n47932, n47933, n47934, n47935, n47936, n47937, n47938,
         n47939, n47940, n47941, n47942, n47943, n47944, n47945, n47946,
         n47947, n47948, n47949, n47950, n47951, n47952, n47953, n47954,
         n47955, n47956, n47957, n47958, n47959, n47960, n47961, n47962,
         n47963, n47964, n47965, n47966, n47967, n47968, n47969, n47970,
         n47971, n47972, n47973, n47974, n47975, n47976, n47977, n47978,
         n47979, n47980, n47981, n47982, n47983, n47984, n47985, n47986,
         n47987, n47988, n47989, n47990, n47991, n47992, n47993, n47994,
         n47995, n47996, n47997, n47998, n47999, n48000, n48001, n48002,
         n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010,
         n48011, n48012, n48013, n48014, n48015, n48016, n48017, n48018,
         n48019, n48020, n48021, n48022, n48023, n48024, n48025, n48026,
         n48027, n48028, n48029, n48030, n48031, n48032, n48033, n48034,
         n48035, n48036, n48037, n48038, n48039, n48040, n48041, n48042,
         n48043, n48044, n48045, n48046, n48047, n48048, n48049, n48050,
         n48051, n48052, n48053, n48054, n48055, n48056, n48057, n48058,
         n48059, n48060, n48061, n48062, n48063, n48064, n48065, n48066,
         n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074,
         n48075, n48076, n48077, n48078, n48079, n48080, n48081, n48082,
         n48083, n48084, n48085, n48086, n48087, n48088, n48089, n48090,
         n48091, n48092, n48093, n48094, n48095, n48096, n48097, n48098,
         n48099, n48100, n48101, n48102, n48103, n48104, n48105, n48106,
         n48107, n48108, n48109, n48110, n48111, n48112, n48113, n48114,
         n48115, n48116, n48117, n48118, n48119, n48120, n48121, n48122,
         n48123, n48124, n48125, n48126, n48127, n48128, n48129, n48130,
         n48131, n48132, n48133, n48134, n48135, n48136, n48137, n48138,
         n48139, n48140, n48141, n48142, n48143, n48144, n48145, n48146,
         n48147, n48148, n48149, n48150, n48151, n48152, n48153, n48154,
         n48155, n48156, n48157, n48158, n48159, n48160, n48161, n48162,
         n48163, n48164, n48165, n48166, n48167, n48168, n48169, n48170,
         n48171, n48172, n48173, n48174, n48175, n48176, n48177, n48178,
         n48179, n48180, n48181, n48182, n48183, n48184, n48185, n48186,
         n48187, n48188, n48189, n48190, n48191, n48192, n48193, n48194,
         n48195, n48196, n48197, n48198, n48199, n48200, n48201, n48202,
         n48203, n48204, n48205, n48206, n48207, n48208, n48209, n48210,
         n48211, n48212, n48213, n48214, n48215, n48216, n48217, n48218,
         n48219, n48220, n48221, n48222, n48223, n48224, n48225, n48226,
         n48227, n48228, n48229, n48230, n48231, n48232, n48233, n48234,
         n48235, n48236, n48237, n48238, n48239, n48240, n48241, n48242,
         n48243, n48244, n48245, n48246, n48247, n48248, n48249, n48250,
         n48251, n48252, n48253, n48254, n48255, n48256, n48257, n48258,
         n48259, n48260, n48261, n48262, n48263, n48264, n48265, n48266,
         n48267, n48268, n48269, n48270, n48271, n48272, n48273, n48274,
         n48275, n48276, n48277, n48278, n48279, n48280, n48281, n48282,
         n48283, n48284, n48285, n48286, n48287, n48288, n48289, n48290,
         n48291, n48292, n48293, n48294, n48295, n48296, n48297, n48298,
         n48299, n48300, n48301, n48302, n48303, n48304, n48305, n48306,
         n48307, n48308, n48309, n48310, n48311, n48312, n48313, n48314,
         n48315, n48316, n48317, n48318, n48319, n48320, n48321, n48322,
         n48323, n48324, n48325, n48326, n48327, n48328, n48329, n48330,
         n48331, n48332, n48333, n48334, n48335, n48336, n48337, n48338,
         n48339, n48340, n48341, n48342, n48343, n48344, n48345, n48346,
         n48347, n48348, n48349, n48350, n48351, n48352, n48353, n48354,
         n48355, n48356, n48357, n48358, n48359, n48360, n48361, n48362,
         n48363, n48364, n48365, n48366, n48367, n48368, n48369, n48370,
         n48371, n48372, n48373, n48374, n48375, n48376, n48377, n48378,
         n48379, n48380, n48381, n48382, n48383, n48384, n48385, n48386,
         n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394,
         n48395, n48396, n48397, n48398, n48399, n48400, n48401, n48402,
         n48403, n48404, n48405, n48406, n48407, n48408, n48409, n48410,
         n48411, n48412, n48413, n48414, n48415, n48416, n48417, n48418,
         n48419, n48420, n48421, n48422, n48423, n48424, n48425, n48426,
         n48427, n48428, n48429, n48430, n48431, n48432, n48433, n48434,
         n48435, n48436, n48437, n48438, n48439, n48440, n48441, n48442,
         n48443, n48444, n48445, n48446, n48447, n48448, n48449, n48450,
         n48451, n48452, n48453, n48454, n48455, n48456, n48457, n48458,
         n48459, n48460, n48461, n48462, n48463, n48464, n48465, n48466,
         n48467, n48468, n48469, n48470, n48471, n48472, n48473, n48474,
         n48475, n48476, n48477, n48478, n48479, n48480, n48481, n48482,
         n48483, n48484, n48485, n48486, n48487, n48488, n48489, n48490,
         n48491, n48492, n48493, n48494, n48495, n48496, n48497, n48498,
         n48499, n48500, n48501, n48502, n48503, n48504, n48505, n48506,
         n48507, n48508, n48509, n48510, n48511, n48512, n48513, n48514,
         n48515, n48516, n48517, n48518, n48519, n48520, n48521, n48522,
         n48523, n48524, n48525, n48526, n48527, n48528, n48529, n48530,
         n48531, n48532, n48533, n48534, n48535, n48536, n48537, n48538,
         n48539, n48540, n48541, n48542, n48543, n48544, n48545, n48546,
         n48547, n48548, n48549, n48550, n48551, n48552, n48553, n48554,
         n48555, n48556, n48557, n48558, n48559, n48560, n48561, n48562,
         n48563, n48564, n48565, n48566, n48567, n48568, n48569, n48570,
         n48571, n48572, n48573, n48574, n48575, n48576, n48577, n48578,
         n48579, n48580, n48581, n48582, n48583, n48584, n48585, n48586,
         n48587, n48588, n48589, n48590, n48591, n48592, n48593, n48594,
         n48595, n48596, n48597, n48598, n48599, n48600, n48601, n48602,
         n48603, n48604, n48605, n48606, n48607, n48608, n48609, n48610,
         n48611, n48612, n48613, n48614, n48615, n48616, n48617, n48618,
         n48619, n48620, n48621, n48622, n48623, n48624, n48625, n48626,
         n48627, n48628, n48629, n48630, n48631, n48632, n48633, n48634,
         n48635, n48636, n48637, n48638, n48639, n48640, n48641, n48642,
         n48643, n48644, n48645, n48646, n48647, n48648, n48649, n48650,
         n48651, n48652, n48653, n48654, n48655, n48656, n48657, n48658,
         n48659, n48660, n48661, n48662, n48663, n48664, n48665, n48666,
         n48667, n48668, n48669, n48670, n48671, n48672, n48673, n48674,
         n48675, n48676, n48677, n48678, n48679, n48680, n48681, n48682,
         n48683, n48684, n48685, n48686, n48687, n48688, n48689, n48690,
         n48691, n48692, n48693, n48694, n48695, n48696, n48697, n48698,
         n48699, n48700, n48701, n48702, n48703, n48704, n48705, n48706,
         n48707, n48708, n48709, n48710, n48711, n48712, n48713, n48714,
         n48715, n48716, n48717, n48718, n48719, n48720, n48721, n48722,
         n48723, n48724, n48725, n48726, n48727, n48728, n48729, n48730,
         n48731, n48732, n48733, n48734, n48735, n48736, n48737, n48738,
         n48739, n48740, n48741, n48742, n48743, n48744, n48745, n48746,
         n48747, n48748, n48749, n48750, n48751, n48752, n48753, n48754,
         n48755, n48756, n48757, n48758, n48759, n48760, n48761, n48762,
         n48763, n48764, n48765, n48766, n48767, n48768, n48769, n48770,
         n48771, n48772, n48773, n48774, n48775, n48776, n48777, n48778,
         n48779, n48780, n48781, n48782, n48783, n48784, n48785, n48786,
         n48787, n48788, n48789, n48790, n48791, n48792, n48793, n48794,
         n48795, n48796, n48797, n48798, n48799, n48800, n48801, n48802,
         n48803, n48804, n48805, n48806, n48807, n48808, n48809, n48810,
         n48811, n48812, n48813, n48814, n48815, n48816, n48817, n48818,
         n48819, n48820, n48821, n48822, n48823, n48824, n48825, n48826,
         n48827, n48828, n48829, n48830, n48831, n48832, n48833, n48834,
         n48835, n48836, n48837, n48838, n48839, n48840, n48841, n48842,
         n48843, n48844, n48845, n48846, n48847, n48848, n48849, n48850,
         n48851, n48852, n48853, n48854, n48855, n48856, n48857, n48858,
         n48859, n48860, n48861, n48862, n48863, n48864, n48865, n48866,
         n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874,
         n48875, n48876, n48877, n48878, n48879, n48880, n48881, n48882,
         n48883, n48884, n48885, n48886, n48887, n48888, n48889, n48890,
         n48891, n48892, n48893, n48894, n48895, n48896, n48897, n48898,
         n48899, n48900, n48901, n48902, n48903, n48904, n48905, n48906,
         n48907, n48908, n48909, n48910, n48911, n48912, n48913, n48914,
         n48915, n48916, n48917, n48918, n48919, n48920, n48921, n48922,
         n48923, n48924, n48925, n48926, n48927, n48928, n48929, n48930,
         n48931, n48932, n48933, n48934, n48935, n48936, n48937, n48938,
         n48939, n48940, n48941, n48942, n48943, n48944, n48945, n48946,
         n48947, n48948, n48949, n48950, n48951, n48952, n48953, n48954,
         n48955, n48956, n48957, n48958, n48959, n48960, n48961, n48962,
         n48963, n48964, n48965, n48966, n48967, n48968, n48969, n48970,
         n48971, n48972, n48973, n48974, n48975, n48976, n48977, n48978,
         n48979, n48980, n48981, n48982, n48983, n48984, n48985, n48986,
         n48987, n48988, n48989, n48990, n48991, n48992, n48993, n48994,
         n48995, n48996, n48997, n48998, n48999, n49000, n49001, n49002,
         n49003, n49004, n49005, n49006, n49007, n49008, n49009, n49010,
         n49011, n49012, n49013, n49014, n49015, n49016, n49017, n49018,
         n49019, n49020, n49021, n49022, n49023, n49024, n49025, n49026,
         n49027, n49028, n49029, n49030, n49031, n49032, n49033, n49034,
         n49035, n49036, n49037, n49038, n49039, n49040, n49041, n49042,
         n49043, n49044, n49045, n49046, n49047, n49048, n49049, n49050,
         n49051, n49052, n49053, n49054, n49055, n49056, n49057, n49058,
         n49059, n49060, n49061, n49062, n49063, n49064, n49065, n49066,
         n49067, n49068, n49069, n49070, n49071, n49072, n49073, n49074,
         n49075, n49076, n49077, n49078, n49079, n49080, n49081, n49082,
         n49083, n49084, n49085, n49086, n49087, n49088, n49089, n49090,
         n49091, n49092, n49093, n49094, n49095, n49096, n49097, n49098,
         n49099, n49100, n49101, n49102, n49103, n49104, n49105, n49106,
         n49107, n49108, n49109, n49110, n49111, n49112, n49113, n49114,
         n49115, n49116, n49117, n49118, n49119, n49120, n49121, n49122,
         n49123, n49124, n49125, n49126, n49127, n49128, n49129, n49130,
         n49131, n49132, n49133, n49134, n49135, n49136, n49137, n49138,
         n49139, n49140, n49141, n49142, n49143, n49144, n49145, n49146,
         n49147, n49148, n49149, n49150, n49151, n49152, n49153, n49154,
         n49155, n49156, n49157, n49158, n49159, n49160, n49161, n49162,
         n49163, n49164, n49165, n49166, n49167, n49168, n49169, n49170,
         n49171, n49172, n49173, n49174, n49175, n49176, n49177, n49178,
         n49179, n49180, n49181, n49182, n49183, n49184, n49185, n49186,
         n49187, n49188, n49189, n49190, n49191, n49192, n49193, n49194,
         n49195, n49196, n49197, n49198, n49199, n49200, n49201, n49202,
         n49203, n49204, n49205, n49206, n49207, n49208, n49209, n49210,
         n49211, n49212, n49213, n49214, n49215, n49216, n49217, n49218,
         n49219, n49220, n49221, n49222, n49223, n49224, n49225, n49226,
         n49227, n49228, n49229, n49230, n49231, n49232, n49233, n49234,
         n49235, n49236, n49237, n49238, n49239, n49240, n49241, n49242,
         n49243, n49244, n49245, n49246, n49247, n49248, n49249, n49250,
         n49251, n49252, n49253, n49254, n49255, n49256, n49257, n49258,
         n49259, n49260, n49261, n49262, n49263, n49264, n49265, n49266,
         n49267, n49268, n49269, n49270, n49271, n49272, n49273, n49274,
         n49275, n49276, n49277, n49278, n49279, n49280, n49281, n49282,
         n49283, n49284, n49285, n49286, n49287, n49288, n49289, n49290,
         n49291, n49292, n49293, n49294, n49295, n49296, n49297, n49298,
         n49299, n49300, n49301, n49302, n49303, n49304, n49305, n49306,
         n49307, n49308, n49309, n49310, n49311, n49312, n49313, n49314,
         n49315, n49316, n49317, n49318, n49319, n49320, n49321, n49322,
         n49323, n49324, n49325, n49326, n49327, n49328, n49329, n49330,
         n49331, n49332, n49333, n49334, n49335, n49336, n49337, n49338,
         n49339, n49340, n49341, n49342, n49343, n49344, n49345, n49346,
         n49347, n49348, n49349, n49350, n49351, n49352, n49353, n49354,
         n49355, n49356, n49357, n49358, n49359, n49360, n49361, n49362,
         n49363, n49364, n49365, n49366, n49367, n49368, n49369, n49370,
         n49371, n49372, n49373, n49374, n49375, n49376, n49377, n49378,
         n49379, n49380, n49381, n49382, n49383, n49384, n49385, n49386,
         n49387, n49388, n49389, n49390, n49391, n49392, n49393, n49394,
         n49395, n49396, n49397, n49398, n49399, n49400, n49401, n49402,
         n49403, n49404, n49405, n49406, n49407, n49408, n49409, n49410,
         n49411, n49412, n49413, n49414, n49415, n49416, n49417, n49418,
         n49419, n49420, n49421, n49422, n49423, n49424, n49425, n49426,
         n49427, n49428, n49429, n49430, n49431, n49432, n49433, n49434,
         n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442,
         n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450,
         n49451, n49452, n49453, n49454, n49455, n49456, n49457, n49458,
         n49459, n49460, n49461, n49462, n49463, n49464, n49465, n49466,
         n49467, n49468, n49469, n49470, n49471, n49472, n49473, n49474,
         n49475, n49476, n49477, n49478, n49479, n49480, n49481, n49482,
         n49483, n49484, n49485, n49486, n49487, n49488, n49489, n49490,
         n49491, n49492, n49493, n49494, n49495, n49496, n49497, n49498,
         n49499, n49500, n49501, n49502, n49503, n49504, n49505, n49506,
         n49507, n49508, n49509, n49510, n49511, n49512, n49513, n49514,
         n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522,
         n49523, n49524, n49525, n49526, n49527, n49528, n49529, n49530,
         n49531, n49532, n49533, n49534, n49535, n49536, n49537, n49538,
         n49539, n49540, n49541, n49542, n49543, n49544, n49545, n49546,
         n49547, n49548, n49549, n49550, n49551, n49552, n49553, n49554,
         n49555, n49556, n49557, n49558, n49559, n49560, n49561, n49562,
         n49563, n49564, n49565, n49566, n49567, n49568, n49569, n49570,
         n49571, n49572, n49573, n49574, n49575, n49576, n49577, n49578,
         n49579, n49580, n49581, n49582, n49583, n49584, n49585, n49586,
         n49587, n49588, n49589, n49590, n49591, n49592, n49593, n49594,
         n49595, n49596, n49597, n49598, n49599, n49600, n49601, n49602,
         n49603, n49604, n49605, n49606, n49607, n49608, n49609, n49610,
         n49611, n49612, n49613, n49614, n49615, n49616, n49617, n49618,
         n49619, n49620, n49621, n49622, n49623, n49624, n49625, n49626,
         n49627, n49628, n49629, n49630, n49631, n49632, n49633, n49634,
         n49635, n49636, n49637, n49638, n49639, n49640, n49641, n49642,
         n49643, n49644, n49645, n49646, n49647, n49648, n49649, n49650,
         n49651, n49652, n49653, n49654, n49655, n49656, n49657, n49658,
         n49659, n49660, n49661, n49662, n49663, n49664, n49665, n49666,
         n49667, n49668, n49669, n49670, n49671, n49672, n49673, n49674,
         n49675, n49676, n49677, n49678, n49679, n49680, n49681, n49682,
         n49683, n49684, n49685, n49686, n49687, n49688, n49689, n49690,
         n49691, n49692, n49693, n49694, n49695, n49696, n49697, n49698,
         n49699, n49700, n49701, n49702, n49703, n49704, n49705, n49706,
         n49707, n49708, n49709, n49710, n49711, n49712, n49713, n49714,
         n49715, n49716, n49717, n49718, n49719, n49720, n49721, n49722,
         n49723, n49724, n49725, n49726, n49727, n49728, n49729, n49730,
         n49731, n49732, n49733, n49734, n49735, n49736, n49737, n49738,
         n49739, n49740, n49741, n49742, n49743, n49744, n49745, n49746,
         n49747, n49748, n49749, n49750, n49751, n49752, n49753, n49754,
         n49755, n49756, n49757, n49758, n49759, n49760, n49761, n49762,
         n49763, n49764, n49765, n49766, n49767, n49768, n49769, n49770,
         n49771, n49772, n49773, n49774, n49775, n49776, n49777, n49778,
         n49779, n49780, n49781, n49782, n49783, n49784, n49785, n49786,
         n49787, n49788, n49789, n49790, n49791, n49792, n49793, n49794,
         n49795, n49796, n49797, n49798, n49799, n49800, n49801, n49802,
         n49803, n49804, n49805, n49806, n49807, n49808, n49809, n49810,
         n49811, n49812, n49813, n49814, n49815, n49816, n49817, n49818,
         n49819, n49820, n49821, n49822, n49823, n49824, n49825, n49826,
         n49827, n49828, n49829, n49830, n49831, n49832, n49833, n49834,
         n49835, n49836, n49837, n49838, n49839, n49840, n49841, n49842,
         n49843, n49844, n49845, n49846, n49847, n49848, n49849, n49850,
         n49851, n49852, n49853, n49854, n49855, n49856, n49857, n49858,
         n49859, n49860, n49861, n49862, n49863, n49864, n49865, n49866,
         n49867, n49868, n49869, n49870, n49871, n49872, n49873, n49874,
         n49875, n49876, n49877, n49878, n49879, n49880, n49881, n49882,
         n49883, n49884, n49885, n49886, n49887, n49888, n49889, n49890,
         n49891, n49892, n49893, n49894, n49895, n49896, n49897, n49898,
         n49899, n49900, n49901, n49902, n49903, n49904, n49905, n49906,
         n49907, n49908, n49909, n49910, n49911, n49912, n49913, n49914,
         n49915, n49916, n49917, n49918, n49919, n49920, n49921, n49922,
         n49923, n49924, n49925, n49926, n49927, n49928, n49929, n49930,
         n49931, n49932, n49933, n49934, n49935, n49936, n49937, n49938,
         n49939, n49940, n49941, n49942, n49943, n49944, n49945, n49946,
         n49947, n49948, n49949, n49950, n49951, n49952, n49953, n49954,
         n49955, n49956, n49957, n49958, n49959, n49960, n49961, n49962,
         n49963, n49964, n49965, n49966, n49967, n49968, n49969, n49970,
         n49971, n49972, n49973, n49974, n49975, n49976, n49977, n49978,
         n49979, n49980, n49981, n49982, n49983, n49984, n49985, n49986,
         n49987, n49988, n49989, n49990, n49991, n49992, n49993, n49994,
         n49995, n49996, n49997, n49998, n49999, n50000, n50001, n50002,
         n50003, n50004, n50005, n50006, n50007, n50008, n50009, n50010,
         n50011, n50012, n50013, n50014, n50015, n50016, n50017, n50018,
         n50019, n50020, n50021, n50022, n50023, n50024, n50025, n50026,
         n50027, n50028, n50029, n50030, n50031, n50032, n50033, n50034,
         n50035, n50036, n50037, n50038, n50039, n50040, n50041, n50042,
         n50043, n50044, n50045, n50046, n50047, n50048, n50049, n50050,
         n50051, n50052, n50053, n50054, n50055, n50056, n50057, n50058,
         n50059, n50060, n50061, n50062, n50063, n50064, n50065, n50066,
         n50067, n50068, n50069, n50070, n50071, n50072, n50073, n50074,
         n50075, n50076, n50077, n50078, n50079, n50080, n50081, n50082,
         n50083, n50084, n50085, n50086, n50087, n50088, n50089, n50090,
         n50091, n50092, n50093, n50094, n50095, n50096, n50097, n50098,
         n50099, n50100, n50101, n50102, n50103, n50104, n50105, n50106,
         n50107, n50108, n50109, n50110, n50111, n50112, n50113, n50114,
         n50115, n50116, n50117, n50118, n50119, n50120, n50121, n50122,
         n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130,
         n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138,
         n50139, n50140, n50141, n50142, n50143, n50144, n50145, n50146,
         n50147, n50148, n50149, n50150, n50151, n50152, n50153, n50154,
         n50155, n50156, n50157, n50158, n50159, n50160, n50161, n50162,
         n50163, n50164, n50165, n50166, n50167, n50168, n50169, n50170,
         n50171, n50172, n50173, n50174, n50175, n50176, n50177, n50178,
         n50179, n50180, n50181, n50182, n50183, n50184, n50185, n50186,
         n50187, n50188, n50189, n50190, n50191, n50192, n50193, n50194,
         n50195, n50196, n50197, n50198, n50199, n50200, n50201, n50202,
         n50203, n50204, n50205, n50206, n50207, n50208, n50209, n50210,
         n50211, n50212, n50213, n50214, n50215, n50216, n50217, n50218,
         n50219, n50220, n50221, n50222, n50223, n50224, n50225, n50226,
         n50227, n50228, n50229, n50230, n50231, n50232, n50233, n50234,
         n50235, n50236, n50237, n50238, n50239, n50240, n50241, n50242,
         n50243, n50244, n50245, n50246, n50247, n50248, n50249, n50250,
         n50251, n50252, n50253, n50254, n50255, n50256, n50257, n50258,
         n50259, n50260, n50261, n50262, n50263, n50264, n50265, n50266,
         n50267, n50268, n50269, n50270, n50271, n50272, n50273, n50274,
         n50275, n50276, n50277, n50278, n50279, n50280, n50281, n50282,
         n50283, n50284, n50285, n50286, n50287, n50288, n50289, n50290,
         n50291, n50292, n50293, n50294, n50295, n50296, n50297, n50298,
         n50299, n50300, n50301, n50302, n50303, n50304, n50305, n50306,
         n50307, n50308, n50309, n50310, n50311, n50312, n50313, n50314,
         n50315, n50316, n50317, n50318, n50319, n50320, n50321, n50322,
         n50323, n50324, n50325, n50326, n50327, n50328, n50329, n50330,
         n50331, n50332, n50333, n50334, n50335, n50336, n50337, n50338,
         n50339, n50340, n50341, n50342, n50343, n50344, n50345, n50346,
         n50347, n50348, n50349, n50350, n50351, n50352, n50353, n50354,
         n50355, n50356, n50357, n50358, n50359, n50360, n50361, n50362,
         n50363, n50364, n50365, n50366, n50367, n50368, n50369, n50370,
         n50371, n50372, n50373, n50374, n50375, n50376, n50377, n50378,
         n50379, n50380, n50381, n50382, n50383, n50384, n50385, n50386,
         n50387, n50388, n50389, n50390, n50391, n50392, n50393, n50394,
         n50395, n50396, n50397, n50398, n50399, n50400, n50401, n50402,
         n50403, n50404, n50405, n50406, n50407, n50408, n50409, n50410,
         n50411, n50412, n50413, n50414, n50415, n50416, n50417, n50418,
         n50419, n50420, n50421, n50422, n50423, n50424, n50425, n50426,
         n50427, n50428, n50429, n50430, n50431, n50432, n50433, n50434,
         n50435, n50436, n50437, n50438, n50439, n50440, n50441, n50442,
         n50443, n50444, n50445, n50446, n50447, n50448, n50449, n50450,
         n50451, n50452, n50453, n50454, n50455, n50456, n50457, n50458,
         n50459, n50460, n50461, n50462, n50463, n50464, n50465, n50466,
         n50467, n50468, n50469, n50470, n50471, n50472, n50473, n50474,
         n50475, n50476, n50477, n50478, n50479, n50480, n50481, n50482,
         n50483, n50484, n50485, n50486, n50487, n50488, n50489, n50490,
         n50491, n50492, n50493, n50494, n50495, n50496, n50497, n50498,
         n50499, n50500, n50501, n50502, n50503, n50504, n50505, n50506,
         n50507, n50508, n50509, n50510, n50511, n50512, n50513, n50514,
         n50515, n50516, n50517, n50518, n50519, n50520, n50521, n50522,
         n50523, n50524, n50525, n50526, n50527, n50528, n50529, n50530,
         n50531, n50532, n50533, n50534, n50535, n50536, n50537, n50538,
         n50539, n50540, n50541, n50542, n50543, n50544, n50545, n50546,
         n50547, n50548, n50549, n50550, n50551, n50552, n50553, n50554,
         n50555, n50556, n50557, n50558, n50559, n50560, n50561, n50562,
         n50563, n50564, n50565, n50566, n50567, n50568, n50569, n50570,
         n50571, n50572, n50573, n50574, n50575, n50576, n50577, n50578,
         n50579, n50580, n50581, n50582, n50583, n50584, n50585, n50586,
         n50587, n50588, n50589, n50590, n50591, n50592, n50593, n50594,
         n50595, n50596, n50597, n50598, n50599, n50600, n50601, n50602,
         n50603, n50604, n50605, n50606, n50607, n50608, n50609, n50610,
         n50611, n50612, n50613, n50614, n50615, n50616, n50617, n50618,
         n50619, n50620, n50621, n50622, n50623, n50624, n50625, n50626,
         n50627, n50628, n50629, n50630, n50631, n50632, n50633, n50634,
         n50635, n50636, n50637, n50638, n50639, n50640, n50641, n50642,
         n50643, n50644, n50645, n50646, n50647, n50648, n50649, n50650,
         n50651, n50652, n50653, n50654, n50655, n50656, n50657, n50658,
         n50659, n50660, n50661, n50662, n50663, n50664, n50665, n50666,
         n50667, n50668, n50669, n50670, n50671, n50672, n50673, n50674,
         n50675, n50676, n50677, n50678, n50679, n50680, n50681, n50682,
         n50683, n50684, n50685, n50686, n50687, n50688, n50689, n50690,
         n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50698,
         n50699, n50700, n50701, n50702, n50703, n50704, n50705, n50706,
         n50707, n50708, n50709, n50710, n50711, n50712, n50713, n50714,
         n50715, n50716, n50717, n50718, n50719, n50720, n50721, n50722,
         n50723, n50724, n50725, n50726, n50727, n50728, n50729, n50730,
         n50731, n50732, n50733, n50734, n50735, n50736, n50737, n50738,
         n50739, n50740, n50741, n50742, n50743, n50744, n50745, n50746,
         n50747, n50748, n50749, n50750, n50751, n50752, n50753, n50754,
         n50755, n50756, n50757, n50758, n50759, n50760, n50761, n50762,
         n50763, n50764, n50765, n50766, n50767, n50768, n50769, n50770,
         n50771, n50772, n50773, n50774, n50775, n50776, n50777, n50778,
         n50779, n50780, n50781, n50782, n50783, n50784, n50785, n50786,
         n50787, n50788, n50789, n50790, n50791, n50792, n50793, n50794,
         n50795, n50796, n50797, n50798, n50799, n50800, n50801, n50802,
         n50803, n50804, n50805, n50806, n50807, n50808, n50809, n50810,
         n50811, n50812, n50813, n50814, n50815, n50816, n50817, n50818,
         n50819, n50820, n50821, n50822, n50823, n50824, n50825, n50826,
         n50827, n50828, n50829, n50830, n50831, n50832, n50833, n50834,
         n50835, n50836, n50837, n50838, n50839, n50840, n50841, n50842,
         n50843, n50844, n50845, n50846, n50847, n50848, n50849, n50850,
         n50851, n50852, n50853, n50854, n50855, n50856, n50857, n50858,
         n50859, n50860, n50861, n50862, n50863, n50864, n50865, n50866,
         n50867, n50868, n50869, n50870, n50871, n50872, n50873, n50874,
         n50875, n50876, n50877, n50878, n50879, n50880, n50881, n50882,
         n50883, n50884, n50885, n50886, n50887, n50888, n50889, n50890,
         n50891, n50892, n50893, n50894, n50895, n50896, n50897, n50898,
         n50899, n50900, n50901, n50902, n50903, n50904, n50905, n50906,
         n50907, n50908, n50909, n50910, n50911, n50912, n50913, n50914,
         n50915, n50916, n50917, n50918, n50919, n50920, n50921, n50922,
         n50923, n50924, n50925, n50926, n50927, n50928, n50929, n50930,
         n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938,
         n50939, n50940, n50941, n50942, n50943, n50944, n50945, n50946,
         n50947, n50948, n50949, n50950, n50951, n50952, n50953, n50954,
         n50955, n50956, n50957, n50958, n50959, n50960, n50961, n50962,
         n50963, n50964, n50965, n50966, n50967, n50968, n50969, n50970,
         n50971, n50972, n50973, n50974, n50975, n50976, n50977, n50978,
         n50979, n50980, n50981, n50982, n50983, n50984, n50985, n50986,
         n50987, n50988, n50989, n50990, n50991, n50992, n50993, n50994,
         n50995, n50996, n50997, n50998, n50999, n51000, n51001, n51002,
         n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010,
         n51011, n51012, n51013, n51014, n51015, n51016, n51017, n51018,
         n51019, n51020, n51021, n51022, n51023, n51024, n51025, n51026,
         n51027, n51028, n51029, n51030, n51031, n51032, n51033, n51034,
         n51035, n51036, n51037, n51038, n51039, n51040, n51041, n51042,
         n51043, n51044, n51045, n51046, n51047, n51048, n51049, n51050,
         n51051, n51052, n51053, n51054, n51055, n51056, n51057, n51058,
         n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066,
         n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074,
         n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082,
         n51083, n51084, n51085, n51086, n51087, n51088, n51089, n51090,
         n51091, n51092, n51093, n51094, n51095, n51096, n51097, n51098,
         n51099, n51100, n51101, n51102, n51103, n51104, n51105, n51106,
         n51107, n51108, n51109, n51110, n51111, n51112, n51113, n51114,
         n51115, n51116, n51117, n51118, n51119, n51120, n51121, n51122,
         n51123, n51124, n51125, n51126, n51127, n51128, n51129, n51130,
         n51131, n51132, n51133, n51134, n51135, n51136, n51137, n51138,
         n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146,
         n51147, n51148, n51149, n51150, n51151, n51152, n51153, n51154,
         n51155, n51156, n51157, n51158, n51159, n51160, n51161, n51162,
         n51163, n51164, n51165, n51166, n51167, n51168, n51169, n51170,
         n51171, n51172, n51173, n51174, n51175, n51176, n51177, n51178,
         n51179, n51180, n51181, n51182, n51183, n51184, n51185, n51186,
         n51187, n51188, n51189, n51190, n51191, n51192, n51193, n51194,
         n51195, n51196, n51197, n51198, n51199, n51200, n51201, n51202,
         n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210,
         n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218,
         n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226,
         n51227, n51228, n51229, n51230, n51231, n51232, n51233, n51234,
         n51235, n51236, n51237, n51238, n51239, n51240, n51241, n51242,
         n51243, n51244, n51245, n51246, n51247, n51248, n51249, n51250,
         n51251, n51252, n51253, n51254, n51255, n51256, n51257, n51258,
         n51259, n51260, n51261, n51262, n51263, n51264, n51265, n51266,
         n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274,
         n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282,
         n51283, n51284, n51285, n51286, n51287, n51288, n51289, n51290,
         n51291, n51292, n51293, n51294, n51295, n51296, n51297, n51298,
         n51299, n51300, n51301, n51302, n51303, n51304, n51305, n51306,
         n51307, n51308, n51309, n51310, n51311, n51312, n51313, n51314,
         n51315, n51316, n51317, n51318, n51319, n51320, n51321, n51322,
         n51323, n51324, n51325, n51326, n51327, n51328, n51329, n51330,
         n51331, n51332, n51333, n51334, n51335, n51336, n51337, n51338,
         n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346,
         n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354,
         n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362,
         n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370,
         n51371, n51372, n51373, n51374, n51375, n51376, n51377, n51378,
         n51379, n51380, n51381, n51382, n51383, n51384, n51385, n51386,
         n51387, n51388, n51389, n51390, n51391, n51392, n51393, n51394,
         n51395, n51396, n51397, n51398, n51399, n51400, n51401, n51402,
         n51403, n51404, n51405, n51406, n51407, n51408, n51409, n51410,
         n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418,
         n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426,
         n51427, n51428, n51429, n51430, n51431, n51432, n51433, n51434,
         n51435, n51436, n51437, n51438, n51439, n51440, n51441, n51442,
         n51443, n51444, n51445, n51446, n51447, n51448, n51449, n51450,
         n51451, n51452, n51453, n51454, n51455, n51456, n51457, n51458,
         n51459, n51460, n51461, n51462, n51463, n51464, n51465, n51466,
         n51467, n51468, n51469, n51470, n51471, n51472, n51473, n51474,
         n51475, n51476, n51477, n51478, n51479, n51480, n51481, n51482,
         n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490,
         n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498,
         n51499, n51500, n51501, n51502, n51503, n51504, n51505, n51506,
         n51507, n51508, n51509, n51510, n51511, n51512, n51513, n51514,
         n51515, n51516, n51517, n51518, n51519, n51520, n51521, n51522,
         n51523, n51524, n51525, n51526, n51527, n51528, n51529, n51530,
         n51531, n51532, n51533, n51534, n51535, n51536, n51537, n51538,
         n51539, n51540, n51541, n51542, n51543, n51544, n51545, n51546,
         n51547, n51548, n51549, n51550, n51551, n51552, n51553, n51554,
         n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562,
         n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51570,
         n51571, n51572, n51573, n51574, n51575, n51576, n51577, n51578,
         n51579, n51580, n51581, n51582, n51583, n51584, n51585, n51586,
         n51587, n51588, n51589, n51590, n51591, n51592, n51593, n51594,
         n51595, n51596, n51597, n51598, n51599, n51600, n51601, n51602,
         n51603, n51604, n51605, n51606, n51607, n51608, n51609, n51610,
         n51611, n51612, n51613, n51614, n51615, n51616, n51617, n51618,
         n51619, n51620, n51621, n51622, n51623, n51624, n51625, n51626,
         n51627, n51628, n51629, n51630, n51631, n51632, n51633, n51634,
         n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642,
         n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650,
         n51651, n51652, n51653, n51654, n51655, n51656, n51657, n51658,
         n51659, n51660, n51661, n51662, n51663, n51664, n51665, n51666,
         n51667, n51668, n51669, n51670, n51671, n51672, n51673, n51674,
         n51675, n51676, n51677, n51678, n51679, n51680, n51681, n51682,
         n51683, n51684, n51685, n51686, n51687, n51688, n51689, n51690,
         n51691, n51692, n51693, n51694, n51695, n51696, n51697, n51698,
         n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706,
         n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714,
         n51715, n51716, n51717, n51718, n51719, n51720, n51721, n51722,
         n51723, n51724, n51725, n51726, n51727, n51728, n51729, n51730,
         n51731, n51732, n51733, n51734, n51735, n51736, n51737, n51738,
         n51739, n51740, n51741, n51742, n51743, n51744, n51745, n51746,
         n51747, n51748, n51749, n51750, n51751, n51752, n51753, n51754,
         n51755, n51756, n51757, n51758, n51759, n51760, n51761, n51762,
         n51763, n51764, n51765, n51766, n51767, n51768, n51769, n51770,
         n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778,
         n51779, n51780, n51781, n51782, n51783, n51784, n51785, n51786,
         n51787, n51788, n51789, n51790, n51791, n51792, n51793, n51794,
         n51795, n51796, n51797, n51798, n51799, n51800, n51801, n51802,
         n51803, n51804, n51805, n51806, n51807, n51808, n51809, n51810,
         n51811, n51812, n51813, n51814, n51815, n51816, n51817, n51818,
         n51819, n51820, n51821, n51822, n51823, n51824, n51825, n51826,
         n51827, n51828, n51829, n51830, n51831, n51832, n51833, n51834,
         n51835, n51836, n51837, n51838, n51839, n51840, n51841, n51842,
         n51843, n51844, n51845, n51846, n51847, n51848, n51849, n51850,
         n51851, n51852, n51853, n51854, n51855, n51856, n51857, n51858,
         n51859, n51860, n51861, n51862, n51863, n51864, n51865, n51866,
         n51867, n51868, n51869, n51870, n51871, n51872, n51873, n51874,
         n51875, n51876, n51877, n51878, n51879, n51880, n51881, n51882,
         n51883, n51884, n51885, n51886, n51887, n51888, n51889, n51890,
         n51891, n51892, n51893, n51894, n51895, n51896, n51897, n51898,
         n51899, n51900, n51901, n51902, n51903, n51904, n51905, n51906,
         n51907, n51908, n51909, n51910, n51911, n51912, n51913, n51914,
         n51915, n51916, n51917, n51918, n51919, n51920, n51921, n51922,
         n51923, n51924, n51925, n51926, n51927, n51928, n51929, n51930,
         n51931, n51932, n51933, n51934, n51935, n51936, n51937, n51938,
         n51939, n51940, n51941, n51942, n51943, n51944, n51945, n51946,
         n51947, n51948, n51949, n51950, n51951, n51952, n51953, n51954,
         n51955, n51956, n51957, n51958, n51959, n51960, n51961, n51962,
         n51963, n51964, n51965, n51966, n51967, n51968, n51969, n51970,
         n51971, n51972, n51973, n51974, n51975, n51976, n51977, n51978,
         n51979, n51980, n51981, n51982, n51983, n51984, n51985, n51986,
         n51987, n51988, n51989, n51990, n51991, n51992, n51993, n51994,
         n51995, n51996, n51997, n51998, n51999, n52000, n52001, n52002,
         n52003, n52004, n52005, n52006, n52007, n52008, n52009, n52010,
         n52011, n52012, n52013, n52014, n52015, n52016, n52017, n52018,
         n52019, n52020, n52021, n52022, n52023, n52024, n52025, n52026,
         n52027, n52028, n52029, n52030, n52031, n52032, n52033, n52034,
         n52035, n52036, n52037, n52038, n52039, n52040, n52041, n52042,
         n52043, n52044, n52045, n52046, n52047, n52048, n52049, n52050,
         n52051, n52052, n52053, n52054, n52055, n52056, n52057, n52058,
         n52059, n52060, n52061, n52062, n52063, n52064, n52065, n52066,
         n52067, n52068, n52069, n52070, n52071, n52072, n52073, n52074,
         n52075, n52076, n52077, n52078, n52079, n52080, n52081, n52082,
         n52083, n52084, n52085, n52086, n52087, n52088, n52089, n52090,
         n52091, n52092, n52093, n52094, n52095, n52096, n52097, n52098,
         n52099, n52100, n52101, n52102, n52103, n52104, n52105, n52106,
         n52107, n52108, n52109, n52110, n52111, n52112, n52113, n52114,
         n52115, n52116, n52117, n52118, n52119, n52120, n52121, n52122,
         n52123, n52124, n52125, n52126, n52127, n52128, n52129, n52130,
         n52131, n52132, n52133, n52134, n52135, n52136, n52137, n52138,
         n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146,
         n52147, n52148, n52149, n52150, n52151, n52152, n52153, n52154,
         n52155, n52156, n52157, n52158, n52159, n52160, n52161, n52162,
         n52163, n52164, n52165, n52166, n52167, n52168, n52169, n52170,
         n52171, n52172, n52173, n52174, n52175, n52176, n52177, n52178,
         n52179, n52180, n52181, n52182, n52183, n52184, n52185, n52186,
         n52187, n52188, n52189, n52190, n52191, n52192, n52193, n52194,
         n52195, n52196, n52197, n52198, n52199, n52200, n52201, n52202,
         n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210,
         n52211, n52212, n52213, n52214, n52215, n52216, n52217, n52218,
         n52219, n52220, n52221, n52222, n52223, n52224, n52225, n52226,
         n52227, n52228, n52229, n52230, n52231, n52232, n52233, n52234,
         n52235, n52236, n52237, n52238, n52239, n52240, n52241, n52242,
         n52243, n52244, n52245, n52246, n52247, n52248, n52249, n52250,
         n52251, n52252, n52253, n52254, n52255, n52256, n52257, n52258,
         n52259, n52260, n52261, n52262, n52263, n52264, n52265, n52266,
         n52267, n52268, n52269, n52270, n52271, n52272, n52273, n52274,
         n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282,
         n52283, n52284, n52285, n52286, n52287, n52288, n52289, n52290,
         n52291, n52292, n52293, n52294, n52295, n52296, n52297, n52298,
         n52299, n52300, n52301, n52302, n52303, n52304, n52305, n52306,
         n52307, n52308, n52309, n52310, n52311, n52312, n52313, n52314,
         n52315, n52316, n52317, n52318, n52319, n52320, n52321, n52322,
         n52323, n52324, n52325, n52326, n52327, n52328, n52329, n52330,
         n52331, n52332, n52333, n52334, n52335, n52336, n52337, n52338,
         n52339, n52340, n52341, n52342, n52343, n52344, n52345, n52346,
         n52347, n52348, n52349, n52350, n52351, n52352, n52353, n52354,
         n52355, n52356, n52357, n52358, n52359, n52360, n52361, n52362,
         n52363, n52364, n52365, n52366, n52367, n52368, n52369, n52370,
         n52371, n52372, n52373, n52374, n52375, n52376, n52377, n52378,
         n52379, n52380, n52381, n52382, n52383, n52384, n52385, n52386,
         n52387, n52388, n52389, n52390, n52391, n52392, n52393, n52394,
         n52395, n52396, n52397, n52398, n52399, n52400, n52401, n52402,
         n52403, n52404, n52405, n52406, n52407, n52408, n52409, n52410,
         n52411, n52412, n52413, n52414, n52415, n52416, n52417, n52418,
         n52419, n52420, n52421, n52422, n52423, n52424, n52425, n52426,
         n52427, n52428, n52429, n52430, n52431, n52432, n52433, n52434,
         n52435, n52436, n52437, n52438, n52439, n52440, n52441, n52442,
         n52443, n52444, n52445, n52446, n52447, n52448, n52449, n52450,
         n52451, n52452, n52453, n52454, n52455, n52456, n52457, n52458,
         n52459, n52460, n52461, n52462, n52463, n52464, n52465, n52466,
         n52467, n52468, n52469, n52470, n52471, n52472, n52473, n52474,
         n52475, n52476, n52477, n52478, n52479, n52480, n52481, n52482,
         n52483, n52484, n52485, n52486, n52487, n52488, n52489, n52490,
         n52491, n52492, n52493, n52494, n52495, n52496, n52497, n52498,
         n52499, n52500, n52501, n52502, n52503, n52504, n52505, n52506,
         n52507, n52508, n52509, n52510, n52511, n52512, n52513, n52514,
         n52515, n52516, n52517, n52518, n52519, n52520, n52521, n52522,
         n52523, n52524, n52525, n52526, n52527, n52528, n52529, n52530,
         n52531, n52532, n52533, n52534, n52535, n52536, n52537, n52538,
         n52539, n52540, n52541, n52542, n52543, n52544, n52545, n52546,
         n52547, n52548, n52549, n52550, n52551, n52552, n52553, n52554,
         n52555, n52556, n52557, n52558, n52559, n52560, n52561, n52562,
         n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570,
         n52571, n52572, n52573, n52574, n52575, n52576, n52577, n52578,
         n52579, n52580, n52581, n52582, n52583, n52584, n52585, n52586,
         n52587, n52588, n52589, n52590, n52591, n52592, n52593, n52594,
         n52595, n52596, n52597, n52598, n52599, n52600, n52601, n52602,
         n52603, n52604, n52605, n52606, n52607, n52608, n52609, n52610,
         n52611, n52612, n52613, n52614, n52615, n52616, n52617, n52618,
         n52619, n52620, n52621, n52622, n52623, n52624, n52625, n52626,
         n52627, n52628, n52629, n52630, n52631, n52632, n52633, n52634,
         n52635, n52636, n52637, n52638, n52639, n52640, n52641, n52642,
         n52643, n52644, n52645, n52646, n52647, n52648, n52649, n52650,
         n52651, n52652, n52653, n52654, n52655, n52656, n52657, n52658,
         n52659, n52660, n52661, n52662, n52663, n52664, n52665, n52666,
         n52667, n52668, n52669, n52670, n52671, n52672, n52673, n52674,
         n52675, n52676, n52677, n52678, n52679, n52680, n52681, n52682,
         n52683, n52684, n52685, n52686, n52687, n52688, n52689, n52690,
         n52691, n52692, n52693, n52694, n52695, n52696, n52697, n52698,
         n52699, n52700, n52701, n52702, n52703, n52704, n52705, n52706,
         n52707, n52708, n52709, n52710, n52711, n52712, n52713, n52714,
         n52715, n52716, n52717, n52718, n52719, n52720, n52721, n52722,
         n52723, n52724, n52725, n52726, n52727, n52728, n52729, n52730,
         n52731, n52732, n52733, n52734, n52735, n52736, n52737, n52738,
         n52739, n52740, n52741, n52742, n52743, n52744, n52745, n52746,
         n52747, n52748, n52749, n52750, n52751, n52752, n52753, n52754,
         n52755, n52756, n52757, n52758, n52759, n52760, n52761, n52762,
         n52763, n52764, n52765, n52766, n52767, n52768, n52769, n52770,
         n52771, n52772, n52773, n52774, n52775, n52776, n52777, n52778,
         n52779, n52780, n52781, n52782, n52783, n52784, n52785, n52786,
         n52787, n52788, n52789, n52790, n52791, n52792, n52793, n52794,
         n52795, n52796, n52797, n52798, n52799, n52800, n52801, n52802,
         n52803, n52804, n52805, n52806, n52807, n52808, n52809, n52810,
         n52811, n52812, n52813, n52814, n52815, n52816, n52817, n52818,
         n52819, n52820, n52821, n52822, n52823, n52824, n52825, n52826,
         n52827, n52828, n52829, n52830, n52831, n52832, n52833, n52834,
         n52835, n52836, n52837, n52838, n52839, n52840, n52841, n52842,
         n52843, n52844, n52845, n52846, n52847, n52848, n52849, n52850,
         n52851, n52852, n52853, n52854, n52855, n52856, n52857, n52858,
         n52859, n52860, n52861, n52862, n52863, n52864, n52865, n52866,
         n52867, n52868, n52869, n52870, n52871, n52872, n52873, n52874,
         n52875, n52876, n52877, n52878, n52879, n52880, n52881, n52882,
         n52883, n52884, n52885, n52886, n52887, n52888, n52889, n52890,
         n52891, n52892, n52893, n52894, n52895, n52896, n52897, n52898,
         n52899, n52900, n52901, n52902, n52903, n52904, n52905, n52906,
         n52907, n52908, n52909, n52910, n52911, n52912, n52913, n52914,
         n52915, n52916, n52917, n52918, n52919, n52920, n52921, n52922,
         n52923, n52924, n52925, n52926, n52927, n52928, n52929, n52930,
         n52931, n52932, n52933, n52934, n52935, n52936, n52937, n52938,
         n52939, n52940, n52941, n52942, n52943, n52944, n52945, n52946,
         n52947, n52948, n52949, n52950, n52951, n52952, n52953, n52954,
         n52955, n52956, n52957, n52958, n52959, n52960, n52961, n52962,
         n52963, n52964, n52965, n52966, n52967, n52968, n52969, n52970,
         n52971, n52972, n52973, n52974, n52975, n52976, n52977, n52978,
         n52979, n52980, n52981, n52982, n52983, n52984, n52985, n52986,
         n52987, n52988, n52989, n52990, n52991, n52992, n52993, n52994,
         n52995, n52996, n52997, n52998, n52999, n53000, n53001, n53002,
         n53003, n53004, n53005, n53006, n53007, n53008, n53009, n53010,
         n53011, n53012, n53013, n53014, n53015, n53016, n53017, n53018,
         n53019, n53020, n53021, n53022, n53023, n53024, n53025, n53026,
         n53027, n53028, n53029, n53030, n53031, n53032, n53033, n53034,
         n53035, n53036, n53037, n53038, n53039, n53040, n53041, n53042,
         n53043, n53044, n53045, n53046, n53047, n53048, n53049, n53050,
         n53051, n53052, n53053, n53054, n53055, n53056, n53057, n53058,
         n53059, n53060, n53061, n53062, n53063, n53064, n53065, n53066,
         n53067, n53068, n53069, n53070, n53071, n53072, n53073, n53074,
         n53075, n53076, n53077, n53078, n53079, n53080, n53081, n53082,
         n53083, n53084, n53085, n53086, n53087, n53088, n53089, n53090,
         n53091, n53092, n53093, n53094, n53095, n53096, n53097, n53098,
         n53099, n53100, n53101, n53102, n53103, n53104, n53105, n53106,
         n53107, n53108, n53109, n53110, n53111, n53112, n53113, n53114,
         n53115, n53116, n53117, n53118, n53119, n53120, n53121, n53122,
         n53123, n53124, n53125, n53126, n53127, n53128, n53129, n53130,
         n53131, n53132, n53133, n53134, n53135, n53136, n53137, n53138,
         n53139, n53140, n53141, n53142, n53143, n53144, n53145, n53146,
         n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154,
         n53155, n53156, n53157, n53158, n53159, n53160, n53161, n53162,
         n53163, n53164, n53165, n53166, n53167, n53168, n53169, n53170,
         n53171, n53172, n53173, n53174, n53175, n53176, n53177, n53178,
         n53179, n53180, n53181, n53182, n53183, n53184, n53185, n53186,
         n53187, n53188, n53189, n53190, n53191, n53192, n53193, n53194,
         n53195, n53196, n53197, n53198, n53199, n53200, n53201, n53202,
         n53203, n53204, n53205, n53206, n53207, n53208, n53209, n53210,
         n53211, n53212, n53213, n53214, n53215, n53216, n53217, n53218,
         n53219, n53220, n53221, n53222, n53223, n53224, n53225, n53226,
         n53227, n53228, n53229, n53230, n53231, n53232, n53233, n53234,
         n53235, n53236, n53237, n53238, n53239, n53240, n53241, n53242,
         n53243, n53244, n53245, n53246, n53247, n53248, n53249, n53250,
         n53251, n53252, n53253, n53254, n53255, n53256, n53257, n53258,
         n53259, n53260, n53261, n53262, n53263, n53264, n53265, n53266,
         n53267, n53268, n53269, n53270, n53271, n53272, n53273, n53274,
         n53275, n53276, n53277, n53278, n53279, n53280, n53281, n53282,
         n53283, n53284, n53285, n53286, n53287, n53288, n53289, n53290,
         n53291, n53292, n53293, n53294, n53295, n53296, n53297, n53298,
         n53299, n53300, n53301, n53302, n53303, n53304, n53305, n53306,
         n53307, n53308, n53309, n53310, n53311, n53312, n53313, n53314,
         n53315, n53316, n53317, n53318, n53319, n53320, n53321, n53322,
         n53323, n53324, n53325, n53326, n53327, n53328, n53329, n53330,
         n53331, n53332, n53333, n53334, n53335, n53336, n53337, n53338,
         n53339, n53340, n53341, n53342, n53343, n53344, n53345, n53346,
         n53347, n53348, n53349, n53350, n53351, n53352, n53353, n53354,
         n53355, n53356, n53357, n53358, n53359, n53360, n53361, n53362,
         n53363, n53364, n53365, n53366, n53367, n53368, n53369, n53370,
         n53371, n53372, n53373, n53374, n53375, n53376, n53377, n53378,
         n53379, n53380, n53381, n53382, n53383, n53384, n53385, n53386,
         n53387, n53388, n53389, n53390, n53391, n53392, n53393, n53394,
         n53395, n53396, n53397, n53398, n53399, n53400, n53401, n53402,
         n53403, n53404, n53405, n53406, n53407, n53408, n53409, n53410,
         n53411, n53412, n53413, n53414, n53415, n53416, n53417, n53418,
         n53419, n53420, n53421, n53422, n53423, n53424, n53425, n53426,
         n53427, n53428, n53429, n53430, n53431, n53432, n53433, n53434,
         n53435, n53436, n53437, n53438, n53439, n53440, n53441, n53442,
         n53443, n53444, n53445, n53446, n53447, n53448, n53449, n53450,
         n53451, n53452, n53453, n53454, n53455, n53456, n53457, n53458,
         n53459, n53460, n53461, n53462, n53463, n53464, n53465, n53466,
         n53467, n53468, n53469, n53470, n53471, n53472, n53473, n53474,
         n53475, n53476, n53477, n53478, n53479, n53480, n53481, n53482,
         n53483, n53484, n53485, n53486, n53487, n53488, n53489, n53490,
         n53491, n53492, n53493, n53494, n53495, n53496, n53497, n53498,
         n53499, n53500, n53501, n53502, n53503, n53504, n53505, n53506,
         n53507, n53508, n53509, n53510, n53511, n53512, n53513, n53514,
         n53515, n53516, n53517, n53518, n53519, n53520, n53521, n53522,
         n53523, n53524, n53525, n53526, n53527, n53528, n53529, n53530,
         n53531, n53532, n53533, n53534, n53535, n53536, n53537, n53538,
         n53539, n53540, n53541, n53542, n53543, n53544, n53545, n53546,
         n53547, n53548, n53549, n53550, n53551, n53552, n53553, n53554,
         n53555, n53556, n53557, n53558, n53559, n53560, n53561, n53562,
         n53563, n53564, n53565, n53566, n53567, n53568, n53569, n53570,
         n53571, n53572, n53573, n53574, n53575, n53576, n53577, n53578,
         n53579, n53580, n53581, n53582, n53583, n53584, n53585, n53586,
         n53587, n53588, n53589, n53590, n53591, n53592, n53593, n53594,
         n53595, n53596, n53597, n53598, n53599, n53600, n53601, n53602,
         n53603, n53604, n53605, n53606, n53607, n53608, n53609, n53610,
         n53611, n53612, n53613, n53614, n53615, n53616, n53617, n53618,
         n53619, n53620, n53621, n53622, n53623, n53624, n53625, n53626,
         n53627, n53628, n53629, n53630, n53631, n53632, n53633, n53634,
         n53635, n53636, n53637, n53638, n53639, n53640, n53641, n53642,
         n53643, n53644, n53645, n53646, n53647, n53648, n53649, n53650,
         n53651, n53652, n53653, n53654, n53655, n53656, n53657, n53658,
         n53659, n53660, n53661, n53662, n53663, n53664, n53665, n53666,
         n53667, n53668, n53669, n53670, n53671, n53672, n53673, n53674,
         n53675, n53676, n53677, n53678, n53679, n53680, n53681, n53682,
         n53683, n53684, n53685, n53686, n53687, n53688, n53689, n53690,
         n53691, n53692, n53693, n53694, n53695, n53696, n53697, n53698,
         n53699, n53700, n53701, n53702, n53703, n53704, n53705, n53706,
         n53707, n53708, n53709, n53710, n53711, n53712, n53713, n53714,
         n53715, n53716, n53717, n53718, n53719, n53720, n53721, n53722,
         n53723, n53724, n53725, n53726, n53727, n53728, n53729, n53730,
         n53731, n53732, n53733, n53734, n53735, n53736, n53737, n53738,
         n53739, n53740, n53741, n53742, n53743, n53744, n53745, n53746,
         n53747, n53748, n53749, n53750, n53751, n53752, n53753, n53754,
         n53755, n53756, n53757, n53758, n53759, n53760, n53761, n53762,
         n53763, n53764, n53765, n53766, n53767, n53768, n53769, n53770,
         n53771, n53772, n53773, n53774, n53775, n53776, n53777, n53778,
         n53779, n53780, n53781, n53782, n53783, n53784, n53785, n53786,
         n53787, n53788, n53789, n53790, n53791, n53792, n53793, n53794,
         n53795, n53796, n53797, n53798, n53799, n53800, n53801, n53802,
         n53803, n53804, n53805, n53806, n53807, n53808, n53809, n53810,
         n53811, n53812, n53813, n53814, n53815, n53816, n53817, n53818,
         n53819, n53820, n53821, n53822, n53823, n53824, n53825, n53826,
         n53827, n53828, n53829, n53830, n53831, n53832, n53833, n53834,
         n53835, n53836, n53837, n53838, n53839, n53840, n53841, n53842,
         n53843, n53844, n53845, n53846, n53847, n53848, n53849, n53850,
         n53851, n53852, n53853, n53854, n53855, n53856, n53857, n53858,
         n53859, n53860, n53861, n53862, n53863, n53864, n53865, n53866,
         n53867, n53868, n53869, n53870, n53871, n53872, n53873, n53874,
         n53875, n53876, n53877, n53878, n53879, n53880, n53881, n53882,
         n53883, n53884, n53885, n53886, n53887, n53888, n53889, n53890,
         n53891, n53892, n53893, n53894, n53895, n53896, n53897, n53898,
         n53899, n53900, n53901, n53902, n53903, n53904, n53905, n53906,
         n53907, n53908, n53909, n53910, n53911, n53912, n53913, n53914,
         n53915, n53916, n53917, n53918, n53919, n53920, n53921, n53922,
         n53923, n53924, n53925, n53926, n53927, n53928, n53929, n53930,
         n53931, n53932, n53933, n53934, n53935, n53936, n53937, n53938,
         n53939, n53940, n53941, n53942, n53943, n53944, n53945, n53946,
         n53947, n53948, n53949, n53950, n53951, n53952, n53953, n53954,
         n53955, n53956, n53957, n53958, n53959, n53960, n53961, n53962,
         n53963, n53964, n53965, n53966, n53967, n53968, n53969, n53970,
         n53971, n53972, n53973, n53974, n53975, n53976, n53977, n53978,
         n53979, n53980, n53981, n53982, n53983, n53984, n53985, n53986,
         n53987, n53988, n53989, n53990, n53991, n53992, n53993, n53994,
         n53995, n53996, n53997, n53998, n53999, n54000, n54001, n54002,
         n54003, n54004, n54005, n54006, n54007, n54008, n54009, n54010,
         n54011, n54012, n54013, n54014, n54015, n54016, n54017, n54018,
         n54019, n54020, n54021, n54022, n54023, n54024, n54025, n54026,
         n54027, n54028, n54029, n54030, n54031, n54032, n54033, n54034,
         n54035, n54036, n54037, n54038, n54039, n54040, n54041, n54042,
         n54043, n54044, n54045, n54046, n54047, n54048, n54049, n54050,
         n54051, n54052, n54053, n54054, n54055, n54056, n54057, n54058,
         n54059, n54060, n54061, n54062, n54063, n54064, n54065, n54066,
         n54067, n54068, n54069, n54070, n54071, n54072, n54073, n54074,
         n54075, n54076, n54077, n54078, n54079, n54080, n54081, n54082,
         n54083, n54084, n54085, n54086, n54087, n54088, n54089, n54090,
         n54091, n54092, n54093, n54094, n54095, n54096, n54097, n54098,
         n54099, n54100, n54101, n54102, n54103, n54104, n54105, n54106,
         n54107, n54108, n54109, n54110, n54111, n54112, n54113, n54114,
         n54115, n54116, n54117, n54118, n54119, n54120, n54121, n54122,
         n54123, n54124, n54125, n54126, n54127, n54128, n54129, n54130,
         n54131, n54132, n54133, n54134, n54135, n54136, n54137, n54138,
         n54139, n54140, n54141, n54142, n54143, n54144, n54145, n54146,
         n54147, n54148, n54149, n54150, n54151, n54152, n54153, n54154,
         n54155, n54156, n54157, n54158, n54159, n54160, n54161, n54162,
         n54163, n54164, n54165, n54166, n54167, n54168, n54169, n54170,
         n54171, n54172, n54173, n54174, n54175, n54176, n54177, n54178,
         n54179, n54180, n54181, n54182, n54183, n54184, n54185, n54186,
         n54187, n54188, n54189, n54190, n54191, n54192, n54193, n54194,
         n54195, n54196, n54197, n54198, n54199, n54200, n54201, n54202,
         n54203, n54204, n54205, n54206, n54207, n54208, n54209, n54210,
         n54211, n54212, n54213, n54214, n54215, n54216, n54217, n54218,
         n54219, n54220, n54221, n54222, n54223, n54224, n54225, n54226,
         n54227, n54228, n54229, n54230, n54231, n54232, n54233, n54234,
         n54235, n54236, n54237, n54238, n54239, n54240, n54241, n54242,
         n54243, n54244, n54245, n54246, n54247, n54248, n54249, n54250,
         n54251, n54252, n54253, n54254, n54255, n54256, n54257, n54258,
         n54259, n54260, n54261, n54262, n54263, n54264, n54265, n54266,
         n54267, n54268, n54269, n54270, n54271, n54272, n54273, n54274,
         n54275, n54276, n54277, n54278, n54279, n54280, n54281, n54282,
         n54283, n54284, n54285, n54286, n54287, n54288, n54289, n54290,
         n54291, n54292, n54293, n54294, n54295, n54296, n54297, n54298,
         n54299, n54300, n54301, n54302, n54303, n54304, n54305, n54306,
         n54307, n54308, n54309, n54310, n54311, n54312, n54313, n54314,
         n54315, n54316, n54317, n54318, n54319, n54320, n54321, n54322,
         n54323, n54324, n54325, n54326, n54327, n54328, n54329, n54330,
         n54331, n54332, n54333, n54334, n54335, n54336, n54337, n54338,
         n54339, n54340, n54341, n54342, n54343, n54344, n54345, n54346,
         n54347, n54348, n54349, n54350, n54351, n54352, n54353, n54354,
         n54355, n54356, n54357, n54358, n54359, n54360, n54361, n54362,
         n54363, n54364, n54365, n54366, n54367, n54368, n54369, n54370,
         n54371, n54372, n54373, n54374, n54375, n54376, n54377, n54378,
         n54379, n54380, n54381, n54382, n54383, n54384, n54385, n54386,
         n54387, n54388, n54389, n54390, n54391, n54392, n54393, n54394,
         n54395, n54396, n54397, n54398, n54399, n54400, n54401, n54402,
         n54403, n54404, n54405, n54406, n54407, n54408, n54409, n54410,
         n54411, n54412, n54413, n54414, n54415, n54416, n54417, n54418,
         n54419, n54420, n54421, n54422, n54423, n54424, n54425, n54426,
         n54427, n54428, n54429, n54430, n54431, n54432, n54433, n54434,
         n54435, n54436, n54437, n54438, n54439, n54440, n54441, n54442,
         n54443, n54444, n54445, n54446, n54447, n54448, n54449, n54450,
         n54451, n54452, n54453, n54454, n54455, n54456, n54457, n54458,
         n54459, n54460, n54461, n54462, n54463, n54464, n54465, n54466,
         n54467, n54468, n54469, n54470, n54471, n54472, n54473, n54474,
         n54475, n54476, n54477, n54478, n54479, n54480, n54481, n54482,
         n54483, n54484, n54485, n54486, n54487, n54488, n54489, n54490,
         n54491, n54492, n54493, n54494, n54495, n54496, n54497, n54498,
         n54499, n54500, n54501, n54502, n54503, n54504, n54505, n54506,
         n54507, n54508, n54509, n54510, n54511, n54512, n54513, n54514,
         n54515, n54516, n54517, n54518, n54519, n54520, n54521, n54522,
         n54523, n54524, n54525, n54526, n54527, n54528, n54529, n54530,
         n54531, n54532, n54533, n54534, n54535, n54536, n54537, n54538,
         n54539, n54540, n54541, n54542, n54543, n54544, n54545, n54546,
         n54547, n54548, n54549, n54550, n54551, n54552, n54553, n54554,
         n54555, n54556, n54557, n54558, n54559, n54560, n54561, n54562,
         n54563, n54564, n54565, n54566, n54567, n54568, n54569, n54570,
         n54571, n54572, n54573, n54574, n54575, n54576, n54577, n54578,
         n54579, n54580, n54581, n54582, n54583, n54584, n54585, n54586,
         n54587, n54588, n54589, n54590, n54591, n54592, n54593, n54594,
         n54595, n54596, n54597, n54598, n54599, n54600, n54601, n54602,
         n54603, n54604, n54605, n54606, n54607, n54608, n54609, n54610,
         n54611, n54612, n54613, n54614, n54615, n54616, n54617, n54618,
         n54619, n54620, n54621, n54622, n54623, n54624, n54625, n54626,
         n54627, n54628, n54629, n54630, n54631, n54632, n54633, n54634,
         n54635, n54636, n54637, n54638, n54639, n54640, n54641, n54642,
         n54643, n54644, n54645, n54646, n54647, n54648, n54649, n54650,
         n54651, n54652, n54653, n54654, n54655, n54656, n54657, n54658,
         n54659, n54660, n54661, n54662, n54663, n54664, n54665, n54666,
         n54667, n54668, n54669, n54670, n54671, n54672, n54673, n54674,
         n54675, n54676, n54677, n54678, n54679, n54680, n54681, n54682,
         n54683, n54684, n54685, n54686, n54687, n54688, n54689, n54690,
         n54691, n54692, n54693, n54694, n54695, n54696, n54697, n54698,
         n54699, n54700, n54701, n54702, n54703, n54704, n54705, n54706,
         n54707, n54708, n54709, n54710, n54711, n54712, n54713, n54714,
         n54715, n54716, n54717, n54718, n54719, n54720, n54721, n54722,
         n54723, n54724, n54725, n54726, n54727, n54728, n54729, n54730,
         n54731, n54732, n54733, n54734, n54735, n54736, n54737, n54738,
         n54739, n54740, n54741, n54742, n54743, n54744, n54745, n54746,
         n54747, n54748, n54749, n54750, n54751, n54752, n54753, n54754,
         n54755, n54756, n54757, n54758, n54759, n54760, n54761, n54762,
         n54763, n54764, n54765, n54766, n54767, n54768, n54769, n54770,
         n54771, n54772, n54773, n54774, n54775, n54776, n54777, n54778,
         n54779, n54780, n54781, n54782, n54783, n54784, n54785, n54786,
         n54787, n54788, n54789, n54790, n54791, n54792, n54793, n54794,
         n54795, n54796, n54797, n54798, n54799, n54800, n54801, n54802,
         n54803, n54804, n54805, n54806, n54807, n54808, n54809, n54810,
         n54811, n54812, n54813, n54814, n54815, n54816, n54817, n54818,
         n54819, n54820, n54821, n54822, n54823, n54824, n54825, n54826,
         n54827, n54828, n54829, n54830, n54831, n54832, n54833, n54834,
         n54835, n54836, n54837, n54838, n54839, n54840, n54841, n54842,
         n54843, n54844, n54845, n54846, n54847, n54848, n54849, n54850,
         n54851, n54852, n54853, n54854, n54855, n54856, n54857, n54858,
         n54859, n54860, n54861, n54862, n54863, n54864, n54865, n54866,
         n54867, n54868, n54869, n54870, n54871, n54872, n54873, n54874,
         n54875, n54876, n54877, n54878, n54879, n54880, n54881, n54882,
         n54883, n54884, n54885, n54886, n54887, n54888, n54889, n54890,
         n54891, n54892, n54893, n54894, n54895, n54896, n54897, n54898,
         n54899, n54900, n54901, n54902, n54903, n54904, n54905, n54906,
         n54907, n54908, n54909, n54910, n54911, n54912, n54913, n54914,
         n54915, n54916, n54917, n54918, n54919, n54920, n54921, n54922,
         n54923, n54924, n54925, n54926, n54927, n54928, n54929, n54930,
         n54931, n54932, n54933, n54934, n54935, n54936, n54937, n54938,
         n54939, n54940, n54941, n54942, n54943, n54944, n54945, n54946,
         n54947, n54948, n54949, n54950, n54951, n54952, n54953, n54954,
         n54955, n54956, n54957, n54958, n54959, n54960, n54961, n54962,
         n54963, n54964, n54965, n54966, n54967, n54968, n54969, n54970,
         n54971, n54972, n54973, n54974, n54975, n54976, n54977, n54978,
         n54979, n54980, n54981, n54982, n54983, n54984, n54985, n54986,
         n54987, n54988, n54989, n54990, n54991, n54992, n54993, n54994,
         n54995, n54996, n54997, n54998, n54999, n55000, n55001, n55002,
         n55003, n55004, n55005, n55006, n55007, n55008, n55009, n55010,
         n55011, n55012, n55013, n55014, n55015, n55016, n55017, n55018,
         n55019, n55020, n55021, n55022, n55023, n55024, n55025, n55026,
         n55027, n55028, n55029, n55030, n55031, n55032, n55033, n55034,
         n55035, n55036, n55037, n55038, n55039, n55040, n55041, n55042,
         n55043, n55044, n55045, n55046, n55047, n55048, n55049, n55050,
         n55051, n55052, n55053, n55054, n55055, n55056, n55057, n55058,
         n55059, n55060, n55061, n55062, n55063, n55064, n55065, n55066,
         n55067, n55068, n55069, n55070, n55071, n55072, n55073, n55074,
         n55075, n55076, n55077, n55078, n55079, n55080, n55081, n55082,
         n55083, n55084, n55085, n55086, n55087, n55088, n55089, n55090,
         n55091, n55092, n55093, n55094, n55095, n55096, n55097, n55098,
         n55099, n55100, n55101, n55102, n55103, n55104, n55105, n55106,
         n55107, n55108, n55109, n55110, n55111, n55112, n55113, n55114,
         n55115, n55116, n55117, n55118, n55119, n55120, n55121, n55122,
         n55123, n55124, n55125, n55126, n55127, n55128, n55129, n55130,
         n55131, n55132, n55133, n55134, n55135, n55136, n55137, n55138,
         n55139, n55140, n55141, n55142, n55143, n55144, n55145, n55146,
         n55147, n55148, n55149, n55150, n55151, n55152, n55153, n55154,
         n55155, n55156, n55157, n55158, n55159, n55160, n55161, n55162,
         n55163, n55164, n55165, n55166, n55167, n55168, n55169, n55170,
         n55171, n55172, n55173, n55174, n55175, n55176, n55177, n55178,
         n55179, n55180, n55181, n55182, n55183, n55184, n55185, n55186,
         n55187, n55188, n55189, n55190, n55191, n55192, n55193, n55194,
         n55195, n55196, n55197, n55198, n55199, n55200, n55201, n55202,
         n55203, n55204, n55205, n55206, n55207, n55208, n55209, n55210,
         n55211, n55212, n55213, n55214, n55215, n55216, n55217, n55218,
         n55219, n55220, n55221, n55222, n55223, n55224, n55225, n55226,
         n55227, n55228, n55229, n55230, n55231, n55232, n55233, n55234,
         n55235, n55236, n55237, n55238, n55239, n55240, n55241, n55242,
         n55243, n55244, n55245, n55246, n55247, n55248, n55249, n55250,
         n55251, n55252, n55253, n55254, n55255, n55256, n55257, n55258,
         n55259, n55260, n55261, n55262, n55263, n55264, n55265, n55266,
         n55267, n55268, n55269, n55270, n55271, n55272, n55273, n55274,
         n55275, n55276, n55277, n55278, n55279, n55280, n55281, n55282,
         n55283, n55284, n55285, n55286, n55287, n55288, n55289, n55290,
         n55291, n55292, n55293, n55294, n55295, n55296, n55297, n55298,
         n55299, n55300, n55301, n55302, n55303, n55304, n55305, n55306,
         n55307, n55308, n55309, n55310, n55311, n55312, n55313, n55314,
         n55315, n55316, n55317, n55318, n55319, n55320, n55321, n55322,
         n55323, n55324, n55325, n55326, n55327, n55328, n55329, n55330,
         n55331, n55332, n55333, n55334, n55335, n55336, n55337, n55338,
         n55339, n55340, n55341, n55342, n55343, n55344, n55345, n55346,
         n55347, n55348, n55349, n55350, n55351, n55352, n55353, n55354,
         n55355, n55356, n55357, n55358, n55359, n55360, n55361, n55362,
         n55363, n55364, n55365, n55366, n55367, n55368, n55369, n55370,
         n55371, n55372, n55373, n55374, n55375, n55376, n55377, n55378,
         n55379, n55380, n55381, n55382, n55383, n55384, n55385, n55386,
         n55387, n55388, n55389, n55390, n55391, n55392, n55393, n55394,
         n55395, n55396, n55397, n55398, n55399, n55400, n55401, n55402,
         n55403, n55404, n55405, n55406, n55407, n55408, n55409, n55410,
         n55411, n55412, n55413, n55414, n55415, n55416, n55417, n55418,
         n55419, n55420, n55421, n55422, n55423, n55424, n55425, n55426,
         n55427, n55428, n55429, n55430, n55431, n55432, n55433, n55434,
         n55435, n55436, n55437, n55438, n55439, n55440, n55441, n55442,
         n55443, n55444, n55445, n55446, n55447, n55448, n55449, n55450,
         n55451, n55452, n55453, n55454, n55455, n55456, n55457, n55458,
         n55459, n55460, n55461, n55462, n55463, n55464, n55465, n55466,
         n55467, n55468, n55469, n55470, n55471, n55472, n55473, n55474,
         n55475, n55476, n55477, n55478, n55479, n55480, n55481, n55482,
         n55483, n55484, n55485, n55486, n55487, n55488, n55489, n55490,
         n55491, n55492, n55493, n55494, n55495, n55496, n55497, n55498,
         n55499, n55500, n55501, n55502, n55503, n55504, n55505, n55506,
         n55507, n55508, n55509, n55510, n55511, n55512, n55513, n55514,
         n55515, n55516, n55517, n55518, n55519, n55520, n55521, n55522,
         n55523, n55524, n55525, n55526, n55527, n55528, n55529, n55530,
         n55531, n55532, n55533, n55534, n55535, n55536, n55537, n55538,
         n55539, n55540, n55541, n55542, n55543, n55544, n55545, n55546,
         n55547, n55548, n55549, n55550, n55551, n55552, n55553, n55554,
         n55555, n55556, n55557, n55558, n55559, n55560, n55561, n55562,
         n55563, n55564, n55565, n55566, n55567, n55568, n55569, n55570,
         n55571, n55572, n55573, n55574, n55575, n55576, n55577, n55578,
         n55579, n55580, n55581, n55582, n55583, n55584, n55585, n55586,
         n55587, n55588, n55589, n55590, n55591, n55592, n55593, n55594,
         n55595, n55596, n55597, n55598, n55599, n55600, n55601, n55602,
         n55603, n55604, n55605, n55606, n55607, n55608, n55609, n55610,
         n55611, n55612, n55613, n55614, n55615, n55616, n55617, n55618,
         n55619, n55620, n55621, n55622, n55623, n55624, n55625, n55626,
         n55627, n55628, n55629, n55630, n55631, n55632, n55633, n55634,
         n55635, n55636, n55637, n55638, n55639, n55640, n55641, n55642,
         n55643, n55644, n55645, n55646, n55647, n55648, n55649, n55650,
         n55651, n55652, n55653, n55654, n55655, n55656, n55657, n55658,
         n55659, n55660, n55661, n55662, n55663, n55664, n55665, n55666,
         n55667, n55668, n55669, n55670, n55671, n55672, n55673, n55674,
         n55675, n55676, n55677, n55678, n55679, n55680, n55681, n55682,
         n55683, n55684, n55685, n55686, n55687, n55688, n55689, n55690,
         n55691, n55692, n55693, n55694, n55695, n55696, n55697, n55698,
         n55699, n55700, n55701, n55702, n55703, n55704, n55705, n55706,
         n55707, n55708, n55709, n55710, n55711, n55712, n55713, n55714,
         n55715, n55716, n55717, n55718, n55719, n55720, n55721, n55722,
         n55723, n55724, n55725, n55726, n55727, n55728, n55729, n55730,
         n55731, n55732, n55733, n55734, n55735, n55736, n55737, n55738,
         n55739, n55740, n55741, n55742, n55743, n55744, n55745, n55746,
         n55747, n55748, n55749, n55750, n55751, n55752, n55753, n55754,
         n55755, n55756, n55757, n55758, n55759, n55760, n55761, n55762,
         n55763, n55764, n55765, n55766, n55767, n55768, n55769, n55770,
         n55771, n55772, n55773, n55774, n55775, n55776, n55777, n55778,
         n55779, n55780, n55781, n55782, n55783, n55784, n55785, n55786,
         n55787, n55788, n55789, n55790, n55791, n55792, n55793, n55794,
         n55795, n55796, n55797, n55798, n55799, n55800, n55801, n55802,
         n55803, n55804, n55805, n55806, n55807, n55808, n55809, n55810,
         n55811, n55812, n55813, n55814, n55815, n55816, n55817, n55818,
         n55819, n55820, n55821, n55822, n55823, n55824, n55825, n55826,
         n55827, n55828, n55829, n55830, n55831, n55832, n55833, n55834,
         n55835, n55836, n55837, n55838, n55839, n55840, n55841, n55842,
         n55843, n55844, n55845, n55846, n55847, n55848, n55849, n55850,
         n55851, n55852, n55853, n55854, n55855, n55856, n55857, n55858,
         n55859, n55860, n55861, n55862, n55863, n55864, n55865, n55866,
         n55867, n55868, n55869, n55870, n55871, n55872, n55873, n55874,
         n55875, n55876, n55877, n55878, n55879, n55880, n55881, n55882,
         n55883, n55884, n55885, n55886, n55887, n55888, n55889, n55890,
         n55891, n55892, n55893, n55894, n55895, n55896, n55897, n55898,
         n55899, n55900, n55901, n55902, n55903, n55904, n55905, n55906,
         n55907, n55908, n55909, n55910, n55911, n55912, n55913, n55914,
         n55915, n55916, n55917, n55918, n55919, n55920, n55921, n55922,
         n55923, n55924, n55925, n55926, n55927, n55928, n55929, n55930,
         n55931, n55932, n55933, n55934, n55935, n55936, n55937, n55938,
         n55939, n55940, n55941, n55942, n55943, n55944, n55945, n55946,
         n55947, n55948, n55949, n55950, n55951, n55952, n55953, n55954,
         n55955, n55956, n55957, n55958, n55959, n55960, n55961, n55962,
         n55963, n55964, n55965, n55966, n55967, n55968, n55969, n55970,
         n55971, n55972, n55973, n55974, n55975, n55976, n55977, n55978,
         n55979, n55980, n55981, n55982, n55983, n55984, n55985, n55986,
         n55987, n55988, n55989, n55990, n55991, n55992, n55993, n55994,
         n55995, n55996, n55997, n55998, n55999, n56000, n56001, n56002,
         n56003, n56004, n56005, n56006, n56007, n56008, n56009, n56010,
         n56011, n56012, n56013, n56014, n56015, n56016, n56017, n56018,
         n56019, n56020, n56021, n56022, n56023, n56024, n56025, n56026,
         n56027, n56028, n56029, n56030, n56031, n56032, n56033, n56034,
         n56035, n56036, n56037, n56038, n56039, n56040, n56041, n56042,
         n56043, n56044, n56045, n56046, n56047, n56048, n56049, n56050,
         n56051, n56052, n56053, n56054, n56055, n56056, n56057, n56058,
         n56059, n56060, n56061, n56062, n56063, n56064, n56065, n56066,
         n56067, n56068, n56069, n56070, n56071, n56072, n56073, n56074,
         n56075, n56076, n56077, n56078, n56079, n56080, n56081, n56082,
         n56083, n56084, n56085, n56086, n56087, n56088, n56089, n56090,
         n56091, n56092, n56093, n56094, n56095, n56096, n56097, n56098,
         n56099, n56100, n56101, n56102, n56103, n56104, n56105, n56106,
         n56107, n56108, n56109, n56110, n56111, n56112, n56113, n56114,
         n56115, n56116, n56117, n56118, n56119, n56120, n56121, n56122,
         n56123, n56124, n56125, n56126, n56127, n56128, n56129, n56130,
         n56131, n56132, n56133, n56134, n56135, n56136, n56137, n56138,
         n56139, n56140, n56141, n56142, n56143, n56144, n56145, n56146,
         n56147, n56148, n56149, n56150, n56151, n56152, n56153, n56154,
         n56155, n56156, n56157, n56158, n56159, n56160, n56161, n56162,
         n56163, n56164, n56165, n56166, n56167, n56168, n56169, n56170,
         n56171, n56172, n56173, n56174, n56175, n56176, n56177, n56178,
         n56179, n56180, n56181, n56182, n56183, n56184, n56185, n56186,
         n56187, n56188, n56189, n56190, n56191, n56192, n56193, n56194,
         n56195, n56196, n56197, n56198, n56199, n56200, n56201, n56202,
         n56203, n56204, n56205, n56206, n56207, n56208, n56209, n56210,
         n56211, n56212, n56213, n56214, n56215, n56216, n56217, n56218,
         n56219, n56220, n56221, n56222, n56223, n56224, n56225, n56226,
         n56227, n56228, n56229, n56230, n56231, n56232, n56233, n56234,
         n56235, n56236, n56237, n56238, n56239, n56240, n56241, n56242,
         n56243, n56244, n56245, n56246, n56247, n56248, n56249, n56250,
         n56251, n56252, n56253, n56254, n56255, n56256, n56257, n56258,
         n56259, n56260, n56261, n56262, n56263, n56264, n56265, n56266,
         n56267, n56268, n56269, n56270, n56271, n56272, n56273, n56274,
         n56275, n56276, n56277, n56278, n56279, n56280, n56281, n56282,
         n56283, n56284, n56285, n56286, n56287, n56288, n56289, n56290,
         n56291, n56292, n56293, n56294, n56295, n56296, n56297, n56298,
         n56299, n56300, n56301, n56302, n56303, n56304, n56305, n56306,
         n56307, n56308, n56309, n56310, n56311, n56312, n56313, n56314,
         n56315, n56316, n56317, n56318, n56319, n56320, n56321, n56322,
         n56323, n56324, n56325, n56326, n56327, n56328, n56329, n56330,
         n56331, n56332, n56333, n56334, n56335, n56336, n56337, n56338,
         n56339, n56340, n56341, n56342, n56343, n56344, n56345, n56346,
         n56347, n56348, n56349, n56350, n56351, n56352, n56353, n56354,
         n56355, n56356, n56357, n56358, n56359, n56360, n56361, n56362,
         n56363, n56364, n56365, n56366, n56367, n56368, n56369, n56370,
         n56371, n56372, n56373, n56374, n56375, n56376, n56377, n56378,
         n56379, n56380, n56381, n56382, n56383, n56384, n56385, n56386,
         n56387, n56388, n56389, n56390, n56391, n56392, n56393, n56394,
         n56395, n56396, n56397, n56398, n56399, n56400, n56401, n56402,
         n56403, n56404, n56405, n56406, n56407, n56408, n56409, n56410,
         n56411, n56412, n56413, n56414, n56415, n56416, n56417, n56418,
         n56419, n56420, n56421, n56422, n56423, n56424, n56425, n56426,
         n56427, n56428, n56429, n56430, n56431, n56432, n56433, n56434,
         n56435, n56436, n56437, n56438, n56439, n56440, n56441, n56442,
         n56443, n56444, n56445, n56446, n56447, n56448, n56449, n56450,
         n56451, n56452, n56453, n56454, n56455, n56456, n56457, n56458,
         n56459, n56460, n56461, n56462, n56463, n56464, n56465, n56466,
         n56467, n56468, n56469, n56470, n56471, n56472, n56473, n56474,
         n56475, n56476, n56477, n56478, n56479, n56480, n56481, n56482,
         n56483, n56484, n56485, n56486, n56487, n56488, n56489, n56490,
         n56491, n56492, n56493, n56494, n56495, n56496, n56497, n56498,
         n56499, n56500, n56501, n56502, n56503, n56504, n56505, n56506,
         n56507, n56508, n56509, n56510, n56511, n56512, n56513, n56514,
         n56515, n56516, n56517, n56518, n56519, n56520, n56521, n56522,
         n56523, n56524, n56525, n56526, n56527, n56528, n56529, n56530,
         n56531, n56532, n56533, n56534, n56535, n56536, n56537, n56538,
         n56539, n56540, n56541, n56542, n56543, n56544, n56545, n56546,
         n56547, n56548, n56549, n56550, n56551, n56552, n56553, n56554,
         n56555, n56556, n56557, n56558, n56559, n56560, n56561, n56562,
         n56563, n56564, n56565, n56566, n56567, n56568, n56569, n56570,
         n56571, n56572, n56573, n56574, n56575, n56576, n56577, n56578,
         n56579, n56580, n56581, n56582, n56583, n56584, n56585, n56586,
         n56587, n56588, n56589, n56590, n56591, n56592, n56593, n56594,
         n56595, n56596, n56597, n56598, n56599, n56600, n56601, n56602,
         n56603, n56604, n56605, n56606, n56607, n56608, n56609, n56610,
         n56611, n56612, n56613, n56614, n56615, n56616, n56617, n56618,
         n56619, n56620, n56621, n56622, n56623, n56624, n56625, n56626,
         n56627, n56628, n56629, n56630, n56631, n56632, n56633, n56634,
         n56635, n56636, n56637, n56638, n56639, n56640, n56641, n56642,
         n56643, n56644, n56645, n56646, n56647, n56648, n56649, n56650,
         n56651, n56652, n56653, n56654, n56655, n56656, n56657, n56658,
         n56659, n56660, n56661, n56662, n56663, n56664, n56665, n56666,
         n56667, n56668, n56669, n56670, n56671, n56672, n56673, n56674,
         n56675, n56676, n56677, n56678, n56679, n56680, n56681, n56682,
         n56683, n56684, n56685, n56686, n56687, n56688, n56689, n56690,
         n56691, n56692, n56693, n56694, n56695, n56696, n56697, n56698,
         n56699, n56700, n56701, n56702, n56703, n56704, n56705, n56706,
         n56707, n56708, n56709, n56710, n56711, n56712, n56713, n56714,
         n56715, n56716, n56717, n56718, n56719, n56720, n56721, n56722,
         n56723, n56724, n56725, n56726, n56727, n56728, n56729, n56730,
         n56731, n56732, n56733, n56734, n56735, n56736, n56737, n56738,
         n56739, n56740, n56741, n56742, n56743, n56744, n56745, n56746,
         n56747, n56748, n56749, n56750, n56751, n56752, n56753, n56754,
         n56755, n56756, n56757, n56758, n56759, n56760, n56761, n56762,
         n56763, n56764, n56765, n56766, n56767, n56768, n56769, n56770,
         n56771, n56772, n56773, n56774, n56775, n56776, n56777, n56778,
         n56779, n56780, n56781, n56782, n56783, n56784, n56785, n56786,
         n56787, n56788, n56789, n56790, n56791, n56792, n56793, n56794,
         n56795, n56796, n56797, n56798, n56799, n56800, n56801, n56802,
         n56803, n56804, n56805, n56806, n56807, n56808, n56809, n56810,
         n56811, n56812, n56813, n56814, n56815, n56816, n56817, n56818,
         n56819, n56820, n56821, n56822, n56823, n56824, n56825, n56826,
         n56827, n56828, n56829, n56830, n56831, n56832, n56833, n56834,
         n56835, n56836, n56837, n56838, n56839, n56840, n56841, n56842,
         n56843, n56844, n56845, n56846, n56847, n56848, n56849, n56850,
         n56851, n56852, n56853, n56854, n56855, n56856, n56857, n56858,
         n56859, n56860, n56861, n56862, n56863, n56864, n56865, n56866,
         n56867, n56868, n56869, n56870, n56871, n56872, n56873, n56874,
         n56875, n56876, n56877, n56878, n56879, n56880, n56881, n56882,
         n56883, n56884, n56885, n56886, n56887, n56888, n56889, n56890,
         n56891, n56892, n56893, n56894, n56895, n56896, n56897, n56898,
         n56899, n56900, n56901, n56902, n56903, n56904, n56905, n56906,
         n56907, n56908, n56909, n56910, n56911, n56912, n56913, n56914,
         n56915, n56916, n56917, n56918, n56919, n56920, n56921, n56922,
         n56923, n56924, n56925, n56926, n56927, n56928, n56929, n56930,
         n56931, n56932, n56933, n56934, n56935, n56936, n56937, n56938,
         n56939, n56940, n56941, n56942, n56943, n56944, n56945, n56946,
         n56947, n56948, n56949, n56950, n56951, n56952, n56953, n56954,
         n56955, n56956, n56957, n56958, n56959, n56960, n56961, n56962,
         n56963, n56964, n56965, n56966, n56967, n56968, n56969, n56970,
         n56971, n56972, n56973, n56974, n56975, n56976, n56977, n56978,
         n56979, n56980, n56981, n56982, n56983, n56984, n56985, n56986,
         n56987, n56988, n56989, n56990, n56991, n56992, n56993, n56994,
         n56995, n56996, n56997, n56998, n56999, n57000, n57001, n57002,
         n57003, n57004, n57005, n57006, n57007, n57008, n57009, n57010,
         n57011, n57012, n57013, n57014, n57015, n57016, n57017, n57018,
         n57019, n57020, n57021, n57022, n57023, n57024, n57025, n57026,
         n57027, n57028, n57029, n57030, n57031, n57032, n57033, n57034,
         n57035, n57036, n57037, n57038, n57039, n57040, n57041, n57042,
         n57043, n57044, n57045, n57046, n57047, n57048, n57049, n57050,
         n57051, n57052, n57053, n57054, n57055, n57056, n57057, n57058,
         n57059, n57060, n57061, n57062, n57063, n57064, n57065, n57066,
         n57067, n57068, n57069, n57070, n57071, n57072, n57073, n57074,
         n57075, n57076, n57077, n57078, n57079, n57080, n57081, n57082,
         n57083, n57084, n57085, n57086, n57087, n57088, n57089, n57090,
         n57091, n57092, n57093, n57094, n57095, n57096, n57097, n57098,
         n57099, n57100, n57101, n57102, n57103, n57104, n57105, n57106,
         n57107, n57108, n57109, n57110, n57111, n57112, n57113, n57114,
         n57115, n57116, n57117, n57118, n57119, n57120, n57121, n57122,
         n57123, n57124, n57125, n57126, n57127, n57128, n57129, n57130,
         n57131, n57132, n57133, n57134, n57135, n57136, n57137, n57138,
         n57139, n57140, n57141, n57142, n57143, n57144, n57145, n57146,
         n57147, n57148, n57149, n57150, n57151, n57152, n57153, n57154,
         n57155, n57156, n57157, n57158, n57159, n57160, n57161, n57162,
         n57163, n57164, n57165, n57166, n57167, n57168, n57169, n57170,
         n57171, n57172, n57173, n57174, n57175, n57176, n57177, n57178,
         n57179, n57180, n57181, n57182, n57183, n57184, n57185, n57186,
         n57187, n57188, n57189, n57190, n57191, n57192, n57193, n57194,
         n57195, n57196, n57197, n57198, n57199, n57200, n57201, n57202,
         n57203, n57204, n57205, n57206, n57207, n57208, n57209, n57210,
         n57211, n57212, n57213, n57214, n57215, n57216, n57217, n57218,
         n57219, n57220, n57221, n57222, n57223, n57224, n57225, n57226,
         n57227, n57228, n57229, n57230, n57231, n57232, n57233, n57234,
         n57235, n57236, n57237, n57238, n57239, n57240, n57241, n57242,
         n57243, n57244, n57245, n57246, n57247, n57248, n57249, n57250,
         n57251, n57252, n57253, n57254, n57255, n57256, n57257, n57258,
         n57259, n57260, n57261, n57262, n57263, n57264, n57265, n57266,
         n57267, n57268, n57269, n57270, n57271, n57272, n57273, n57274,
         n57275, n57276, n57277, n57278, n57279, n57280, n57281, n57282,
         n57283, n57284, n57285, n57286, n57287, n57288, n57289, n57290,
         n57291, n57292, n57293, n57294, n57295, n57296, n57297, n57298,
         n57299, n57300, n57301, n57302, n57303, n57304, n57305, n57306,
         n57307, n57308, n57309, n57310, n57311, n57312, n57313, n57314,
         n57315, n57316, n57317, n57318, n57319, n57320, n57321, n57322,
         n57323, n57324, n57325, n57326, n57327, n57328, n57329, n57330,
         n57331, n57332, n57333, n57334, n57335, n57336, n57337, n57338,
         n57339, n57340, n57341, n57342, n57343, n57344, n57345, n57346,
         n57347, n57348, n57349, n57350, n57351, n57352, n57353, n57354,
         n57355, n57356, n57357, n57358, n57359, n57360, n57361, n57362,
         n57363, n57364, n57365, n57366, n57367, n57368, n57369, n57370,
         n57371, n57372, n57373, n57374, n57375, n57376, n57377, n57378,
         n57379, n57380, n57381, n57382, n57383, n57384, n57385, n57386,
         n57387, n57388, n57389, n57390, n57391, n57392, n57393, n57394,
         n57395, n57396, n57397, n57398, n57399, n57400, n57401, n57402,
         n57403, n57404, n57405, n57406, n57407, n57408, n57409, n57410,
         n57411, n57412, n57413, n57414, n57415, n57416, n57417, n57418,
         n57419, n57420, n57421, n57422, n57423, n57424, n57425, n57426,
         n57427, n57428, n57429, n57430, n57431, n57432, n57433, n57434,
         n57435, n57436, n57437, n57438, n57439, n57440, n57441, n57442,
         n57443, n57444, n57445, n57446, n57447, n57448, n57449, n57450,
         n57451, n57452, n57453, n57454, n57455, n57456, n57457, n57458,
         n57459, n57460, n57461, n57462, n57463, n57464, n57465, n57466,
         n57467, n57468, n57469, n57470, n57471, n57472, n57473, n57474,
         n57475, n57476, n57477, n57478, n57479, n57480, n57481, n57482,
         n57483, n57484, n57485, n57486, n57487, n57488, n57489, n57490,
         n57491, n57492, n57493, n57494, n57495, n57496, n57497, n57498,
         n57499, n57500, n57501, n57502, n57503, n57504, n57505, n57506,
         n57507, n57508, n57509, n57510, n57511, n57512, n57513, n57514,
         n57515, n57516, n57517, n57518, n57519, n57520, n57521, n57522,
         n57523, n57524, n57525, n57526, n57527, n57528, n57529, n57530,
         n57531, n57532, n57533, n57534, n57535, n57536, n57537, n57538,
         n57539, n57540, n57541, n57542, n57543, n57544, n57545, n57546,
         n57547, n57548, n57549, n57550, n57551, n57552, n57553, n57554,
         n57555, n57556, n57557, n57558, n57559, n57560, n57561, n57562,
         n57563, n57564, n57565, n57566, n57567, n57568, n57569, n57570,
         n57571, n57572, n57573, n57574, n57575, n57576, n57577, n57578,
         n57579, n57580, n57581, n57582, n57583, n57584, n57585, n57586,
         n57587, n57588, n57589, n57590, n57591, n57592, n57593, n57594,
         n57595, n57596, n57597, n57598, n57599, n57600, n57601, n57602,
         n57603, n57604, n57605, n57606, n57607, n57608, n57609, n57610,
         n57611, n57612, n57613, n57614, n57615, n57616, n57617, n57618,
         n57619, n57620, n57621, n57622, n57623, n57624, n57625, n57626,
         n57627, n57628, n57629, n57630, n57631, n57632, n57633, n57634,
         n57635, n57636, n57637, n57638, n57639, n57640, n57641, n57642,
         n57643, n57644, n57645, n57646, n57647, n57648, n57649, n57650,
         n57651, n57652, n57653, n57654, n57655, n57656, n57657, n57658,
         n57659, n57660, n57661, n57662, n57663, n57664, n57665, n57666,
         n57667, n57668, n57669, n57670, n57671, n57672, n57673, n57674,
         n57675, n57676, n57677, n57678, n57679, n57680, n57681, n57682,
         n57683, n57684, n57685, n57686, n57687, n57688, n57689, n57690,
         n57691, n57692, n57693, n57694, n57695, n57696, n57697, n57698,
         n57699, n57700, n57701, n57702, n57703, n57704, n57705, n57706,
         n57707, n57708, n57709, n57710, n57711, n57712, n57713, n57714,
         n57715, n57716, n57717, n57718, n57719, n57720, n57721, n57722,
         n57723, n57724, n57725, n57726, n57727, n57728, n57729, n57730,
         n57731, n57732, n57733, n57734, n57735, n57736, n57737, n57738,
         n57739, n57740, n57741, n57742, n57743, n57744, n57745, n57746,
         n57747, n57748, n57749, n57750, n57751, n57752, n57753, n57754,
         n57755, n57756, n57757, n57758, n57759, n57760, n57761, n57762,
         n57763, n57764, n57765, n57766, n57767, n57768, n57769, n57770,
         n57771, n57772, n57773, n57774, n57775, n57776, n57777, n57778,
         n57779, n57780, n57781, n57782, n57783, n57784, n57785, n57786,
         n57787, n57788, n57789, n57790, n57791, n57792, n57793, n57794,
         n57795, n57796, n57797, n57798, n57799, n57800, n57801, n57802,
         n57803, n57804, n57805, n57806, n57807, n57808, n57809, n57810,
         n57811, n57812, n57813, n57814, n57815, n57816, n57817, n57818,
         n57819, n57820, n57821, n57822, n57823, n57824, n57825, n57826,
         n57827, n57828, n57829, n57830, n57831, n57832, n57833, n57834,
         n57835, n57836, n57837, n57838, n57839, n57840, n57841, n57842,
         n57843, n57844, n57845, n57846, n57847, n57848, n57849, n57850,
         n57851, n57852, n57853, n57854, n57855, n57856, n57857, n57858,
         n57859, n57860, n57861, n57862, n57863, n57864, n57865, n57866,
         n57867, n57868, n57869, n57870, n57871, n57872, n57873, n57874,
         n57875, n57876, n57877, n57878, n57879, n57880, n57881, n57882,
         n57883, n57884, n57885, n57886, n57887, n57888, n57889, n57890,
         n57891, n57892, n57893, n57894, n57895, n57896, n57897, n57898,
         n57899, n57900, n57901, n57902, n57903, n57904, n57905, n57906,
         n57907, n57908, n57909, n57910, n57911, n57912, n57913, n57914,
         n57915, n57916, n57917, n57918, n57919, n57920, n57921, n57922,
         n57923, n57924, n57925, n57926, n57927, n57928, n57929, n57930,
         n57931, n57932, n57933, n57934, n57935, n57936, n57937, n57938,
         n57939, n57940, n57941, n57942, n57943, n57944, n57945, n57946,
         n57947, n57948, n57949, n57950, n57951, n57952, n57953, n57954,
         n57955, n57956, n57957, n57958, n57959, n57960, n57961, n57962,
         n57963, n57964, n57965, n57966, n57967, n57968, n57969, n57970,
         n57971, n57972, n57973, n57974, n57975, n57976, n57977, n57978,
         n57979, n57980, n57981, n57982, n57983, n57984, n57985, n57986,
         n57987, n57988, n57989, n57990, n57991, n57992, n57993, n57994,
         n57995, n57996, n57997, n57998, n57999, n58000, n58001, n58002,
         n58003, n58004, n58005, n58006, n58007, n58008, n58009, n58010,
         n58011, n58012, n58013, n58014, n58015, n58016, n58017, n58018,
         n58019, n58020, n58021, n58022, n58023, n58024, n58025, n58026,
         n58027, n58028, n58029, n58030, n58031, n58032, n58033, n58034,
         n58035, n58036, n58037, n58038, n58039, n58040, n58041, n58042,
         n58043, n58044, n58045, n58046, n58047, n58048, n58049, n58050,
         n58051, n58052, n58053, n58054, n58055, n58056, n58057, n58058,
         n58059, n58060, n58061, n58062, n58063, n58064, n58065, n58066,
         n58067, n58068, n58069, n58070, n58071, n58072, n58073, n58074,
         n58075, n58076, n58077, n58078, n58079, n58080, n58081, n58082,
         n58083, n58084, n58085, n58086, n58087, n58088, n58089, n58090,
         n58091, n58092, n58093, n58094, n58095, n58096, n58097, n58098,
         n58099, n58100, n58101, n58102, n58103, n58104, n58105, n58106,
         n58107, n58108, n58109, n58110, n58111, n58112, n58113, n58114,
         n58115, n58116, n58117, n58118, n58119, n58120, n58121, n58122,
         n58123, n58124, n58125, n58126, n58127, n58128, n58129, n58130,
         n58131, n58132, n58133, n58134, n58135, n58136, n58137, n58138,
         n58139, n58140, n58141, n58142, n58143, n58144, n58145, n58146,
         n58147, n58148, n58149, n58150, n58151, n58152, n58153, n58154,
         n58155, n58156, n58157, n58158, n58159, n58160, n58161, n58162,
         n58163, n58164, n58165, n58166, n58167, n58168, n58169, n58170,
         n58171, n58172, n58173, n58174, n58175, n58176, n58177, n58178,
         n58179, n58180, n58181, n58182, n58183, n58184, n58185, n58186,
         n58187, n58188, n58189, n58190, n58191, n58192, n58193, n58194,
         n58195, n58196, n58197, n58198, n58199, n58200, n58201, n58202,
         n58203, n58204, n58205, n58206, n58207, n58208, n58209, n58210,
         n58211, n58212, n58213, n58214, n58215, n58216, n58217, n58218,
         n58219, n58220, n58221, n58222, n58223, n58224, n58225, n58226,
         n58227, n58228, n58229, n58230, n58231, n58232, n58233, n58234,
         n58235, n58236, n58237, n58238, n58239, n58240, n58241, n58242,
         n58243, n58244, n58245, n58246, n58247, n58248, n58249, n58250,
         n58251, n58252, n58253, n58254, n58255, n58256, n58257, n58258,
         n58259, n58260, n58261, n58262, n58263, n58264, n58265, n58266,
         n58267, n58268, n58269, n58270, n58271, n58272, n58273, n58274,
         n58275, n58276, n58277, n58278, n58279, n58280, n58281, n58282,
         n58283, n58284, n58285, n58286, n58287, n58288, n58289, n58290,
         n58291, n58292, n58293, n58294, n58295, n58296, n58297, n58298,
         n58299, n58300, n58301, n58302, n58303, n58304, n58305, n58306,
         n58307, n58308, n58309, n58310, n58311, n58312, n58313, n58314,
         n58315, n58316, n58317, n58318, n58319, n58320, n58321, n58322,
         n58323, n58324, n58325, n58326, n58327, n58328, n58329, n58330,
         n58331, n58332, n58333, n58334, n58335, n58336, n58337, n58338,
         n58339, n58340, n58341, n58342, n58343, n58344, n58345, n58346,
         n58347, n58348, n58349, n58350, n58351, n58352, n58353, n58354,
         n58355, n58356, n58357, n58358, n58359, n58360, n58361, n58362,
         n58363, n58364, n58365, n58366, n58367, n58368, n58369, n58370,
         n58371, n58372, n58373, n58374, n58375, n58376, n58377, n58378,
         n58379, n58380, n58381, n58382, n58383, n58384, n58385, n58386,
         n58387, n58388, n58389, n58390, n58391, n58392, n58393, n58394,
         n58395, n58396, n58397, n58398, n58399, n58400, n58401, n58402,
         n58403, n58404, n58405, n58406, n58407, n58408, n58409, n58410,
         n58411, n58412, n58413, n58414, n58415, n58416, n58417, n58418,
         n58419, n58420, n58421, n58422, n58423, n58424, n58425, n58426,
         n58427, n58428, n58429, n58430, n58431, n58432, n58433, n58434,
         n58435, n58436, n58437, n58438, n58439, n58440, n58441, n58442,
         n58443, n58444, n58445, n58446, n58447, n58448, n58449, n58450,
         n58451, n58452, n58453, n58454, n58455, n58456, n58457, n58458,
         n58459, n58460, n58461, n58462, n58463, n58464, n58465, n58466,
         n58467, n58468, n58469, n58470, n58471, n58472, n58473, n58474,
         n58475, n58476, n58477, n58478, n58479, n58480, n58481, n58482,
         n58483, n58484, n58485, n58486, n58487, n58488, n58489, n58490,
         n58491, n58492, n58493, n58494, n58495, n58496, n58497, n58498,
         n58499, n58500, n58501, n58502, n58503, n58504, n58505, n58506,
         n58507, n58508, n58509, n58510, n58511, n58512, n58513, n58514,
         n58515, n58516, n58517, n58518, n58519, n58520, n58521, n58522,
         n58523, n58524, n58525, n58526, n58527, n58528, n58529, n58530,
         n58531, n58532, n58533, n58534, n58535, n58536, n58537, n58538,
         n58539, n58540, n58541, n58542, n58543, n58544, n58545, n58546,
         n58547, n58548, n58549, n58550, n58551, n58552, n58553, n58554,
         n58555, n58556, n58557, n58558, n58559, n58560, n58561, n58562,
         n58563, n58564, n58565, n58566, n58567, n58568, n58569, n58570,
         n58571, n58572, n58573, n58574, n58575, n58576, n58577, n58578,
         n58579, n58580, n58581, n58582, n58583, n58584, n58585, n58586,
         n58587, n58588, n58589, n58590, n58591, n58592, n58593, n58594,
         n58595, n58596, n58597, n58598, n58599, n58600, n58601, n58602,
         n58603, n58604, n58605, n58606, n58607, n58608, n58609, n58610,
         n58611, n58612, n58613, n58614, n58615, n58616, n58617, n58618,
         n58619, n58620, n58621, n58622, n58623, n58624, n58625, n58626,
         n58627, n58628, n58629, n58630, n58631, n58632, n58633, n58634,
         n58635, n58636, n58637, n58638, n58639, n58640, n58641, n58642,
         n58643, n58644, n58645, n58646;

  IV U35632 ( .A(n42713), .Z(n24435) );
  IV U35633 ( .A(n42714), .Z(n24436) );
  NOR U35634 ( .A(n42713), .B(n24436), .Z(n24437) );
  NOR U35635 ( .A(n42714), .B(n24435), .Z(n24438) );
  NOR U35636 ( .A(n42712), .B(n24438), .Z(n24439) );
  NOR U35637 ( .A(n24437), .B(n24439), .Z(n45817) );
  IV U35638 ( .A(n45820), .Z(n24440) );
  IV U35639 ( .A(n45821), .Z(n24441) );
  NOR U35640 ( .A(n45820), .B(n24441), .Z(n24442) );
  NOR U35641 ( .A(n45821), .B(n24440), .Z(n24443) );
  NOR U35642 ( .A(n45819), .B(n24443), .Z(n24444) );
  NOR U35643 ( .A(n24442), .B(n24444), .Z(n24445) );
  NOR U35644 ( .A(n45818), .B(n45817), .Z(n24446) );
  NOR U35645 ( .A(n24446), .B(n24445), .Z(n49365) );
  NOR U35646 ( .A(n49361), .B(n49360), .Z(n24447) );
  NOR U35647 ( .A(n49362), .B(n24447), .Z(n24448) );
  NOR U35648 ( .A(n49364), .B(n49363), .Z(n24449) );
  NOR U35649 ( .A(n49365), .B(n24449), .Z(n24450) );
  NOR U35650 ( .A(n24448), .B(n24450), .Z(n53189) );
  NOR U35651 ( .A(n56271), .B(n56270), .Z(n24451) );
  NOR U35652 ( .A(n56272), .B(n24451), .Z(n24452) );
  NOR U35653 ( .A(n56273), .B(n24452), .Z(n56274) );
  IV U35654 ( .A(n42341), .Z(n24453) );
  NOR U35655 ( .A(n42340), .B(n24453), .Z(n24454) );
  NOR U35656 ( .A(n42341), .B(n45465), .Z(n24455) );
  NOR U35657 ( .A(n42339), .B(n24455), .Z(n24456) );
  NOR U35658 ( .A(n24454), .B(n24456), .Z(n24457) );
  XOR U35659 ( .A(n45466), .B(n24457), .Z(n45450) );
  IV U35660 ( .A(n43353), .Z(n24458) );
  NOR U35661 ( .A(n38724), .B(n24458), .Z(n24459) );
  NOR U35662 ( .A(n42086), .B(n24459), .Z(n24460) );
  XOR U35663 ( .A(n43345), .B(n43343), .Z(n24461) );
  XOR U35664 ( .A(n24462), .B(n24461), .Z(n42075) );
  IV U35665 ( .A(n24460), .Z(n24462) );
  IV U35666 ( .A(n52633), .Z(n24463) );
  NOR U35667 ( .A(n52633), .B(n52634), .Z(n24464) );
  NOR U35668 ( .A(n53757), .B(n24463), .Z(n24465) );
  NOR U35669 ( .A(n52635), .B(n24465), .Z(n24466) );
  NOR U35670 ( .A(n24464), .B(n24466), .Z(n56952) );
  NOR U35671 ( .A(n54169), .B(n54168), .Z(n24467) );
  NOR U35672 ( .A(n54170), .B(n24467), .Z(n24468) );
  IV U35673 ( .A(n24468), .Z(n57530) );
  IV U35674 ( .A(n44879), .Z(n24469) );
  XOR U35675 ( .A(n44880), .B(n24469), .Z(n24470) );
  IV U35676 ( .A(n44878), .Z(n24471) );
  NOR U35677 ( .A(n24470), .B(n24471), .Z(n24472) );
  IV U35678 ( .A(n44880), .Z(n24473) );
  NOR U35679 ( .A(n24473), .B(n24469), .Z(n24474) );
  NOR U35680 ( .A(n24472), .B(n24474), .Z(n48293) );
  IV U35681 ( .A(n51803), .Z(n24475) );
  IV U35682 ( .A(n51804), .Z(n24476) );
  IV U35683 ( .A(n51805), .Z(n24477) );
  XOR U35684 ( .A(n51805), .B(n24475), .Z(n24478) );
  NOR U35685 ( .A(n24478), .B(n24476), .Z(n24479) );
  NOR U35686 ( .A(n24477), .B(n24475), .Z(n24480) );
  NOR U35687 ( .A(n24479), .B(n24480), .Z(n57897) );
  NOR U35688 ( .A(n54585), .B(n54584), .Z(n24481) );
  NOR U35689 ( .A(n54586), .B(n24481), .Z(n24482) );
  IV U35690 ( .A(n24482), .Z(n55139) );
  NOR U35691 ( .A(n51572), .B(n51573), .Z(n24483) );
  NOR U35692 ( .A(n51574), .B(n24483), .Z(n24484) );
  IV U35693 ( .A(n24484), .Z(n58196) );
  NOR U35694 ( .A(n51390), .B(n51389), .Z(n24485) );
  NOR U35695 ( .A(n51391), .B(n24485), .Z(n24486) );
  IV U35696 ( .A(n24486), .Z(n58510) );
  XOR U35697 ( .A(x[1023]), .B(y[1023]), .Z(n24487) );
  IV U35698 ( .A(n24487), .Z(n54929) );
  XOR U35699 ( .A(x[1022]), .B(y[1022]), .Z(n54893) );
  XOR U35700 ( .A(x[1021]), .B(y[1021]), .Z(n51321) );
  XOR U35701 ( .A(x[1020]), .B(y[1020]), .Z(n51312) );
  XOR U35702 ( .A(x[1019]), .B(y[1019]), .Z(n51278) );
  XOR U35703 ( .A(x[1018]), .B(y[1018]), .Z(n51240) );
  XOR U35704 ( .A(x[1017]), .B(y[1017]), .Z(n51224) );
  XOR U35705 ( .A(x[1016]), .B(y[1016]), .Z(n47753) );
  XOR U35706 ( .A(x[1015]), .B(y[1015]), .Z(n47736) );
  XOR U35707 ( .A(x[1014]), .B(y[1014]), .Z(n44408) );
  XOR U35708 ( .A(x[1013]), .B(y[1013]), .Z(n44372) );
  XOR U35709 ( .A(x[1012]), .B(y[1012]), .Z(n44349) );
  XOR U35710 ( .A(x[1011]), .B(y[1011]), .Z(n34426) );
  XOR U35711 ( .A(x[1010]), .B(y[1010]), .Z(n34420) );
  XOR U35712 ( .A(x[1009]), .B(y[1009]), .Z(n34404) );
  XOR U35713 ( .A(x[1008]), .B(y[1008]), .Z(n34399) );
  XOR U35714 ( .A(x[1007]), .B(y[1007]), .Z(n34391) );
  XOR U35715 ( .A(x[1006]), .B(y[1006]), .Z(n34387) );
  XOR U35716 ( .A(x[1005]), .B(y[1005]), .Z(n34373) );
  XOR U35717 ( .A(x[1004]), .B(y[1004]), .Z(n31266) );
  XOR U35718 ( .A(x[1003]), .B(y[1003]), .Z(n31259) );
  XOR U35719 ( .A(x[1002]), .B(y[1002]), .Z(n31250) );
  XOR U35720 ( .A(x[1001]), .B(y[1001]), .Z(n31244) );
  XOR U35721 ( .A(x[1000]), .B(y[1000]), .Z(n28115) );
  XOR U35722 ( .A(x[999]), .B(y[999]), .Z(n24491) );
  XOR U35723 ( .A(x[998]), .B(y[998]), .Z(n28110) );
  XOR U35724 ( .A(x[997]), .B(y[997]), .Z(n28107) );
  XOR U35725 ( .A(x[996]), .B(y[996]), .Z(n28103) );
  XOR U35726 ( .A(x[995]), .B(y[995]), .Z(n28100) );
  XOR U35727 ( .A(x[994]), .B(y[994]), .Z(n24494) );
  XOR U35728 ( .A(x[993]), .B(y[993]), .Z(n28096) );
  XOR U35729 ( .A(x[992]), .B(y[992]), .Z(n28093) );
  XOR U35730 ( .A(x[991]), .B(y[991]), .Z(n28089) );
  XOR U35731 ( .A(x[990]), .B(y[990]), .Z(n28086) );
  XOR U35732 ( .A(x[989]), .B(y[989]), .Z(n24497) );
  XOR U35733 ( .A(x[988]), .B(y[988]), .Z(n28083) );
  XOR U35734 ( .A(x[987]), .B(y[987]), .Z(n28080) );
  XOR U35735 ( .A(x[986]), .B(y[986]), .Z(n28076) );
  XOR U35736 ( .A(x[985]), .B(y[985]), .Z(n28073) );
  XOR U35737 ( .A(x[984]), .B(y[984]), .Z(n24500) );
  XOR U35738 ( .A(x[983]), .B(y[983]), .Z(n24506) );
  XOR U35739 ( .A(x[982]), .B(y[982]), .Z(n24503) );
  XOR U35740 ( .A(x[981]), .B(y[981]), .Z(n24512) );
  XOR U35741 ( .A(x[980]), .B(y[980]), .Z(n24509) );
  XOR U35742 ( .A(x[979]), .B(y[979]), .Z(n24518) );
  XOR U35743 ( .A(x[978]), .B(y[978]), .Z(n24515) );
  XOR U35744 ( .A(x[977]), .B(y[977]), .Z(n28068) );
  XOR U35745 ( .A(x[976]), .B(y[976]), .Z(n28065) );
  XOR U35746 ( .A(x[975]), .B(y[975]), .Z(n24524) );
  XOR U35747 ( .A(x[974]), .B(y[974]), .Z(n24521) );
  XOR U35748 ( .A(x[973]), .B(y[973]), .Z(n24527) );
  XOR U35749 ( .A(x[972]), .B(y[972]), .Z(n24533) );
  XOR U35750 ( .A(x[971]), .B(y[971]), .Z(n24530) );
  XOR U35751 ( .A(x[970]), .B(y[970]), .Z(n24539) );
  XOR U35752 ( .A(x[969]), .B(y[969]), .Z(n24536) );
  XOR U35753 ( .A(x[968]), .B(y[968]), .Z(n24546) );
  XOR U35754 ( .A(x[967]), .B(y[967]), .Z(n24543) );
  XOR U35755 ( .A(x[966]), .B(y[966]), .Z(n24552) );
  XOR U35756 ( .A(x[965]), .B(y[965]), .Z(n24549) );
  XOR U35757 ( .A(x[964]), .B(y[964]), .Z(n24555) );
  XOR U35758 ( .A(x[963]), .B(y[963]), .Z(n24561) );
  XOR U35759 ( .A(x[962]), .B(y[962]), .Z(n24558) );
  XOR U35760 ( .A(x[961]), .B(y[961]), .Z(n24567) );
  XOR U35761 ( .A(x[960]), .B(y[960]), .Z(n24564) );
  XOR U35762 ( .A(x[959]), .B(y[959]), .Z(n28057) );
  XOR U35763 ( .A(x[958]), .B(y[958]), .Z(n28054) );
  XOR U35764 ( .A(x[957]), .B(y[957]), .Z(n24573) );
  XOR U35765 ( .A(x[956]), .B(y[956]), .Z(n24570) );
  XOR U35766 ( .A(x[955]), .B(y[955]), .Z(n28050) );
  XOR U35767 ( .A(x[954]), .B(y[954]), .Z(n28047) );
  XOR U35768 ( .A(x[953]), .B(y[953]), .Z(n24580) );
  XOR U35769 ( .A(x[952]), .B(y[952]), .Z(n24577) );
  XOR U35770 ( .A(x[951]), .B(y[951]), .Z(n24583) );
  XOR U35771 ( .A(x[950]), .B(y[950]), .Z(n24589) );
  XOR U35772 ( .A(x[949]), .B(y[949]), .Z(n24586) );
  XOR U35773 ( .A(x[948]), .B(y[948]), .Z(n24595) );
  XOR U35774 ( .A(x[947]), .B(y[947]), .Z(n24592) );
  XOR U35775 ( .A(x[946]), .B(y[946]), .Z(n24598) );
  XOR U35776 ( .A(x[945]), .B(y[945]), .Z(n24604) );
  XOR U35777 ( .A(x[944]), .B(y[944]), .Z(n24601) );
  XOR U35778 ( .A(x[943]), .B(y[943]), .Z(n24610) );
  XOR U35779 ( .A(x[942]), .B(y[942]), .Z(n24607) );
  XOR U35780 ( .A(x[941]), .B(y[941]), .Z(n24613) );
  XOR U35781 ( .A(x[940]), .B(y[940]), .Z(n28040) );
  XOR U35782 ( .A(x[939]), .B(y[939]), .Z(n28037) );
  XOR U35783 ( .A(x[938]), .B(y[938]), .Z(n28033) );
  XOR U35784 ( .A(x[937]), .B(y[937]), .Z(n28030) );
  XOR U35785 ( .A(x[936]), .B(y[936]), .Z(n28026) );
  XOR U35786 ( .A(x[935]), .B(y[935]), .Z(n28023) );
  XOR U35787 ( .A(x[934]), .B(y[934]), .Z(n24619) );
  XOR U35788 ( .A(x[933]), .B(y[933]), .Z(n24616) );
  XOR U35789 ( .A(x[932]), .B(y[932]), .Z(n24625) );
  XOR U35790 ( .A(x[931]), .B(y[931]), .Z(n24622) );
  XOR U35791 ( .A(x[930]), .B(y[930]), .Z(n24631) );
  XOR U35792 ( .A(x[929]), .B(y[929]), .Z(n24628) );
  XOR U35793 ( .A(x[928]), .B(y[928]), .Z(n24637) );
  XOR U35794 ( .A(x[927]), .B(y[927]), .Z(n24634) );
  XOR U35795 ( .A(x[926]), .B(y[926]), .Z(n28001) );
  XOR U35796 ( .A(x[925]), .B(y[925]), .Z(n24640) );
  XOR U35797 ( .A(x[924]), .B(y[924]), .Z(n28004) );
  XOR U35798 ( .A(x[923]), .B(y[923]), .Z(n27996) );
  XOR U35799 ( .A(x[922]), .B(y[922]), .Z(n27993) );
  XOR U35800 ( .A(x[921]), .B(y[921]), .Z(n24646) );
  XOR U35801 ( .A(x[920]), .B(y[920]), .Z(n24643) );
  XOR U35802 ( .A(x[919]), .B(y[919]), .Z(n27989) );
  XOR U35803 ( .A(x[918]), .B(y[918]), .Z(n27986) );
  XOR U35804 ( .A(x[917]), .B(y[917]), .Z(n24653) );
  XOR U35805 ( .A(x[916]), .B(y[916]), .Z(n24650) );
  XOR U35806 ( .A(x[915]), .B(y[915]), .Z(n24656) );
  XOR U35807 ( .A(x[914]), .B(y[914]), .Z(n24662) );
  XOR U35808 ( .A(x[913]), .B(y[913]), .Z(n24659) );
  XOR U35809 ( .A(x[912]), .B(y[912]), .Z(n24668) );
  XOR U35810 ( .A(x[911]), .B(y[911]), .Z(n24665) );
  XOR U35811 ( .A(x[910]), .B(y[910]), .Z(n24671) );
  XOR U35812 ( .A(x[909]), .B(y[909]), .Z(n27981) );
  XOR U35813 ( .A(x[908]), .B(y[908]), .Z(n27978) );
  XOR U35814 ( .A(x[907]), .B(y[907]), .Z(n24677) );
  XOR U35815 ( .A(x[906]), .B(y[906]), .Z(n24674) );
  XOR U35816 ( .A(x[905]), .B(y[905]), .Z(n24680) );
  XOR U35817 ( .A(x[904]), .B(y[904]), .Z(n27973) );
  XOR U35818 ( .A(x[903]), .B(y[903]), .Z(n27970) );
  XOR U35819 ( .A(x[902]), .B(y[902]), .Z(n24686) );
  XOR U35820 ( .A(x[901]), .B(y[901]), .Z(n24683) );
  XOR U35821 ( .A(x[900]), .B(y[900]), .Z(n24692) );
  XOR U35822 ( .A(x[899]), .B(y[899]), .Z(n24689) );
  XOR U35823 ( .A(x[898]), .B(y[898]), .Z(n27965) );
  XOR U35824 ( .A(x[897]), .B(y[897]), .Z(n27962) );
  XOR U35825 ( .A(x[896]), .B(y[896]), .Z(n24695) );
  XOR U35826 ( .A(x[895]), .B(y[895]), .Z(n27958) );
  XOR U35827 ( .A(x[894]), .B(y[894]), .Z(n27955) );
  XOR U35828 ( .A(x[893]), .B(y[893]), .Z(n24701) );
  XOR U35829 ( .A(x[892]), .B(y[892]), .Z(n24698) );
  XOR U35830 ( .A(x[891]), .B(y[891]), .Z(n24705) );
  XOR U35831 ( .A(x[890]), .B(y[890]), .Z(n27952) );
  XOR U35832 ( .A(x[889]), .B(y[889]), .Z(n27949) );
  XOR U35833 ( .A(x[888]), .B(y[888]), .Z(n24711) );
  XOR U35834 ( .A(x[887]), .B(y[887]), .Z(n24708) );
  XOR U35835 ( .A(x[886]), .B(y[886]), .Z(n27945) );
  XOR U35836 ( .A(x[885]), .B(y[885]), .Z(n27942) );
  XOR U35837 ( .A(x[884]), .B(y[884]), .Z(n24717) );
  XOR U35838 ( .A(x[883]), .B(y[883]), .Z(n24714) );
  XOR U35839 ( .A(x[882]), .B(y[882]), .Z(n27939) );
  XOR U35840 ( .A(x[881]), .B(y[881]), .Z(n27936) );
  XOR U35841 ( .A(x[880]), .B(y[880]), .Z(n24720) );
  XOR U35842 ( .A(x[879]), .B(y[879]), .Z(n27929) );
  XOR U35843 ( .A(x[878]), .B(y[878]), .Z(n24723) );
  XOR U35844 ( .A(x[877]), .B(y[877]), .Z(n24729) );
  XOR U35845 ( .A(x[876]), .B(y[876]), .Z(n24726) );
  XOR U35846 ( .A(x[875]), .B(y[875]), .Z(n24735) );
  XOR U35847 ( .A(x[874]), .B(y[874]), .Z(n24732) );
  XOR U35848 ( .A(x[873]), .B(y[873]), .Z(n24738) );
  XOR U35849 ( .A(x[872]), .B(y[872]), .Z(n24744) );
  XOR U35850 ( .A(x[871]), .B(y[871]), .Z(n24741) );
  XOR U35851 ( .A(x[870]), .B(y[870]), .Z(n24750) );
  XOR U35852 ( .A(x[869]), .B(y[869]), .Z(n24747) );
  XOR U35853 ( .A(x[868]), .B(y[868]), .Z(n24753) );
  XOR U35854 ( .A(x[867]), .B(y[867]), .Z(n24759) );
  XOR U35855 ( .A(x[866]), .B(y[866]), .Z(n24756) );
  XOR U35856 ( .A(x[865]), .B(y[865]), .Z(n24765) );
  XOR U35857 ( .A(x[864]), .B(y[864]), .Z(n24762) );
  XOR U35858 ( .A(x[863]), .B(y[863]), .Z(n27918) );
  XOR U35859 ( .A(x[862]), .B(y[862]), .Z(n27915) );
  XOR U35860 ( .A(x[861]), .B(y[861]), .Z(n24771) );
  XOR U35861 ( .A(x[860]), .B(y[860]), .Z(n24768) );
  XOR U35862 ( .A(x[859]), .B(y[859]), .Z(n24777) );
  XOR U35863 ( .A(x[858]), .B(y[858]), .Z(n24774) );
  XOR U35864 ( .A(x[857]), .B(y[857]), .Z(n24783) );
  XOR U35865 ( .A(x[856]), .B(y[856]), .Z(n24780) );
  XOR U35866 ( .A(x[855]), .B(y[855]), .Z(n24789) );
  XOR U35867 ( .A(x[854]), .B(y[854]), .Z(n24786) );
  XOR U35868 ( .A(x[853]), .B(y[853]), .Z(n27910) );
  XOR U35869 ( .A(x[852]), .B(y[852]), .Z(n27907) );
  XOR U35870 ( .A(x[851]), .B(y[851]), .Z(n24792) );
  XOR U35871 ( .A(x[850]), .B(y[850]), .Z(n27901) );
  XOR U35872 ( .A(x[849]), .B(y[849]), .Z(n24795) );
  XOR U35873 ( .A(x[848]), .B(y[848]), .Z(n27894) );
  XOR U35874 ( .A(x[847]), .B(y[847]), .Z(n27891) );
  XOR U35875 ( .A(x[846]), .B(y[846]), .Z(n24801) );
  XOR U35876 ( .A(x[845]), .B(y[845]), .Z(n24798) );
  XOR U35877 ( .A(x[844]), .B(y[844]), .Z(n24807) );
  XOR U35878 ( .A(x[843]), .B(y[843]), .Z(n24804) );
  XOR U35879 ( .A(x[842]), .B(y[842]), .Z(n27886) );
  XOR U35880 ( .A(x[841]), .B(y[841]), .Z(n27883) );
  XOR U35881 ( .A(x[840]), .B(y[840]), .Z(n27879) );
  XOR U35882 ( .A(x[839]), .B(y[839]), .Z(n27876) );
  XOR U35883 ( .A(x[838]), .B(y[838]), .Z(n27872) );
  XOR U35884 ( .A(x[837]), .B(y[837]), .Z(n27869) );
  XOR U35885 ( .A(x[836]), .B(y[836]), .Z(n27865) );
  XOR U35886 ( .A(x[835]), .B(y[835]), .Z(n27862) );
  XOR U35887 ( .A(x[834]), .B(y[834]), .Z(n27858) );
  XOR U35888 ( .A(x[833]), .B(y[833]), .Z(n27855) );
  XOR U35889 ( .A(x[832]), .B(y[832]), .Z(n27851) );
  XOR U35890 ( .A(x[831]), .B(y[831]), .Z(n27848) );
  XOR U35891 ( .A(x[830]), .B(y[830]), .Z(n24810) );
  XOR U35892 ( .A(x[829]), .B(y[829]), .Z(n24816) );
  XOR U35893 ( .A(x[828]), .B(y[828]), .Z(n24813) );
  XOR U35894 ( .A(x[827]), .B(y[827]), .Z(n27843) );
  XOR U35895 ( .A(x[826]), .B(y[826]), .Z(n27840) );
  XOR U35896 ( .A(x[825]), .B(y[825]), .Z(n27837) );
  XOR U35897 ( .A(x[824]), .B(y[824]), .Z(n27834) );
  XOR U35898 ( .A(x[823]), .B(y[823]), .Z(n27830) );
  XOR U35899 ( .A(x[822]), .B(y[822]), .Z(n27827) );
  XOR U35900 ( .A(x[821]), .B(y[821]), .Z(n24822) );
  XOR U35901 ( .A(x[820]), .B(y[820]), .Z(n24819) );
  XOR U35902 ( .A(x[819]), .B(y[819]), .Z(n27822) );
  XOR U35903 ( .A(x[818]), .B(y[818]), .Z(n27819) );
  XOR U35904 ( .A(x[817]), .B(y[817]), .Z(n27815) );
  XOR U35905 ( .A(x[816]), .B(y[816]), .Z(n27812) );
  XOR U35906 ( .A(x[815]), .B(y[815]), .Z(n27808) );
  XOR U35907 ( .A(x[814]), .B(y[814]), .Z(n27805) );
  XOR U35908 ( .A(x[813]), .B(y[813]), .Z(n24828) );
  XOR U35909 ( .A(x[812]), .B(y[812]), .Z(n24825) );
  XOR U35910 ( .A(x[811]), .B(y[811]), .Z(n27801) );
  XOR U35911 ( .A(x[810]), .B(y[810]), .Z(n27798) );
  XOR U35912 ( .A(x[809]), .B(y[809]), .Z(n24834) );
  XOR U35913 ( .A(x[808]), .B(y[808]), .Z(n24831) );
  XOR U35914 ( .A(x[807]), .B(y[807]), .Z(n27793) );
  XOR U35915 ( .A(x[806]), .B(y[806]), .Z(n27790) );
  XOR U35916 ( .A(x[805]), .B(y[805]), .Z(n24840) );
  XOR U35917 ( .A(x[804]), .B(y[804]), .Z(n24837) );
  XOR U35918 ( .A(x[803]), .B(y[803]), .Z(n27786) );
  XOR U35919 ( .A(x[802]), .B(y[802]), .Z(n27783) );
  XOR U35920 ( .A(x[801]), .B(y[801]), .Z(n27779) );
  XOR U35921 ( .A(x[800]), .B(y[800]), .Z(n27776) );
  XOR U35922 ( .A(x[799]), .B(y[799]), .Z(n24846) );
  XOR U35923 ( .A(x[798]), .B(y[798]), .Z(n24843) );
  XOR U35924 ( .A(x[797]), .B(y[797]), .Z(n24852) );
  XOR U35925 ( .A(x[796]), .B(y[796]), .Z(n24849) );
  XOR U35926 ( .A(x[795]), .B(y[795]), .Z(n24855) );
  XOR U35927 ( .A(x[794]), .B(y[794]), .Z(n24861) );
  XOR U35928 ( .A(x[793]), .B(y[793]), .Z(n24858) );
  XOR U35929 ( .A(x[792]), .B(y[792]), .Z(n24867) );
  XOR U35930 ( .A(x[791]), .B(y[791]), .Z(n24864) );
  XOR U35931 ( .A(x[790]), .B(y[790]), .Z(n27768) );
  XOR U35932 ( .A(x[789]), .B(y[789]), .Z(n27765) );
  XOR U35933 ( .A(x[788]), .B(y[788]), .Z(n24873) );
  XOR U35934 ( .A(x[787]), .B(y[787]), .Z(n24870) );
  XOR U35935 ( .A(x[786]), .B(y[786]), .Z(n27761) );
  XOR U35936 ( .A(x[785]), .B(y[785]), .Z(n27758) );
  XOR U35937 ( .A(x[784]), .B(y[784]), .Z(n24876) );
  XOR U35938 ( .A(x[783]), .B(y[783]), .Z(n27754) );
  XOR U35939 ( .A(x[782]), .B(y[782]), .Z(n27751) );
  XOR U35940 ( .A(x[781]), .B(y[781]), .Z(n27747) );
  XOR U35941 ( .A(x[780]), .B(y[780]), .Z(n27744) );
  XOR U35942 ( .A(x[779]), .B(y[779]), .Z(n24882) );
  XOR U35943 ( .A(x[778]), .B(y[778]), .Z(n24879) );
  XOR U35944 ( .A(x[777]), .B(y[777]), .Z(n24888) );
  XOR U35945 ( .A(x[776]), .B(y[776]), .Z(n24885) );
  XOR U35946 ( .A(x[775]), .B(y[775]), .Z(n24891) );
  XOR U35947 ( .A(x[774]), .B(y[774]), .Z(n27740) );
  XOR U35948 ( .A(x[773]), .B(y[773]), .Z(n27737) );
  XOR U35949 ( .A(x[772]), .B(y[772]), .Z(n24897) );
  XOR U35950 ( .A(x[771]), .B(y[771]), .Z(n24894) );
  XOR U35951 ( .A(x[770]), .B(y[770]), .Z(n24903) );
  XOR U35952 ( .A(x[769]), .B(y[769]), .Z(n24900) );
  XOR U35953 ( .A(x[768]), .B(y[768]), .Z(n24909) );
  XOR U35954 ( .A(x[767]), .B(y[767]), .Z(n24906) );
  XOR U35955 ( .A(x[766]), .B(y[766]), .Z(n24915) );
  XOR U35956 ( .A(x[765]), .B(y[765]), .Z(n24912) );
  XOR U35957 ( .A(x[764]), .B(y[764]), .Z(n27731) );
  XOR U35958 ( .A(x[763]), .B(y[763]), .Z(n27728) );
  XOR U35959 ( .A(x[762]), .B(y[762]), .Z(n24919) );
  XOR U35960 ( .A(x[761]), .B(y[761]), .Z(n27724) );
  XOR U35961 ( .A(x[760]), .B(y[760]), .Z(n27721) );
  XOR U35962 ( .A(x[759]), .B(y[759]), .Z(n27717) );
  XOR U35963 ( .A(x[758]), .B(y[758]), .Z(n27714) );
  XOR U35964 ( .A(x[757]), .B(y[757]), .Z(n24925) );
  XOR U35965 ( .A(x[756]), .B(y[756]), .Z(n24922) );
  XOR U35966 ( .A(x[755]), .B(y[755]), .Z(n27709) );
  XOR U35967 ( .A(x[754]), .B(y[754]), .Z(n27706) );
  XOR U35968 ( .A(x[753]), .B(y[753]), .Z(n24931) );
  XOR U35969 ( .A(x[752]), .B(y[752]), .Z(n24928) );
  XOR U35970 ( .A(x[751]), .B(y[751]), .Z(n24934) );
  XOR U35971 ( .A(x[750]), .B(y[750]), .Z(n27700) );
  XOR U35972 ( .A(x[749]), .B(y[749]), .Z(n27697) );
  XOR U35973 ( .A(x[748]), .B(y[748]), .Z(n24940) );
  XOR U35974 ( .A(x[747]), .B(y[747]), .Z(n24937) );
  XOR U35975 ( .A(x[746]), .B(y[746]), .Z(n27693) );
  XOR U35976 ( .A(x[745]), .B(y[745]), .Z(n27690) );
  XOR U35977 ( .A(x[744]), .B(y[744]), .Z(n24943) );
  XOR U35978 ( .A(x[743]), .B(y[743]), .Z(n24949) );
  XOR U35979 ( .A(x[742]), .B(y[742]), .Z(n24946) );
  XOR U35980 ( .A(x[741]), .B(y[741]), .Z(n24953) );
  XOR U35981 ( .A(x[740]), .B(y[740]), .Z(n27686) );
  XOR U35982 ( .A(x[739]), .B(y[739]), .Z(n27683) );
  XOR U35983 ( .A(x[738]), .B(y[738]), .Z(n24959) );
  XOR U35984 ( .A(x[737]), .B(y[737]), .Z(n24956) );
  XOR U35985 ( .A(x[736]), .B(y[736]), .Z(n24962) );
  XOR U35986 ( .A(x[735]), .B(y[735]), .Z(n27679) );
  XOR U35987 ( .A(x[734]), .B(y[734]), .Z(n27676) );
  XOR U35988 ( .A(x[733]), .B(y[733]), .Z(n24968) );
  XOR U35989 ( .A(x[732]), .B(y[732]), .Z(n24965) );
  XOR U35990 ( .A(x[731]), .B(y[731]), .Z(n24974) );
  XOR U35991 ( .A(x[730]), .B(y[730]), .Z(n24971) );
  XOR U35992 ( .A(x[729]), .B(y[729]), .Z(n24980) );
  XOR U35993 ( .A(x[728]), .B(y[728]), .Z(n24977) );
  XOR U35994 ( .A(x[727]), .B(y[727]), .Z(n24983) );
  XOR U35995 ( .A(x[726]), .B(y[726]), .Z(n27662) );
  XOR U35996 ( .A(x[725]), .B(y[725]), .Z(n24986) );
  XOR U35997 ( .A(x[724]), .B(y[724]), .Z(n27654) );
  XOR U35998 ( .A(x[723]), .B(y[723]), .Z(n24989) );
  XOR U35999 ( .A(x[722]), .B(y[722]), .Z(n24992) );
  XOR U36000 ( .A(x[721]), .B(y[721]), .Z(n24998) );
  XOR U36001 ( .A(x[720]), .B(y[720]), .Z(n24995) );
  XOR U36002 ( .A(x[719]), .B(y[719]), .Z(n27641) );
  XOR U36003 ( .A(x[718]), .B(y[718]), .Z(n27638) );
  XOR U36004 ( .A(x[717]), .B(y[717]), .Z(n25004) );
  XOR U36005 ( .A(x[716]), .B(y[716]), .Z(n25001) );
  XOR U36006 ( .A(x[715]), .B(y[715]), .Z(n27634) );
  XOR U36007 ( .A(x[714]), .B(y[714]), .Z(n27631) );
  XOR U36008 ( .A(x[713]), .B(y[713]), .Z(n27627) );
  XOR U36009 ( .A(x[712]), .B(y[712]), .Z(n27624) );
  XOR U36010 ( .A(x[711]), .B(y[711]), .Z(n25007) );
  XOR U36011 ( .A(x[710]), .B(y[710]), .Z(n27620) );
  XOR U36012 ( .A(x[709]), .B(y[709]), .Z(n27617) );
  XOR U36013 ( .A(x[708]), .B(y[708]), .Z(n25010) );
  XOR U36014 ( .A(x[707]), .B(y[707]), .Z(n25013) );
  XOR U36015 ( .A(x[706]), .B(y[706]), .Z(n27606) );
  XOR U36016 ( .A(x[705]), .B(y[705]), .Z(n25016) );
  XOR U36017 ( .A(x[704]), .B(y[704]), .Z(n27600) );
  XOR U36018 ( .A(x[703]), .B(y[703]), .Z(n27597) );
  XOR U36019 ( .A(x[702]), .B(y[702]), .Z(n25022) );
  XOR U36020 ( .A(x[701]), .B(y[701]), .Z(n25019) );
  XOR U36021 ( .A(x[700]), .B(y[700]), .Z(n25028) );
  XOR U36022 ( .A(x[699]), .B(y[699]), .Z(n25025) );
  XOR U36023 ( .A(x[698]), .B(y[698]), .Z(n27585) );
  XOR U36024 ( .A(x[697]), .B(y[697]), .Z(n25031) );
  XOR U36025 ( .A(x[696]), .B(y[696]), .Z(n27588) );
  XOR U36026 ( .A(x[695]), .B(y[695]), .Z(n27582) );
  XOR U36027 ( .A(x[694]), .B(y[694]), .Z(n27579) );
  XOR U36028 ( .A(x[693]), .B(y[693]), .Z(n25035) );
  XOR U36029 ( .A(x[692]), .B(y[692]), .Z(n27567) );
  XOR U36030 ( .A(x[691]), .B(y[691]), .Z(n27561) );
  XOR U36031 ( .A(x[690]), .B(y[690]), .Z(n27558) );
  XOR U36032 ( .A(x[689]), .B(y[689]), .Z(n27555) );
  XOR U36033 ( .A(x[688]), .B(y[688]), .Z(n27552) );
  XOR U36034 ( .A(x[687]), .B(y[687]), .Z(n27548) );
  XOR U36035 ( .A(x[686]), .B(y[686]), .Z(n27545) );
  XOR U36036 ( .A(x[685]), .B(y[685]), .Z(n25038) );
  XOR U36037 ( .A(x[684]), .B(y[684]), .Z(n27542) );
  XOR U36038 ( .A(x[683]), .B(y[683]), .Z(n27539) );
  XOR U36039 ( .A(x[682]), .B(y[682]), .Z(n27535) );
  XOR U36040 ( .A(x[681]), .B(y[681]), .Z(n27532) );
  XOR U36041 ( .A(x[680]), .B(y[680]), .Z(n25041) );
  XOR U36042 ( .A(x[679]), .B(y[679]), .Z(n27529) );
  XOR U36043 ( .A(x[678]), .B(y[678]), .Z(n27526) );
  XOR U36044 ( .A(x[677]), .B(y[677]), .Z(n27522) );
  XOR U36045 ( .A(x[676]), .B(y[676]), .Z(n27519) );
  XOR U36046 ( .A(x[675]), .B(y[675]), .Z(n25044) );
  XOR U36047 ( .A(x[674]), .B(y[674]), .Z(n27516) );
  XOR U36048 ( .A(x[673]), .B(y[673]), .Z(n27513) );
  XOR U36049 ( .A(x[672]), .B(y[672]), .Z(n27509) );
  XOR U36050 ( .A(x[671]), .B(y[671]), .Z(n27506) );
  XOR U36051 ( .A(x[670]), .B(y[670]), .Z(n25047) );
  XOR U36052 ( .A(x[669]), .B(y[669]), .Z(n27503) );
  XOR U36053 ( .A(x[668]), .B(y[668]), .Z(n27500) );
  XOR U36054 ( .A(x[667]), .B(y[667]), .Z(n27496) );
  XOR U36055 ( .A(x[666]), .B(y[666]), .Z(n27493) );
  XOR U36056 ( .A(x[665]), .B(y[665]), .Z(n25053) );
  XOR U36057 ( .A(x[664]), .B(y[664]), .Z(n25050) );
  XOR U36058 ( .A(x[663]), .B(y[663]), .Z(n25059) );
  XOR U36059 ( .A(x[662]), .B(y[662]), .Z(n25056) );
  XOR U36060 ( .A(x[661]), .B(y[661]), .Z(n27489) );
  XOR U36061 ( .A(x[660]), .B(y[660]), .Z(n27486) );
  XOR U36062 ( .A(x[659]), .B(y[659]), .Z(n27482) );
  XOR U36063 ( .A(x[658]), .B(y[658]), .Z(n27479) );
  XOR U36064 ( .A(x[657]), .B(y[657]), .Z(n27475) );
  XOR U36065 ( .A(x[656]), .B(y[656]), .Z(n27472) );
  XOR U36066 ( .A(x[655]), .B(y[655]), .Z(n27468) );
  XOR U36067 ( .A(x[654]), .B(y[654]), .Z(n27465) );
  XOR U36068 ( .A(x[653]), .B(y[653]), .Z(n27461) );
  XOR U36069 ( .A(x[652]), .B(y[652]), .Z(n27458) );
  XOR U36070 ( .A(x[651]), .B(y[651]), .Z(n27454) );
  XOR U36071 ( .A(x[650]), .B(y[650]), .Z(n27451) );
  XOR U36072 ( .A(x[649]), .B(y[649]), .Z(n25065) );
  XOR U36073 ( .A(x[648]), .B(y[648]), .Z(n25062) );
  XOR U36074 ( .A(x[647]), .B(y[647]), .Z(n27447) );
  XOR U36075 ( .A(x[646]), .B(y[646]), .Z(n27444) );
  XOR U36076 ( .A(x[645]), .B(y[645]), .Z(n27440) );
  XOR U36077 ( .A(x[644]), .B(y[644]), .Z(n27437) );
  XOR U36078 ( .A(x[643]), .B(y[643]), .Z(n27433) );
  XOR U36079 ( .A(x[642]), .B(y[642]), .Z(n27430) );
  XOR U36080 ( .A(x[641]), .B(y[641]), .Z(n25071) );
  XOR U36081 ( .A(x[640]), .B(y[640]), .Z(n25068) );
  XOR U36082 ( .A(x[639]), .B(y[639]), .Z(n25077) );
  XOR U36083 ( .A(x[638]), .B(y[638]), .Z(n25074) );
  XOR U36084 ( .A(x[637]), .B(y[637]), .Z(n25083) );
  XOR U36085 ( .A(x[636]), .B(y[636]), .Z(n25080) );
  XOR U36086 ( .A(x[635]), .B(y[635]), .Z(n27424) );
  XOR U36087 ( .A(x[634]), .B(y[634]), .Z(n25086) );
  XOR U36088 ( .A(x[633]), .B(y[633]), .Z(n27416) );
  XOR U36089 ( .A(x[632]), .B(y[632]), .Z(n27413) );
  XOR U36090 ( .A(x[631]), .B(y[631]), .Z(n27409) );
  XOR U36091 ( .A(x[630]), .B(y[630]), .Z(n27406) );
  XOR U36092 ( .A(x[629]), .B(y[629]), .Z(n25092) );
  XOR U36093 ( .A(x[628]), .B(y[628]), .Z(n25089) );
  XOR U36094 ( .A(x[627]), .B(y[627]), .Z(n25098) );
  XOR U36095 ( .A(x[626]), .B(y[626]), .Z(n25095) );
  XOR U36096 ( .A(x[625]), .B(y[625]), .Z(n27402) );
  XOR U36097 ( .A(x[624]), .B(y[624]), .Z(n27399) );
  XOR U36098 ( .A(x[623]), .B(y[623]), .Z(n25105) );
  XOR U36099 ( .A(x[622]), .B(y[622]), .Z(n25102) );
  XOR U36100 ( .A(x[621]), .B(y[621]), .Z(n27394) );
  XOR U36101 ( .A(x[620]), .B(y[620]), .Z(n27391) );
  XOR U36102 ( .A(x[619]), .B(y[619]), .Z(n27387) );
  XOR U36103 ( .A(x[618]), .B(y[618]), .Z(n27384) );
  XOR U36104 ( .A(x[617]), .B(y[617]), .Z(n25111) );
  XOR U36105 ( .A(x[616]), .B(y[616]), .Z(n25108) );
  XOR U36106 ( .A(x[615]), .B(y[615]), .Z(n25117) );
  XOR U36107 ( .A(x[614]), .B(y[614]), .Z(n25114) );
  XOR U36108 ( .A(x[613]), .B(y[613]), .Z(n27372) );
  XOR U36109 ( .A(x[612]), .B(y[612]), .Z(n25120) );
  XOR U36110 ( .A(x[611]), .B(y[611]), .Z(n27375) );
  XOR U36111 ( .A(x[610]), .B(y[610]), .Z(n27369) );
  XOR U36112 ( .A(x[609]), .B(y[609]), .Z(n27366) );
  XOR U36113 ( .A(x[608]), .B(y[608]), .Z(n27355) );
  XOR U36114 ( .A(x[607]), .B(y[607]), .Z(n25124) );
  XOR U36115 ( .A(x[606]), .B(y[606]), .Z(n27358) );
  XOR U36116 ( .A(x[605]), .B(y[605]), .Z(n27352) );
  XOR U36117 ( .A(x[604]), .B(y[604]), .Z(n27349) );
  XOR U36118 ( .A(x[603]), .B(y[603]), .Z(n25131) );
  XOR U36119 ( .A(x[602]), .B(y[602]), .Z(n25128) );
  XOR U36120 ( .A(x[601]), .B(y[601]), .Z(n27346) );
  XOR U36121 ( .A(x[600]), .B(y[600]), .Z(n27343) );
  XOR U36122 ( .A(x[599]), .B(y[599]), .Z(n25137) );
  XOR U36123 ( .A(x[598]), .B(y[598]), .Z(n25134) );
  XOR U36124 ( .A(x[597]), .B(y[597]), .Z(n25143) );
  XOR U36125 ( .A(x[596]), .B(y[596]), .Z(n25140) );
  XOR U36126 ( .A(x[595]), .B(y[595]), .Z(n27338) );
  XOR U36127 ( .A(x[594]), .B(y[594]), .Z(n27335) );
  XOR U36128 ( .A(x[593]), .B(y[593]), .Z(n25149) );
  XOR U36129 ( .A(x[592]), .B(y[592]), .Z(n25146) );
  XOR U36130 ( .A(x[591]), .B(y[591]), .Z(n25155) );
  XOR U36131 ( .A(x[590]), .B(y[590]), .Z(n25152) );
  XOR U36132 ( .A(x[589]), .B(y[589]), .Z(n25158) );
  XOR U36133 ( .A(x[588]), .B(y[588]), .Z(n27329) );
  XOR U36134 ( .A(x[587]), .B(y[587]), .Z(n27326) );
  XOR U36135 ( .A(x[586]), .B(y[586]), .Z(n25164) );
  XOR U36136 ( .A(x[585]), .B(y[585]), .Z(n25161) );
  XOR U36137 ( .A(x[584]), .B(y[584]), .Z(n25167) );
  XOR U36138 ( .A(x[583]), .B(y[583]), .Z(n25173) );
  XOR U36139 ( .A(x[582]), .B(y[582]), .Z(n25170) );
  XOR U36140 ( .A(x[581]), .B(y[581]), .Z(n27320) );
  XOR U36141 ( .A(x[580]), .B(y[580]), .Z(n27317) );
  XOR U36142 ( .A(x[579]), .B(y[579]), .Z(n25176) );
  XOR U36143 ( .A(x[578]), .B(y[578]), .Z(n27305) );
  XOR U36144 ( .A(x[577]), .B(y[577]), .Z(n25179) );
  XOR U36145 ( .A(x[576]), .B(y[576]), .Z(n27301) );
  XOR U36146 ( .A(x[575]), .B(y[575]), .Z(n27298) );
  XOR U36147 ( .A(x[574]), .B(y[574]), .Z(n25182) );
  XOR U36148 ( .A(x[573]), .B(y[573]), .Z(n27291) );
  XOR U36149 ( .A(x[572]), .B(y[572]), .Z(n25185) );
  XOR U36150 ( .A(x[571]), .B(y[571]), .Z(n27285) );
  XOR U36151 ( .A(x[570]), .B(y[570]), .Z(n27282) );
  XOR U36152 ( .A(x[569]), .B(y[569]), .Z(n25191) );
  XOR U36153 ( .A(x[568]), .B(y[568]), .Z(n25188) );
  XOR U36154 ( .A(x[567]), .B(y[567]), .Z(n25197) );
  XOR U36155 ( .A(x[566]), .B(y[566]), .Z(n25194) );
  XOR U36156 ( .A(x[565]), .B(y[565]), .Z(n25203) );
  XOR U36157 ( .A(x[564]), .B(y[564]), .Z(n25200) );
  XOR U36158 ( .A(x[563]), .B(y[563]), .Z(n25206) );
  XOR U36159 ( .A(x[562]), .B(y[562]), .Z(n25212) );
  XOR U36160 ( .A(x[561]), .B(y[561]), .Z(n25209) );
  XOR U36161 ( .A(x[560]), .B(y[560]), .Z(n27275) );
  XOR U36162 ( .A(x[559]), .B(y[559]), .Z(n27272) );
  XOR U36163 ( .A(x[558]), .B(y[558]), .Z(n27268) );
  XOR U36164 ( .A(x[557]), .B(y[557]), .Z(n27265) );
  XOR U36165 ( .A(x[556]), .B(y[556]), .Z(n27261) );
  XOR U36166 ( .A(x[555]), .B(y[555]), .Z(n27258) );
  XOR U36167 ( .A(x[554]), .B(y[554]), .Z(n27254) );
  XOR U36168 ( .A(x[553]), .B(y[553]), .Z(n27251) );
  XOR U36169 ( .A(x[552]), .B(y[552]), .Z(n25215) );
  XOR U36170 ( .A(x[551]), .B(y[551]), .Z(n25221) );
  XOR U36171 ( .A(x[550]), .B(y[550]), .Z(n25218) );
  XOR U36172 ( .A(x[549]), .B(y[549]), .Z(n27246) );
  XOR U36173 ( .A(x[548]), .B(y[548]), .Z(n27243) );
  XOR U36174 ( .A(x[547]), .B(y[547]), .Z(n25228) );
  XOR U36175 ( .A(x[546]), .B(y[546]), .Z(n25225) );
  XOR U36176 ( .A(x[545]), .B(y[545]), .Z(n27239) );
  XOR U36177 ( .A(x[544]), .B(y[544]), .Z(n27236) );
  XOR U36178 ( .A(x[543]), .B(y[543]), .Z(n27232) );
  XOR U36179 ( .A(x[542]), .B(y[542]), .Z(n27229) );
  XOR U36180 ( .A(x[541]), .B(y[541]), .Z(n25231) );
  XOR U36181 ( .A(x[540]), .B(y[540]), .Z(n27217) );
  XOR U36182 ( .A(x[539]), .B(y[539]), .Z(n25234) );
  XOR U36183 ( .A(x[538]), .B(y[538]), .Z(n27220) );
  XOR U36184 ( .A(x[537]), .B(y[537]), .Z(n25238) );
  XOR U36185 ( .A(x[536]), .B(y[536]), .Z(n27211) );
  XOR U36186 ( .A(x[535]), .B(y[535]), .Z(n27208) );
  XOR U36187 ( .A(x[534]), .B(y[534]), .Z(n25244) );
  XOR U36188 ( .A(x[533]), .B(y[533]), .Z(n25241) );
  XOR U36189 ( .A(x[532]), .B(y[532]), .Z(n25250) );
  XOR U36190 ( .A(x[531]), .B(y[531]), .Z(n25247) );
  XOR U36191 ( .A(x[530]), .B(y[530]), .Z(n27203) );
  XOR U36192 ( .A(x[529]), .B(y[529]), .Z(n27200) );
  XOR U36193 ( .A(x[528]), .B(y[528]), .Z(n25256) );
  XOR U36194 ( .A(x[527]), .B(y[527]), .Z(n25253) );
  XOR U36195 ( .A(x[526]), .B(y[526]), .Z(n27196) );
  XOR U36196 ( .A(x[525]), .B(y[525]), .Z(n27193) );
  XOR U36197 ( .A(x[524]), .B(y[524]), .Z(n27189) );
  XOR U36198 ( .A(x[523]), .B(y[523]), .Z(n27186) );
  XOR U36199 ( .A(x[522]), .B(y[522]), .Z(n25259) );
  XOR U36200 ( .A(x[521]), .B(y[521]), .Z(n27182) );
  XOR U36201 ( .A(x[520]), .B(y[520]), .Z(n27179) );
  XOR U36202 ( .A(x[519]), .B(y[519]), .Z(n27175) );
  XOR U36203 ( .A(x[518]), .B(y[518]), .Z(n27172) );
  XOR U36204 ( .A(x[517]), .B(y[517]), .Z(n25262) );
  XOR U36205 ( .A(x[516]), .B(y[516]), .Z(n25268) );
  XOR U36206 ( .A(x[515]), .B(y[515]), .Z(n25265) );
  XOR U36207 ( .A(x[514]), .B(y[514]), .Z(n25272) );
  XOR U36208 ( .A(x[513]), .B(y[513]), .Z(n27167) );
  XOR U36209 ( .A(x[512]), .B(y[512]), .Z(n27164) );
  XOR U36210 ( .A(x[511]), .B(y[511]), .Z(n25278) );
  XOR U36211 ( .A(x[510]), .B(y[510]), .Z(n25275) );
  XOR U36212 ( .A(x[509]), .B(y[509]), .Z(n27152) );
  XOR U36213 ( .A(x[508]), .B(y[508]), .Z(n25281) );
  XOR U36214 ( .A(x[507]), .B(y[507]), .Z(n27155) );
  XOR U36215 ( .A(x[506]), .B(y[506]), .Z(n25288) );
  XOR U36216 ( .A(x[505]), .B(y[505]), .Z(n25285) );
  XOR U36217 ( .A(x[504]), .B(y[504]), .Z(n27148) );
  XOR U36218 ( .A(x[503]), .B(y[503]), .Z(n27145) );
  XOR U36219 ( .A(x[502]), .B(y[502]), .Z(n27141) );
  XOR U36220 ( .A(x[501]), .B(y[501]), .Z(n27138) );
  XOR U36221 ( .A(x[500]), .B(y[500]), .Z(n27134) );
  XOR U36222 ( .A(x[499]), .B(y[499]), .Z(n27131) );
  XOR U36223 ( .A(x[498]), .B(y[498]), .Z(n27127) );
  XOR U36224 ( .A(x[497]), .B(y[497]), .Z(n27124) );
  XOR U36225 ( .A(x[496]), .B(y[496]), .Z(n25295) );
  XOR U36226 ( .A(x[495]), .B(y[495]), .Z(n25292) );
  XOR U36227 ( .A(x[494]), .B(y[494]), .Z(n27119) );
  XOR U36228 ( .A(x[493]), .B(y[493]), .Z(n27116) );
  XOR U36229 ( .A(x[492]), .B(y[492]), .Z(n25301) );
  XOR U36230 ( .A(x[491]), .B(y[491]), .Z(n25298) );
  XOR U36231 ( .A(x[490]), .B(y[490]), .Z(n27111) );
  XOR U36232 ( .A(x[489]), .B(y[489]), .Z(n27108) );
  XOR U36233 ( .A(x[488]), .B(y[488]), .Z(n25307) );
  XOR U36234 ( .A(x[487]), .B(y[487]), .Z(n25304) );
  XOR U36235 ( .A(x[486]), .B(y[486]), .Z(n27104) );
  XOR U36236 ( .A(x[485]), .B(y[485]), .Z(n27101) );
  XOR U36237 ( .A(x[484]), .B(y[484]), .Z(n25313) );
  XOR U36238 ( .A(x[483]), .B(y[483]), .Z(n25310) );
  XOR U36239 ( .A(x[482]), .B(y[482]), .Z(n25316) );
  XOR U36240 ( .A(x[481]), .B(y[481]), .Z(n27089) );
  XOR U36241 ( .A(x[480]), .B(y[480]), .Z(n27086) );
  XOR U36242 ( .A(x[479]), .B(y[479]), .Z(n27082) );
  XOR U36243 ( .A(x[478]), .B(y[478]), .Z(n27079) );
  XOR U36244 ( .A(x[477]), .B(y[477]), .Z(n25323) );
  XOR U36245 ( .A(x[476]), .B(y[476]), .Z(n25320) );
  XOR U36246 ( .A(x[475]), .B(y[475]), .Z(n25326) );
  XOR U36247 ( .A(x[474]), .B(y[474]), .Z(n25329) );
  XOR U36248 ( .A(x[473]), .B(y[473]), .Z(n27064) );
  XOR U36249 ( .A(x[472]), .B(y[472]), .Z(n25332) );
  XOR U36250 ( .A(x[471]), .B(y[471]), .Z(n25338) );
  XOR U36251 ( .A(x[470]), .B(y[470]), .Z(n25335) );
  XOR U36252 ( .A(x[469]), .B(y[469]), .Z(n25344) );
  XOR U36253 ( .A(x[468]), .B(y[468]), .Z(n25341) );
  XOR U36254 ( .A(x[467]), .B(y[467]), .Z(n25347) );
  XOR U36255 ( .A(x[466]), .B(y[466]), .Z(n27055) );
  XOR U36256 ( .A(x[465]), .B(y[465]), .Z(n25350) );
  XOR U36257 ( .A(x[464]), .B(y[464]), .Z(n27049) );
  XOR U36258 ( .A(x[463]), .B(y[463]), .Z(n27046) );
  XOR U36259 ( .A(x[462]), .B(y[462]), .Z(n25356) );
  XOR U36260 ( .A(x[461]), .B(y[461]), .Z(n25353) );
  XOR U36261 ( .A(x[460]), .B(y[460]), .Z(n25362) );
  XOR U36262 ( .A(x[459]), .B(y[459]), .Z(n25359) );
  XOR U36263 ( .A(x[458]), .B(y[458]), .Z(n25368) );
  XOR U36264 ( .A(x[457]), .B(y[457]), .Z(n25365) );
  XOR U36265 ( .A(x[456]), .B(y[456]), .Z(n27040) );
  XOR U36266 ( .A(x[455]), .B(y[455]), .Z(n27037) );
  XOR U36267 ( .A(x[454]), .B(y[454]), .Z(n27033) );
  XOR U36268 ( .A(x[453]), .B(y[453]), .Z(n27030) );
  XOR U36269 ( .A(x[452]), .B(y[452]), .Z(n27026) );
  XOR U36270 ( .A(x[451]), .B(y[451]), .Z(n27023) );
  XOR U36271 ( .A(x[450]), .B(y[450]), .Z(n25374) );
  XOR U36272 ( .A(x[449]), .B(y[449]), .Z(n25371) );
  XOR U36273 ( .A(x[448]), .B(y[448]), .Z(n25377) );
  XOR U36274 ( .A(x[447]), .B(y[447]), .Z(n27009) );
  XOR U36275 ( .A(x[446]), .B(y[446]), .Z(n25380) );
  XOR U36276 ( .A(x[445]), .B(y[445]), .Z(n26995) );
  XOR U36277 ( .A(x[444]), .B(y[444]), .Z(n26990) );
  XOR U36278 ( .A(x[443]), .B(y[443]), .Z(n26987) );
  XOR U36279 ( .A(x[442]), .B(y[442]), .Z(n25386) );
  XOR U36280 ( .A(x[441]), .B(y[441]), .Z(n25383) );
  XOR U36281 ( .A(x[440]), .B(y[440]), .Z(n25392) );
  XOR U36282 ( .A(x[439]), .B(y[439]), .Z(n25389) );
  XOR U36283 ( .A(x[438]), .B(y[438]), .Z(n26982) );
  XOR U36284 ( .A(x[437]), .B(y[437]), .Z(n26979) );
  XOR U36285 ( .A(x[436]), .B(y[436]), .Z(n26975) );
  XOR U36286 ( .A(x[435]), .B(y[435]), .Z(n26972) );
  XOR U36287 ( .A(x[434]), .B(y[434]), .Z(n26968) );
  XOR U36288 ( .A(x[433]), .B(y[433]), .Z(n26965) );
  XOR U36289 ( .A(x[432]), .B(y[432]), .Z(n25395) );
  XOR U36290 ( .A(x[431]), .B(y[431]), .Z(n26953) );
  XOR U36291 ( .A(x[430]), .B(y[430]), .Z(n25398) );
  XOR U36292 ( .A(x[429]), .B(y[429]), .Z(n26956) );
  XOR U36293 ( .A(x[428]), .B(y[428]), .Z(n26949) );
  XOR U36294 ( .A(x[427]), .B(y[427]), .Z(n26946) );
  XOR U36295 ( .A(x[426]), .B(y[426]), .Z(n25405) );
  XOR U36296 ( .A(x[425]), .B(y[425]), .Z(n25402) );
  XOR U36297 ( .A(x[424]), .B(y[424]), .Z(n26942) );
  XOR U36298 ( .A(x[423]), .B(y[423]), .Z(n26939) );
  XOR U36299 ( .A(x[422]), .B(y[422]), .Z(n25411) );
  XOR U36300 ( .A(x[421]), .B(y[421]), .Z(n25408) );
  XOR U36301 ( .A(x[420]), .B(y[420]), .Z(n25414) );
  XOR U36302 ( .A(x[419]), .B(y[419]), .Z(n26929) );
  XOR U36303 ( .A(x[418]), .B(y[418]), .Z(n26926) );
  XOR U36304 ( .A(x[417]), .B(y[417]), .Z(n26922) );
  XOR U36305 ( .A(x[416]), .B(y[416]), .Z(n26919) );
  XOR U36306 ( .A(x[415]), .B(y[415]), .Z(n25417) );
  XOR U36307 ( .A(x[414]), .B(y[414]), .Z(n26907) );
  XOR U36308 ( .A(x[413]), .B(y[413]), .Z(n25423) );
  XOR U36309 ( .A(x[412]), .B(y[412]), .Z(n25420) );
  XOR U36310 ( .A(x[411]), .B(y[411]), .Z(n26901) );
  XOR U36311 ( .A(x[410]), .B(y[410]), .Z(n26898) );
  XOR U36312 ( .A(x[409]), .B(y[409]), .Z(n25426) );
  XOR U36313 ( .A(x[408]), .B(y[408]), .Z(n25429) );
  XOR U36314 ( .A(x[407]), .B(y[407]), .Z(n26884) );
  XOR U36315 ( .A(x[406]), .B(y[406]), .Z(n25432) );
  XOR U36316 ( .A(x[405]), .B(y[405]), .Z(n25435) );
  XOR U36317 ( .A(x[404]), .B(y[404]), .Z(n25441) );
  XOR U36318 ( .A(x[403]), .B(y[403]), .Z(n25438) );
  XOR U36319 ( .A(x[402]), .B(y[402]), .Z(n25447) );
  XOR U36320 ( .A(x[401]), .B(y[401]), .Z(n25444) );
  XOR U36321 ( .A(x[400]), .B(y[400]), .Z(n25450) );
  XOR U36322 ( .A(x[399]), .B(y[399]), .Z(n26878) );
  XOR U36323 ( .A(x[398]), .B(y[398]), .Z(n26875) );
  XOR U36324 ( .A(x[397]), .B(y[397]), .Z(n25456) );
  XOR U36325 ( .A(x[396]), .B(y[396]), .Z(n25453) );
  XOR U36326 ( .A(x[395]), .B(y[395]), .Z(n25462) );
  XOR U36327 ( .A(x[394]), .B(y[394]), .Z(n25459) );
  XOR U36328 ( .A(x[393]), .B(y[393]), .Z(n26871) );
  XOR U36329 ( .A(x[392]), .B(y[392]), .Z(n26868) );
  XOR U36330 ( .A(x[391]), .B(y[391]), .Z(n26864) );
  XOR U36331 ( .A(x[390]), .B(y[390]), .Z(n26861) );
  XOR U36332 ( .A(x[389]), .B(y[389]), .Z(n26858) );
  XOR U36333 ( .A(x[388]), .B(y[388]), .Z(n26855) );
  XOR U36334 ( .A(x[387]), .B(y[387]), .Z(n26851) );
  XOR U36335 ( .A(x[386]), .B(y[386]), .Z(n26848) );
  XOR U36336 ( .A(x[385]), .B(y[385]), .Z(n25465) );
  XOR U36337 ( .A(x[384]), .B(y[384]), .Z(n26844) );
  XOR U36338 ( .A(x[383]), .B(y[383]), .Z(n26841) );
  XOR U36339 ( .A(x[382]), .B(y[382]), .Z(n26837) );
  XOR U36340 ( .A(x[381]), .B(y[381]), .Z(n26834) );
  XOR U36341 ( .A(x[380]), .B(y[380]), .Z(n25468) );
  XOR U36342 ( .A(x[379]), .B(y[379]), .Z(n25474) );
  XOR U36343 ( .A(x[378]), .B(y[378]), .Z(n25471) );
  XOR U36344 ( .A(x[377]), .B(y[377]), .Z(n26830) );
  XOR U36345 ( .A(x[376]), .B(y[376]), .Z(n26827) );
  XOR U36346 ( .A(x[375]), .B(y[375]), .Z(n26824) );
  XOR U36347 ( .A(x[374]), .B(y[374]), .Z(n26821) );
  XOR U36348 ( .A(x[373]), .B(y[373]), .Z(n26817) );
  XOR U36349 ( .A(x[372]), .B(y[372]), .Z(n26814) );
  XOR U36350 ( .A(x[371]), .B(y[371]), .Z(n36821) );
  XOR U36351 ( .A(x[370]), .B(y[370]), .Z(n25478) );
  IV U36352 ( .A(x[369]), .Z(n24488) );
  XOR U36353 ( .A(n24488), .B(y[369]), .Z(n25487) );
  XOR U36354 ( .A(x[368]), .B(y[368]), .Z(n25483) );
  XOR U36355 ( .A(x[367]), .B(y[367]), .Z(n25489) );
  XOR U36356 ( .A(x[366]), .B(y[366]), .Z(n25495) );
  XOR U36357 ( .A(x[365]), .B(y[365]), .Z(n25492) );
  XOR U36358 ( .A(x[364]), .B(y[364]), .Z(n26809) );
  XOR U36359 ( .A(x[363]), .B(y[363]), .Z(n26806) );
  XOR U36360 ( .A(x[362]), .B(y[362]), .Z(n25498) );
  XOR U36361 ( .A(x[361]), .B(y[361]), .Z(n26802) );
  XOR U36362 ( .A(x[360]), .B(y[360]), .Z(n26799) );
  XOR U36363 ( .A(x[359]), .B(y[359]), .Z(n26785) );
  XOR U36364 ( .A(x[358]), .B(y[358]), .Z(n26782) );
  XOR U36365 ( .A(x[357]), .B(y[357]), .Z(n25504) );
  XOR U36366 ( .A(x[356]), .B(y[356]), .Z(n25501) );
  XOR U36367 ( .A(x[355]), .B(y[355]), .Z(n26778) );
  XOR U36368 ( .A(x[354]), .B(y[354]), .Z(n26775) );
  XOR U36369 ( .A(x[353]), .B(y[353]), .Z(n25510) );
  XOR U36370 ( .A(x[352]), .B(y[352]), .Z(n25507) );
  XOR U36371 ( .A(x[351]), .B(y[351]), .Z(n26771) );
  XOR U36372 ( .A(x[350]), .B(y[350]), .Z(n26768) );
  XOR U36373 ( .A(x[349]), .B(y[349]), .Z(n25517) );
  XOR U36374 ( .A(x[348]), .B(y[348]), .Z(n25514) );
  XOR U36375 ( .A(x[347]), .B(y[347]), .Z(n25523) );
  XOR U36376 ( .A(x[346]), .B(y[346]), .Z(n25520) );
  XOR U36377 ( .A(x[345]), .B(y[345]), .Z(n25529) );
  XOR U36378 ( .A(x[344]), .B(y[344]), .Z(n25526) );
  XOR U36379 ( .A(x[343]), .B(y[343]), .Z(n25532) );
  XOR U36380 ( .A(x[342]), .B(y[342]), .Z(n26762) );
  XOR U36381 ( .A(x[341]), .B(y[341]), .Z(n26759) );
  XOR U36382 ( .A(x[340]), .B(y[340]), .Z(n26755) );
  XOR U36383 ( .A(x[339]), .B(y[339]), .Z(n26752) );
  XOR U36384 ( .A(x[338]), .B(y[338]), .Z(n26748) );
  XOR U36385 ( .A(x[337]), .B(y[337]), .Z(n26745) );
  XOR U36386 ( .A(x[336]), .B(y[336]), .Z(n25535) );
  XOR U36387 ( .A(x[335]), .B(y[335]), .Z(n25541) );
  XOR U36388 ( .A(x[334]), .B(y[334]), .Z(n25538) );
  XOR U36389 ( .A(x[333]), .B(y[333]), .Z(n25547) );
  XOR U36390 ( .A(x[332]), .B(y[332]), .Z(n25544) );
  XOR U36391 ( .A(x[331]), .B(y[331]), .Z(n25554) );
  XOR U36392 ( .A(x[330]), .B(y[330]), .Z(n25551) );
  XOR U36393 ( .A(x[329]), .B(y[329]), .Z(n25560) );
  XOR U36394 ( .A(x[328]), .B(y[328]), .Z(n25557) );
  XOR U36395 ( .A(x[327]), .B(y[327]), .Z(n25566) );
  XOR U36396 ( .A(x[326]), .B(y[326]), .Z(n25563) );
  XOR U36397 ( .A(x[325]), .B(y[325]), .Z(n25572) );
  XOR U36398 ( .A(x[324]), .B(y[324]), .Z(n25569) );
  XOR U36399 ( .A(x[323]), .B(y[323]), .Z(n25578) );
  XOR U36400 ( .A(x[322]), .B(y[322]), .Z(n25575) );
  XOR U36401 ( .A(x[321]), .B(y[321]), .Z(n26725) );
  XOR U36402 ( .A(x[320]), .B(y[320]), .Z(n25581) );
  XOR U36403 ( .A(x[319]), .B(y[319]), .Z(n26728) );
  XOR U36404 ( .A(x[318]), .B(y[318]), .Z(n25585) );
  XOR U36405 ( .A(x[317]), .B(y[317]), .Z(n25591) );
  XOR U36406 ( .A(x[316]), .B(y[316]), .Z(n25588) );
  XOR U36407 ( .A(x[315]), .B(y[315]), .Z(n25597) );
  XOR U36408 ( .A(x[314]), .B(y[314]), .Z(n25594) );
  XOR U36409 ( .A(x[313]), .B(y[313]), .Z(n25603) );
  XOR U36410 ( .A(x[312]), .B(y[312]), .Z(n25600) );
  XOR U36411 ( .A(x[311]), .B(y[311]), .Z(n25606) );
  XOR U36412 ( .A(x[310]), .B(y[310]), .Z(n25612) );
  XOR U36413 ( .A(x[309]), .B(y[309]), .Z(n25609) );
  XOR U36414 ( .A(x[308]), .B(y[308]), .Z(n25618) );
  XOR U36415 ( .A(x[307]), .B(y[307]), .Z(n25615) );
  XOR U36416 ( .A(x[306]), .B(y[306]), .Z(n25621) );
  XOR U36417 ( .A(x[305]), .B(y[305]), .Z(n25627) );
  XOR U36418 ( .A(x[304]), .B(y[304]), .Z(n25624) );
  XOR U36419 ( .A(x[303]), .B(y[303]), .Z(n25633) );
  XOR U36420 ( .A(x[302]), .B(y[302]), .Z(n25630) );
  XOR U36421 ( .A(x[301]), .B(y[301]), .Z(n25636) );
  XOR U36422 ( .A(x[300]), .B(y[300]), .Z(n26710) );
  XOR U36423 ( .A(x[299]), .B(y[299]), .Z(n26707) );
  XOR U36424 ( .A(x[298]), .B(y[298]), .Z(n26703) );
  XOR U36425 ( .A(x[297]), .B(y[297]), .Z(n26700) );
  XOR U36426 ( .A(x[296]), .B(y[296]), .Z(n26696) );
  XOR U36427 ( .A(x[295]), .B(y[295]), .Z(n26693) );
  XOR U36428 ( .A(x[294]), .B(y[294]), .Z(n25639) );
  XOR U36429 ( .A(x[293]), .B(y[293]), .Z(n25645) );
  XOR U36430 ( .A(x[292]), .B(y[292]), .Z(n25642) );
  XOR U36431 ( .A(x[291]), .B(y[291]), .Z(n25651) );
  XOR U36432 ( .A(x[290]), .B(y[290]), .Z(n25648) );
  XOR U36433 ( .A(x[289]), .B(y[289]), .Z(n25657) );
  XOR U36434 ( .A(x[288]), .B(y[288]), .Z(n25654) );
  XOR U36435 ( .A(x[287]), .B(y[287]), .Z(n26688) );
  XOR U36436 ( .A(x[286]), .B(y[286]), .Z(n26685) );
  XOR U36437 ( .A(x[285]), .B(y[285]), .Z(n25663) );
  XOR U36438 ( .A(x[284]), .B(y[284]), .Z(n25660) );
  XOR U36439 ( .A(x[283]), .B(y[283]), .Z(n25669) );
  XOR U36440 ( .A(x[282]), .B(y[282]), .Z(n25666) );
  XOR U36441 ( .A(x[281]), .B(y[281]), .Z(n25675) );
  XOR U36442 ( .A(x[280]), .B(y[280]), .Z(n25672) );
  XOR U36443 ( .A(x[279]), .B(y[279]), .Z(n25679) );
  XOR U36444 ( .A(x[278]), .B(y[278]), .Z(n25685) );
  XOR U36445 ( .A(x[277]), .B(y[277]), .Z(n25682) );
  XOR U36446 ( .A(x[276]), .B(y[276]), .Z(n26678) );
  XOR U36447 ( .A(x[275]), .B(y[275]), .Z(n26675) );
  XOR U36448 ( .A(x[274]), .B(y[274]), .Z(n25688) );
  XOR U36449 ( .A(x[273]), .B(y[273]), .Z(n26667) );
  XOR U36450 ( .A(x[272]), .B(y[272]), .Z(n26664) );
  XOR U36451 ( .A(x[271]), .B(y[271]), .Z(n26660) );
  XOR U36452 ( .A(x[270]), .B(y[270]), .Z(n26657) );
  XOR U36453 ( .A(x[269]), .B(y[269]), .Z(n26653) );
  XOR U36454 ( .A(x[268]), .B(y[268]), .Z(n26650) );
  XOR U36455 ( .A(x[267]), .B(y[267]), .Z(n25691) );
  XOR U36456 ( .A(x[266]), .B(y[266]), .Z(n26638) );
  XOR U36457 ( .A(x[265]), .B(y[265]), .Z(n25698) );
  XOR U36458 ( .A(x[264]), .B(y[264]), .Z(n25695) );
  XOR U36459 ( .A(x[263]), .B(y[263]), .Z(n26632) );
  XOR U36460 ( .A(x[262]), .B(y[262]), .Z(n26629) );
  XOR U36461 ( .A(x[261]), .B(y[261]), .Z(n25704) );
  XOR U36462 ( .A(x[260]), .B(y[260]), .Z(n25701) );
  XOR U36463 ( .A(x[259]), .B(y[259]), .Z(n26625) );
  XOR U36464 ( .A(x[258]), .B(y[258]), .Z(n26622) );
  XOR U36465 ( .A(x[257]), .B(y[257]), .Z(n25710) );
  XOR U36466 ( .A(x[256]), .B(y[256]), .Z(n25707) );
  XOR U36467 ( .A(x[255]), .B(y[255]), .Z(n25713) );
  XOR U36468 ( .A(x[254]), .B(y[254]), .Z(n25719) );
  XOR U36469 ( .A(x[253]), .B(y[253]), .Z(n25716) );
  XOR U36470 ( .A(x[252]), .B(y[252]), .Z(n25725) );
  XOR U36471 ( .A(x[251]), .B(y[251]), .Z(n25722) );
  XOR U36472 ( .A(x[250]), .B(y[250]), .Z(n25728) );
  XOR U36473 ( .A(x[249]), .B(y[249]), .Z(n25734) );
  XOR U36474 ( .A(x[248]), .B(y[248]), .Z(n25731) );
  XOR U36475 ( .A(x[247]), .B(y[247]), .Z(n25740) );
  XOR U36476 ( .A(x[246]), .B(y[246]), .Z(n25737) );
  XOR U36477 ( .A(x[245]), .B(y[245]), .Z(n26617) );
  XOR U36478 ( .A(x[244]), .B(y[244]), .Z(n26614) );
  XOR U36479 ( .A(x[243]), .B(y[243]), .Z(n25747) );
  XOR U36480 ( .A(x[242]), .B(y[242]), .Z(n25744) );
  XOR U36481 ( .A(x[241]), .B(y[241]), .Z(n26610) );
  XOR U36482 ( .A(x[240]), .B(y[240]), .Z(n26607) );
  XOR U36483 ( .A(x[239]), .B(y[239]), .Z(n25753) );
  XOR U36484 ( .A(x[238]), .B(y[238]), .Z(n25750) );
  XOR U36485 ( .A(x[237]), .B(y[237]), .Z(n25759) );
  XOR U36486 ( .A(x[236]), .B(y[236]), .Z(n25756) );
  XOR U36487 ( .A(x[235]), .B(y[235]), .Z(n25763) );
  XOR U36488 ( .A(x[234]), .B(y[234]), .Z(n26604) );
  XOR U36489 ( .A(x[233]), .B(y[233]), .Z(n26601) );
  XOR U36490 ( .A(x[232]), .B(y[232]), .Z(n26597) );
  XOR U36491 ( .A(x[231]), .B(y[231]), .Z(n26594) );
  XOR U36492 ( .A(x[230]), .B(y[230]), .Z(n25766) );
  XOR U36493 ( .A(x[229]), .B(y[229]), .Z(n25773) );
  XOR U36494 ( .A(x[228]), .B(y[228]), .Z(n25770) );
  XOR U36495 ( .A(x[227]), .B(y[227]), .Z(n25779) );
  XOR U36496 ( .A(x[226]), .B(y[226]), .Z(n25776) );
  XOR U36497 ( .A(x[225]), .B(y[225]), .Z(n26589) );
  XOR U36498 ( .A(x[224]), .B(y[224]), .Z(n26586) );
  XOR U36499 ( .A(x[223]), .B(y[223]), .Z(n25782) );
  XOR U36500 ( .A(x[222]), .B(y[222]), .Z(n26580) );
  XOR U36501 ( .A(x[221]), .B(y[221]), .Z(n25785) );
  XOR U36502 ( .A(x[220]), .B(y[220]), .Z(n26574) );
  XOR U36503 ( .A(x[219]), .B(y[219]), .Z(n26571) );
  XOR U36504 ( .A(x[218]), .B(y[218]), .Z(n25788) );
  XOR U36505 ( .A(x[217]), .B(y[217]), .Z(n25795) );
  XOR U36506 ( .A(x[216]), .B(y[216]), .Z(n25792) );
  XOR U36507 ( .A(x[215]), .B(y[215]), .Z(n26566) );
  XOR U36508 ( .A(x[214]), .B(y[214]), .Z(n26563) );
  XOR U36509 ( .A(x[213]), .B(y[213]), .Z(n25798) );
  XOR U36510 ( .A(x[212]), .B(y[212]), .Z(n25804) );
  XOR U36511 ( .A(x[211]), .B(y[211]), .Z(n25801) );
  XOR U36512 ( .A(x[210]), .B(y[210]), .Z(n25808) );
  XOR U36513 ( .A(x[209]), .B(y[209]), .Z(n25814) );
  XOR U36514 ( .A(x[208]), .B(y[208]), .Z(n25811) );
  XOR U36515 ( .A(x[207]), .B(y[207]), .Z(n26558) );
  XOR U36516 ( .A(x[206]), .B(y[206]), .Z(n26555) );
  XOR U36517 ( .A(x[205]), .B(y[205]), .Z(n26551) );
  XOR U36518 ( .A(x[204]), .B(y[204]), .Z(n26548) );
  XOR U36519 ( .A(x[203]), .B(y[203]), .Z(n25820) );
  XOR U36520 ( .A(x[202]), .B(y[202]), .Z(n25817) );
  XOR U36521 ( .A(x[201]), .B(y[201]), .Z(n26545) );
  XOR U36522 ( .A(x[200]), .B(y[200]), .Z(n26542) );
  XOR U36523 ( .A(x[199]), .B(y[199]), .Z(n25826) );
  XOR U36524 ( .A(x[198]), .B(y[198]), .Z(n25823) );
  XOR U36525 ( .A(x[197]), .B(y[197]), .Z(n26538) );
  XOR U36526 ( .A(x[196]), .B(y[196]), .Z(n26535) );
  XOR U36527 ( .A(x[195]), .B(y[195]), .Z(n25832) );
  XOR U36528 ( .A(x[194]), .B(y[194]), .Z(n25829) );
  XOR U36529 ( .A(x[193]), .B(y[193]), .Z(n26531) );
  XOR U36530 ( .A(x[192]), .B(y[192]), .Z(n26528) );
  XOR U36531 ( .A(x[191]), .B(y[191]), .Z(n25835) );
  XOR U36532 ( .A(x[190]), .B(y[190]), .Z(n26522) );
  XOR U36533 ( .A(x[189]), .B(y[189]), .Z(n25838) );
  XOR U36534 ( .A(x[188]), .B(y[188]), .Z(n26516) );
  XOR U36535 ( .A(x[187]), .B(y[187]), .Z(n26513) );
  XOR U36536 ( .A(x[186]), .B(y[186]), .Z(n25841) );
  XOR U36537 ( .A(x[185]), .B(y[185]), .Z(n26509) );
  XOR U36538 ( .A(x[184]), .B(y[184]), .Z(n26506) );
  XOR U36539 ( .A(x[183]), .B(y[183]), .Z(n26502) );
  XOR U36540 ( .A(x[182]), .B(y[182]), .Z(n26499) );
  XOR U36541 ( .A(x[181]), .B(y[181]), .Z(n25848) );
  XOR U36542 ( .A(x[180]), .B(y[180]), .Z(n25845) );
  XOR U36543 ( .A(x[179]), .B(y[179]), .Z(n26494) );
  XOR U36544 ( .A(x[178]), .B(y[178]), .Z(n26491) );
  XOR U36545 ( .A(x[177]), .B(y[177]), .Z(n25854) );
  XOR U36546 ( .A(x[176]), .B(y[176]), .Z(n25851) );
  XOR U36547 ( .A(x[175]), .B(y[175]), .Z(n25860) );
  XOR U36548 ( .A(x[174]), .B(y[174]), .Z(n25857) );
  XOR U36549 ( .A(x[173]), .B(y[173]), .Z(n25866) );
  XOR U36550 ( .A(x[172]), .B(y[172]), .Z(n25863) );
  XOR U36551 ( .A(x[171]), .B(y[171]), .Z(n25873) );
  XOR U36552 ( .A(x[170]), .B(y[170]), .Z(n25870) );
  XOR U36553 ( .A(x[169]), .B(y[169]), .Z(n25877) );
  XOR U36554 ( .A(x[168]), .B(y[168]), .Z(n25883) );
  XOR U36555 ( .A(x[167]), .B(y[167]), .Z(n25880) );
  XOR U36556 ( .A(x[166]), .B(y[166]), .Z(n25887) );
  XOR U36557 ( .A(x[165]), .B(y[165]), .Z(n26485) );
  XOR U36558 ( .A(x[164]), .B(y[164]), .Z(n26482) );
  XOR U36559 ( .A(x[163]), .B(y[163]), .Z(n26478) );
  XOR U36560 ( .A(x[162]), .B(y[162]), .Z(n26475) );
  XOR U36561 ( .A(x[161]), .B(y[161]), .Z(n26471) );
  XOR U36562 ( .A(x[160]), .B(y[160]), .Z(n26468) );
  XOR U36563 ( .A(x[159]), .B(y[159]), .Z(n25890) );
  XOR U36564 ( .A(x[158]), .B(y[158]), .Z(n26464) );
  XOR U36565 ( .A(x[157]), .B(y[157]), .Z(n26461) );
  XOR U36566 ( .A(x[156]), .B(y[156]), .Z(n26457) );
  XOR U36567 ( .A(x[155]), .B(y[155]), .Z(n26454) );
  XOR U36568 ( .A(x[154]), .B(y[154]), .Z(n25894) );
  XOR U36569 ( .A(x[153]), .B(y[153]), .Z(n26450) );
  XOR U36570 ( .A(x[152]), .B(y[152]), .Z(n26447) );
  XOR U36571 ( .A(x[151]), .B(y[151]), .Z(n26443) );
  XOR U36572 ( .A(x[150]), .B(y[150]), .Z(n26440) );
  XOR U36573 ( .A(x[149]), .B(y[149]), .Z(n25900) );
  XOR U36574 ( .A(x[148]), .B(y[148]), .Z(n25897) );
  XOR U36575 ( .A(x[147]), .B(y[147]), .Z(n26437) );
  XOR U36576 ( .A(x[146]), .B(y[146]), .Z(n26434) );
  XOR U36577 ( .A(x[145]), .B(y[145]), .Z(n25906) );
  XOR U36578 ( .A(x[144]), .B(y[144]), .Z(n25903) );
  XOR U36579 ( .A(x[143]), .B(y[143]), .Z(n25909) );
  XOR U36580 ( .A(x[142]), .B(y[142]), .Z(n26430) );
  XOR U36581 ( .A(x[141]), .B(y[141]), .Z(n26427) );
  XOR U36582 ( .A(x[140]), .B(y[140]), .Z(n25915) );
  XOR U36583 ( .A(x[139]), .B(y[139]), .Z(n25912) );
  XOR U36584 ( .A(x[138]), .B(y[138]), .Z(n25918) );
  XOR U36585 ( .A(x[137]), .B(y[137]), .Z(n26415) );
  XOR U36586 ( .A(x[136]), .B(y[136]), .Z(n26402) );
  XOR U36587 ( .A(x[135]), .B(y[135]), .Z(n25921) );
  XOR U36588 ( .A(x[134]), .B(y[134]), .Z(n25924) );
  XOR U36589 ( .A(x[133]), .B(y[133]), .Z(n25930) );
  XOR U36590 ( .A(x[132]), .B(y[132]), .Z(n25927) );
  XOR U36591 ( .A(x[131]), .B(y[131]), .Z(n25936) );
  XOR U36592 ( .A(x[130]), .B(y[130]), .Z(n25933) );
  XOR U36593 ( .A(x[129]), .B(y[129]), .Z(n25943) );
  XOR U36594 ( .A(x[128]), .B(y[128]), .Z(n25940) );
  XOR U36595 ( .A(x[127]), .B(y[127]), .Z(n25946) );
  XOR U36596 ( .A(x[126]), .B(y[126]), .Z(n26391) );
  XOR U36597 ( .A(x[125]), .B(y[125]), .Z(n26388) );
  XOR U36598 ( .A(x[124]), .B(y[124]), .Z(n25952) );
  XOR U36599 ( .A(x[123]), .B(y[123]), .Z(n25949) );
  XOR U36600 ( .A(x[122]), .B(y[122]), .Z(n25955) );
  XOR U36601 ( .A(x[121]), .B(y[121]), .Z(n26383) );
  XOR U36602 ( .A(x[120]), .B(y[120]), .Z(n26380) );
  XOR U36603 ( .A(x[119]), .B(y[119]), .Z(n26376) );
  XOR U36604 ( .A(x[118]), .B(y[118]), .Z(n26373) );
  XOR U36605 ( .A(x[117]), .B(y[117]), .Z(n26369) );
  XOR U36606 ( .A(x[116]), .B(y[116]), .Z(n26366) );
  XOR U36607 ( .A(x[115]), .B(y[115]), .Z(n25961) );
  XOR U36608 ( .A(x[114]), .B(y[114]), .Z(n25958) );
  XOR U36609 ( .A(x[113]), .B(y[113]), .Z(n25967) );
  XOR U36610 ( .A(x[112]), .B(y[112]), .Z(n25964) );
  XOR U36611 ( .A(x[111]), .B(y[111]), .Z(n25973) );
  XOR U36612 ( .A(x[110]), .B(y[110]), .Z(n25970) );
  XOR U36613 ( .A(x[109]), .B(y[109]), .Z(n25979) );
  XOR U36614 ( .A(x[108]), .B(y[108]), .Z(n25976) );
  XOR U36615 ( .A(x[107]), .B(y[107]), .Z(n25985) );
  XOR U36616 ( .A(x[106]), .B(y[106]), .Z(n25982) );
  XOR U36617 ( .A(x[105]), .B(y[105]), .Z(n25988) );
  XOR U36618 ( .A(x[104]), .B(y[104]), .Z(n36005) );
  XOR U36619 ( .A(x[103]), .B(y[103]), .Z(n25992) );
  IV U36620 ( .A(x[102]), .Z(n24489) );
  XOR U36621 ( .A(n24489), .B(y[102]), .Z(n26000) );
  XOR U36622 ( .A(x[101]), .B(y[101]), .Z(n25997) );
  XOR U36623 ( .A(x[100]), .B(y[100]), .Z(n26360) );
  XOR U36624 ( .A(x[99]), .B(y[99]), .Z(n26357) );
  XOR U36625 ( .A(x[98]), .B(y[98]), .Z(n26350) );
  XOR U36626 ( .A(x[97]), .B(y[97]), .Z(n26002) );
  XOR U36627 ( .A(x[96]), .B(y[96]), .Z(n26346) );
  XOR U36628 ( .A(x[95]), .B(y[95]), .Z(n26343) );
  XOR U36629 ( .A(x[94]), .B(y[94]), .Z(n26339) );
  XOR U36630 ( .A(x[93]), .B(y[93]), .Z(n26336) );
  XOR U36631 ( .A(x[92]), .B(y[92]), .Z(n26008) );
  XOR U36632 ( .A(x[91]), .B(y[91]), .Z(n26005) );
  XOR U36633 ( .A(x[90]), .B(y[90]), .Z(n26011) );
  XOR U36634 ( .A(x[89]), .B(y[89]), .Z(n26321) );
  XOR U36635 ( .A(x[88]), .B(y[88]), .Z(n26017) );
  XOR U36636 ( .A(x[87]), .B(y[87]), .Z(n26014) );
  XOR U36637 ( .A(x[86]), .B(y[86]), .Z(n26316) );
  XOR U36638 ( .A(x[85]), .B(y[85]), .Z(n26313) );
  XOR U36639 ( .A(x[84]), .B(y[84]), .Z(n26023) );
  XOR U36640 ( .A(x[83]), .B(y[83]), .Z(n26020) );
  XOR U36641 ( .A(x[82]), .B(y[82]), .Z(n26309) );
  XOR U36642 ( .A(x[81]), .B(y[81]), .Z(n26306) );
  XOR U36643 ( .A(x[80]), .B(y[80]), .Z(n26029) );
  XOR U36644 ( .A(x[79]), .B(y[79]), .Z(n26026) );
  XOR U36645 ( .A(x[78]), .B(y[78]), .Z(n26032) );
  XOR U36646 ( .A(x[77]), .B(y[77]), .Z(n26038) );
  XOR U36647 ( .A(x[76]), .B(y[76]), .Z(n26035) );
  XOR U36648 ( .A(x[75]), .B(y[75]), .Z(n26044) );
  XOR U36649 ( .A(x[74]), .B(y[74]), .Z(n26041) );
  XOR U36650 ( .A(x[73]), .B(y[73]), .Z(n26047) );
  XOR U36651 ( .A(x[72]), .B(y[72]), .Z(n26300) );
  XOR U36652 ( .A(x[71]), .B(y[71]), .Z(n26297) );
  XOR U36653 ( .A(x[70]), .B(y[70]), .Z(n26053) );
  XOR U36654 ( .A(x[69]), .B(y[69]), .Z(n26050) );
  XOR U36655 ( .A(x[68]), .B(y[68]), .Z(n26293) );
  XOR U36656 ( .A(x[67]), .B(y[67]), .Z(n26290) );
  XOR U36657 ( .A(x[66]), .B(y[66]), .Z(n26279) );
  XOR U36658 ( .A(x[65]), .B(y[65]), .Z(n26057) );
  XOR U36659 ( .A(x[64]), .B(y[64]), .Z(n26282) );
  XOR U36660 ( .A(x[63]), .B(y[63]), .Z(n26275) );
  XOR U36661 ( .A(x[62]), .B(y[62]), .Z(n26272) );
  XOR U36662 ( .A(x[61]), .B(y[61]), .Z(n26268) );
  XOR U36663 ( .A(x[60]), .B(y[60]), .Z(n26265) );
  XOR U36664 ( .A(x[59]), .B(y[59]), .Z(n26261) );
  XOR U36665 ( .A(x[58]), .B(y[58]), .Z(n26258) );
  XOR U36666 ( .A(x[57]), .B(y[57]), .Z(n26064) );
  XOR U36667 ( .A(x[56]), .B(y[56]), .Z(n26061) );
  XOR U36668 ( .A(x[55]), .B(y[55]), .Z(n26070) );
  XOR U36669 ( .A(x[54]), .B(y[54]), .Z(n26067) );
  XOR U36670 ( .A(x[53]), .B(y[53]), .Z(n26076) );
  XOR U36671 ( .A(x[52]), .B(y[52]), .Z(n26073) );
  XOR U36672 ( .A(x[51]), .B(y[51]), .Z(n26254) );
  XOR U36673 ( .A(x[50]), .B(y[50]), .Z(n26251) );
  XOR U36674 ( .A(x[49]), .B(y[49]), .Z(n26082) );
  XOR U36675 ( .A(x[48]), .B(y[48]), .Z(n26079) );
  XOR U36676 ( .A(x[47]), .B(y[47]), .Z(n26247) );
  XOR U36677 ( .A(x[46]), .B(y[46]), .Z(n26244) );
  XOR U36678 ( .A(x[45]), .B(y[45]), .Z(n26088) );
  XOR U36679 ( .A(x[44]), .B(y[44]), .Z(n26085) );
  XOR U36680 ( .A(x[43]), .B(y[43]), .Z(n26241) );
  XOR U36681 ( .A(x[42]), .B(y[42]), .Z(n26238) );
  XOR U36682 ( .A(x[41]), .B(y[41]), .Z(n26234) );
  XOR U36683 ( .A(x[40]), .B(y[40]), .Z(n26231) );
  XOR U36684 ( .A(x[39]), .B(y[39]), .Z(n26091) );
  XOR U36685 ( .A(x[38]), .B(y[38]), .Z(n26097) );
  XOR U36686 ( .A(x[37]), .B(y[37]), .Z(n26094) );
  XOR U36687 ( .A(x[36]), .B(y[36]), .Z(n26225) );
  XOR U36688 ( .A(x[35]), .B(y[35]), .Z(n26222) );
  XOR U36689 ( .A(x[34]), .B(y[34]), .Z(n26218) );
  XOR U36690 ( .A(x[33]), .B(y[33]), .Z(n26215) );
  XOR U36691 ( .A(x[32]), .B(y[32]), .Z(n26212) );
  XOR U36692 ( .A(x[31]), .B(y[31]), .Z(n26209) );
  XOR U36693 ( .A(x[30]), .B(y[30]), .Z(n26205) );
  XOR U36694 ( .A(x[29]), .B(y[29]), .Z(n26202) );
  XOR U36695 ( .A(x[28]), .B(y[28]), .Z(n26100) );
  XOR U36696 ( .A(x[27]), .B(y[27]), .Z(n26198) );
  XOR U36697 ( .A(x[26]), .B(y[26]), .Z(n26195) );
  XOR U36698 ( .A(x[25]), .B(y[25]), .Z(n26191) );
  XOR U36699 ( .A(x[24]), .B(y[24]), .Z(n26188) );
  XOR U36700 ( .A(x[23]), .B(y[23]), .Z(n26184) );
  XOR U36701 ( .A(x[22]), .B(y[22]), .Z(n26181) );
  XOR U36702 ( .A(x[21]), .B(y[21]), .Z(n26177) );
  XOR U36703 ( .A(x[20]), .B(y[20]), .Z(n26174) );
  XOR U36704 ( .A(x[19]), .B(y[19]), .Z(n26103) );
  XOR U36705 ( .A(x[18]), .B(y[18]), .Z(n26170) );
  XOR U36706 ( .A(x[17]), .B(y[17]), .Z(n26167) );
  XOR U36707 ( .A(x[16]), .B(y[16]), .Z(n26163) );
  XOR U36708 ( .A(x[15]), .B(y[15]), .Z(n26160) );
  XOR U36709 ( .A(x[14]), .B(y[14]), .Z(n26109) );
  XOR U36710 ( .A(x[13]), .B(y[13]), .Z(n26106) );
  XOR U36711 ( .A(x[12]), .B(y[12]), .Z(n26112) );
  XOR U36712 ( .A(x[11]), .B(y[11]), .Z(n26118) );
  XOR U36713 ( .A(x[10]), .B(y[10]), .Z(n26115) );
  XOR U36714 ( .A(x[9]), .B(y[9]), .Z(n26124) );
  XOR U36715 ( .A(x[8]), .B(y[8]), .Z(n26121) );
  XOR U36716 ( .A(x[7]), .B(y[7]), .Z(n26151) );
  XOR U36717 ( .A(x[6]), .B(y[6]), .Z(n26148) );
  XOR U36718 ( .A(x[5]), .B(y[5]), .Z(n26127) );
  XOR U36719 ( .A(x[4]), .B(y[4]), .Z(n26130) );
  XOR U36720 ( .A(y[3]), .B(x[3]), .Z(n26133) );
  XOR U36721 ( .A(x[2]), .B(y[2]), .Z(n26141) );
  XOR U36722 ( .A(x[1]), .B(y[1]), .Z(n26137) );
  XOR U36723 ( .A(y[0]), .B(x[0]), .Z(n24490) );
  IV U36724 ( .A(n24490), .Z(n26138) );
  XOR U36725 ( .A(n26137), .B(n26138), .Z(n26142) );
  XOR U36726 ( .A(n26141), .B(n26142), .Z(n26134) );
  XOR U36727 ( .A(n26133), .B(n26134), .Z(n26132) );
  XOR U36728 ( .A(n26130), .B(n26132), .Z(n26129) );
  XOR U36729 ( .A(n26127), .B(n26129), .Z(n26149) );
  XOR U36730 ( .A(n26148), .B(n26149), .Z(n26152) );
  XOR U36731 ( .A(n26151), .B(n26152), .Z(n26123) );
  XOR U36732 ( .A(n26121), .B(n26123), .Z(n26125) );
  XOR U36733 ( .A(n26124), .B(n26125), .Z(n26116) );
  XOR U36734 ( .A(n26115), .B(n26116), .Z(n26119) );
  XOR U36735 ( .A(n26118), .B(n26119), .Z(n26113) );
  XOR U36736 ( .A(n26112), .B(n26113), .Z(n26107) );
  XOR U36737 ( .A(n26106), .B(n26107), .Z(n26111) );
  XOR U36738 ( .A(n26109), .B(n26111), .Z(n26162) );
  XOR U36739 ( .A(n26160), .B(n26162), .Z(n26165) );
  XOR U36740 ( .A(n26163), .B(n26165), .Z(n26169) );
  XOR U36741 ( .A(n26167), .B(n26169), .Z(n26172) );
  XOR U36742 ( .A(n26170), .B(n26172), .Z(n26105) );
  XOR U36743 ( .A(n26103), .B(n26105), .Z(n26175) );
  XOR U36744 ( .A(n26174), .B(n26175), .Z(n26179) );
  XOR U36745 ( .A(n26177), .B(n26179), .Z(n26183) );
  XOR U36746 ( .A(n26181), .B(n26183), .Z(n26186) );
  XOR U36747 ( .A(n26184), .B(n26186), .Z(n26189) );
  XOR U36748 ( .A(n26188), .B(n26189), .Z(n26192) );
  XOR U36749 ( .A(n26191), .B(n26192), .Z(n26197) );
  XOR U36750 ( .A(n26195), .B(n26197), .Z(n26200) );
  XOR U36751 ( .A(n26198), .B(n26200), .Z(n26101) );
  XOR U36752 ( .A(n26100), .B(n26101), .Z(n26203) );
  XOR U36753 ( .A(n26202), .B(n26203), .Z(n26207) );
  XOR U36754 ( .A(n26205), .B(n26207), .Z(n26211) );
  XOR U36755 ( .A(n26209), .B(n26211), .Z(n26213) );
  XOR U36756 ( .A(n26212), .B(n26213), .Z(n26216) );
  XOR U36757 ( .A(n26215), .B(n26216), .Z(n26220) );
  XOR U36758 ( .A(n26218), .B(n26220), .Z(n26224) );
  XOR U36759 ( .A(n26222), .B(n26224), .Z(n26227) );
  XOR U36760 ( .A(n26225), .B(n26227), .Z(n26096) );
  XOR U36761 ( .A(n26094), .B(n26096), .Z(n26099) );
  XOR U36762 ( .A(n26097), .B(n26099), .Z(n26093) );
  XOR U36763 ( .A(n26091), .B(n26093), .Z(n26232) );
  XOR U36764 ( .A(n26231), .B(n26232), .Z(n26235) );
  XOR U36765 ( .A(n26234), .B(n26235), .Z(n26240) );
  XOR U36766 ( .A(n26238), .B(n26240), .Z(n26242) );
  XOR U36767 ( .A(n26241), .B(n26242), .Z(n26086) );
  XOR U36768 ( .A(n26085), .B(n26086), .Z(n26090) );
  XOR U36769 ( .A(n26088), .B(n26090), .Z(n26246) );
  XOR U36770 ( .A(n26244), .B(n26246), .Z(n26249) );
  XOR U36771 ( .A(n26247), .B(n26249), .Z(n26080) );
  XOR U36772 ( .A(n26079), .B(n26080), .Z(n26084) );
  XOR U36773 ( .A(n26082), .B(n26084), .Z(n26252) );
  XOR U36774 ( .A(n26251), .B(n26252), .Z(n26256) );
  XOR U36775 ( .A(n26254), .B(n26256), .Z(n26074) );
  XOR U36776 ( .A(n26073), .B(n26074), .Z(n26078) );
  XOR U36777 ( .A(n26076), .B(n26078), .Z(n26069) );
  XOR U36778 ( .A(n26067), .B(n26069), .Z(n26072) );
  XOR U36779 ( .A(n26070), .B(n26072), .Z(n26063) );
  XOR U36780 ( .A(n26061), .B(n26063), .Z(n26066) );
  XOR U36781 ( .A(n26064), .B(n26066), .Z(n26260) );
  XOR U36782 ( .A(n26258), .B(n26260), .Z(n26263) );
  XOR U36783 ( .A(n26261), .B(n26263), .Z(n26267) );
  XOR U36784 ( .A(n26265), .B(n26267), .Z(n26270) );
  XOR U36785 ( .A(n26268), .B(n26270), .Z(n26274) );
  XOR U36786 ( .A(n26272), .B(n26274), .Z(n26277) );
  XOR U36787 ( .A(n26275), .B(n26277), .Z(n26283) );
  XOR U36788 ( .A(n26282), .B(n26283), .Z(n26059) );
  XOR U36789 ( .A(n26057), .B(n26059), .Z(n26281) );
  XOR U36790 ( .A(n26279), .B(n26281), .Z(n26292) );
  XOR U36791 ( .A(n26290), .B(n26292), .Z(n26294) );
  XOR U36792 ( .A(n26293), .B(n26294), .Z(n26051) );
  XOR U36793 ( .A(n26050), .B(n26051), .Z(n26055) );
  XOR U36794 ( .A(n26053), .B(n26055), .Z(n26298) );
  XOR U36795 ( .A(n26297), .B(n26298), .Z(n26301) );
  XOR U36796 ( .A(n26300), .B(n26301), .Z(n26048) );
  XOR U36797 ( .A(n26047), .B(n26048), .Z(n26043) );
  XOR U36798 ( .A(n26041), .B(n26043), .Z(n26046) );
  XOR U36799 ( .A(n26044), .B(n26046), .Z(n26036) );
  XOR U36800 ( .A(n26035), .B(n26036), .Z(n26039) );
  XOR U36801 ( .A(n26038), .B(n26039), .Z(n26034) );
  XOR U36802 ( .A(n26032), .B(n26034), .Z(n26027) );
  XOR U36803 ( .A(n26026), .B(n26027), .Z(n26030) );
  XOR U36804 ( .A(n26029), .B(n26030), .Z(n26307) );
  XOR U36805 ( .A(n26306), .B(n26307), .Z(n26311) );
  XOR U36806 ( .A(n26309), .B(n26311), .Z(n26022) );
  XOR U36807 ( .A(n26020), .B(n26022), .Z(n26024) );
  XOR U36808 ( .A(n26023), .B(n26024), .Z(n26315) );
  XOR U36809 ( .A(n26313), .B(n26315), .Z(n26318) );
  XOR U36810 ( .A(n26316), .B(n26318), .Z(n26016) );
  XOR U36811 ( .A(n26014), .B(n26016), .Z(n26019) );
  XOR U36812 ( .A(n26017), .B(n26019), .Z(n26323) );
  XOR U36813 ( .A(n26321), .B(n26323), .Z(n26012) );
  XOR U36814 ( .A(n26011), .B(n26012), .Z(n26006) );
  XOR U36815 ( .A(n26005), .B(n26006), .Z(n26010) );
  XOR U36816 ( .A(n26008), .B(n26010), .Z(n26338) );
  XOR U36817 ( .A(n26336), .B(n26338), .Z(n26341) );
  XOR U36818 ( .A(n26339), .B(n26341), .Z(n26345) );
  XOR U36819 ( .A(n26343), .B(n26345), .Z(n26347) );
  XOR U36820 ( .A(n26346), .B(n26347), .Z(n26004) );
  XOR U36821 ( .A(n26002), .B(n26004), .Z(n26352) );
  XOR U36822 ( .A(n26350), .B(n26352), .Z(n26358) );
  XOR U36823 ( .A(n26357), .B(n26358), .Z(n26361) );
  XOR U36824 ( .A(n26360), .B(n26361), .Z(n25999) );
  XOR U36825 ( .A(n25997), .B(n25999), .Z(n26001) );
  XOR U36826 ( .A(n26000), .B(n26001), .Z(n25991) );
  IV U36827 ( .A(n25991), .Z(n25993) );
  XOR U36828 ( .A(n25992), .B(n25993), .Z(n36006) );
  XOR U36829 ( .A(n36005), .B(n36006), .Z(n25990) );
  XOR U36830 ( .A(n25988), .B(n25990), .Z(n25984) );
  XOR U36831 ( .A(n25982), .B(n25984), .Z(n25987) );
  XOR U36832 ( .A(n25985), .B(n25987), .Z(n25977) );
  XOR U36833 ( .A(n25976), .B(n25977), .Z(n25981) );
  XOR U36834 ( .A(n25979), .B(n25981), .Z(n25972) );
  XOR U36835 ( .A(n25970), .B(n25972), .Z(n25975) );
  XOR U36836 ( .A(n25973), .B(n25975), .Z(n25965) );
  XOR U36837 ( .A(n25964), .B(n25965), .Z(n25968) );
  XOR U36838 ( .A(n25967), .B(n25968), .Z(n25960) );
  XOR U36839 ( .A(n25958), .B(n25960), .Z(n25963) );
  XOR U36840 ( .A(n25961), .B(n25963), .Z(n26368) );
  XOR U36841 ( .A(n26366), .B(n26368), .Z(n26371) );
  XOR U36842 ( .A(n26369), .B(n26371), .Z(n26375) );
  XOR U36843 ( .A(n26373), .B(n26375), .Z(n26378) );
  XOR U36844 ( .A(n26376), .B(n26378), .Z(n26381) );
  XOR U36845 ( .A(n26380), .B(n26381), .Z(n26384) );
  XOR U36846 ( .A(n26383), .B(n26384), .Z(n25956) );
  XOR U36847 ( .A(n25955), .B(n25956), .Z(n25950) );
  XOR U36848 ( .A(n25949), .B(n25950), .Z(n25953) );
  XOR U36849 ( .A(n25952), .B(n25953), .Z(n26390) );
  XOR U36850 ( .A(n26388), .B(n26390), .Z(n26393) );
  XOR U36851 ( .A(n26391), .B(n26393), .Z(n25948) );
  XOR U36852 ( .A(n25946), .B(n25948), .Z(n25941) );
  XOR U36853 ( .A(n25940), .B(n25941), .Z(n25945) );
  XOR U36854 ( .A(n25943), .B(n25945), .Z(n25935) );
  XOR U36855 ( .A(n25933), .B(n25935), .Z(n25937) );
  XOR U36856 ( .A(n25936), .B(n25937), .Z(n25928) );
  XOR U36857 ( .A(n25927), .B(n25928), .Z(n25931) );
  XOR U36858 ( .A(n25930), .B(n25931), .Z(n25926) );
  XOR U36859 ( .A(n25924), .B(n25926), .Z(n25923) );
  XOR U36860 ( .A(n25921), .B(n25923), .Z(n26403) );
  XOR U36861 ( .A(n26402), .B(n26403), .Z(n26416) );
  XOR U36862 ( .A(n26415), .B(n26416), .Z(n25920) );
  XOR U36863 ( .A(n25918), .B(n25920), .Z(n25914) );
  XOR U36864 ( .A(n25912), .B(n25914), .Z(n25916) );
  XOR U36865 ( .A(n25915), .B(n25916), .Z(n26429) );
  XOR U36866 ( .A(n26427), .B(n26429), .Z(n26432) );
  XOR U36867 ( .A(n26430), .B(n26432), .Z(n25910) );
  XOR U36868 ( .A(n25909), .B(n25910), .Z(n25904) );
  XOR U36869 ( .A(n25903), .B(n25904), .Z(n25907) );
  XOR U36870 ( .A(n25906), .B(n25907), .Z(n26436) );
  XOR U36871 ( .A(n26434), .B(n26436), .Z(n26439) );
  XOR U36872 ( .A(n26437), .B(n26439), .Z(n25899) );
  XOR U36873 ( .A(n25897), .B(n25899), .Z(n25902) );
  XOR U36874 ( .A(n25900), .B(n25902), .Z(n26442) );
  XOR U36875 ( .A(n26440), .B(n26442), .Z(n26445) );
  XOR U36876 ( .A(n26443), .B(n26445), .Z(n26448) );
  XOR U36877 ( .A(n26447), .B(n26448), .Z(n26452) );
  XOR U36878 ( .A(n26450), .B(n26452), .Z(n25896) );
  XOR U36879 ( .A(n25894), .B(n25896), .Z(n26455) );
  XOR U36880 ( .A(n26454), .B(n26455), .Z(n26458) );
  XOR U36881 ( .A(n26457), .B(n26458), .Z(n26463) );
  XOR U36882 ( .A(n26461), .B(n26463), .Z(n26465) );
  XOR U36883 ( .A(n26464), .B(n26465), .Z(n25892) );
  XOR U36884 ( .A(n25890), .B(n25892), .Z(n26470) );
  XOR U36885 ( .A(n26468), .B(n26470), .Z(n26473) );
  XOR U36886 ( .A(n26471), .B(n26473), .Z(n26476) );
  XOR U36887 ( .A(n26475), .B(n26476), .Z(n26480) );
  XOR U36888 ( .A(n26478), .B(n26480), .Z(n26483) );
  XOR U36889 ( .A(n26482), .B(n26483), .Z(n26487) );
  XOR U36890 ( .A(n26485), .B(n26487), .Z(n25889) );
  XOR U36891 ( .A(n25887), .B(n25889), .Z(n25881) );
  XOR U36892 ( .A(n25880), .B(n25881), .Z(n25884) );
  XOR U36893 ( .A(n25883), .B(n25884), .Z(n25879) );
  XOR U36894 ( .A(n25877), .B(n25879), .Z(n25871) );
  XOR U36895 ( .A(n25870), .B(n25871), .Z(n25875) );
  XOR U36896 ( .A(n25873), .B(n25875), .Z(n25864) );
  XOR U36897 ( .A(n25863), .B(n25864), .Z(n25868) );
  XOR U36898 ( .A(n25866), .B(n25868), .Z(n25859) );
  XOR U36899 ( .A(n25857), .B(n25859), .Z(n25861) );
  XOR U36900 ( .A(n25860), .B(n25861), .Z(n25852) );
  XOR U36901 ( .A(n25851), .B(n25852), .Z(n25855) );
  XOR U36902 ( .A(n25854), .B(n25855), .Z(n26493) );
  XOR U36903 ( .A(n26491), .B(n26493), .Z(n26496) );
  XOR U36904 ( .A(n26494), .B(n26496), .Z(n25846) );
  XOR U36905 ( .A(n25845), .B(n25846), .Z(n25850) );
  XOR U36906 ( .A(n25848), .B(n25850), .Z(n26501) );
  XOR U36907 ( .A(n26499), .B(n26501), .Z(n26504) );
  XOR U36908 ( .A(n26502), .B(n26504), .Z(n26507) );
  XOR U36909 ( .A(n26506), .B(n26507), .Z(n26511) );
  XOR U36910 ( .A(n26509), .B(n26511), .Z(n25842) );
  XOR U36911 ( .A(n25841), .B(n25842), .Z(n26514) );
  XOR U36912 ( .A(n26513), .B(n26514), .Z(n26518) );
  XOR U36913 ( .A(n26516), .B(n26518), .Z(n25840) );
  XOR U36914 ( .A(n25838), .B(n25840), .Z(n26524) );
  XOR U36915 ( .A(n26522), .B(n26524), .Z(n25837) );
  XOR U36916 ( .A(n25835), .B(n25837), .Z(n26529) );
  XOR U36917 ( .A(n26528), .B(n26529), .Z(n26533) );
  XOR U36918 ( .A(n26531), .B(n26533), .Z(n25831) );
  XOR U36919 ( .A(n25829), .B(n25831), .Z(n25834) );
  XOR U36920 ( .A(n25832), .B(n25834), .Z(n26537) );
  XOR U36921 ( .A(n26535), .B(n26537), .Z(n26540) );
  XOR U36922 ( .A(n26538), .B(n26540), .Z(n25824) );
  XOR U36923 ( .A(n25823), .B(n25824), .Z(n25828) );
  XOR U36924 ( .A(n25826), .B(n25828), .Z(n26543) );
  XOR U36925 ( .A(n26542), .B(n26543), .Z(n26546) );
  XOR U36926 ( .A(n26545), .B(n26546), .Z(n25819) );
  XOR U36927 ( .A(n25817), .B(n25819), .Z(n25822) );
  XOR U36928 ( .A(n25820), .B(n25822), .Z(n26549) );
  XOR U36929 ( .A(n26548), .B(n26549), .Z(n26552) );
  XOR U36930 ( .A(n26551), .B(n26552), .Z(n26557) );
  XOR U36931 ( .A(n26555), .B(n26557), .Z(n26560) );
  XOR U36932 ( .A(n26558), .B(n26560), .Z(n25813) );
  XOR U36933 ( .A(n25811), .B(n25813), .Z(n25816) );
  XOR U36934 ( .A(n25814), .B(n25816), .Z(n25810) );
  XOR U36935 ( .A(n25808), .B(n25810), .Z(n25803) );
  XOR U36936 ( .A(n25801), .B(n25803), .Z(n25805) );
  XOR U36937 ( .A(n25804), .B(n25805), .Z(n25800) );
  XOR U36938 ( .A(n25798), .B(n25800), .Z(n26565) );
  XOR U36939 ( .A(n26563), .B(n26565), .Z(n26568) );
  XOR U36940 ( .A(n26566), .B(n26568), .Z(n25793) );
  XOR U36941 ( .A(n25792), .B(n25793), .Z(n25796) );
  XOR U36942 ( .A(n25795), .B(n25796), .Z(n25790) );
  XOR U36943 ( .A(n25788), .B(n25790), .Z(n26573) );
  XOR U36944 ( .A(n26571), .B(n26573), .Z(n26575) );
  XOR U36945 ( .A(n26574), .B(n26575), .Z(n25787) );
  XOR U36946 ( .A(n25785), .B(n25787), .Z(n26582) );
  XOR U36947 ( .A(n26580), .B(n26582), .Z(n25784) );
  XOR U36948 ( .A(n25782), .B(n25784), .Z(n26587) );
  XOR U36949 ( .A(n26586), .B(n26587), .Z(n26591) );
  XOR U36950 ( .A(n26589), .B(n26591), .Z(n25778) );
  XOR U36951 ( .A(n25776), .B(n25778), .Z(n25780) );
  XOR U36952 ( .A(n25779), .B(n25780), .Z(n25771) );
  XOR U36953 ( .A(n25770), .B(n25771), .Z(n25774) );
  XOR U36954 ( .A(n25773), .B(n25774), .Z(n25768) );
  XOR U36955 ( .A(n25766), .B(n25768), .Z(n26595) );
  XOR U36956 ( .A(n26594), .B(n26595), .Z(n26598) );
  XOR U36957 ( .A(n26597), .B(n26598), .Z(n26602) );
  XOR U36958 ( .A(n26601), .B(n26602), .Z(n26606) );
  XOR U36959 ( .A(n26604), .B(n26606), .Z(n25765) );
  XOR U36960 ( .A(n25763), .B(n25765), .Z(n25757) );
  XOR U36961 ( .A(n25756), .B(n25757), .Z(n25761) );
  XOR U36962 ( .A(n25759), .B(n25761), .Z(n25752) );
  XOR U36963 ( .A(n25750), .B(n25752), .Z(n25754) );
  XOR U36964 ( .A(n25753), .B(n25754), .Z(n26608) );
  XOR U36965 ( .A(n26607), .B(n26608), .Z(n26611) );
  XOR U36966 ( .A(n26610), .B(n26611), .Z(n25746) );
  XOR U36967 ( .A(n25744), .B(n25746), .Z(n25749) );
  XOR U36968 ( .A(n25747), .B(n25749), .Z(n26615) );
  XOR U36969 ( .A(n26614), .B(n26615), .Z(n26619) );
  XOR U36970 ( .A(n26617), .B(n26619), .Z(n25739) );
  XOR U36971 ( .A(n25737), .B(n25739), .Z(n25742) );
  XOR U36972 ( .A(n25740), .B(n25742), .Z(n25732) );
  XOR U36973 ( .A(n25731), .B(n25732), .Z(n25736) );
  XOR U36974 ( .A(n25734), .B(n25736), .Z(n25730) );
  XOR U36975 ( .A(n25728), .B(n25730), .Z(n25724) );
  XOR U36976 ( .A(n25722), .B(n25724), .Z(n25726) );
  XOR U36977 ( .A(n25725), .B(n25726), .Z(n25718) );
  XOR U36978 ( .A(n25716), .B(n25718), .Z(n25721) );
  XOR U36979 ( .A(n25719), .B(n25721), .Z(n25715) );
  XOR U36980 ( .A(n25713), .B(n25715), .Z(n25708) );
  XOR U36981 ( .A(n25707), .B(n25708), .Z(n25712) );
  XOR U36982 ( .A(n25710), .B(n25712), .Z(n26624) );
  XOR U36983 ( .A(n26622), .B(n26624), .Z(n26626) );
  XOR U36984 ( .A(n26625), .B(n26626), .Z(n25702) );
  XOR U36985 ( .A(n25701), .B(n25702), .Z(n25706) );
  XOR U36986 ( .A(n25704), .B(n25706), .Z(n26630) );
  XOR U36987 ( .A(n26629), .B(n26630), .Z(n26634) );
  XOR U36988 ( .A(n26632), .B(n26634), .Z(n25696) );
  XOR U36989 ( .A(n25695), .B(n25696), .Z(n25700) );
  XOR U36990 ( .A(n25698), .B(n25700), .Z(n26640) );
  XOR U36991 ( .A(n26638), .B(n26640), .Z(n25693) );
  XOR U36992 ( .A(n25691), .B(n25693), .Z(n26652) );
  XOR U36993 ( .A(n26650), .B(n26652), .Z(n26655) );
  XOR U36994 ( .A(n26653), .B(n26655), .Z(n26658) );
  XOR U36995 ( .A(n26657), .B(n26658), .Z(n26662) );
  XOR U36996 ( .A(n26660), .B(n26662), .Z(n26665) );
  XOR U36997 ( .A(n26664), .B(n26665), .Z(n26668) );
  XOR U36998 ( .A(n26667), .B(n26668), .Z(n25690) );
  XOR U36999 ( .A(n25688), .B(n25690), .Z(n26676) );
  XOR U37000 ( .A(n26675), .B(n26676), .Z(n26679) );
  XOR U37001 ( .A(n26678), .B(n26679), .Z(n25684) );
  XOR U37002 ( .A(n25682), .B(n25684), .Z(n25687) );
  XOR U37003 ( .A(n25685), .B(n25687), .Z(n25681) );
  XOR U37004 ( .A(n25679), .B(n25681), .Z(n25673) );
  XOR U37005 ( .A(n25672), .B(n25673), .Z(n25676) );
  XOR U37006 ( .A(n25675), .B(n25676), .Z(n25668) );
  XOR U37007 ( .A(n25666), .B(n25668), .Z(n25671) );
  XOR U37008 ( .A(n25669), .B(n25671), .Z(n25661) );
  XOR U37009 ( .A(n25660), .B(n25661), .Z(n25665) );
  XOR U37010 ( .A(n25663), .B(n25665), .Z(n26686) );
  XOR U37011 ( .A(n26685), .B(n26686), .Z(n26690) );
  XOR U37012 ( .A(n26688), .B(n26690), .Z(n25656) );
  XOR U37013 ( .A(n25654), .B(n25656), .Z(n25659) );
  XOR U37014 ( .A(n25657), .B(n25659), .Z(n25649) );
  XOR U37015 ( .A(n25648), .B(n25649), .Z(n25653) );
  XOR U37016 ( .A(n25651), .B(n25653), .Z(n25644) );
  XOR U37017 ( .A(n25642), .B(n25644), .Z(n25647) );
  XOR U37018 ( .A(n25645), .B(n25647), .Z(n25641) );
  XOR U37019 ( .A(n25639), .B(n25641), .Z(n26694) );
  XOR U37020 ( .A(n26693), .B(n26694), .Z(n26697) );
  XOR U37021 ( .A(n26696), .B(n26697), .Z(n26701) );
  XOR U37022 ( .A(n26700), .B(n26701), .Z(n26705) );
  XOR U37023 ( .A(n26703), .B(n26705), .Z(n26709) );
  XOR U37024 ( .A(n26707), .B(n26709), .Z(n26711) );
  XOR U37025 ( .A(n26710), .B(n26711), .Z(n25638) );
  XOR U37026 ( .A(n25636), .B(n25638), .Z(n25632) );
  XOR U37027 ( .A(n25630), .B(n25632), .Z(n25635) );
  XOR U37028 ( .A(n25633), .B(n25635), .Z(n25625) );
  XOR U37029 ( .A(n25624), .B(n25625), .Z(n25628) );
  XOR U37030 ( .A(n25627), .B(n25628), .Z(n25623) );
  XOR U37031 ( .A(n25621), .B(n25623), .Z(n25617) );
  XOR U37032 ( .A(n25615), .B(n25617), .Z(n25619) );
  XOR U37033 ( .A(n25618), .B(n25619), .Z(n25611) );
  XOR U37034 ( .A(n25609), .B(n25611), .Z(n25614) );
  XOR U37035 ( .A(n25612), .B(n25614), .Z(n25607) );
  XOR U37036 ( .A(n25606), .B(n25607), .Z(n25601) );
  XOR U37037 ( .A(n25600), .B(n25601), .Z(n25605) );
  XOR U37038 ( .A(n25603), .B(n25605), .Z(n25596) );
  XOR U37039 ( .A(n25594), .B(n25596), .Z(n25598) );
  XOR U37040 ( .A(n25597), .B(n25598), .Z(n25589) );
  XOR U37041 ( .A(n25588), .B(n25589), .Z(n25593) );
  XOR U37042 ( .A(n25591), .B(n25593), .Z(n25586) );
  XOR U37043 ( .A(n25585), .B(n25586), .Z(n26730) );
  XOR U37044 ( .A(n26728), .B(n26730), .Z(n25582) );
  XOR U37045 ( .A(n25581), .B(n25582), .Z(n26727) );
  XOR U37046 ( .A(n26725), .B(n26727), .Z(n25577) );
  XOR U37047 ( .A(n25575), .B(n25577), .Z(n25580) );
  XOR U37048 ( .A(n25578), .B(n25580), .Z(n25570) );
  XOR U37049 ( .A(n25569), .B(n25570), .Z(n25574) );
  XOR U37050 ( .A(n25572), .B(n25574), .Z(n25565) );
  XOR U37051 ( .A(n25563), .B(n25565), .Z(n25568) );
  XOR U37052 ( .A(n25566), .B(n25568), .Z(n25558) );
  XOR U37053 ( .A(n25557), .B(n25558), .Z(n25561) );
  XOR U37054 ( .A(n25560), .B(n25561), .Z(n25553) );
  XOR U37055 ( .A(n25551), .B(n25553), .Z(n25556) );
  XOR U37056 ( .A(n25554), .B(n25556), .Z(n25545) );
  XOR U37057 ( .A(n25544), .B(n25545), .Z(n25549) );
  XOR U37058 ( .A(n25547), .B(n25549), .Z(n25540) );
  XOR U37059 ( .A(n25538), .B(n25540), .Z(n25542) );
  XOR U37060 ( .A(n25541), .B(n25542), .Z(n25536) );
  XOR U37061 ( .A(n25535), .B(n25536), .Z(n26746) );
  XOR U37062 ( .A(n26745), .B(n26746), .Z(n26750) );
  XOR U37063 ( .A(n26748), .B(n26750), .Z(n26754) );
  XOR U37064 ( .A(n26752), .B(n26754), .Z(n26756) );
  XOR U37065 ( .A(n26755), .B(n26756), .Z(n26761) );
  XOR U37066 ( .A(n26759), .B(n26761), .Z(n26763) );
  XOR U37067 ( .A(n26762), .B(n26763), .Z(n25534) );
  XOR U37068 ( .A(n25532), .B(n25534), .Z(n25527) );
  XOR U37069 ( .A(n25526), .B(n25527), .Z(n25530) );
  XOR U37070 ( .A(n25529), .B(n25530), .Z(n25521) );
  XOR U37071 ( .A(n25520), .B(n25521), .Z(n25525) );
  XOR U37072 ( .A(n25523), .B(n25525), .Z(n25515) );
  XOR U37073 ( .A(n25514), .B(n25515), .Z(n25519) );
  XOR U37074 ( .A(n25517), .B(n25519), .Z(n26770) );
  XOR U37075 ( .A(n26768), .B(n26770), .Z(n26772) );
  XOR U37076 ( .A(n26771), .B(n26772), .Z(n25508) );
  XOR U37077 ( .A(n25507), .B(n25508), .Z(n25512) );
  XOR U37078 ( .A(n25510), .B(n25512), .Z(n26777) );
  XOR U37079 ( .A(n26775), .B(n26777), .Z(n26779) );
  XOR U37080 ( .A(n26778), .B(n26779), .Z(n25502) );
  XOR U37081 ( .A(n25501), .B(n25502), .Z(n25506) );
  XOR U37082 ( .A(n25504), .B(n25506), .Z(n26784) );
  XOR U37083 ( .A(n26782), .B(n26784), .Z(n26787) );
  XOR U37084 ( .A(n26785), .B(n26787), .Z(n26800) );
  XOR U37085 ( .A(n26799), .B(n26800), .Z(n26803) );
  XOR U37086 ( .A(n26802), .B(n26803), .Z(n25500) );
  XOR U37087 ( .A(n25498), .B(n25500), .Z(n26808) );
  XOR U37088 ( .A(n26806), .B(n26808), .Z(n26810) );
  XOR U37089 ( .A(n26809), .B(n26810), .Z(n25494) );
  XOR U37090 ( .A(n25492), .B(n25494), .Z(n25497) );
  XOR U37091 ( .A(n25495), .B(n25497), .Z(n25490) );
  XOR U37092 ( .A(n25489), .B(n25490), .Z(n25484) );
  XOR U37093 ( .A(n25483), .B(n25484), .Z(n25486) );
  XOR U37094 ( .A(n25487), .B(n25486), .Z(n25477) );
  IV U37095 ( .A(n25477), .Z(n25480) );
  XOR U37096 ( .A(n25478), .B(n25480), .Z(n36823) );
  XOR U37097 ( .A(n36821), .B(n36823), .Z(n26816) );
  XOR U37098 ( .A(n26814), .B(n26816), .Z(n26819) );
  XOR U37099 ( .A(n26817), .B(n26819), .Z(n26823) );
  XOR U37100 ( .A(n26821), .B(n26823), .Z(n26826) );
  XOR U37101 ( .A(n26824), .B(n26826), .Z(n26828) );
  XOR U37102 ( .A(n26827), .B(n26828), .Z(n26832) );
  XOR U37103 ( .A(n26830), .B(n26832), .Z(n25473) );
  XOR U37104 ( .A(n25471), .B(n25473), .Z(n25475) );
  XOR U37105 ( .A(n25474), .B(n25475), .Z(n25469) );
  XOR U37106 ( .A(n25468), .B(n25469), .Z(n26836) );
  XOR U37107 ( .A(n26834), .B(n26836), .Z(n26839) );
  XOR U37108 ( .A(n26837), .B(n26839), .Z(n26842) );
  XOR U37109 ( .A(n26841), .B(n26842), .Z(n26845) );
  XOR U37110 ( .A(n26844), .B(n26845), .Z(n25467) );
  XOR U37111 ( .A(n25465), .B(n25467), .Z(n26850) );
  XOR U37112 ( .A(n26848), .B(n26850), .Z(n26852) );
  XOR U37113 ( .A(n26851), .B(n26852), .Z(n26856) );
  XOR U37114 ( .A(n26855), .B(n26856), .Z(n26859) );
  XOR U37115 ( .A(n26858), .B(n26859), .Z(n26863) );
  XOR U37116 ( .A(n26861), .B(n26863), .Z(n26866) );
  XOR U37117 ( .A(n26864), .B(n26866), .Z(n26869) );
  XOR U37118 ( .A(n26868), .B(n26869), .Z(n26873) );
  XOR U37119 ( .A(n26871), .B(n26873), .Z(n25461) );
  XOR U37120 ( .A(n25459), .B(n25461), .Z(n25463) );
  XOR U37121 ( .A(n25462), .B(n25463), .Z(n25454) );
  XOR U37122 ( .A(n25453), .B(n25454), .Z(n25458) );
  XOR U37123 ( .A(n25456), .B(n25458), .Z(n26876) );
  XOR U37124 ( .A(n26875), .B(n26876), .Z(n26880) );
  XOR U37125 ( .A(n26878), .B(n26880), .Z(n25451) );
  XOR U37126 ( .A(n25450), .B(n25451), .Z(n25445) );
  XOR U37127 ( .A(n25444), .B(n25445), .Z(n25449) );
  XOR U37128 ( .A(n25447), .B(n25449), .Z(n25440) );
  XOR U37129 ( .A(n25438), .B(n25440), .Z(n25442) );
  XOR U37130 ( .A(n25441), .B(n25442), .Z(n25437) );
  XOR U37131 ( .A(n25435), .B(n25437), .Z(n25434) );
  XOR U37132 ( .A(n25432), .B(n25434), .Z(n26885) );
  XOR U37133 ( .A(n26884), .B(n26885), .Z(n25430) );
  XOR U37134 ( .A(n25429), .B(n25430), .Z(n25428) );
  XOR U37135 ( .A(n25426), .B(n25428), .Z(n26900) );
  XOR U37136 ( .A(n26898), .B(n26900), .Z(n26903) );
  XOR U37137 ( .A(n26901), .B(n26903), .Z(n25422) );
  XOR U37138 ( .A(n25420), .B(n25422), .Z(n25425) );
  XOR U37139 ( .A(n25423), .B(n25425), .Z(n26909) );
  XOR U37140 ( .A(n26907), .B(n26909), .Z(n25419) );
  XOR U37141 ( .A(n25417), .B(n25419), .Z(n26920) );
  XOR U37142 ( .A(n26919), .B(n26920), .Z(n26923) );
  XOR U37143 ( .A(n26922), .B(n26923), .Z(n26928) );
  XOR U37144 ( .A(n26926), .B(n26928), .Z(n26931) );
  XOR U37145 ( .A(n26929), .B(n26931), .Z(n25415) );
  XOR U37146 ( .A(n25414), .B(n25415), .Z(n25409) );
  XOR U37147 ( .A(n25408), .B(n25409), .Z(n25413) );
  XOR U37148 ( .A(n25411), .B(n25413), .Z(n26940) );
  XOR U37149 ( .A(n26939), .B(n26940), .Z(n26943) );
  XOR U37150 ( .A(n26942), .B(n26943), .Z(n25403) );
  XOR U37151 ( .A(n25402), .B(n25403), .Z(n25407) );
  XOR U37152 ( .A(n25405), .B(n25407), .Z(n26948) );
  XOR U37153 ( .A(n26946), .B(n26948), .Z(n26950) );
  XOR U37154 ( .A(n26949), .B(n26950), .Z(n26958) );
  XOR U37155 ( .A(n26956), .B(n26958), .Z(n25400) );
  XOR U37156 ( .A(n25398), .B(n25400), .Z(n26955) );
  XOR U37157 ( .A(n26953), .B(n26955), .Z(n25396) );
  XOR U37158 ( .A(n25395), .B(n25396), .Z(n26966) );
  XOR U37159 ( .A(n26965), .B(n26966), .Z(n26970) );
  XOR U37160 ( .A(n26968), .B(n26970), .Z(n26973) );
  XOR U37161 ( .A(n26972), .B(n26973), .Z(n26976) );
  XOR U37162 ( .A(n26975), .B(n26976), .Z(n26980) );
  XOR U37163 ( .A(n26979), .B(n26980), .Z(n26984) );
  XOR U37164 ( .A(n26982), .B(n26984), .Z(n25390) );
  XOR U37165 ( .A(n25389), .B(n25390), .Z(n25393) );
  XOR U37166 ( .A(n25392), .B(n25393), .Z(n25384) );
  XOR U37167 ( .A(n25383), .B(n25384), .Z(n25388) );
  XOR U37168 ( .A(n25386), .B(n25388), .Z(n26989) );
  XOR U37169 ( .A(n26987), .B(n26989), .Z(n26991) );
  XOR U37170 ( .A(n26990), .B(n26991), .Z(n26997) );
  XOR U37171 ( .A(n26995), .B(n26997), .Z(n25382) );
  XOR U37172 ( .A(n25380), .B(n25382), .Z(n27011) );
  XOR U37173 ( .A(n27009), .B(n27011), .Z(n25378) );
  XOR U37174 ( .A(n25377), .B(n25378), .Z(n25372) );
  XOR U37175 ( .A(n25371), .B(n25372), .Z(n25376) );
  XOR U37176 ( .A(n25374), .B(n25376), .Z(n27024) );
  XOR U37177 ( .A(n27023), .B(n27024), .Z(n27027) );
  XOR U37178 ( .A(n27026), .B(n27027), .Z(n27031) );
  XOR U37179 ( .A(n27030), .B(n27031), .Z(n27035) );
  XOR U37180 ( .A(n27033), .B(n27035), .Z(n27039) );
  XOR U37181 ( .A(n27037), .B(n27039), .Z(n27041) );
  XOR U37182 ( .A(n27040), .B(n27041), .Z(n25366) );
  XOR U37183 ( .A(n25365), .B(n25366), .Z(n25370) );
  XOR U37184 ( .A(n25368), .B(n25370), .Z(n25361) );
  XOR U37185 ( .A(n25359), .B(n25361), .Z(n25364) );
  XOR U37186 ( .A(n25362), .B(n25364), .Z(n25355) );
  XOR U37187 ( .A(n25353), .B(n25355), .Z(n25358) );
  XOR U37188 ( .A(n25356), .B(n25358), .Z(n27047) );
  XOR U37189 ( .A(n27046), .B(n27047), .Z(n27050) );
  XOR U37190 ( .A(n27049), .B(n27050), .Z(n25351) );
  XOR U37191 ( .A(n25350), .B(n25351), .Z(n27057) );
  XOR U37192 ( .A(n27055), .B(n27057), .Z(n25348) );
  XOR U37193 ( .A(n25347), .B(n25348), .Z(n25342) );
  XOR U37194 ( .A(n25341), .B(n25342), .Z(n25346) );
  XOR U37195 ( .A(n25344), .B(n25346), .Z(n25337) );
  XOR U37196 ( .A(n25335), .B(n25337), .Z(n25340) );
  XOR U37197 ( .A(n25338), .B(n25340), .Z(n25334) );
  XOR U37198 ( .A(n25332), .B(n25334), .Z(n27066) );
  XOR U37199 ( .A(n27064), .B(n27066), .Z(n25330) );
  XOR U37200 ( .A(n25329), .B(n25330), .Z(n25328) );
  XOR U37201 ( .A(n25326), .B(n25328), .Z(n25322) );
  XOR U37202 ( .A(n25320), .B(n25322), .Z(n25325) );
  XOR U37203 ( .A(n25323), .B(n25325), .Z(n27081) );
  XOR U37204 ( .A(n27079), .B(n27081), .Z(n27084) );
  XOR U37205 ( .A(n27082), .B(n27084), .Z(n27088) );
  XOR U37206 ( .A(n27086), .B(n27088), .Z(n27090) );
  XOR U37207 ( .A(n27089), .B(n27090), .Z(n25317) );
  XOR U37208 ( .A(n25316), .B(n25317), .Z(n25312) );
  XOR U37209 ( .A(n25310), .B(n25312), .Z(n25315) );
  XOR U37210 ( .A(n25313), .B(n25315), .Z(n27103) );
  XOR U37211 ( .A(n27101), .B(n27103), .Z(n27106) );
  XOR U37212 ( .A(n27104), .B(n27106), .Z(n25306) );
  XOR U37213 ( .A(n25304), .B(n25306), .Z(n25308) );
  XOR U37214 ( .A(n25307), .B(n25308), .Z(n27110) );
  XOR U37215 ( .A(n27108), .B(n27110), .Z(n27113) );
  XOR U37216 ( .A(n27111), .B(n27113), .Z(n25300) );
  XOR U37217 ( .A(n25298), .B(n25300), .Z(n25302) );
  XOR U37218 ( .A(n25301), .B(n25302), .Z(n27118) );
  XOR U37219 ( .A(n27116), .B(n27118), .Z(n27121) );
  XOR U37220 ( .A(n27119), .B(n27121), .Z(n25294) );
  XOR U37221 ( .A(n25292), .B(n25294), .Z(n25297) );
  XOR U37222 ( .A(n25295), .B(n25297), .Z(n27125) );
  XOR U37223 ( .A(n27124), .B(n27125), .Z(n27128) );
  XOR U37224 ( .A(n27127), .B(n27128), .Z(n27133) );
  XOR U37225 ( .A(n27131), .B(n27133), .Z(n27136) );
  XOR U37226 ( .A(n27134), .B(n27136), .Z(n27140) );
  XOR U37227 ( .A(n27138), .B(n27140), .Z(n27143) );
  XOR U37228 ( .A(n27141), .B(n27143), .Z(n27146) );
  XOR U37229 ( .A(n27145), .B(n27146), .Z(n27149) );
  XOR U37230 ( .A(n27148), .B(n27149), .Z(n25287) );
  XOR U37231 ( .A(n25285), .B(n25287), .Z(n25290) );
  XOR U37232 ( .A(n25288), .B(n25290), .Z(n27157) );
  XOR U37233 ( .A(n27155), .B(n27157), .Z(n25282) );
  XOR U37234 ( .A(n25281), .B(n25282), .Z(n27154) );
  XOR U37235 ( .A(n27152), .B(n27154), .Z(n25277) );
  XOR U37236 ( .A(n25275), .B(n25277), .Z(n25280) );
  XOR U37237 ( .A(n25278), .B(n25280), .Z(n27165) );
  XOR U37238 ( .A(n27164), .B(n27165), .Z(n27168) );
  XOR U37239 ( .A(n27167), .B(n27168), .Z(n25274) );
  XOR U37240 ( .A(n25272), .B(n25274), .Z(n25267) );
  XOR U37241 ( .A(n25265), .B(n25267), .Z(n25269) );
  XOR U37242 ( .A(n25268), .B(n25269), .Z(n25263) );
  XOR U37243 ( .A(n25262), .B(n25263), .Z(n27174) );
  XOR U37244 ( .A(n27172), .B(n27174), .Z(n27177) );
  XOR U37245 ( .A(n27175), .B(n27177), .Z(n27180) );
  XOR U37246 ( .A(n27179), .B(n27180), .Z(n27183) );
  XOR U37247 ( .A(n27182), .B(n27183), .Z(n25261) );
  XOR U37248 ( .A(n25259), .B(n25261), .Z(n27187) );
  XOR U37249 ( .A(n27186), .B(n27187), .Z(n27190) );
  XOR U37250 ( .A(n27189), .B(n27190), .Z(n27194) );
  XOR U37251 ( .A(n27193), .B(n27194), .Z(n27198) );
  XOR U37252 ( .A(n27196), .B(n27198), .Z(n25254) );
  XOR U37253 ( .A(n25253), .B(n25254), .Z(n25257) );
  XOR U37254 ( .A(n25256), .B(n25257), .Z(n27201) );
  XOR U37255 ( .A(n27200), .B(n27201), .Z(n27205) );
  XOR U37256 ( .A(n27203), .B(n27205), .Z(n25249) );
  XOR U37257 ( .A(n25247), .B(n25249), .Z(n25251) );
  XOR U37258 ( .A(n25250), .B(n25251), .Z(n25242) );
  XOR U37259 ( .A(n25241), .B(n25242), .Z(n25246) );
  XOR U37260 ( .A(n25244), .B(n25246), .Z(n27209) );
  XOR U37261 ( .A(n27208), .B(n27209), .Z(n27212) );
  XOR U37262 ( .A(n27211), .B(n27212), .Z(n25240) );
  XOR U37263 ( .A(n25238), .B(n25240), .Z(n27222) );
  XOR U37264 ( .A(n27220), .B(n27222), .Z(n25235) );
  XOR U37265 ( .A(n25234), .B(n25235), .Z(n27218) );
  XOR U37266 ( .A(n27217), .B(n27218), .Z(n25233) );
  XOR U37267 ( .A(n25231), .B(n25233), .Z(n27231) );
  XOR U37268 ( .A(n27229), .B(n27231), .Z(n27234) );
  XOR U37269 ( .A(n27232), .B(n27234), .Z(n27237) );
  XOR U37270 ( .A(n27236), .B(n27237), .Z(n27240) );
  XOR U37271 ( .A(n27239), .B(n27240), .Z(n25227) );
  XOR U37272 ( .A(n25225), .B(n25227), .Z(n25230) );
  XOR U37273 ( .A(n25228), .B(n25230), .Z(n27244) );
  XOR U37274 ( .A(n27243), .B(n27244), .Z(n27248) );
  XOR U37275 ( .A(n27246), .B(n27248), .Z(n25219) );
  XOR U37276 ( .A(n25218), .B(n25219), .Z(n25223) );
  XOR U37277 ( .A(n25221), .B(n25223), .Z(n25216) );
  XOR U37278 ( .A(n25215), .B(n25216), .Z(n27252) );
  XOR U37279 ( .A(n27251), .B(n27252), .Z(n27256) );
  XOR U37280 ( .A(n27254), .B(n27256), .Z(n27260) );
  XOR U37281 ( .A(n27258), .B(n27260), .Z(n27262) );
  XOR U37282 ( .A(n27261), .B(n27262), .Z(n27267) );
  XOR U37283 ( .A(n27265), .B(n27267), .Z(n27270) );
  XOR U37284 ( .A(n27268), .B(n27270), .Z(n27273) );
  XOR U37285 ( .A(n27272), .B(n27273), .Z(n27276) );
  XOR U37286 ( .A(n27275), .B(n27276), .Z(n25210) );
  XOR U37287 ( .A(n25209), .B(n25210), .Z(n25214) );
  XOR U37288 ( .A(n25212), .B(n25214), .Z(n25208) );
  XOR U37289 ( .A(n25206), .B(n25208), .Z(n25202) );
  XOR U37290 ( .A(n25200), .B(n25202), .Z(n25205) );
  XOR U37291 ( .A(n25203), .B(n25205), .Z(n25196) );
  XOR U37292 ( .A(n25194), .B(n25196), .Z(n25199) );
  XOR U37293 ( .A(n25197), .B(n25199), .Z(n25189) );
  XOR U37294 ( .A(n25188), .B(n25189), .Z(n25192) );
  XOR U37295 ( .A(n25191), .B(n25192), .Z(n27284) );
  XOR U37296 ( .A(n27282), .B(n27284), .Z(n27287) );
  XOR U37297 ( .A(n27285), .B(n27287), .Z(n25186) );
  XOR U37298 ( .A(n25185), .B(n25186), .Z(n27293) );
  XOR U37299 ( .A(n27291), .B(n27293), .Z(n25184) );
  XOR U37300 ( .A(n25182), .B(n25184), .Z(n27299) );
  XOR U37301 ( .A(n27298), .B(n27299), .Z(n27302) );
  XOR U37302 ( .A(n27301), .B(n27302), .Z(n25181) );
  XOR U37303 ( .A(n25179), .B(n25181), .Z(n27307) );
  XOR U37304 ( .A(n27305), .B(n27307), .Z(n25178) );
  XOR U37305 ( .A(n25176), .B(n25178), .Z(n27318) );
  XOR U37306 ( .A(n27317), .B(n27318), .Z(n27321) );
  XOR U37307 ( .A(n27320), .B(n27321), .Z(n25172) );
  XOR U37308 ( .A(n25170), .B(n25172), .Z(n25175) );
  XOR U37309 ( .A(n25173), .B(n25175), .Z(n25168) );
  XOR U37310 ( .A(n25167), .B(n25168), .Z(n25163) );
  XOR U37311 ( .A(n25161), .B(n25163), .Z(n25166) );
  XOR U37312 ( .A(n25164), .B(n25166), .Z(n27327) );
  XOR U37313 ( .A(n27326), .B(n27327), .Z(n27330) );
  XOR U37314 ( .A(n27329), .B(n27330), .Z(n25160) );
  XOR U37315 ( .A(n25158), .B(n25160), .Z(n25154) );
  XOR U37316 ( .A(n25152), .B(n25154), .Z(n25157) );
  XOR U37317 ( .A(n25155), .B(n25157), .Z(n25147) );
  XOR U37318 ( .A(n25146), .B(n25147), .Z(n25150) );
  XOR U37319 ( .A(n25149), .B(n25150), .Z(n27337) );
  XOR U37320 ( .A(n27335), .B(n27337), .Z(n27340) );
  XOR U37321 ( .A(n27338), .B(n27340), .Z(n25142) );
  XOR U37322 ( .A(n25140), .B(n25142), .Z(n25145) );
  XOR U37323 ( .A(n25143), .B(n25145), .Z(n25135) );
  XOR U37324 ( .A(n25134), .B(n25135), .Z(n25139) );
  XOR U37325 ( .A(n25137), .B(n25139), .Z(n27344) );
  XOR U37326 ( .A(n27343), .B(n27344), .Z(n27348) );
  XOR U37327 ( .A(n27346), .B(n27348), .Z(n25129) );
  XOR U37328 ( .A(n25128), .B(n25129), .Z(n25133) );
  XOR U37329 ( .A(n25131), .B(n25133), .Z(n27350) );
  XOR U37330 ( .A(n27349), .B(n27350), .Z(n27354) );
  XOR U37331 ( .A(n27352), .B(n27354), .Z(n27360) );
  XOR U37332 ( .A(n27358), .B(n27360), .Z(n25126) );
  XOR U37333 ( .A(n25124), .B(n25126), .Z(n27356) );
  XOR U37334 ( .A(n27355), .B(n27356), .Z(n27367) );
  XOR U37335 ( .A(n27366), .B(n27367), .Z(n27371) );
  XOR U37336 ( .A(n27369), .B(n27371), .Z(n27377) );
  XOR U37337 ( .A(n27375), .B(n27377), .Z(n25121) );
  XOR U37338 ( .A(n25120), .B(n25121), .Z(n27374) );
  XOR U37339 ( .A(n27372), .B(n27374), .Z(n25116) );
  XOR U37340 ( .A(n25114), .B(n25116), .Z(n25119) );
  XOR U37341 ( .A(n25117), .B(n25119), .Z(n25109) );
  XOR U37342 ( .A(n25108), .B(n25109), .Z(n25113) );
  XOR U37343 ( .A(n25111), .B(n25113), .Z(n27385) );
  XOR U37344 ( .A(n27384), .B(n27385), .Z(n27389) );
  XOR U37345 ( .A(n27387), .B(n27389), .Z(n27392) );
  XOR U37346 ( .A(n27391), .B(n27392), .Z(n27396) );
  XOR U37347 ( .A(n27394), .B(n27396), .Z(n25104) );
  XOR U37348 ( .A(n25102), .B(n25104), .Z(n25106) );
  XOR U37349 ( .A(n25105), .B(n25106), .Z(n27400) );
  XOR U37350 ( .A(n27399), .B(n27400), .Z(n27403) );
  XOR U37351 ( .A(n27402), .B(n27403), .Z(n25097) );
  XOR U37352 ( .A(n25095), .B(n25097), .Z(n25100) );
  XOR U37353 ( .A(n25098), .B(n25100), .Z(n25090) );
  XOR U37354 ( .A(n25089), .B(n25090), .Z(n25094) );
  XOR U37355 ( .A(n25092), .B(n25094), .Z(n27408) );
  XOR U37356 ( .A(n27406), .B(n27408), .Z(n27410) );
  XOR U37357 ( .A(n27409), .B(n27410), .Z(n27414) );
  XOR U37358 ( .A(n27413), .B(n27414), .Z(n27417) );
  XOR U37359 ( .A(n27416), .B(n27417), .Z(n25088) );
  XOR U37360 ( .A(n25086), .B(n25088), .Z(n27426) );
  XOR U37361 ( .A(n27424), .B(n27426), .Z(n25081) );
  XOR U37362 ( .A(n25080), .B(n25081), .Z(n25085) );
  XOR U37363 ( .A(n25083), .B(n25085), .Z(n25076) );
  XOR U37364 ( .A(n25074), .B(n25076), .Z(n25079) );
  XOR U37365 ( .A(n25077), .B(n25079), .Z(n25069) );
  XOR U37366 ( .A(n25068), .B(n25069), .Z(n25072) );
  XOR U37367 ( .A(n25071), .B(n25072), .Z(n27431) );
  XOR U37368 ( .A(n27430), .B(n27431), .Z(n27435) );
  XOR U37369 ( .A(n27433), .B(n27435), .Z(n27438) );
  XOR U37370 ( .A(n27437), .B(n27438), .Z(n27441) );
  XOR U37371 ( .A(n27440), .B(n27441), .Z(n27446) );
  XOR U37372 ( .A(n27444), .B(n27446), .Z(n27449) );
  XOR U37373 ( .A(n27447), .B(n27449), .Z(n25063) );
  XOR U37374 ( .A(n25062), .B(n25063), .Z(n25067) );
  XOR U37375 ( .A(n25065), .B(n25067), .Z(n27453) );
  XOR U37376 ( .A(n27451), .B(n27453), .Z(n27455) );
  XOR U37377 ( .A(n27454), .B(n27455), .Z(n27459) );
  XOR U37378 ( .A(n27458), .B(n27459), .Z(n27463) );
  XOR U37379 ( .A(n27461), .B(n27463), .Z(n27467) );
  XOR U37380 ( .A(n27465), .B(n27467), .Z(n27470) );
  XOR U37381 ( .A(n27468), .B(n27470), .Z(n27473) );
  XOR U37382 ( .A(n27472), .B(n27473), .Z(n27476) );
  XOR U37383 ( .A(n27475), .B(n27476), .Z(n27481) );
  XOR U37384 ( .A(n27479), .B(n27481), .Z(n27484) );
  XOR U37385 ( .A(n27482), .B(n27484), .Z(n27487) );
  XOR U37386 ( .A(n27486), .B(n27487), .Z(n27491) );
  XOR U37387 ( .A(n27489), .B(n27491), .Z(n25058) );
  XOR U37388 ( .A(n25056), .B(n25058), .Z(n25060) );
  XOR U37389 ( .A(n25059), .B(n25060), .Z(n25051) );
  XOR U37390 ( .A(n25050), .B(n25051), .Z(n25055) );
  XOR U37391 ( .A(n25053), .B(n25055), .Z(n27495) );
  XOR U37392 ( .A(n27493), .B(n27495), .Z(n27498) );
  XOR U37393 ( .A(n27496), .B(n27498), .Z(n27502) );
  XOR U37394 ( .A(n27500), .B(n27502), .Z(n27505) );
  XOR U37395 ( .A(n27503), .B(n27505), .Z(n25049) );
  XOR U37396 ( .A(n25047), .B(n25049), .Z(n27508) );
  XOR U37397 ( .A(n27506), .B(n27508), .Z(n27510) );
  XOR U37398 ( .A(n27509), .B(n27510), .Z(n27515) );
  XOR U37399 ( .A(n27513), .B(n27515), .Z(n27518) );
  XOR U37400 ( .A(n27516), .B(n27518), .Z(n25046) );
  XOR U37401 ( .A(n25044), .B(n25046), .Z(n27521) );
  XOR U37402 ( .A(n27519), .B(n27521), .Z(n27524) );
  XOR U37403 ( .A(n27522), .B(n27524), .Z(n27528) );
  XOR U37404 ( .A(n27526), .B(n27528), .Z(n27531) );
  XOR U37405 ( .A(n27529), .B(n27531), .Z(n25042) );
  XOR U37406 ( .A(n25041), .B(n25042), .Z(n27533) );
  XOR U37407 ( .A(n27532), .B(n27533), .Z(n27537) );
  XOR U37408 ( .A(n27535), .B(n27537), .Z(n27541) );
  XOR U37409 ( .A(n27539), .B(n27541), .Z(n27543) );
  XOR U37410 ( .A(n27542), .B(n27543), .Z(n25040) );
  XOR U37411 ( .A(n25038), .B(n25040), .Z(n27547) );
  XOR U37412 ( .A(n27545), .B(n27547), .Z(n27550) );
  XOR U37413 ( .A(n27548), .B(n27550), .Z(n27553) );
  XOR U37414 ( .A(n27552), .B(n27553), .Z(n27556) );
  XOR U37415 ( .A(n27555), .B(n27556), .Z(n27560) );
  XOR U37416 ( .A(n27558), .B(n27560), .Z(n27563) );
  XOR U37417 ( .A(n27561), .B(n27563), .Z(n27568) );
  XOR U37418 ( .A(n27567), .B(n27568), .Z(n25037) );
  XOR U37419 ( .A(n25035), .B(n25037), .Z(n27581) );
  XOR U37420 ( .A(n27579), .B(n27581), .Z(n27583) );
  XOR U37421 ( .A(n27582), .B(n27583), .Z(n27589) );
  XOR U37422 ( .A(n27588), .B(n27589), .Z(n25032) );
  XOR U37423 ( .A(n25031), .B(n25032), .Z(n27587) );
  XOR U37424 ( .A(n27585), .B(n27587), .Z(n25026) );
  XOR U37425 ( .A(n25025), .B(n25026), .Z(n25029) );
  XOR U37426 ( .A(n25028), .B(n25029), .Z(n25021) );
  XOR U37427 ( .A(n25019), .B(n25021), .Z(n25024) );
  XOR U37428 ( .A(n25022), .B(n25024), .Z(n27599) );
  XOR U37429 ( .A(n27597), .B(n27599), .Z(n27601) );
  XOR U37430 ( .A(n27600), .B(n27601), .Z(n25017) );
  XOR U37431 ( .A(n25016), .B(n25017), .Z(n27608) );
  XOR U37432 ( .A(n27606), .B(n27608), .Z(n25015) );
  XOR U37433 ( .A(n25013), .B(n25015), .Z(n25011) );
  XOR U37434 ( .A(n25010), .B(n25011), .Z(n27618) );
  XOR U37435 ( .A(n27617), .B(n27618), .Z(n27622) );
  XOR U37436 ( .A(n27620), .B(n27622), .Z(n25009) );
  XOR U37437 ( .A(n25007), .B(n25009), .Z(n27625) );
  XOR U37438 ( .A(n27624), .B(n27625), .Z(n27629) );
  XOR U37439 ( .A(n27627), .B(n27629), .Z(n27633) );
  XOR U37440 ( .A(n27631), .B(n27633), .Z(n27636) );
  XOR U37441 ( .A(n27634), .B(n27636), .Z(n25002) );
  XOR U37442 ( .A(n25001), .B(n25002), .Z(n25006) );
  XOR U37443 ( .A(n25004), .B(n25006), .Z(n27640) );
  XOR U37444 ( .A(n27638), .B(n27640), .Z(n27643) );
  XOR U37445 ( .A(n27641), .B(n27643), .Z(n24996) );
  XOR U37446 ( .A(n24995), .B(n24996), .Z(n25000) );
  XOR U37447 ( .A(n24998), .B(n25000), .Z(n24994) );
  XOR U37448 ( .A(n24992), .B(n24994), .Z(n24991) );
  XOR U37449 ( .A(n24989), .B(n24991), .Z(n27655) );
  XOR U37450 ( .A(n27654), .B(n27655), .Z(n24988) );
  XOR U37451 ( .A(n24986), .B(n24988), .Z(n27664) );
  XOR U37452 ( .A(n27662), .B(n27664), .Z(n24985) );
  XOR U37453 ( .A(n24983), .B(n24985), .Z(n24978) );
  XOR U37454 ( .A(n24977), .B(n24978), .Z(n24982) );
  XOR U37455 ( .A(n24980), .B(n24982), .Z(n24973) );
  XOR U37456 ( .A(n24971), .B(n24973), .Z(n24976) );
  XOR U37457 ( .A(n24974), .B(n24976), .Z(n24966) );
  XOR U37458 ( .A(n24965), .B(n24966), .Z(n24970) );
  XOR U37459 ( .A(n24968), .B(n24970), .Z(n27678) );
  XOR U37460 ( .A(n27676), .B(n27678), .Z(n27681) );
  XOR U37461 ( .A(n27679), .B(n27681), .Z(n24963) );
  XOR U37462 ( .A(n24962), .B(n24963), .Z(n24957) );
  XOR U37463 ( .A(n24956), .B(n24957), .Z(n24961) );
  XOR U37464 ( .A(n24959), .B(n24961), .Z(n27685) );
  XOR U37465 ( .A(n27683), .B(n27685), .Z(n27687) );
  XOR U37466 ( .A(n27686), .B(n27687), .Z(n24954) );
  XOR U37467 ( .A(n24953), .B(n24954), .Z(n24948) );
  XOR U37468 ( .A(n24946), .B(n24948), .Z(n24950) );
  XOR U37469 ( .A(n24949), .B(n24950), .Z(n24944) );
  XOR U37470 ( .A(n24943), .B(n24944), .Z(n27691) );
  XOR U37471 ( .A(n27690), .B(n27691), .Z(n27695) );
  XOR U37472 ( .A(n27693), .B(n27695), .Z(n24939) );
  XOR U37473 ( .A(n24937), .B(n24939), .Z(n24941) );
  XOR U37474 ( .A(n24940), .B(n24941), .Z(n27699) );
  XOR U37475 ( .A(n27697), .B(n27699), .Z(n27702) );
  XOR U37476 ( .A(n27700), .B(n27702), .Z(n24936) );
  XOR U37477 ( .A(n24934), .B(n24936), .Z(n24929) );
  XOR U37478 ( .A(n24928), .B(n24929), .Z(n24932) );
  XOR U37479 ( .A(n24931), .B(n24932), .Z(n27708) );
  XOR U37480 ( .A(n27706), .B(n27708), .Z(n27711) );
  XOR U37481 ( .A(n27709), .B(n27711), .Z(n24924) );
  XOR U37482 ( .A(n24922), .B(n24924), .Z(n24927) );
  XOR U37483 ( .A(n24925), .B(n24927), .Z(n27716) );
  XOR U37484 ( .A(n27714), .B(n27716), .Z(n27719) );
  XOR U37485 ( .A(n27717), .B(n27719), .Z(n27722) );
  XOR U37486 ( .A(n27721), .B(n27722), .Z(n27725) );
  XOR U37487 ( .A(n27724), .B(n27725), .Z(n24921) );
  XOR U37488 ( .A(n24919), .B(n24921), .Z(n27730) );
  XOR U37489 ( .A(n27728), .B(n27730), .Z(n27732) );
  XOR U37490 ( .A(n27731), .B(n27732), .Z(n24914) );
  XOR U37491 ( .A(n24912), .B(n24914), .Z(n24916) );
  XOR U37492 ( .A(n24915), .B(n24916), .Z(n24908) );
  XOR U37493 ( .A(n24906), .B(n24908), .Z(n24910) );
  XOR U37494 ( .A(n24909), .B(n24910), .Z(n24901) );
  XOR U37495 ( .A(n24900), .B(n24901), .Z(n24905) );
  XOR U37496 ( .A(n24903), .B(n24905), .Z(n24896) );
  XOR U37497 ( .A(n24894), .B(n24896), .Z(n24898) );
  XOR U37498 ( .A(n24897), .B(n24898), .Z(n27739) );
  XOR U37499 ( .A(n27737), .B(n27739), .Z(n27742) );
  XOR U37500 ( .A(n27740), .B(n27742), .Z(n24893) );
  XOR U37501 ( .A(n24891), .B(n24893), .Z(n24886) );
  XOR U37502 ( .A(n24885), .B(n24886), .Z(n24890) );
  XOR U37503 ( .A(n24888), .B(n24890), .Z(n24881) );
  XOR U37504 ( .A(n24879), .B(n24881), .Z(n24884) );
  XOR U37505 ( .A(n24882), .B(n24884), .Z(n27745) );
  XOR U37506 ( .A(n27744), .B(n27745), .Z(n27749) );
  XOR U37507 ( .A(n27747), .B(n27749), .Z(n27753) );
  XOR U37508 ( .A(n27751), .B(n27753), .Z(n27755) );
  XOR U37509 ( .A(n27754), .B(n27755), .Z(n24877) );
  XOR U37510 ( .A(n24876), .B(n24877), .Z(n27759) );
  XOR U37511 ( .A(n27758), .B(n27759), .Z(n27763) );
  XOR U37512 ( .A(n27761), .B(n27763), .Z(n24872) );
  XOR U37513 ( .A(n24870), .B(n24872), .Z(n24874) );
  XOR U37514 ( .A(n24873), .B(n24874), .Z(n27767) );
  XOR U37515 ( .A(n27765), .B(n27767), .Z(n27770) );
  XOR U37516 ( .A(n27768), .B(n27770), .Z(n24866) );
  XOR U37517 ( .A(n24864), .B(n24866), .Z(n24869) );
  XOR U37518 ( .A(n24867), .B(n24869), .Z(n24860) );
  XOR U37519 ( .A(n24858), .B(n24860), .Z(n24862) );
  XOR U37520 ( .A(n24861), .B(n24862), .Z(n24856) );
  XOR U37521 ( .A(n24855), .B(n24856), .Z(n24851) );
  XOR U37522 ( .A(n24849), .B(n24851), .Z(n24854) );
  XOR U37523 ( .A(n24852), .B(n24854), .Z(n24845) );
  XOR U37524 ( .A(n24843), .B(n24845), .Z(n24848) );
  XOR U37525 ( .A(n24846), .B(n24848), .Z(n27777) );
  XOR U37526 ( .A(n27776), .B(n27777), .Z(n27780) );
  XOR U37527 ( .A(n27779), .B(n27780), .Z(n27785) );
  XOR U37528 ( .A(n27783), .B(n27785), .Z(n27788) );
  XOR U37529 ( .A(n27786), .B(n27788), .Z(n24839) );
  XOR U37530 ( .A(n24837), .B(n24839), .Z(n24842) );
  XOR U37531 ( .A(n24840), .B(n24842), .Z(n27791) );
  XOR U37532 ( .A(n27790), .B(n27791), .Z(n27795) );
  XOR U37533 ( .A(n27793), .B(n27795), .Z(n24832) );
  XOR U37534 ( .A(n24831), .B(n24832), .Z(n24835) );
  XOR U37535 ( .A(n24834), .B(n24835), .Z(n27800) );
  XOR U37536 ( .A(n27798), .B(n27800), .Z(n27803) );
  XOR U37537 ( .A(n27801), .B(n27803), .Z(n24826) );
  XOR U37538 ( .A(n24825), .B(n24826), .Z(n24830) );
  XOR U37539 ( .A(n24828), .B(n24830), .Z(n27807) );
  XOR U37540 ( .A(n27805), .B(n27807), .Z(n27809) );
  XOR U37541 ( .A(n27808), .B(n27809), .Z(n27813) );
  XOR U37542 ( .A(n27812), .B(n27813), .Z(n27816) );
  XOR U37543 ( .A(n27815), .B(n27816), .Z(n27821) );
  XOR U37544 ( .A(n27819), .B(n27821), .Z(n27824) );
  XOR U37545 ( .A(n27822), .B(n27824), .Z(n24820) );
  XOR U37546 ( .A(n24819), .B(n24820), .Z(n24824) );
  XOR U37547 ( .A(n24822), .B(n24824), .Z(n27829) );
  XOR U37548 ( .A(n27827), .B(n27829), .Z(n27831) );
  XOR U37549 ( .A(n27830), .B(n27831), .Z(n27835) );
  XOR U37550 ( .A(n27834), .B(n27835), .Z(n27838) );
  XOR U37551 ( .A(n27837), .B(n27838), .Z(n27842) );
  XOR U37552 ( .A(n27840), .B(n27842), .Z(n27844) );
  XOR U37553 ( .A(n27843), .B(n27844), .Z(n24814) );
  XOR U37554 ( .A(n24813), .B(n24814), .Z(n24818) );
  XOR U37555 ( .A(n24816), .B(n24818), .Z(n24811) );
  XOR U37556 ( .A(n24810), .B(n24811), .Z(n27850) );
  XOR U37557 ( .A(n27848), .B(n27850), .Z(n27852) );
  XOR U37558 ( .A(n27851), .B(n27852), .Z(n27856) );
  XOR U37559 ( .A(n27855), .B(n27856), .Z(n27860) );
  XOR U37560 ( .A(n27858), .B(n27860), .Z(n27864) );
  XOR U37561 ( .A(n27862), .B(n27864), .Z(n27866) );
  XOR U37562 ( .A(n27865), .B(n27866), .Z(n27870) );
  XOR U37563 ( .A(n27869), .B(n27870), .Z(n27874) );
  XOR U37564 ( .A(n27872), .B(n27874), .Z(n27878) );
  XOR U37565 ( .A(n27876), .B(n27878), .Z(n27880) );
  XOR U37566 ( .A(n27879), .B(n27880), .Z(n27884) );
  XOR U37567 ( .A(n27883), .B(n27884), .Z(n27888) );
  XOR U37568 ( .A(n27886), .B(n27888), .Z(n24805) );
  XOR U37569 ( .A(n24804), .B(n24805), .Z(n24808) );
  XOR U37570 ( .A(n24807), .B(n24808), .Z(n24800) );
  XOR U37571 ( .A(n24798), .B(n24800), .Z(n24803) );
  XOR U37572 ( .A(n24801), .B(n24803), .Z(n27892) );
  XOR U37573 ( .A(n27891), .B(n27892), .Z(n27895) );
  XOR U37574 ( .A(n27894), .B(n27895), .Z(n24796) );
  XOR U37575 ( .A(n24795), .B(n24796), .Z(n27903) );
  XOR U37576 ( .A(n27901), .B(n27903), .Z(n24794) );
  XOR U37577 ( .A(n24792), .B(n24794), .Z(n27908) );
  XOR U37578 ( .A(n27907), .B(n27908), .Z(n27912) );
  XOR U37579 ( .A(n27910), .B(n27912), .Z(n24788) );
  XOR U37580 ( .A(n24786), .B(n24788), .Z(n24790) );
  XOR U37581 ( .A(n24789), .B(n24790), .Z(n24781) );
  XOR U37582 ( .A(n24780), .B(n24781), .Z(n24784) );
  XOR U37583 ( .A(n24783), .B(n24784), .Z(n24776) );
  XOR U37584 ( .A(n24774), .B(n24776), .Z(n24779) );
  XOR U37585 ( .A(n24777), .B(n24779), .Z(n24769) );
  XOR U37586 ( .A(n24768), .B(n24769), .Z(n24773) );
  XOR U37587 ( .A(n24771), .B(n24773), .Z(n27917) );
  XOR U37588 ( .A(n27915), .B(n27917), .Z(n27920) );
  XOR U37589 ( .A(n27918), .B(n27920), .Z(n24763) );
  XOR U37590 ( .A(n24762), .B(n24763), .Z(n24767) );
  XOR U37591 ( .A(n24765), .B(n24767), .Z(n24757) );
  XOR U37592 ( .A(n24756), .B(n24757), .Z(n24761) );
  XOR U37593 ( .A(n24759), .B(n24761), .Z(n24754) );
  XOR U37594 ( .A(n24753), .B(n24754), .Z(n24748) );
  XOR U37595 ( .A(n24747), .B(n24748), .Z(n24752) );
  XOR U37596 ( .A(n24750), .B(n24752), .Z(n24743) );
  XOR U37597 ( .A(n24741), .B(n24743), .Z(n24745) );
  XOR U37598 ( .A(n24744), .B(n24745), .Z(n24739) );
  XOR U37599 ( .A(n24738), .B(n24739), .Z(n24734) );
  XOR U37600 ( .A(n24732), .B(n24734), .Z(n24737) );
  XOR U37601 ( .A(n24735), .B(n24737), .Z(n24727) );
  XOR U37602 ( .A(n24726), .B(n24727), .Z(n24731) );
  XOR U37603 ( .A(n24729), .B(n24731), .Z(n24724) );
  XOR U37604 ( .A(n24723), .B(n24724), .Z(n27931) );
  XOR U37605 ( .A(n27929), .B(n27931), .Z(n24721) );
  XOR U37606 ( .A(n24720), .B(n24721), .Z(n27937) );
  XOR U37607 ( .A(n27936), .B(n27937), .Z(n27941) );
  XOR U37608 ( .A(n27939), .B(n27941), .Z(n24716) );
  XOR U37609 ( .A(n24714), .B(n24716), .Z(n24718) );
  XOR U37610 ( .A(n24717), .B(n24718), .Z(n27944) );
  XOR U37611 ( .A(n27942), .B(n27944), .Z(n27946) );
  XOR U37612 ( .A(n27945), .B(n27946), .Z(n24709) );
  XOR U37613 ( .A(n24708), .B(n24709), .Z(n24712) );
  XOR U37614 ( .A(n24711), .B(n24712), .Z(n27950) );
  XOR U37615 ( .A(n27949), .B(n27950), .Z(n27954) );
  XOR U37616 ( .A(n27952), .B(n27954), .Z(n24707) );
  XOR U37617 ( .A(n24705), .B(n24707), .Z(n24699) );
  XOR U37618 ( .A(n24698), .B(n24699), .Z(n24703) );
  XOR U37619 ( .A(n24701), .B(n24703), .Z(n27957) );
  XOR U37620 ( .A(n27955), .B(n27957), .Z(n27960) );
  XOR U37621 ( .A(n27958), .B(n27960), .Z(n24696) );
  XOR U37622 ( .A(n24695), .B(n24696), .Z(n27963) );
  XOR U37623 ( .A(n27962), .B(n27963), .Z(n27967) );
  XOR U37624 ( .A(n27965), .B(n27967), .Z(n24691) );
  XOR U37625 ( .A(n24689), .B(n24691), .Z(n24693) );
  XOR U37626 ( .A(n24692), .B(n24693), .Z(n24684) );
  XOR U37627 ( .A(n24683), .B(n24684), .Z(n24688) );
  XOR U37628 ( .A(n24686), .B(n24688), .Z(n27972) );
  XOR U37629 ( .A(n27970), .B(n27972), .Z(n27974) );
  XOR U37630 ( .A(n27973), .B(n27974), .Z(n24681) );
  XOR U37631 ( .A(n24680), .B(n24681), .Z(n24676) );
  XOR U37632 ( .A(n24674), .B(n24676), .Z(n24679) );
  XOR U37633 ( .A(n24677), .B(n24679), .Z(n27979) );
  XOR U37634 ( .A(n27978), .B(n27979), .Z(n27982) );
  XOR U37635 ( .A(n27981), .B(n27982), .Z(n24673) );
  XOR U37636 ( .A(n24671), .B(n24673), .Z(n24667) );
  XOR U37637 ( .A(n24665), .B(n24667), .Z(n24669) );
  XOR U37638 ( .A(n24668), .B(n24669), .Z(n24660) );
  XOR U37639 ( .A(n24659), .B(n24660), .Z(n24664) );
  XOR U37640 ( .A(n24662), .B(n24664), .Z(n24658) );
  XOR U37641 ( .A(n24656), .B(n24658), .Z(n24651) );
  XOR U37642 ( .A(n24650), .B(n24651), .Z(n24655) );
  XOR U37643 ( .A(n24653), .B(n24655), .Z(n27988) );
  XOR U37644 ( .A(n27986), .B(n27988), .Z(n27991) );
  XOR U37645 ( .A(n27989), .B(n27991), .Z(n24644) );
  XOR U37646 ( .A(n24643), .B(n24644), .Z(n24647) );
  XOR U37647 ( .A(n24646), .B(n24647), .Z(n27995) );
  XOR U37648 ( .A(n27993), .B(n27995), .Z(n27998) );
  XOR U37649 ( .A(n27996), .B(n27998), .Z(n28005) );
  XOR U37650 ( .A(n28004), .B(n28005), .Z(n24642) );
  XOR U37651 ( .A(n24640), .B(n24642), .Z(n28003) );
  XOR U37652 ( .A(n28001), .B(n28003), .Z(n24636) );
  XOR U37653 ( .A(n24634), .B(n24636), .Z(n24638) );
  XOR U37654 ( .A(n24637), .B(n24638), .Z(n24629) );
  XOR U37655 ( .A(n24628), .B(n24629), .Z(n24633) );
  XOR U37656 ( .A(n24631), .B(n24633), .Z(n24624) );
  XOR U37657 ( .A(n24622), .B(n24624), .Z(n24626) );
  XOR U37658 ( .A(n24625), .B(n24626), .Z(n24617) );
  XOR U37659 ( .A(n24616), .B(n24617), .Z(n24621) );
  XOR U37660 ( .A(n24619), .B(n24621), .Z(n28025) );
  XOR U37661 ( .A(n28023), .B(n28025), .Z(n28027) );
  XOR U37662 ( .A(n28026), .B(n28027), .Z(n28031) );
  XOR U37663 ( .A(n28030), .B(n28031), .Z(n28035) );
  XOR U37664 ( .A(n28033), .B(n28035), .Z(n28039) );
  XOR U37665 ( .A(n28037), .B(n28039), .Z(n28041) );
  XOR U37666 ( .A(n28040), .B(n28041), .Z(n24615) );
  XOR U37667 ( .A(n24613), .B(n24615), .Z(n24609) );
  XOR U37668 ( .A(n24607), .B(n24609), .Z(n24612) );
  XOR U37669 ( .A(n24610), .B(n24612), .Z(n24602) );
  XOR U37670 ( .A(n24601), .B(n24602), .Z(n24606) );
  XOR U37671 ( .A(n24604), .B(n24606), .Z(n24600) );
  XOR U37672 ( .A(n24598), .B(n24600), .Z(n24594) );
  XOR U37673 ( .A(n24592), .B(n24594), .Z(n24596) );
  XOR U37674 ( .A(n24595), .B(n24596), .Z(n24588) );
  XOR U37675 ( .A(n24586), .B(n24588), .Z(n24591) );
  XOR U37676 ( .A(n24589), .B(n24591), .Z(n24585) );
  XOR U37677 ( .A(n24583), .B(n24585), .Z(n24578) );
  XOR U37678 ( .A(n24577), .B(n24578), .Z(n24581) );
  XOR U37679 ( .A(n24580), .B(n24581), .Z(n28049) );
  XOR U37680 ( .A(n28047), .B(n28049), .Z(n28052) );
  XOR U37681 ( .A(n28050), .B(n28052), .Z(n24571) );
  XOR U37682 ( .A(n24570), .B(n24571), .Z(n24575) );
  XOR U37683 ( .A(n24573), .B(n24575), .Z(n28056) );
  XOR U37684 ( .A(n28054), .B(n28056), .Z(n28059) );
  XOR U37685 ( .A(n28057), .B(n28059), .Z(n24566) );
  XOR U37686 ( .A(n24564), .B(n24566), .Z(n24569) );
  XOR U37687 ( .A(n24567), .B(n24569), .Z(n24560) );
  XOR U37688 ( .A(n24558), .B(n24560), .Z(n24562) );
  XOR U37689 ( .A(n24561), .B(n24562), .Z(n24556) );
  XOR U37690 ( .A(n24555), .B(n24556), .Z(n24550) );
  XOR U37691 ( .A(n24549), .B(n24550), .Z(n24554) );
  XOR U37692 ( .A(n24552), .B(n24554), .Z(n24544) );
  XOR U37693 ( .A(n24543), .B(n24544), .Z(n24547) );
  XOR U37694 ( .A(n24546), .B(n24547), .Z(n24538) );
  XOR U37695 ( .A(n24536), .B(n24538), .Z(n24541) );
  XOR U37696 ( .A(n24539), .B(n24541), .Z(n24531) );
  XOR U37697 ( .A(n24530), .B(n24531), .Z(n24534) );
  XOR U37698 ( .A(n24533), .B(n24534), .Z(n24529) );
  XOR U37699 ( .A(n24527), .B(n24529), .Z(n24522) );
  XOR U37700 ( .A(n24521), .B(n24522), .Z(n24526) );
  XOR U37701 ( .A(n24524), .B(n24526), .Z(n28066) );
  XOR U37702 ( .A(n28065), .B(n28066), .Z(n28069) );
  XOR U37703 ( .A(n28068), .B(n28069), .Z(n24517) );
  XOR U37704 ( .A(n24515), .B(n24517), .Z(n24520) );
  XOR U37705 ( .A(n24518), .B(n24520), .Z(n24510) );
  XOR U37706 ( .A(n24509), .B(n24510), .Z(n24514) );
  XOR U37707 ( .A(n24512), .B(n24514), .Z(n24505) );
  XOR U37708 ( .A(n24503), .B(n24505), .Z(n24507) );
  XOR U37709 ( .A(n24506), .B(n24507), .Z(n24501) );
  XOR U37710 ( .A(n24500), .B(n24501), .Z(n28074) );
  XOR U37711 ( .A(n28073), .B(n28074), .Z(n28078) );
  XOR U37712 ( .A(n28076), .B(n28078), .Z(n28082) );
  XOR U37713 ( .A(n28080), .B(n28082), .Z(n28084) );
  XOR U37714 ( .A(n28083), .B(n28084), .Z(n24499) );
  XOR U37715 ( .A(n24497), .B(n24499), .Z(n28088) );
  XOR U37716 ( .A(n28086), .B(n28088), .Z(n28090) );
  XOR U37717 ( .A(n28089), .B(n28090), .Z(n28094) );
  XOR U37718 ( .A(n28093), .B(n28094), .Z(n28097) );
  XOR U37719 ( .A(n28096), .B(n28097), .Z(n24496) );
  XOR U37720 ( .A(n24494), .B(n24496), .Z(n28102) );
  XOR U37721 ( .A(n28100), .B(n28102), .Z(n28104) );
  XOR U37722 ( .A(n28103), .B(n28104), .Z(n28108) );
  XOR U37723 ( .A(n28107), .B(n28108), .Z(n28112) );
  XOR U37724 ( .A(n28110), .B(n28112), .Z(n24493) );
  XOR U37725 ( .A(n24491), .B(n24493), .Z(n28116) );
  XOR U37726 ( .A(n28115), .B(n28116), .Z(n31246) );
  XOR U37727 ( .A(n31244), .B(n31246), .Z(n31251) );
  XOR U37728 ( .A(n31250), .B(n31251), .Z(n31260) );
  XOR U37729 ( .A(n31259), .B(n31260), .Z(n31267) );
  XOR U37730 ( .A(n31266), .B(n31267), .Z(n34374) );
  XOR U37731 ( .A(n34373), .B(n34374), .Z(n34388) );
  XOR U37732 ( .A(n34387), .B(n34388), .Z(n34392) );
  XOR U37733 ( .A(n34391), .B(n34392), .Z(n34400) );
  XOR U37734 ( .A(n34399), .B(n34400), .Z(n34405) );
  XOR U37735 ( .A(n34404), .B(n34405), .Z(n34421) );
  XOR U37736 ( .A(n34420), .B(n34421), .Z(n34427) );
  XOR U37737 ( .A(n34426), .B(n34427), .Z(n44350) );
  XOR U37738 ( .A(n44349), .B(n44350), .Z(n44373) );
  XOR U37739 ( .A(n44372), .B(n44373), .Z(n44409) );
  XOR U37740 ( .A(n44408), .B(n44409), .Z(n47737) );
  XOR U37741 ( .A(n47736), .B(n47737), .Z(n47754) );
  XOR U37742 ( .A(n47753), .B(n47754), .Z(n51225) );
  XOR U37743 ( .A(n51224), .B(n51225), .Z(n51241) );
  XOR U37744 ( .A(n51240), .B(n51241), .Z(n51279) );
  XOR U37745 ( .A(n51278), .B(n51279), .Z(n51313) );
  XOR U37746 ( .A(n51312), .B(n51313), .Z(n51322) );
  XOR U37747 ( .A(n51321), .B(n51322), .Z(n54894) );
  XOR U37748 ( .A(n54893), .B(n54894), .Z(n54928) );
  XOR U37749 ( .A(n54929), .B(n54928), .Z(o[0]) );
  IV U37750 ( .A(n24491), .Z(n24492) );
  NOR U37751 ( .A(n24493), .B(n24492), .Z(n31248) );
  IV U37752 ( .A(n31248), .Z(n28114) );
  IV U37753 ( .A(n24494), .Z(n24495) );
  NOR U37754 ( .A(n24496), .B(n24495), .Z(n31229) );
  IV U37755 ( .A(n24497), .Z(n24498) );
  NOR U37756 ( .A(n24499), .B(n24498), .Z(n28138) );
  IV U37757 ( .A(n24500), .Z(n24502) );
  NOR U37758 ( .A(n24502), .B(n24501), .Z(n28148) );
  IV U37759 ( .A(n24503), .Z(n24504) );
  NOR U37760 ( .A(n24505), .B(n24504), .Z(n37849) );
  IV U37761 ( .A(n24506), .Z(n24508) );
  NOR U37762 ( .A(n24508), .B(n24507), .Z(n37844) );
  NOR U37763 ( .A(n37849), .B(n37844), .Z(n34334) );
  IV U37764 ( .A(n34334), .Z(n28153) );
  IV U37765 ( .A(n24509), .Z(n24511) );
  NOR U37766 ( .A(n24511), .B(n24510), .Z(n31303) );
  IV U37767 ( .A(n24512), .Z(n24513) );
  NOR U37768 ( .A(n24514), .B(n24513), .Z(n31296) );
  NOR U37769 ( .A(n31303), .B(n31296), .Z(n28151) );
  IV U37770 ( .A(n24515), .Z(n24516) );
  NOR U37771 ( .A(n24517), .B(n24516), .Z(n28161) );
  IV U37772 ( .A(n24518), .Z(n24519) );
  NOR U37773 ( .A(n24520), .B(n24519), .Z(n28159) );
  NOR U37774 ( .A(n28161), .B(n28159), .Z(n28072) );
  IV U37775 ( .A(n24521), .Z(n24523) );
  NOR U37776 ( .A(n24523), .B(n24522), .Z(n28167) );
  IV U37777 ( .A(n24524), .Z(n24525) );
  NOR U37778 ( .A(n24526), .B(n24525), .Z(n31221) );
  NOR U37779 ( .A(n28167), .B(n31221), .Z(n28064) );
  IV U37780 ( .A(n24527), .Z(n24528) );
  NOR U37781 ( .A(n24529), .B(n24528), .Z(n28171) );
  IV U37782 ( .A(n24530), .Z(n24532) );
  NOR U37783 ( .A(n24532), .B(n24531), .Z(n31321) );
  IV U37784 ( .A(n24533), .Z(n24535) );
  NOR U37785 ( .A(n24535), .B(n24534), .Z(n31314) );
  NOR U37786 ( .A(n31321), .B(n31314), .Z(n28170) );
  IV U37787 ( .A(n24536), .Z(n24537) );
  NOR U37788 ( .A(n24538), .B(n24537), .Z(n34317) );
  IV U37789 ( .A(n24539), .Z(n24540) );
  NOR U37790 ( .A(n24541), .B(n24540), .Z(n24542) );
  NOR U37791 ( .A(n34317), .B(n24542), .Z(n31215) );
  IV U37792 ( .A(n31215), .Z(n28063) );
  IV U37793 ( .A(n24543), .Z(n24545) );
  NOR U37794 ( .A(n24545), .B(n24544), .Z(n34299) );
  IV U37795 ( .A(n24546), .Z(n24548) );
  NOR U37796 ( .A(n24548), .B(n24547), .Z(n34308) );
  NOR U37797 ( .A(n34299), .B(n34308), .Z(n31214) );
  IV U37798 ( .A(n24549), .Z(n24551) );
  NOR U37799 ( .A(n24551), .B(n24550), .Z(n28176) );
  IV U37800 ( .A(n24552), .Z(n24553) );
  NOR U37801 ( .A(n24554), .B(n24553), .Z(n28178) );
  NOR U37802 ( .A(n28176), .B(n28178), .Z(n28062) );
  IV U37803 ( .A(n24555), .Z(n24557) );
  NOR U37804 ( .A(n24557), .B(n24556), .Z(n31196) );
  IV U37805 ( .A(n24558), .Z(n24559) );
  NOR U37806 ( .A(n24560), .B(n24559), .Z(n31182) );
  IV U37807 ( .A(n24561), .Z(n24563) );
  NOR U37808 ( .A(n24563), .B(n24562), .Z(n31191) );
  NOR U37809 ( .A(n31182), .B(n31191), .Z(n28061) );
  IV U37810 ( .A(n24564), .Z(n24565) );
  NOR U37811 ( .A(n24566), .B(n24565), .Z(n31177) );
  IV U37812 ( .A(n24567), .Z(n24568) );
  NOR U37813 ( .A(n24569), .B(n24568), .Z(n31185) );
  NOR U37814 ( .A(n31177), .B(n31185), .Z(n28060) );
  IV U37815 ( .A(n24570), .Z(n24572) );
  NOR U37816 ( .A(n24572), .B(n24571), .Z(n34280) );
  IV U37817 ( .A(n24573), .Z(n24574) );
  NOR U37818 ( .A(n24575), .B(n24574), .Z(n24576) );
  NOR U37819 ( .A(n34280), .B(n24576), .Z(n28181) );
  IV U37820 ( .A(n24577), .Z(n24579) );
  NOR U37821 ( .A(n24579), .B(n24578), .Z(n28184) );
  IV U37822 ( .A(n24580), .Z(n24582) );
  NOR U37823 ( .A(n24582), .B(n24581), .Z(n28182) );
  NOR U37824 ( .A(n28184), .B(n28182), .Z(n28046) );
  IV U37825 ( .A(n24583), .Z(n24584) );
  NOR U37826 ( .A(n24585), .B(n24584), .Z(n31158) );
  IV U37827 ( .A(n24586), .Z(n24587) );
  NOR U37828 ( .A(n24588), .B(n24587), .Z(n34256) );
  IV U37829 ( .A(n24589), .Z(n24590) );
  NOR U37830 ( .A(n24591), .B(n24590), .Z(n31346) );
  NOR U37831 ( .A(n34256), .B(n31346), .Z(n31157) );
  IV U37832 ( .A(n24592), .Z(n24593) );
  NOR U37833 ( .A(n24594), .B(n24593), .Z(n28192) );
  IV U37834 ( .A(n24595), .Z(n24597) );
  NOR U37835 ( .A(n24597), .B(n24596), .Z(n28187) );
  NOR U37836 ( .A(n28192), .B(n28187), .Z(n28045) );
  IV U37837 ( .A(n24598), .Z(n24599) );
  NOR U37838 ( .A(n24600), .B(n24599), .Z(n28190) );
  IV U37839 ( .A(n24601), .Z(n24603) );
  NOR U37840 ( .A(n24603), .B(n24602), .Z(n31351) );
  IV U37841 ( .A(n24604), .Z(n24605) );
  NOR U37842 ( .A(n24606), .B(n24605), .Z(n34249) );
  NOR U37843 ( .A(n31351), .B(n34249), .Z(n28196) );
  IV U37844 ( .A(n24607), .Z(n24608) );
  NOR U37845 ( .A(n24609), .B(n24608), .Z(n28203) );
  IV U37846 ( .A(n24610), .Z(n24611) );
  NOR U37847 ( .A(n24612), .B(n24611), .Z(n28197) );
  NOR U37848 ( .A(n28203), .B(n28197), .Z(n28044) );
  IV U37849 ( .A(n24613), .Z(n24614) );
  NOR U37850 ( .A(n24615), .B(n24614), .Z(n28201) );
  IV U37851 ( .A(n24616), .Z(n24618) );
  NOR U37852 ( .A(n24618), .B(n24617), .Z(n31377) );
  IV U37853 ( .A(n24619), .Z(n24620) );
  NOR U37854 ( .A(n24621), .B(n24620), .Z(n31371) );
  NOR U37855 ( .A(n31377), .B(n31371), .Z(n31139) );
  IV U37856 ( .A(n24622), .Z(n24623) );
  NOR U37857 ( .A(n24624), .B(n24623), .Z(n37736) );
  IV U37858 ( .A(n24625), .Z(n24627) );
  NOR U37859 ( .A(n24627), .B(n24626), .Z(n34527) );
  NOR U37860 ( .A(n37736), .B(n34527), .Z(n31138) );
  IV U37861 ( .A(n24628), .Z(n24630) );
  NOR U37862 ( .A(n24630), .B(n24629), .Z(n37720) );
  IV U37863 ( .A(n24631), .Z(n24632) );
  NOR U37864 ( .A(n24633), .B(n24632), .Z(n37732) );
  NOR U37865 ( .A(n37720), .B(n37732), .Z(n31126) );
  IV U37866 ( .A(n24634), .Z(n24635) );
  NOR U37867 ( .A(n24636), .B(n24635), .Z(n34535) );
  IV U37868 ( .A(n24637), .Z(n24639) );
  NOR U37869 ( .A(n24639), .B(n24638), .Z(n37728) );
  NOR U37870 ( .A(n34535), .B(n37728), .Z(n31131) );
  IV U37871 ( .A(n24640), .Z(n24641) );
  NOR U37872 ( .A(n24642), .B(n24641), .Z(n28017) );
  IV U37873 ( .A(n28017), .Z(n28000) );
  IV U37874 ( .A(n24643), .Z(n24645) );
  NOR U37875 ( .A(n24645), .B(n24644), .Z(n37712) );
  IV U37876 ( .A(n24646), .Z(n24648) );
  NOR U37877 ( .A(n24648), .B(n24647), .Z(n24649) );
  NOR U37878 ( .A(n37712), .B(n24649), .Z(n31115) );
  IV U37879 ( .A(n24650), .Z(n24652) );
  NOR U37880 ( .A(n24652), .B(n24651), .Z(n31392) );
  IV U37881 ( .A(n24653), .Z(n24654) );
  NOR U37882 ( .A(n24655), .B(n24654), .Z(n31388) );
  NOR U37883 ( .A(n31392), .B(n31388), .Z(n31102) );
  IV U37884 ( .A(n24656), .Z(n24657) );
  NOR U37885 ( .A(n24658), .B(n24657), .Z(n31094) );
  IV U37886 ( .A(n24659), .Z(n24661) );
  NOR U37887 ( .A(n24661), .B(n24660), .Z(n34206) );
  IV U37888 ( .A(n24662), .Z(n24663) );
  NOR U37889 ( .A(n24664), .B(n24663), .Z(n31399) );
  NOR U37890 ( .A(n34206), .B(n31399), .Z(n31093) );
  IV U37891 ( .A(n24665), .Z(n24666) );
  NOR U37892 ( .A(n24667), .B(n24666), .Z(n31085) );
  IV U37893 ( .A(n24668), .Z(n24670) );
  NOR U37894 ( .A(n24670), .B(n24669), .Z(n31088) );
  NOR U37895 ( .A(n31085), .B(n31088), .Z(n27985) );
  IV U37896 ( .A(n24671), .Z(n24672) );
  NOR U37897 ( .A(n24673), .B(n24672), .Z(n31079) );
  IV U37898 ( .A(n24674), .Z(n24675) );
  NOR U37899 ( .A(n24676), .B(n24675), .Z(n28215) );
  IV U37900 ( .A(n24677), .Z(n24678) );
  NOR U37901 ( .A(n24679), .B(n24678), .Z(n31075) );
  NOR U37902 ( .A(n28215), .B(n31075), .Z(n27977) );
  IV U37903 ( .A(n24680), .Z(n24682) );
  NOR U37904 ( .A(n24682), .B(n24681), .Z(n28218) );
  IV U37905 ( .A(n24683), .Z(n24685) );
  NOR U37906 ( .A(n24685), .B(n24684), .Z(n31419) );
  IV U37907 ( .A(n24686), .Z(n24687) );
  NOR U37908 ( .A(n24688), .B(n24687), .Z(n31414) );
  NOR U37909 ( .A(n31419), .B(n31414), .Z(n28221) );
  IV U37910 ( .A(n24689), .Z(n24690) );
  NOR U37911 ( .A(n24691), .B(n24690), .Z(n28229) );
  IV U37912 ( .A(n24692), .Z(n24694) );
  NOR U37913 ( .A(n24694), .B(n24693), .Z(n28227) );
  NOR U37914 ( .A(n28229), .B(n28227), .Z(n27969) );
  IV U37915 ( .A(n24695), .Z(n24697) );
  NOR U37916 ( .A(n24697), .B(n24696), .Z(n28237) );
  IV U37917 ( .A(n24698), .Z(n24700) );
  NOR U37918 ( .A(n24700), .B(n24699), .Z(n34187) );
  IV U37919 ( .A(n24701), .Z(n24702) );
  NOR U37920 ( .A(n24703), .B(n24702), .Z(n24704) );
  NOR U37921 ( .A(n34187), .B(n24704), .Z(n31032) );
  IV U37922 ( .A(n24705), .Z(n24706) );
  NOR U37923 ( .A(n24707), .B(n24706), .Z(n28243) );
  IV U37924 ( .A(n24708), .Z(n24710) );
  NOR U37925 ( .A(n24710), .B(n24709), .Z(n28251) );
  IV U37926 ( .A(n24711), .Z(n24713) );
  NOR U37927 ( .A(n24713), .B(n24712), .Z(n28247) );
  NOR U37928 ( .A(n28251), .B(n28247), .Z(n27948) );
  IV U37929 ( .A(n24714), .Z(n24715) );
  NOR U37930 ( .A(n24716), .B(n24715), .Z(n34607) );
  IV U37931 ( .A(n24717), .Z(n24719) );
  NOR U37932 ( .A(n24719), .B(n24718), .Z(n34602) );
  NOR U37933 ( .A(n34607), .B(n34602), .Z(n34179) );
  IV U37934 ( .A(n24720), .Z(n24722) );
  NOR U37935 ( .A(n24722), .B(n24721), .Z(n27934) );
  IV U37936 ( .A(n27934), .Z(n27928) );
  IV U37937 ( .A(n24723), .Z(n24725) );
  NOR U37938 ( .A(n24725), .B(n24724), .Z(n31005) );
  IV U37939 ( .A(n24726), .Z(n24728) );
  NOR U37940 ( .A(n24728), .B(n24727), .Z(n30988) );
  IV U37941 ( .A(n24729), .Z(n24730) );
  NOR U37942 ( .A(n24731), .B(n24730), .Z(n28255) );
  NOR U37943 ( .A(n30988), .B(n28255), .Z(n27926) );
  IV U37944 ( .A(n24732), .Z(n24733) );
  NOR U37945 ( .A(n24734), .B(n24733), .Z(n28260) );
  IV U37946 ( .A(n24735), .Z(n24736) );
  NOR U37947 ( .A(n24737), .B(n24736), .Z(n28257) );
  NOR U37948 ( .A(n28260), .B(n28257), .Z(n27925) );
  IV U37949 ( .A(n24738), .Z(n24740) );
  NOR U37950 ( .A(n24740), .B(n24739), .Z(n28264) );
  IV U37951 ( .A(n24741), .Z(n24742) );
  NOR U37952 ( .A(n24743), .B(n24742), .Z(n31472) );
  IV U37953 ( .A(n24744), .Z(n24746) );
  NOR U37954 ( .A(n24746), .B(n24745), .Z(n31468) );
  NOR U37955 ( .A(n31472), .B(n31468), .Z(n28263) );
  IV U37956 ( .A(n24747), .Z(n24749) );
  NOR U37957 ( .A(n24749), .B(n24748), .Z(n30971) );
  IV U37958 ( .A(n24750), .Z(n24751) );
  NOR U37959 ( .A(n24752), .B(n24751), .Z(n28268) );
  NOR U37960 ( .A(n30971), .B(n28268), .Z(n27924) );
  IV U37961 ( .A(n24753), .Z(n24755) );
  NOR U37962 ( .A(n24755), .B(n24754), .Z(n30969) );
  IV U37963 ( .A(n24756), .Z(n24758) );
  NOR U37964 ( .A(n24758), .B(n24757), .Z(n34639) );
  IV U37965 ( .A(n24759), .Z(n24760) );
  NOR U37966 ( .A(n24761), .B(n24760), .Z(n34634) );
  NOR U37967 ( .A(n34639), .B(n34634), .Z(n30976) );
  IV U37968 ( .A(n24762), .Z(n24764) );
  NOR U37969 ( .A(n24764), .B(n24763), .Z(n30962) );
  IV U37970 ( .A(n24765), .Z(n24766) );
  NOR U37971 ( .A(n24767), .B(n24766), .Z(n28271) );
  NOR U37972 ( .A(n30962), .B(n28271), .Z(n27922) );
  IV U37973 ( .A(n24768), .Z(n24770) );
  NOR U37974 ( .A(n24770), .B(n24769), .Z(n34662) );
  IV U37975 ( .A(n24771), .Z(n24772) );
  NOR U37976 ( .A(n24773), .B(n24772), .Z(n34654) );
  NOR U37977 ( .A(n34662), .B(n34654), .Z(n30952) );
  IV U37978 ( .A(n24774), .Z(n24775) );
  NOR U37979 ( .A(n24776), .B(n24775), .Z(n34673) );
  IV U37980 ( .A(n24777), .Z(n24778) );
  NOR U37981 ( .A(n24779), .B(n24778), .Z(n34665) );
  NOR U37982 ( .A(n34673), .B(n34665), .Z(n28277) );
  IV U37983 ( .A(n24780), .Z(n24782) );
  NOR U37984 ( .A(n24782), .B(n24781), .Z(n37608) );
  IV U37985 ( .A(n24783), .Z(n24785) );
  NOR U37986 ( .A(n24785), .B(n24784), .Z(n34676) );
  NOR U37987 ( .A(n37608), .B(n34676), .Z(n30946) );
  IV U37988 ( .A(n24786), .Z(n24787) );
  NOR U37989 ( .A(n24788), .B(n24787), .Z(n30936) );
  IV U37990 ( .A(n24789), .Z(n24791) );
  NOR U37991 ( .A(n24791), .B(n24790), .Z(n28278) );
  NOR U37992 ( .A(n30936), .B(n28278), .Z(n27914) );
  IV U37993 ( .A(n24792), .Z(n24793) );
  NOR U37994 ( .A(n24794), .B(n24793), .Z(n27905) );
  IV U37995 ( .A(n27905), .Z(n27900) );
  IV U37996 ( .A(n24795), .Z(n24797) );
  NOR U37997 ( .A(n24797), .B(n24796), .Z(n28288) );
  IV U37998 ( .A(n24798), .Z(n24799) );
  NOR U37999 ( .A(n24800), .B(n24799), .Z(n28297) );
  IV U38000 ( .A(n24801), .Z(n24802) );
  NOR U38001 ( .A(n24803), .B(n24802), .Z(n28293) );
  NOR U38002 ( .A(n28297), .B(n28293), .Z(n27890) );
  IV U38003 ( .A(n24804), .Z(n24806) );
  NOR U38004 ( .A(n24806), .B(n24805), .Z(n31521) );
  IV U38005 ( .A(n24807), .Z(n24809) );
  NOR U38006 ( .A(n24809), .B(n24808), .Z(n31517) );
  NOR U38007 ( .A(n31521), .B(n31517), .Z(n28296) );
  IV U38008 ( .A(n24810), .Z(n24812) );
  NOR U38009 ( .A(n24812), .B(n24811), .Z(n28315) );
  IV U38010 ( .A(n24813), .Z(n24815) );
  NOR U38011 ( .A(n24815), .B(n24814), .Z(n34114) );
  IV U38012 ( .A(n24816), .Z(n24817) );
  NOR U38013 ( .A(n24818), .B(n24817), .Z(n34121) );
  NOR U38014 ( .A(n34114), .B(n34121), .Z(n30892) );
  IV U38015 ( .A(n30892), .Z(n27847) );
  IV U38016 ( .A(n24819), .Z(n24821) );
  NOR U38017 ( .A(n24821), .B(n24820), .Z(n30877) );
  IV U38018 ( .A(n24822), .Z(n24823) );
  NOR U38019 ( .A(n24824), .B(n24823), .Z(n30879) );
  NOR U38020 ( .A(n30877), .B(n30879), .Z(n27826) );
  IV U38021 ( .A(n24825), .Z(n24827) );
  NOR U38022 ( .A(n24827), .B(n24826), .Z(n34745) );
  IV U38023 ( .A(n24828), .Z(n24829) );
  NOR U38024 ( .A(n24830), .B(n24829), .Z(n34740) );
  NOR U38025 ( .A(n34745), .B(n34740), .Z(n30858) );
  IV U38026 ( .A(n24831), .Z(n24833) );
  NOR U38027 ( .A(n24833), .B(n24832), .Z(n30837) );
  IV U38028 ( .A(n24834), .Z(n24836) );
  NOR U38029 ( .A(n24836), .B(n24835), .Z(n30832) );
  NOR U38030 ( .A(n30837), .B(n30832), .Z(n27797) );
  IV U38031 ( .A(n24837), .Z(n24838) );
  NOR U38032 ( .A(n24839), .B(n24838), .Z(n34094) );
  IV U38033 ( .A(n24840), .Z(n24841) );
  NOR U38034 ( .A(n24842), .B(n24841), .Z(n31577) );
  NOR U38035 ( .A(n34094), .B(n31577), .Z(n30827) );
  IV U38036 ( .A(n24843), .Z(n24844) );
  NOR U38037 ( .A(n24845), .B(n24844), .Z(n30817) );
  IV U38038 ( .A(n24846), .Z(n24847) );
  NOR U38039 ( .A(n24848), .B(n24847), .Z(n28342) );
  NOR U38040 ( .A(n30817), .B(n28342), .Z(n27775) );
  IV U38041 ( .A(n24849), .Z(n24850) );
  NOR U38042 ( .A(n24851), .B(n24850), .Z(n30813) );
  IV U38043 ( .A(n24852), .Z(n24853) );
  NOR U38044 ( .A(n24854), .B(n24853), .Z(n30820) );
  NOR U38045 ( .A(n30813), .B(n30820), .Z(n27774) );
  IV U38046 ( .A(n24855), .Z(n24857) );
  NOR U38047 ( .A(n24857), .B(n24856), .Z(n30811) );
  IV U38048 ( .A(n24858), .Z(n24859) );
  NOR U38049 ( .A(n24860), .B(n24859), .Z(n28349) );
  IV U38050 ( .A(n24861), .Z(n24863) );
  NOR U38051 ( .A(n24863), .B(n24862), .Z(n28347) );
  NOR U38052 ( .A(n28349), .B(n28347), .Z(n27772) );
  IV U38053 ( .A(n24864), .Z(n24865) );
  NOR U38054 ( .A(n24866), .B(n24865), .Z(n30806) );
  IV U38055 ( .A(n24867), .Z(n24868) );
  NOR U38056 ( .A(n24869), .B(n24868), .Z(n28352) );
  NOR U38057 ( .A(n30806), .B(n28352), .Z(n27771) );
  IV U38058 ( .A(n24870), .Z(n24871) );
  NOR U38059 ( .A(n24872), .B(n24871), .Z(n31593) );
  IV U38060 ( .A(n24873), .Z(n24875) );
  NOR U38061 ( .A(n24875), .B(n24874), .Z(n31588) );
  NOR U38062 ( .A(n31593), .B(n31588), .Z(n30802) );
  IV U38063 ( .A(n24876), .Z(n24878) );
  NOR U38064 ( .A(n24878), .B(n24877), .Z(n28361) );
  IV U38065 ( .A(n24879), .Z(n24880) );
  NOR U38066 ( .A(n24881), .B(n24880), .Z(n34810) );
  IV U38067 ( .A(n24882), .Z(n24883) );
  NOR U38068 ( .A(n24884), .B(n24883), .Z(n37469) );
  NOR U38069 ( .A(n34810), .B(n37469), .Z(n34061) );
  IV U38070 ( .A(n24885), .Z(n24887) );
  NOR U38071 ( .A(n24887), .B(n24886), .Z(n34046) );
  IV U38072 ( .A(n24888), .Z(n24889) );
  NOR U38073 ( .A(n24890), .B(n24889), .Z(n34053) );
  NOR U38074 ( .A(n34046), .B(n34053), .Z(n30777) );
  IV U38075 ( .A(n24891), .Z(n24892) );
  NOR U38076 ( .A(n24893), .B(n24892), .Z(n28366) );
  IV U38077 ( .A(n24894), .Z(n24895) );
  NOR U38078 ( .A(n24896), .B(n24895), .Z(n28371) );
  IV U38079 ( .A(n24897), .Z(n24899) );
  NOR U38080 ( .A(n24899), .B(n24898), .Z(n30768) );
  NOR U38081 ( .A(n28371), .B(n30768), .Z(n27736) );
  IV U38082 ( .A(n24900), .Z(n24902) );
  NOR U38083 ( .A(n24902), .B(n24901), .Z(n28377) );
  IV U38084 ( .A(n24903), .Z(n24904) );
  NOR U38085 ( .A(n24905), .B(n24904), .Z(n28373) );
  NOR U38086 ( .A(n28377), .B(n28373), .Z(n27735) );
  IV U38087 ( .A(n24906), .Z(n24907) );
  NOR U38088 ( .A(n24908), .B(n24907), .Z(n31623) );
  IV U38089 ( .A(n24909), .Z(n24911) );
  NOR U38090 ( .A(n24911), .B(n24910), .Z(n31614) );
  NOR U38091 ( .A(n31623), .B(n31614), .Z(n28376) );
  IV U38092 ( .A(n24912), .Z(n24913) );
  NOR U38093 ( .A(n24914), .B(n24913), .Z(n31627) );
  IV U38094 ( .A(n24915), .Z(n24917) );
  NOR U38095 ( .A(n24917), .B(n24916), .Z(n24918) );
  NOR U38096 ( .A(n31627), .B(n24918), .Z(n28382) );
  IV U38097 ( .A(n24919), .Z(n24920) );
  NOR U38098 ( .A(n24921), .B(n24920), .Z(n30751) );
  IV U38099 ( .A(n24922), .Z(n24923) );
  NOR U38100 ( .A(n24924), .B(n24923), .Z(n31646) );
  IV U38101 ( .A(n24925), .Z(n24926) );
  NOR U38102 ( .A(n24927), .B(n24926), .Z(n31639) );
  NOR U38103 ( .A(n31646), .B(n31639), .Z(n30733) );
  IV U38104 ( .A(n24928), .Z(n24930) );
  NOR U38105 ( .A(n24930), .B(n24929), .Z(n30726) );
  IV U38106 ( .A(n24931), .Z(n24933) );
  NOR U38107 ( .A(n24933), .B(n24932), .Z(n28391) );
  NOR U38108 ( .A(n30726), .B(n28391), .Z(n27705) );
  IV U38109 ( .A(n24934), .Z(n24935) );
  NOR U38110 ( .A(n24936), .B(n24935), .Z(n30719) );
  IV U38111 ( .A(n24937), .Z(n24938) );
  NOR U38112 ( .A(n24939), .B(n24938), .Z(n31669) );
  IV U38113 ( .A(n24940), .Z(n24942) );
  NOR U38114 ( .A(n24942), .B(n24941), .Z(n31660) );
  NOR U38115 ( .A(n31669), .B(n31660), .Z(n30708) );
  IV U38116 ( .A(n24943), .Z(n24945) );
  NOR U38117 ( .A(n24945), .B(n24944), .Z(n30698) );
  IV U38118 ( .A(n24946), .Z(n24947) );
  NOR U38119 ( .A(n24948), .B(n24947), .Z(n30689) );
  IV U38120 ( .A(n24949), .Z(n24951) );
  NOR U38121 ( .A(n24951), .B(n24950), .Z(n30694) );
  NOR U38122 ( .A(n30689), .B(n30694), .Z(n24952) );
  IV U38123 ( .A(n24952), .Z(n27689) );
  IV U38124 ( .A(n24953), .Z(n24955) );
  NOR U38125 ( .A(n24955), .B(n24954), .Z(n30687) );
  IV U38126 ( .A(n24956), .Z(n24958) );
  NOR U38127 ( .A(n24958), .B(n24957), .Z(n34863) );
  IV U38128 ( .A(n24959), .Z(n24960) );
  NOR U38129 ( .A(n24961), .B(n24960), .Z(n34856) );
  NOR U38130 ( .A(n34863), .B(n34856), .Z(n30679) );
  IV U38131 ( .A(n24962), .Z(n24964) );
  NOR U38132 ( .A(n24964), .B(n24963), .Z(n28399) );
  IV U38133 ( .A(n24965), .Z(n24967) );
  NOR U38134 ( .A(n24967), .B(n24966), .Z(n30654) );
  IV U38135 ( .A(n24968), .Z(n24969) );
  NOR U38136 ( .A(n24970), .B(n24969), .Z(n30648) );
  NOR U38137 ( .A(n30654), .B(n30648), .Z(n28402) );
  IV U38138 ( .A(n24971), .Z(n24972) );
  NOR U38139 ( .A(n24973), .B(n24972), .Z(n30638) );
  IV U38140 ( .A(n24974), .Z(n24975) );
  NOR U38141 ( .A(n24976), .B(n24975), .Z(n30635) );
  NOR U38142 ( .A(n30638), .B(n30635), .Z(n27675) );
  IV U38143 ( .A(n24977), .Z(n24979) );
  NOR U38144 ( .A(n24979), .B(n24978), .Z(n28403) );
  IV U38145 ( .A(n24980), .Z(n24981) );
  NOR U38146 ( .A(n24982), .B(n24981), .Z(n30641) );
  NOR U38147 ( .A(n28403), .B(n30641), .Z(n27674) );
  IV U38148 ( .A(n24983), .Z(n24984) );
  NOR U38149 ( .A(n24985), .B(n24984), .Z(n27672) );
  IV U38150 ( .A(n27672), .Z(n27661) );
  IV U38151 ( .A(n24986), .Z(n24987) );
  NOR U38152 ( .A(n24988), .B(n24987), .Z(n27658) );
  IV U38153 ( .A(n27658), .Z(n27653) );
  IV U38154 ( .A(n24989), .Z(n24990) );
  NOR U38155 ( .A(n24991), .B(n24990), .Z(n28410) );
  IV U38156 ( .A(n24992), .Z(n24993) );
  NOR U38157 ( .A(n24994), .B(n24993), .Z(n27647) );
  IV U38158 ( .A(n24995), .Z(n24997) );
  NOR U38159 ( .A(n24997), .B(n24996), .Z(n30629) );
  IV U38160 ( .A(n24998), .Z(n24999) );
  NOR U38161 ( .A(n25000), .B(n24999), .Z(n28413) );
  NOR U38162 ( .A(n30629), .B(n28413), .Z(n27645) );
  IV U38163 ( .A(n25001), .Z(n25003) );
  NOR U38164 ( .A(n25003), .B(n25002), .Z(n31719) );
  IV U38165 ( .A(n25004), .Z(n25005) );
  NOR U38166 ( .A(n25006), .B(n25005), .Z(n31715) );
  NOR U38167 ( .A(n31719), .B(n31715), .Z(n30619) );
  IV U38168 ( .A(n25007), .Z(n25008) );
  NOR U38169 ( .A(n25009), .B(n25008), .Z(n30606) );
  IV U38170 ( .A(n25010), .Z(n25012) );
  NOR U38171 ( .A(n25012), .B(n25011), .Z(n27612) );
  IV U38172 ( .A(n25013), .Z(n25014) );
  NOR U38173 ( .A(n25015), .B(n25014), .Z(n27610) );
  IV U38174 ( .A(n27610), .Z(n27605) );
  IV U38175 ( .A(n25016), .Z(n25018) );
  NOR U38176 ( .A(n25018), .B(n25017), .Z(n30592) );
  IV U38177 ( .A(n25019), .Z(n25020) );
  NOR U38178 ( .A(n25021), .B(n25020), .Z(n28423) );
  IV U38179 ( .A(n25022), .Z(n25023) );
  NOR U38180 ( .A(n25024), .B(n25023), .Z(n30582) );
  NOR U38181 ( .A(n28423), .B(n30582), .Z(n27596) );
  IV U38182 ( .A(n25025), .Z(n25027) );
  NOR U38183 ( .A(n25027), .B(n25026), .Z(n33955) );
  IV U38184 ( .A(n25028), .Z(n25030) );
  NOR U38185 ( .A(n25030), .B(n25029), .Z(n31736) );
  NOR U38186 ( .A(n33955), .B(n31736), .Z(n30572) );
  IV U38187 ( .A(n25031), .Z(n25033) );
  NOR U38188 ( .A(n25033), .B(n25032), .Z(n25034) );
  IV U38189 ( .A(n25034), .Z(n27592) );
  IV U38190 ( .A(n25035), .Z(n25036) );
  NOR U38191 ( .A(n25037), .B(n25036), .Z(n27574) );
  IV U38192 ( .A(n27574), .Z(n27566) );
  IV U38193 ( .A(n25038), .Z(n25039) );
  NOR U38194 ( .A(n25040), .B(n25039), .Z(n28439) );
  IV U38195 ( .A(n25041), .Z(n25043) );
  NOR U38196 ( .A(n25043), .B(n25042), .Z(n30539) );
  IV U38197 ( .A(n25044), .Z(n25045) );
  NOR U38198 ( .A(n25046), .B(n25045), .Z(n28446) );
  IV U38199 ( .A(n25047), .Z(n25048) );
  NOR U38200 ( .A(n25049), .B(n25048), .Z(n30513) );
  IV U38201 ( .A(n25050), .Z(n25052) );
  NOR U38202 ( .A(n25052), .B(n25051), .Z(n33900) );
  IV U38203 ( .A(n25053), .Z(n25054) );
  NOR U38204 ( .A(n25055), .B(n25054), .Z(n33905) );
  NOR U38205 ( .A(n33900), .B(n33905), .Z(n28452) );
  IV U38206 ( .A(n25056), .Z(n25057) );
  NOR U38207 ( .A(n25058), .B(n25057), .Z(n30501) );
  IV U38208 ( .A(n25059), .Z(n25061) );
  NOR U38209 ( .A(n25061), .B(n25060), .Z(n30496) );
  NOR U38210 ( .A(n30501), .B(n30496), .Z(n30493) );
  IV U38211 ( .A(n25062), .Z(n25064) );
  NOR U38212 ( .A(n25064), .B(n25063), .Z(n30465) );
  IV U38213 ( .A(n25065), .Z(n25066) );
  NOR U38214 ( .A(n25067), .B(n25066), .Z(n30468) );
  NOR U38215 ( .A(n30465), .B(n30468), .Z(n27450) );
  IV U38216 ( .A(n25068), .Z(n25070) );
  NOR U38217 ( .A(n25070), .B(n25069), .Z(n28498) );
  IV U38218 ( .A(n25071), .Z(n25073) );
  NOR U38219 ( .A(n25073), .B(n25072), .Z(n28491) );
  NOR U38220 ( .A(n28498), .B(n28491), .Z(n27428) );
  IV U38221 ( .A(n25074), .Z(n25075) );
  NOR U38222 ( .A(n25076), .B(n25075), .Z(n31827) );
  IV U38223 ( .A(n25077), .Z(n25078) );
  NOR U38224 ( .A(n25079), .B(n25078), .Z(n33872) );
  NOR U38225 ( .A(n31827), .B(n33872), .Z(n28497) );
  IV U38226 ( .A(n25080), .Z(n25082) );
  NOR U38227 ( .A(n25082), .B(n25081), .Z(n35064) );
  IV U38228 ( .A(n25083), .Z(n25084) );
  NOR U38229 ( .A(n25085), .B(n25084), .Z(n28502) );
  NOR U38230 ( .A(n35064), .B(n28502), .Z(n27427) );
  IV U38231 ( .A(n25086), .Z(n25087) );
  NOR U38232 ( .A(n25088), .B(n25087), .Z(n27421) );
  IV U38233 ( .A(n25089), .Z(n25091) );
  NOR U38234 ( .A(n25091), .B(n25090), .Z(n35088) );
  IV U38235 ( .A(n25092), .Z(n25093) );
  NOR U38236 ( .A(n25094), .B(n25093), .Z(n35081) );
  NOR U38237 ( .A(n35088), .B(n35081), .Z(n30440) );
  IV U38238 ( .A(n25095), .Z(n25096) );
  NOR U38239 ( .A(n25097), .B(n25096), .Z(n40285) );
  IV U38240 ( .A(n25098), .Z(n25099) );
  NOR U38241 ( .A(n25100), .B(n25099), .Z(n25101) );
  NOR U38242 ( .A(n40285), .B(n25101), .Z(n35094) );
  IV U38243 ( .A(n25102), .Z(n25103) );
  NOR U38244 ( .A(n25104), .B(n25103), .Z(n30427) );
  IV U38245 ( .A(n25105), .Z(n25107) );
  NOR U38246 ( .A(n25107), .B(n25106), .Z(n30425) );
  NOR U38247 ( .A(n30427), .B(n30425), .Z(n27398) );
  IV U38248 ( .A(n25108), .Z(n25110) );
  NOR U38249 ( .A(n25110), .B(n25109), .Z(n28523) );
  IV U38250 ( .A(n25111), .Z(n25112) );
  NOR U38251 ( .A(n25113), .B(n25112), .Z(n30408) );
  NOR U38252 ( .A(n28523), .B(n30408), .Z(n27383) );
  IV U38253 ( .A(n25114), .Z(n25115) );
  NOR U38254 ( .A(n25116), .B(n25115), .Z(n37220) );
  IV U38255 ( .A(n25117), .Z(n25118) );
  NOR U38256 ( .A(n25119), .B(n25118), .Z(n35116) );
  NOR U38257 ( .A(n37220), .B(n35116), .Z(n30404) );
  IV U38258 ( .A(n25120), .Z(n25122) );
  NOR U38259 ( .A(n25122), .B(n25121), .Z(n25123) );
  IV U38260 ( .A(n25123), .Z(n27379) );
  IV U38261 ( .A(n25124), .Z(n25125) );
  NOR U38262 ( .A(n25126), .B(n25125), .Z(n25127) );
  IV U38263 ( .A(n25127), .Z(n27362) );
  IV U38264 ( .A(n25128), .Z(n25130) );
  NOR U38265 ( .A(n25130), .B(n25129), .Z(n30379) );
  IV U38266 ( .A(n25131), .Z(n25132) );
  NOR U38267 ( .A(n25133), .B(n25132), .Z(n30384) );
  NOR U38268 ( .A(n30379), .B(n30384), .Z(n31905) );
  IV U38269 ( .A(n25134), .Z(n25136) );
  NOR U38270 ( .A(n25136), .B(n25135), .Z(n28534) );
  IV U38271 ( .A(n25137), .Z(n25138) );
  NOR U38272 ( .A(n25139), .B(n25138), .Z(n28529) );
  NOR U38273 ( .A(n28534), .B(n28529), .Z(n27342) );
  IV U38274 ( .A(n25140), .Z(n25141) );
  NOR U38275 ( .A(n25142), .B(n25141), .Z(n31921) );
  IV U38276 ( .A(n25143), .Z(n25144) );
  NOR U38277 ( .A(n25145), .B(n25144), .Z(n33850) );
  NOR U38278 ( .A(n31921), .B(n33850), .Z(n28533) );
  IV U38279 ( .A(n25146), .Z(n25148) );
  NOR U38280 ( .A(n25148), .B(n25147), .Z(n30362) );
  IV U38281 ( .A(n25149), .Z(n25151) );
  NOR U38282 ( .A(n25151), .B(n25150), .Z(n30365) );
  NOR U38283 ( .A(n30362), .B(n30365), .Z(n27334) );
  IV U38284 ( .A(n25152), .Z(n25153) );
  NOR U38285 ( .A(n25154), .B(n25153), .Z(n28544) );
  IV U38286 ( .A(n25155), .Z(n25156) );
  NOR U38287 ( .A(n25157), .B(n25156), .Z(n30346) );
  NOR U38288 ( .A(n28544), .B(n30346), .Z(n27333) );
  IV U38289 ( .A(n25158), .Z(n25159) );
  NOR U38290 ( .A(n25160), .B(n25159), .Z(n28542) );
  IV U38291 ( .A(n25161), .Z(n25162) );
  NOR U38292 ( .A(n25163), .B(n25162), .Z(n28549) );
  IV U38293 ( .A(n25164), .Z(n25165) );
  NOR U38294 ( .A(n25166), .B(n25165), .Z(n30340) );
  NOR U38295 ( .A(n28549), .B(n30340), .Z(n27325) );
  IV U38296 ( .A(n25167), .Z(n25169) );
  NOR U38297 ( .A(n25169), .B(n25168), .Z(n28552) );
  IV U38298 ( .A(n25170), .Z(n25171) );
  NOR U38299 ( .A(n25172), .B(n25171), .Z(n37142) );
  IV U38300 ( .A(n25173), .Z(n25174) );
  NOR U38301 ( .A(n25175), .B(n25174), .Z(n37152) );
  NOR U38302 ( .A(n37142), .B(n37152), .Z(n33828) );
  IV U38303 ( .A(n25176), .Z(n25177) );
  NOR U38304 ( .A(n25178), .B(n25177), .Z(n27312) );
  IV U38305 ( .A(n25179), .Z(n25180) );
  NOR U38306 ( .A(n25181), .B(n25180), .Z(n30328) );
  IV U38307 ( .A(n25182), .Z(n25183) );
  NOR U38308 ( .A(n25184), .B(n25183), .Z(n27295) );
  IV U38309 ( .A(n27295), .Z(n27290) );
  IV U38310 ( .A(n25185), .Z(n25187) );
  NOR U38311 ( .A(n25187), .B(n25186), .Z(n28568) );
  IV U38312 ( .A(n25188), .Z(n25190) );
  NOR U38313 ( .A(n25190), .B(n25189), .Z(n31948) );
  IV U38314 ( .A(n25191), .Z(n25193) );
  NOR U38315 ( .A(n25193), .B(n25192), .Z(n33799) );
  NOR U38316 ( .A(n31948), .B(n33799), .Z(n30311) );
  IV U38317 ( .A(n25194), .Z(n25195) );
  NOR U38318 ( .A(n25196), .B(n25195), .Z(n30300) );
  IV U38319 ( .A(n25197), .Z(n25198) );
  NOR U38320 ( .A(n25199), .B(n25198), .Z(n28574) );
  NOR U38321 ( .A(n30300), .B(n28574), .Z(n27281) );
  IV U38322 ( .A(n25200), .Z(n25201) );
  NOR U38323 ( .A(n25202), .B(n25201), .Z(n30290) );
  IV U38324 ( .A(n25203), .Z(n25204) );
  NOR U38325 ( .A(n25205), .B(n25204), .Z(n30303) );
  NOR U38326 ( .A(n30290), .B(n30303), .Z(n27280) );
  IV U38327 ( .A(n25206), .Z(n25207) );
  NOR U38328 ( .A(n25208), .B(n25207), .Z(n30293) );
  IV U38329 ( .A(n25209), .Z(n25211) );
  NOR U38330 ( .A(n25211), .B(n25210), .Z(n31969) );
  IV U38331 ( .A(n25212), .Z(n25213) );
  NOR U38332 ( .A(n25214), .B(n25213), .Z(n31965) );
  NOR U38333 ( .A(n31969), .B(n31965), .Z(n30292) );
  IV U38334 ( .A(n25215), .Z(n25217) );
  NOR U38335 ( .A(n25217), .B(n25216), .Z(n28588) );
  IV U38336 ( .A(n25218), .Z(n25220) );
  NOR U38337 ( .A(n25220), .B(n25219), .Z(n38520) );
  IV U38338 ( .A(n25221), .Z(n25222) );
  NOR U38339 ( .A(n25223), .B(n25222), .Z(n25224) );
  NOR U38340 ( .A(n38520), .B(n25224), .Z(n35227) );
  IV U38341 ( .A(n35227), .Z(n27250) );
  IV U38342 ( .A(n25225), .Z(n25226) );
  NOR U38343 ( .A(n25227), .B(n25226), .Z(n33784) );
  IV U38344 ( .A(n25228), .Z(n25229) );
  NOR U38345 ( .A(n25230), .B(n25229), .Z(n31999) );
  NOR U38346 ( .A(n33784), .B(n31999), .Z(n28592) );
  IV U38347 ( .A(n25231), .Z(n25232) );
  NOR U38348 ( .A(n25233), .B(n25232), .Z(n28600) );
  IV U38349 ( .A(n25234), .Z(n25236) );
  NOR U38350 ( .A(n25236), .B(n25235), .Z(n25237) );
  IV U38351 ( .A(n25237), .Z(n27224) );
  IV U38352 ( .A(n25238), .Z(n25239) );
  NOR U38353 ( .A(n25240), .B(n25239), .Z(n28609) );
  IV U38354 ( .A(n25241), .Z(n25243) );
  NOR U38355 ( .A(n25243), .B(n25242), .Z(n32020) );
  IV U38356 ( .A(n25244), .Z(n25245) );
  NOR U38357 ( .A(n25246), .B(n25245), .Z(n33771) );
  NOR U38358 ( .A(n32020), .B(n33771), .Z(n28613) );
  IV U38359 ( .A(n25247), .Z(n25248) );
  NOR U38360 ( .A(n25249), .B(n25248), .Z(n28619) );
  IV U38361 ( .A(n25250), .Z(n25252) );
  NOR U38362 ( .A(n25252), .B(n25251), .Z(n28617) );
  NOR U38363 ( .A(n28619), .B(n28617), .Z(n27207) );
  IV U38364 ( .A(n25253), .Z(n25255) );
  NOR U38365 ( .A(n25255), .B(n25254), .Z(n30235) );
  IV U38366 ( .A(n25256), .Z(n25258) );
  NOR U38367 ( .A(n25258), .B(n25257), .Z(n30231) );
  NOR U38368 ( .A(n30235), .B(n30231), .Z(n30227) );
  IV U38369 ( .A(n25259), .Z(n25260) );
  NOR U38370 ( .A(n25261), .B(n25260), .Z(n28629) );
  IV U38371 ( .A(n25262), .Z(n25264) );
  NOR U38372 ( .A(n25264), .B(n25263), .Z(n28638) );
  IV U38373 ( .A(n25265), .Z(n25266) );
  NOR U38374 ( .A(n25267), .B(n25266), .Z(n28652) );
  IV U38375 ( .A(n25268), .Z(n25270) );
  NOR U38376 ( .A(n25270), .B(n25269), .Z(n28644) );
  NOR U38377 ( .A(n28652), .B(n28644), .Z(n25271) );
  IV U38378 ( .A(n25271), .Z(n27171) );
  IV U38379 ( .A(n25272), .Z(n25273) );
  NOR U38380 ( .A(n25274), .B(n25273), .Z(n28647) );
  IV U38381 ( .A(n25275), .Z(n25276) );
  NOR U38382 ( .A(n25277), .B(n25276), .Z(n33724) );
  IV U38383 ( .A(n25278), .Z(n25279) );
  NOR U38384 ( .A(n25280), .B(n25279), .Z(n33737) );
  NOR U38385 ( .A(n33724), .B(n33737), .Z(n28656) );
  IV U38386 ( .A(n25281), .Z(n25283) );
  NOR U38387 ( .A(n25283), .B(n25282), .Z(n25284) );
  IV U38388 ( .A(n25284), .Z(n27159) );
  IV U38389 ( .A(n25285), .Z(n25286) );
  NOR U38390 ( .A(n25287), .B(n25286), .Z(n33714) );
  IV U38391 ( .A(n25288), .Z(n25289) );
  NOR U38392 ( .A(n25290), .B(n25289), .Z(n25291) );
  NOR U38393 ( .A(n33714), .B(n25291), .Z(n30212) );
  IV U38394 ( .A(n25292), .Z(n25293) );
  NOR U38395 ( .A(n25294), .B(n25293), .Z(n28670) );
  IV U38396 ( .A(n25295), .Z(n25296) );
  NOR U38397 ( .A(n25297), .B(n25296), .Z(n28668) );
  NOR U38398 ( .A(n28670), .B(n28668), .Z(n27123) );
  IV U38399 ( .A(n25298), .Z(n25299) );
  NOR U38400 ( .A(n25300), .B(n25299), .Z(n28675) );
  IV U38401 ( .A(n25301), .Z(n25303) );
  NOR U38402 ( .A(n25303), .B(n25302), .Z(n28673) );
  NOR U38403 ( .A(n28675), .B(n28673), .Z(n27115) );
  IV U38404 ( .A(n25304), .Z(n25305) );
  NOR U38405 ( .A(n25306), .B(n25305), .Z(n30154) );
  IV U38406 ( .A(n25307), .Z(n25309) );
  NOR U38407 ( .A(n25309), .B(n25308), .Z(n30165) );
  NOR U38408 ( .A(n30154), .B(n30165), .Z(n27107) );
  IV U38409 ( .A(n25310), .Z(n25311) );
  NOR U38410 ( .A(n25312), .B(n25311), .Z(n27099) );
  IV U38411 ( .A(n25313), .Z(n25314) );
  NOR U38412 ( .A(n25315), .B(n25314), .Z(n27095) );
  IV U38413 ( .A(n25316), .Z(n25318) );
  NOR U38414 ( .A(n25318), .B(n25317), .Z(n25319) );
  IV U38415 ( .A(n25319), .Z(n28685) );
  IV U38416 ( .A(n25320), .Z(n25321) );
  NOR U38417 ( .A(n25322), .B(n25321), .Z(n30139) );
  IV U38418 ( .A(n25323), .Z(n25324) );
  NOR U38419 ( .A(n25325), .B(n25324), .Z(n28693) );
  NOR U38420 ( .A(n30139), .B(n28693), .Z(n27077) );
  IV U38421 ( .A(n25326), .Z(n25327) );
  NOR U38422 ( .A(n25328), .B(n25327), .Z(n30135) );
  IV U38423 ( .A(n25329), .Z(n25331) );
  NOR U38424 ( .A(n25331), .B(n25330), .Z(n27071) );
  IV U38425 ( .A(n27071), .Z(n27063) );
  IV U38426 ( .A(n25332), .Z(n25333) );
  NOR U38427 ( .A(n25334), .B(n25333), .Z(n28696) );
  IV U38428 ( .A(n25335), .Z(n25336) );
  NOR U38429 ( .A(n25337), .B(n25336), .Z(n32087) );
  IV U38430 ( .A(n25338), .Z(n25339) );
  NOR U38431 ( .A(n25340), .B(n25339), .Z(n33632) );
  NOR U38432 ( .A(n32087), .B(n33632), .Z(n28700) );
  IV U38433 ( .A(n25341), .Z(n25343) );
  NOR U38434 ( .A(n25343), .B(n25342), .Z(n28707) );
  IV U38435 ( .A(n25344), .Z(n25345) );
  NOR U38436 ( .A(n25346), .B(n25345), .Z(n28701) );
  NOR U38437 ( .A(n28707), .B(n28701), .Z(n27061) );
  IV U38438 ( .A(n25347), .Z(n25349) );
  NOR U38439 ( .A(n25349), .B(n25348), .Z(n27059) );
  IV U38440 ( .A(n27059), .Z(n27054) );
  IV U38441 ( .A(n25350), .Z(n25352) );
  NOR U38442 ( .A(n25352), .B(n25351), .Z(n28711) );
  IV U38443 ( .A(n25353), .Z(n25354) );
  NOR U38444 ( .A(n25355), .B(n25354), .Z(n28720) );
  IV U38445 ( .A(n25356), .Z(n25357) );
  NOR U38446 ( .A(n25358), .B(n25357), .Z(n28716) );
  NOR U38447 ( .A(n28720), .B(n28716), .Z(n27045) );
  IV U38448 ( .A(n25359), .Z(n25360) );
  NOR U38449 ( .A(n25361), .B(n25360), .Z(n35405) );
  IV U38450 ( .A(n25362), .Z(n25363) );
  NOR U38451 ( .A(n25364), .B(n25363), .Z(n35393) );
  NOR U38452 ( .A(n35405), .B(n35393), .Z(n30120) );
  IV U38453 ( .A(n25365), .Z(n25367) );
  NOR U38454 ( .A(n25367), .B(n25366), .Z(n28722) );
  IV U38455 ( .A(n25368), .Z(n25369) );
  NOR U38456 ( .A(n25370), .B(n25369), .Z(n30121) );
  NOR U38457 ( .A(n28722), .B(n30121), .Z(n27044) );
  IV U38458 ( .A(n25371), .Z(n25373) );
  NOR U38459 ( .A(n25373), .B(n25372), .Z(n28736) );
  IV U38460 ( .A(n25374), .Z(n25375) );
  NOR U38461 ( .A(n25376), .B(n25375), .Z(n28733) );
  NOR U38462 ( .A(n28736), .B(n28733), .Z(n27022) );
  IV U38463 ( .A(n25377), .Z(n25379) );
  NOR U38464 ( .A(n25379), .B(n25378), .Z(n27017) );
  IV U38465 ( .A(n27017), .Z(n27008) );
  IV U38466 ( .A(n25380), .Z(n25381) );
  NOR U38467 ( .A(n25382), .B(n25381), .Z(n27005) );
  IV U38468 ( .A(n27005), .Z(n26994) );
  IV U38469 ( .A(n25383), .Z(n25385) );
  NOR U38470 ( .A(n25385), .B(n25384), .Z(n28744) );
  IV U38471 ( .A(n25386), .Z(n25387) );
  NOR U38472 ( .A(n25388), .B(n25387), .Z(n30089) );
  NOR U38473 ( .A(n28744), .B(n30089), .Z(n26986) );
  IV U38474 ( .A(n25389), .Z(n25391) );
  NOR U38475 ( .A(n25391), .B(n25390), .Z(n32148) );
  IV U38476 ( .A(n25392), .Z(n25394) );
  NOR U38477 ( .A(n25394), .B(n25393), .Z(n32143) );
  NOR U38478 ( .A(n32148), .B(n32143), .Z(n28743) );
  IV U38479 ( .A(n25395), .Z(n25397) );
  NOR U38480 ( .A(n25397), .B(n25396), .Z(n28764) );
  IV U38481 ( .A(n25398), .Z(n25399) );
  NOR U38482 ( .A(n25400), .B(n25399), .Z(n25401) );
  IV U38483 ( .A(n25401), .Z(n26960) );
  IV U38484 ( .A(n25402), .Z(n25404) );
  NOR U38485 ( .A(n25404), .B(n25403), .Z(n32165) );
  IV U38486 ( .A(n25405), .Z(n25406) );
  NOR U38487 ( .A(n25407), .B(n25406), .Z(n33563) );
  NOR U38488 ( .A(n32165), .B(n33563), .Z(n28775) );
  IV U38489 ( .A(n25408), .Z(n25410) );
  NOR U38490 ( .A(n25410), .B(n25409), .Z(n30056) );
  IV U38491 ( .A(n25411), .Z(n25412) );
  NOR U38492 ( .A(n25413), .B(n25412), .Z(n30052) );
  NOR U38493 ( .A(n30056), .B(n30052), .Z(n26938) );
  IV U38494 ( .A(n25414), .Z(n25416) );
  NOR U38495 ( .A(n25416), .B(n25415), .Z(n26934) );
  IV U38496 ( .A(n25417), .Z(n25418) );
  NOR U38497 ( .A(n25419), .B(n25418), .Z(n26917) );
  IV U38498 ( .A(n26917), .Z(n26906) );
  IV U38499 ( .A(n25420), .Z(n25421) );
  NOR U38500 ( .A(n25422), .B(n25421), .Z(n28778) );
  IV U38501 ( .A(n25423), .Z(n25424) );
  NOR U38502 ( .A(n25425), .B(n25424), .Z(n28780) );
  NOR U38503 ( .A(n28778), .B(n28780), .Z(n26905) );
  IV U38504 ( .A(n25426), .Z(n25427) );
  NOR U38505 ( .A(n25428), .B(n25427), .Z(n30030) );
  IV U38506 ( .A(n25429), .Z(n25431) );
  NOR U38507 ( .A(n25431), .B(n25430), .Z(n26891) );
  IV U38508 ( .A(n26891), .Z(n26883) );
  IV U38509 ( .A(n25432), .Z(n25433) );
  NOR U38510 ( .A(n25434), .B(n25433), .Z(n30012) );
  IV U38511 ( .A(n25435), .Z(n25436) );
  NOR U38512 ( .A(n25437), .B(n25436), .Z(n30015) );
  IV U38513 ( .A(n25438), .Z(n25439) );
  NOR U38514 ( .A(n25440), .B(n25439), .Z(n33532) );
  IV U38515 ( .A(n25441), .Z(n25443) );
  NOR U38516 ( .A(n25443), .B(n25442), .Z(n32202) );
  NOR U38517 ( .A(n33532), .B(n32202), .Z(n28788) );
  IV U38518 ( .A(n25444), .Z(n25446) );
  NOR U38519 ( .A(n25446), .B(n25445), .Z(n30000) );
  IV U38520 ( .A(n25447), .Z(n25448) );
  NOR U38521 ( .A(n25449), .B(n25448), .Z(n28789) );
  NOR U38522 ( .A(n30000), .B(n28789), .Z(n26882) );
  IV U38523 ( .A(n25450), .Z(n25452) );
  NOR U38524 ( .A(n25452), .B(n25451), .Z(n30003) );
  IV U38525 ( .A(n25453), .Z(n25455) );
  NOR U38526 ( .A(n25455), .B(n25454), .Z(n33504) );
  IV U38527 ( .A(n25456), .Z(n25457) );
  NOR U38528 ( .A(n25458), .B(n25457), .Z(n33514) );
  NOR U38529 ( .A(n33504), .B(n33514), .Z(n29996) );
  IV U38530 ( .A(n25459), .Z(n25460) );
  NOR U38531 ( .A(n25461), .B(n25460), .Z(n32213) );
  IV U38532 ( .A(n25462), .Z(n25464) );
  NOR U38533 ( .A(n25464), .B(n25463), .Z(n32206) );
  NOR U38534 ( .A(n32213), .B(n32206), .Z(n29994) );
  IV U38535 ( .A(n25465), .Z(n25466) );
  NOR U38536 ( .A(n25467), .B(n25466), .Z(n28802) );
  IV U38537 ( .A(n25468), .Z(n25470) );
  NOR U38538 ( .A(n25470), .B(n25469), .Z(n29970) );
  IV U38539 ( .A(n25471), .Z(n25472) );
  NOR U38540 ( .A(n25473), .B(n25472), .Z(n29953) );
  IV U38541 ( .A(n25474), .Z(n25476) );
  NOR U38542 ( .A(n25476), .B(n25475), .Z(n28810) );
  NOR U38543 ( .A(n29953), .B(n28810), .Z(n26833) );
  NOR U38544 ( .A(n25477), .B(n25478), .Z(n25482) );
  IV U38545 ( .A(n25478), .Z(n25479) );
  NOR U38546 ( .A(n25480), .B(n25479), .Z(n36814) );
  NOR U38547 ( .A(n36814), .B(n36821), .Z(n25481) );
  NOR U38548 ( .A(n25482), .B(n25481), .Z(n29945) );
  IV U38549 ( .A(n25483), .Z(n25485) );
  NOR U38550 ( .A(n25485), .B(n25484), .Z(n28819) );
  NOR U38551 ( .A(n25487), .B(n25486), .Z(n28815) );
  NOR U38552 ( .A(n28819), .B(n28815), .Z(n25488) );
  IV U38553 ( .A(n25488), .Z(n26813) );
  IV U38554 ( .A(n25489), .Z(n25491) );
  NOR U38555 ( .A(n25491), .B(n25490), .Z(n28821) );
  IV U38556 ( .A(n25492), .Z(n25493) );
  NOR U38557 ( .A(n25494), .B(n25493), .Z(n33473) );
  IV U38558 ( .A(n25495), .Z(n25496) );
  NOR U38559 ( .A(n25497), .B(n25496), .Z(n32277) );
  NOR U38560 ( .A(n33473), .B(n32277), .Z(n28825) );
  IV U38561 ( .A(n25498), .Z(n25499) );
  NOR U38562 ( .A(n25500), .B(n25499), .Z(n28833) );
  IV U38563 ( .A(n25501), .Z(n25503) );
  NOR U38564 ( .A(n25503), .B(n25502), .Z(n29923) );
  IV U38565 ( .A(n25504), .Z(n25505) );
  NOR U38566 ( .A(n25506), .B(n25505), .Z(n29935) );
  NOR U38567 ( .A(n29923), .B(n29935), .Z(n26781) );
  IV U38568 ( .A(n25507), .Z(n25509) );
  NOR U38569 ( .A(n25509), .B(n25508), .Z(n33438) );
  IV U38570 ( .A(n25510), .Z(n25511) );
  NOR U38571 ( .A(n25512), .B(n25511), .Z(n25513) );
  NOR U38572 ( .A(n33438), .B(n25513), .Z(n29925) );
  IV U38573 ( .A(n25514), .Z(n25516) );
  NOR U38574 ( .A(n25516), .B(n25515), .Z(n29906) );
  IV U38575 ( .A(n25517), .Z(n25518) );
  NOR U38576 ( .A(n25519), .B(n25518), .Z(n29917) );
  NOR U38577 ( .A(n29906), .B(n29917), .Z(n26767) );
  IV U38578 ( .A(n25520), .Z(n25522) );
  NOR U38579 ( .A(n25522), .B(n25521), .Z(n33427) );
  IV U38580 ( .A(n25523), .Z(n25524) );
  NOR U38581 ( .A(n25525), .B(n25524), .Z(n32295) );
  NOR U38582 ( .A(n33427), .B(n32295), .Z(n29905) );
  IV U38583 ( .A(n25526), .Z(n25528) );
  NOR U38584 ( .A(n25528), .B(n25527), .Z(n28852) );
  IV U38585 ( .A(n25529), .Z(n25531) );
  NOR U38586 ( .A(n25531), .B(n25530), .Z(n28846) );
  NOR U38587 ( .A(n28852), .B(n28846), .Z(n26766) );
  IV U38588 ( .A(n25532), .Z(n25533) );
  NOR U38589 ( .A(n25534), .B(n25533), .Z(n28850) );
  IV U38590 ( .A(n25535), .Z(n25537) );
  NOR U38591 ( .A(n25537), .B(n25536), .Z(n28863) );
  IV U38592 ( .A(n25538), .Z(n25539) );
  NOR U38593 ( .A(n25540), .B(n25539), .Z(n32309) );
  IV U38594 ( .A(n25541), .Z(n25543) );
  NOR U38595 ( .A(n25543), .B(n25542), .Z(n33410) );
  NOR U38596 ( .A(n32309), .B(n33410), .Z(n29889) );
  IV U38597 ( .A(n25544), .Z(n25546) );
  NOR U38598 ( .A(n25546), .B(n25545), .Z(n32319) );
  IV U38599 ( .A(n25547), .Z(n25548) );
  NOR U38600 ( .A(n25549), .B(n25548), .Z(n25550) );
  NOR U38601 ( .A(n32319), .B(n25550), .Z(n29887) );
  IV U38602 ( .A(n25551), .Z(n25552) );
  NOR U38603 ( .A(n25553), .B(n25552), .Z(n29870) );
  IV U38604 ( .A(n25554), .Z(n25555) );
  NOR U38605 ( .A(n25556), .B(n25555), .Z(n29884) );
  NOR U38606 ( .A(n29870), .B(n29884), .Z(n26744) );
  IV U38607 ( .A(n25557), .Z(n25559) );
  NOR U38608 ( .A(n25559), .B(n25558), .Z(n29874) );
  IV U38609 ( .A(n25560), .Z(n25562) );
  NOR U38610 ( .A(n25562), .B(n25561), .Z(n29876) );
  NOR U38611 ( .A(n29874), .B(n29876), .Z(n26743) );
  IV U38612 ( .A(n25563), .Z(n25564) );
  NOR U38613 ( .A(n25565), .B(n25564), .Z(n35611) );
  IV U38614 ( .A(n25566), .Z(n25567) );
  NOR U38615 ( .A(n25568), .B(n25567), .Z(n35606) );
  NOR U38616 ( .A(n35611), .B(n35606), .Z(n33398) );
  IV U38617 ( .A(n33398), .Z(n28868) );
  IV U38618 ( .A(n25569), .Z(n25571) );
  NOR U38619 ( .A(n25571), .B(n25570), .Z(n33386) );
  IV U38620 ( .A(n25572), .Z(n25573) );
  NOR U38621 ( .A(n25574), .B(n25573), .Z(n33392) );
  NOR U38622 ( .A(n33386), .B(n33392), .Z(n28866) );
  IV U38623 ( .A(n25575), .Z(n25576) );
  NOR U38624 ( .A(n25577), .B(n25576), .Z(n28873) );
  IV U38625 ( .A(n25578), .Z(n25579) );
  NOR U38626 ( .A(n25580), .B(n25579), .Z(n28871) );
  NOR U38627 ( .A(n28873), .B(n28871), .Z(n26742) );
  IV U38628 ( .A(n25581), .Z(n25583) );
  NOR U38629 ( .A(n25583), .B(n25582), .Z(n25584) );
  IV U38630 ( .A(n25584), .Z(n26737) );
  IV U38631 ( .A(n25585), .Z(n25587) );
  NOR U38632 ( .A(n25587), .B(n25586), .Z(n26720) );
  IV U38633 ( .A(n25588), .Z(n25590) );
  NOR U38634 ( .A(n25590), .B(n25589), .Z(n28884) );
  IV U38635 ( .A(n25591), .Z(n25592) );
  NOR U38636 ( .A(n25593), .B(n25592), .Z(n28881) );
  NOR U38637 ( .A(n28884), .B(n28881), .Z(n26719) );
  IV U38638 ( .A(n25594), .Z(n25595) );
  NOR U38639 ( .A(n25596), .B(n25595), .Z(n29857) );
  IV U38640 ( .A(n25597), .Z(n25599) );
  NOR U38641 ( .A(n25599), .B(n25598), .Z(n29861) );
  NOR U38642 ( .A(n29857), .B(n29861), .Z(n26718) );
  IV U38643 ( .A(n25600), .Z(n25602) );
  NOR U38644 ( .A(n25602), .B(n25601), .Z(n29851) );
  IV U38645 ( .A(n25603), .Z(n25604) );
  NOR U38646 ( .A(n25605), .B(n25604), .Z(n28887) );
  NOR U38647 ( .A(n29851), .B(n28887), .Z(n26717) );
  IV U38648 ( .A(n25606), .Z(n25608) );
  NOR U38649 ( .A(n25608), .B(n25607), .Z(n29847) );
  IV U38650 ( .A(n25609), .Z(n25610) );
  NOR U38651 ( .A(n25611), .B(n25610), .Z(n32339) );
  IV U38652 ( .A(n25612), .Z(n25613) );
  NOR U38653 ( .A(n25614), .B(n25613), .Z(n32333) );
  NOR U38654 ( .A(n32339), .B(n32333), .Z(n29846) );
  IV U38655 ( .A(n25615), .Z(n25616) );
  NOR U38656 ( .A(n25617), .B(n25616), .Z(n29842) );
  IV U38657 ( .A(n25618), .Z(n25620) );
  NOR U38658 ( .A(n25620), .B(n25619), .Z(n28890) );
  NOR U38659 ( .A(n29842), .B(n28890), .Z(n26716) );
  IV U38660 ( .A(n25621), .Z(n25622) );
  NOR U38661 ( .A(n25623), .B(n25622), .Z(n28894) );
  IV U38662 ( .A(n25624), .Z(n25626) );
  NOR U38663 ( .A(n25626), .B(n25625), .Z(n28897) );
  IV U38664 ( .A(n25627), .Z(n25629) );
  NOR U38665 ( .A(n25629), .B(n25628), .Z(n28899) );
  NOR U38666 ( .A(n28897), .B(n28899), .Z(n26715) );
  IV U38667 ( .A(n25630), .Z(n25631) );
  NOR U38668 ( .A(n25632), .B(n25631), .Z(n28906) );
  IV U38669 ( .A(n25633), .Z(n25634) );
  NOR U38670 ( .A(n25635), .B(n25634), .Z(n28903) );
  NOR U38671 ( .A(n28906), .B(n28903), .Z(n26714) );
  IV U38672 ( .A(n25636), .Z(n25637) );
  NOR U38673 ( .A(n25638), .B(n25637), .Z(n28908) );
  IV U38674 ( .A(n25639), .Z(n25640) );
  NOR U38675 ( .A(n25641), .B(n25640), .Z(n29803) );
  IV U38676 ( .A(n25642), .Z(n25643) );
  NOR U38677 ( .A(n25644), .B(n25643), .Z(n35681) );
  IV U38678 ( .A(n25645), .Z(n25646) );
  NOR U38679 ( .A(n25647), .B(n25646), .Z(n35675) );
  NOR U38680 ( .A(n35681), .B(n35675), .Z(n29816) );
  IV U38681 ( .A(n29816), .Z(n26692) );
  IV U38682 ( .A(n25648), .Z(n25650) );
  NOR U38683 ( .A(n25650), .B(n25649), .Z(n32368) );
  IV U38684 ( .A(n25651), .Z(n25652) );
  NOR U38685 ( .A(n25653), .B(n25652), .Z(n32364) );
  NOR U38686 ( .A(n32368), .B(n32364), .Z(n29806) );
  IV U38687 ( .A(n25654), .Z(n25655) );
  NOR U38688 ( .A(n25656), .B(n25655), .Z(n28916) );
  IV U38689 ( .A(n25657), .Z(n25658) );
  NOR U38690 ( .A(n25659), .B(n25658), .Z(n28911) );
  NOR U38691 ( .A(n28916), .B(n28911), .Z(n26691) );
  IV U38692 ( .A(n25660), .Z(n25662) );
  NOR U38693 ( .A(n25662), .B(n25661), .Z(n33319) );
  IV U38694 ( .A(n25663), .Z(n25664) );
  NOR U38695 ( .A(n25665), .B(n25664), .Z(n32392) );
  NOR U38696 ( .A(n33319), .B(n32392), .Z(n32378) );
  IV U38697 ( .A(n25666), .Z(n25667) );
  NOR U38698 ( .A(n25668), .B(n25667), .Z(n29784) );
  IV U38699 ( .A(n25669), .Z(n25670) );
  NOR U38700 ( .A(n25671), .B(n25670), .Z(n28920) );
  NOR U38701 ( .A(n29784), .B(n28920), .Z(n26684) );
  IV U38702 ( .A(n25672), .Z(n25674) );
  NOR U38703 ( .A(n25674), .B(n25673), .Z(n29787) );
  IV U38704 ( .A(n25675), .Z(n25677) );
  NOR U38705 ( .A(n25677), .B(n25676), .Z(n29779) );
  NOR U38706 ( .A(n29787), .B(n29779), .Z(n25678) );
  IV U38707 ( .A(n25678), .Z(n26683) );
  IV U38708 ( .A(n25679), .Z(n25680) );
  NOR U38709 ( .A(n25681), .B(n25680), .Z(n29790) );
  IV U38710 ( .A(n25682), .Z(n25683) );
  NOR U38711 ( .A(n25684), .B(n25683), .Z(n33298) );
  IV U38712 ( .A(n25685), .Z(n25686) );
  NOR U38713 ( .A(n25687), .B(n25686), .Z(n33304) );
  NOR U38714 ( .A(n33298), .B(n33304), .Z(n28922) );
  IV U38715 ( .A(n25688), .Z(n25689) );
  NOR U38716 ( .A(n25690), .B(n25689), .Z(n26671) );
  IV U38717 ( .A(n25691), .Z(n25692) );
  NOR U38718 ( .A(n25693), .B(n25692), .Z(n25694) );
  IV U38719 ( .A(n25694), .Z(n26646) );
  IV U38720 ( .A(n25695), .Z(n25697) );
  NOR U38721 ( .A(n25697), .B(n25696), .Z(n29752) );
  IV U38722 ( .A(n25698), .Z(n25699) );
  NOR U38723 ( .A(n25700), .B(n25699), .Z(n29744) );
  NOR U38724 ( .A(n29752), .B(n29744), .Z(n26636) );
  IV U38725 ( .A(n25701), .Z(n25703) );
  NOR U38726 ( .A(n25703), .B(n25702), .Z(n38927) );
  IV U38727 ( .A(n25704), .Z(n25705) );
  NOR U38728 ( .A(n25706), .B(n25705), .Z(n38913) );
  NOR U38729 ( .A(n38927), .B(n38913), .Z(n33278) );
  IV U38730 ( .A(n25707), .Z(n25709) );
  NOR U38731 ( .A(n25709), .B(n25708), .Z(n33254) );
  IV U38732 ( .A(n25710), .Z(n25711) );
  NOR U38733 ( .A(n25712), .B(n25711), .Z(n33270) );
  NOR U38734 ( .A(n33254), .B(n33270), .Z(n29730) );
  IV U38735 ( .A(n25713), .Z(n25714) );
  NOR U38736 ( .A(n25715), .B(n25714), .Z(n28943) );
  IV U38737 ( .A(n25716), .Z(n25717) );
  NOR U38738 ( .A(n25718), .B(n25717), .Z(n32426) );
  IV U38739 ( .A(n25719), .Z(n25720) );
  NOR U38740 ( .A(n25721), .B(n25720), .Z(n33262) );
  NOR U38741 ( .A(n32426), .B(n33262), .Z(n29724) );
  IV U38742 ( .A(n25722), .Z(n25723) );
  NOR U38743 ( .A(n25724), .B(n25723), .Z(n29711) );
  IV U38744 ( .A(n25725), .Z(n25727) );
  NOR U38745 ( .A(n25727), .B(n25726), .Z(n28946) );
  NOR U38746 ( .A(n29711), .B(n28946), .Z(n26621) );
  IV U38747 ( .A(n25728), .Z(n25729) );
  NOR U38748 ( .A(n25730), .B(n25729), .Z(n29709) );
  IV U38749 ( .A(n25731), .Z(n25733) );
  NOR U38750 ( .A(n25733), .B(n25732), .Z(n36609) );
  IV U38751 ( .A(n25734), .Z(n25735) );
  NOR U38752 ( .A(n25736), .B(n25735), .Z(n35755) );
  NOR U38753 ( .A(n36609), .B(n35755), .Z(n28951) );
  IV U38754 ( .A(n25737), .Z(n25738) );
  NOR U38755 ( .A(n25739), .B(n25738), .Z(n39641) );
  IV U38756 ( .A(n25740), .Z(n25741) );
  NOR U38757 ( .A(n25742), .B(n25741), .Z(n25743) );
  NOR U38758 ( .A(n39641), .B(n25743), .Z(n28950) );
  IV U38759 ( .A(n25744), .Z(n25745) );
  NOR U38760 ( .A(n25746), .B(n25745), .Z(n36594) );
  IV U38761 ( .A(n25747), .Z(n25748) );
  NOR U38762 ( .A(n25749), .B(n25748), .Z(n36585) );
  NOR U38763 ( .A(n36594), .B(n36585), .Z(n33242) );
  IV U38764 ( .A(n25750), .Z(n25751) );
  NOR U38765 ( .A(n25752), .B(n25751), .Z(n32441) );
  IV U38766 ( .A(n25753), .Z(n25755) );
  NOR U38767 ( .A(n25755), .B(n25754), .Z(n32436) );
  NOR U38768 ( .A(n32441), .B(n32436), .Z(n29692) );
  IV U38769 ( .A(n25756), .Z(n25758) );
  NOR U38770 ( .A(n25758), .B(n25757), .Z(n33222) );
  IV U38771 ( .A(n25759), .Z(n25760) );
  NOR U38772 ( .A(n25761), .B(n25760), .Z(n25762) );
  NOR U38773 ( .A(n33222), .B(n25762), .Z(n29695) );
  IV U38774 ( .A(n25763), .Z(n25764) );
  NOR U38775 ( .A(n25765), .B(n25764), .Z(n33224) );
  IV U38776 ( .A(n33224), .Z(n28962) );
  IV U38777 ( .A(n25766), .Z(n25767) );
  NOR U38778 ( .A(n25768), .B(n25767), .Z(n25769) );
  IV U38779 ( .A(n25769), .Z(n29677) );
  IV U38780 ( .A(n25770), .Z(n25772) );
  NOR U38781 ( .A(n25772), .B(n25771), .Z(n29672) );
  IV U38782 ( .A(n25773), .Z(n25775) );
  NOR U38783 ( .A(n25775), .B(n25774), .Z(n29679) );
  NOR U38784 ( .A(n29672), .B(n29679), .Z(n26593) );
  IV U38785 ( .A(n25776), .Z(n25777) );
  NOR U38786 ( .A(n25778), .B(n25777), .Z(n32454) );
  IV U38787 ( .A(n25779), .Z(n25781) );
  NOR U38788 ( .A(n25781), .B(n25780), .Z(n32450) );
  NOR U38789 ( .A(n32454), .B(n32450), .Z(n29671) );
  IV U38790 ( .A(n25782), .Z(n25783) );
  NOR U38791 ( .A(n25784), .B(n25783), .Z(n26584) );
  IV U38792 ( .A(n26584), .Z(n26579) );
  IV U38793 ( .A(n25785), .Z(n25786) );
  NOR U38794 ( .A(n25787), .B(n25786), .Z(n28976) );
  IV U38795 ( .A(n25788), .Z(n25789) );
  NOR U38796 ( .A(n25790), .B(n25789), .Z(n25791) );
  IV U38797 ( .A(n25791), .Z(n28985) );
  IV U38798 ( .A(n25792), .Z(n25794) );
  NOR U38799 ( .A(n25794), .B(n25793), .Z(n28989) );
  IV U38800 ( .A(n25795), .Z(n25797) );
  NOR U38801 ( .A(n25797), .B(n25796), .Z(n28992) );
  NOR U38802 ( .A(n28989), .B(n28992), .Z(n26570) );
  IV U38803 ( .A(n25798), .Z(n25799) );
  NOR U38804 ( .A(n25800), .B(n25799), .Z(n29003) );
  IV U38805 ( .A(n25801), .Z(n25802) );
  NOR U38806 ( .A(n25803), .B(n25802), .Z(n29012) );
  IV U38807 ( .A(n25804), .Z(n25806) );
  NOR U38808 ( .A(n25806), .B(n25805), .Z(n29007) );
  NOR U38809 ( .A(n29012), .B(n29007), .Z(n25807) );
  IV U38810 ( .A(n25807), .Z(n26562) );
  IV U38811 ( .A(n25808), .Z(n25809) );
  NOR U38812 ( .A(n25810), .B(n25809), .Z(n29010) );
  IV U38813 ( .A(n25811), .Z(n25812) );
  NOR U38814 ( .A(n25813), .B(n25812), .Z(n32479) );
  IV U38815 ( .A(n25814), .Z(n25815) );
  NOR U38816 ( .A(n25816), .B(n25815), .Z(n32475) );
  NOR U38817 ( .A(n32479), .B(n32475), .Z(n29658) );
  IV U38818 ( .A(n25817), .Z(n25818) );
  NOR U38819 ( .A(n25819), .B(n25818), .Z(n35838) );
  IV U38820 ( .A(n25820), .Z(n25821) );
  NOR U38821 ( .A(n25822), .B(n25821), .Z(n35829) );
  NOR U38822 ( .A(n35838), .B(n35829), .Z(n29644) );
  IV U38823 ( .A(n25823), .Z(n25825) );
  NOR U38824 ( .A(n25825), .B(n25824), .Z(n29633) );
  IV U38825 ( .A(n25826), .Z(n25827) );
  NOR U38826 ( .A(n25828), .B(n25827), .Z(n29637) );
  NOR U38827 ( .A(n29633), .B(n29637), .Z(n26541) );
  IV U38828 ( .A(n25829), .Z(n25830) );
  NOR U38829 ( .A(n25831), .B(n25830), .Z(n33156) );
  IV U38830 ( .A(n25832), .Z(n25833) );
  NOR U38831 ( .A(n25834), .B(n25833), .Z(n33161) );
  NOR U38832 ( .A(n33156), .B(n33161), .Z(n29624) );
  IV U38833 ( .A(n25835), .Z(n25836) );
  NOR U38834 ( .A(n25837), .B(n25836), .Z(n26526) );
  IV U38835 ( .A(n26526), .Z(n26521) );
  IV U38836 ( .A(n25838), .Z(n25839) );
  NOR U38837 ( .A(n25840), .B(n25839), .Z(n29015) );
  IV U38838 ( .A(n25841), .Z(n25843) );
  NOR U38839 ( .A(n25843), .B(n25842), .Z(n25844) );
  IV U38840 ( .A(n25844), .Z(n29024) );
  IV U38841 ( .A(n25845), .Z(n25847) );
  NOR U38842 ( .A(n25847), .B(n25846), .Z(n32515) );
  IV U38843 ( .A(n25848), .Z(n25849) );
  NOR U38844 ( .A(n25850), .B(n25849), .Z(n33119) );
  NOR U38845 ( .A(n32515), .B(n33119), .Z(n29029) );
  IV U38846 ( .A(n25851), .Z(n25853) );
  NOR U38847 ( .A(n25853), .B(n25852), .Z(n29558) );
  IV U38848 ( .A(n25854), .Z(n25856) );
  NOR U38849 ( .A(n25856), .B(n25855), .Z(n29569) );
  NOR U38850 ( .A(n29558), .B(n29569), .Z(n29555) );
  IV U38851 ( .A(n25857), .Z(n25858) );
  NOR U38852 ( .A(n25859), .B(n25858), .Z(n32529) );
  IV U38853 ( .A(n25860), .Z(n25862) );
  NOR U38854 ( .A(n25862), .B(n25861), .Z(n32525) );
  NOR U38855 ( .A(n32529), .B(n32525), .Z(n29559) );
  IV U38856 ( .A(n25863), .Z(n25865) );
  NOR U38857 ( .A(n25865), .B(n25864), .Z(n32536) );
  IV U38858 ( .A(n25866), .Z(n25867) );
  NOR U38859 ( .A(n25868), .B(n25867), .Z(n25869) );
  NOR U38860 ( .A(n32536), .B(n25869), .Z(n29548) );
  IV U38861 ( .A(n25870), .Z(n25872) );
  NOR U38862 ( .A(n25872), .B(n25871), .Z(n33116) );
  IV U38863 ( .A(n25873), .Z(n25874) );
  NOR U38864 ( .A(n25875), .B(n25874), .Z(n25876) );
  NOR U38865 ( .A(n33116), .B(n25876), .Z(n29033) );
  IV U38866 ( .A(n25877), .Z(n25878) );
  NOR U38867 ( .A(n25879), .B(n25878), .Z(n29030) );
  IV U38868 ( .A(n25880), .Z(n25882) );
  NOR U38869 ( .A(n25882), .B(n25881), .Z(n29535) );
  IV U38870 ( .A(n25883), .Z(n25885) );
  NOR U38871 ( .A(n25885), .B(n25884), .Z(n29528) );
  NOR U38872 ( .A(n29535), .B(n29528), .Z(n25886) );
  IV U38873 ( .A(n25886), .Z(n26489) );
  IV U38874 ( .A(n25887), .Z(n25888) );
  NOR U38875 ( .A(n25889), .B(n25888), .Z(n29533) );
  IV U38876 ( .A(n25890), .Z(n25891) );
  NOR U38877 ( .A(n25892), .B(n25891), .Z(n25893) );
  IV U38878 ( .A(n25893), .Z(n29503) );
  IV U38879 ( .A(n25894), .Z(n25895) );
  NOR U38880 ( .A(n25896), .B(n25895), .Z(n29497) );
  IV U38881 ( .A(n29497), .Z(n32572) );
  IV U38882 ( .A(n25897), .Z(n25898) );
  NOR U38883 ( .A(n25899), .B(n25898), .Z(n32590) );
  IV U38884 ( .A(n25900), .Z(n25901) );
  NOR U38885 ( .A(n25902), .B(n25901), .Z(n32585) );
  NOR U38886 ( .A(n32590), .B(n32585), .Z(n29060) );
  IV U38887 ( .A(n25903), .Z(n25905) );
  NOR U38888 ( .A(n25905), .B(n25904), .Z(n33074) );
  IV U38889 ( .A(n25906), .Z(n25908) );
  NOR U38890 ( .A(n25908), .B(n25907), .Z(n32601) );
  NOR U38891 ( .A(n33074), .B(n32601), .Z(n29066) );
  IV U38892 ( .A(n25909), .Z(n25911) );
  NOR U38893 ( .A(n25911), .B(n25910), .Z(n29063) );
  IV U38894 ( .A(n25912), .Z(n25913) );
  NOR U38895 ( .A(n25914), .B(n25913), .Z(n29483) );
  IV U38896 ( .A(n25915), .Z(n25917) );
  NOR U38897 ( .A(n25917), .B(n25916), .Z(n29488) );
  NOR U38898 ( .A(n29483), .B(n29488), .Z(n32610) );
  IV U38899 ( .A(n25918), .Z(n25919) );
  NOR U38900 ( .A(n25920), .B(n25919), .Z(n26424) );
  IV U38901 ( .A(n26424), .Z(n26414) );
  IV U38902 ( .A(n25921), .Z(n25922) );
  NOR U38903 ( .A(n25923), .B(n25922), .Z(n26406) );
  IV U38904 ( .A(n25924), .Z(n25925) );
  NOR U38905 ( .A(n25926), .B(n25925), .Z(n26397) );
  IV U38906 ( .A(n25927), .Z(n25929) );
  NOR U38907 ( .A(n25929), .B(n25928), .Z(n29073) );
  IV U38908 ( .A(n25930), .Z(n25932) );
  NOR U38909 ( .A(n25932), .B(n25931), .Z(n29071) );
  NOR U38910 ( .A(n29073), .B(n29071), .Z(n26396) );
  IV U38911 ( .A(n25933), .Z(n25934) );
  NOR U38912 ( .A(n25935), .B(n25934), .Z(n36412) );
  IV U38913 ( .A(n25936), .Z(n25938) );
  NOR U38914 ( .A(n25938), .B(n25937), .Z(n25939) );
  NOR U38915 ( .A(n36412), .B(n25939), .Z(n35958) );
  IV U38916 ( .A(n25940), .Z(n25942) );
  NOR U38917 ( .A(n25942), .B(n25941), .Z(n29473) );
  IV U38918 ( .A(n25943), .Z(n25944) );
  NOR U38919 ( .A(n25945), .B(n25944), .Z(n29478) );
  NOR U38920 ( .A(n29473), .B(n29478), .Z(n26395) );
  IV U38921 ( .A(n25946), .Z(n25947) );
  NOR U38922 ( .A(n25948), .B(n25947), .Z(n29471) );
  IV U38923 ( .A(n25949), .Z(n25951) );
  NOR U38924 ( .A(n25951), .B(n25950), .Z(n29454) );
  IV U38925 ( .A(n25952), .Z(n25954) );
  NOR U38926 ( .A(n25954), .B(n25953), .Z(n29448) );
  NOR U38927 ( .A(n29454), .B(n29448), .Z(n26387) );
  IV U38928 ( .A(n25955), .Z(n25957) );
  NOR U38929 ( .A(n25957), .B(n25956), .Z(n29452) );
  IV U38930 ( .A(n25958), .Z(n25959) );
  NOR U38931 ( .A(n25960), .B(n25959), .Z(n36366) );
  IV U38932 ( .A(n25961), .Z(n25962) );
  NOR U38933 ( .A(n25963), .B(n25962), .Z(n36375) );
  NOR U38934 ( .A(n36366), .B(n36375), .Z(n33022) );
  IV U38935 ( .A(n25964), .Z(n25966) );
  NOR U38936 ( .A(n25966), .B(n25965), .Z(n33012) );
  IV U38937 ( .A(n25967), .Z(n25969) );
  NOR U38938 ( .A(n25969), .B(n25968), .Z(n32642) );
  NOR U38939 ( .A(n33012), .B(n32642), .Z(n29092) );
  IV U38940 ( .A(n25970), .Z(n25971) );
  NOR U38941 ( .A(n25972), .B(n25971), .Z(n33006) );
  IV U38942 ( .A(n25973), .Z(n25974) );
  NOR U38943 ( .A(n25975), .B(n25974), .Z(n33015) );
  NOR U38944 ( .A(n33006), .B(n33015), .Z(n29436) );
  IV U38945 ( .A(n25976), .Z(n25978) );
  NOR U38946 ( .A(n25978), .B(n25977), .Z(n32646) );
  IV U38947 ( .A(n25979), .Z(n25980) );
  NOR U38948 ( .A(n25981), .B(n25980), .Z(n33003) );
  NOR U38949 ( .A(n32646), .B(n33003), .Z(n29434) );
  IV U38950 ( .A(n25982), .Z(n25983) );
  NOR U38951 ( .A(n25984), .B(n25983), .Z(n29431) );
  IV U38952 ( .A(n25985), .Z(n25986) );
  NOR U38953 ( .A(n25987), .B(n25986), .Z(n29093) );
  NOR U38954 ( .A(n29431), .B(n29093), .Z(n26365) );
  IV U38955 ( .A(n25988), .Z(n25989) );
  NOR U38956 ( .A(n25990), .B(n25989), .Z(n29096) );
  NOR U38957 ( .A(n25992), .B(n25991), .Z(n25996) );
  IV U38958 ( .A(n25992), .Z(n25994) );
  NOR U38959 ( .A(n25994), .B(n25993), .Z(n36016) );
  NOR U38960 ( .A(n36005), .B(n36016), .Z(n25995) );
  NOR U38961 ( .A(n25996), .B(n25995), .Z(n29099) );
  IV U38962 ( .A(n25997), .Z(n25998) );
  NOR U38963 ( .A(n25999), .B(n25998), .Z(n32667) );
  NOR U38964 ( .A(n26001), .B(n26000), .Z(n32663) );
  NOR U38965 ( .A(n32667), .B(n32663), .Z(n29098) );
  IV U38966 ( .A(n26002), .Z(n26003) );
  NOR U38967 ( .A(n26004), .B(n26003), .Z(n29112) );
  IV U38968 ( .A(n26005), .Z(n26007) );
  NOR U38969 ( .A(n26007), .B(n26006), .Z(n36331) );
  IV U38970 ( .A(n26008), .Z(n26009) );
  NOR U38971 ( .A(n26010), .B(n26009), .Z(n36034) );
  NOR U38972 ( .A(n36331), .B(n36034), .Z(n29115) );
  IV U38973 ( .A(n26011), .Z(n26013) );
  NOR U38974 ( .A(n26013), .B(n26012), .Z(n26328) );
  IV U38975 ( .A(n26014), .Z(n26015) );
  NOR U38976 ( .A(n26016), .B(n26015), .Z(n29120) );
  IV U38977 ( .A(n26017), .Z(n26018) );
  NOR U38978 ( .A(n26019), .B(n26018), .Z(n29397) );
  NOR U38979 ( .A(n29120), .B(n29397), .Z(n26319) );
  IV U38980 ( .A(n26020), .Z(n26021) );
  NOR U38981 ( .A(n26022), .B(n26021), .Z(n32978) );
  IV U38982 ( .A(n26023), .Z(n26025) );
  NOR U38983 ( .A(n26025), .B(n26024), .Z(n32693) );
  NOR U38984 ( .A(n32978), .B(n32693), .Z(n29122) );
  IV U38985 ( .A(n26026), .Z(n26028) );
  NOR U38986 ( .A(n26028), .B(n26027), .Z(n29384) );
  IV U38987 ( .A(n26029), .Z(n26031) );
  NOR U38988 ( .A(n26031), .B(n26030), .Z(n29130) );
  NOR U38989 ( .A(n29384), .B(n29130), .Z(n26305) );
  IV U38990 ( .A(n26032), .Z(n26033) );
  NOR U38991 ( .A(n26034), .B(n26033), .Z(n29382) );
  IV U38992 ( .A(n26035), .Z(n26037) );
  NOR U38993 ( .A(n26037), .B(n26036), .Z(n29364) );
  IV U38994 ( .A(n26038), .Z(n26040) );
  NOR U38995 ( .A(n26040), .B(n26039), .Z(n29379) );
  NOR U38996 ( .A(n29364), .B(n29379), .Z(n26304) );
  IV U38997 ( .A(n26041), .Z(n26042) );
  NOR U38998 ( .A(n26043), .B(n26042), .Z(n29135) );
  IV U38999 ( .A(n26044), .Z(n26045) );
  NOR U39000 ( .A(n26046), .B(n26045), .Z(n29368) );
  NOR U39001 ( .A(n29135), .B(n29368), .Z(n26303) );
  IV U39002 ( .A(n26047), .Z(n26049) );
  NOR U39003 ( .A(n26049), .B(n26048), .Z(n29133) );
  IV U39004 ( .A(n26050), .Z(n26052) );
  NOR U39005 ( .A(n26052), .B(n26051), .Z(n36288) );
  IV U39006 ( .A(n26053), .Z(n26054) );
  NOR U39007 ( .A(n26055), .B(n26054), .Z(n26056) );
  NOR U39008 ( .A(n36288), .B(n26056), .Z(n29141) );
  IV U39009 ( .A(n26057), .Z(n26058) );
  NOR U39010 ( .A(n26059), .B(n26058), .Z(n26060) );
  IV U39011 ( .A(n26060), .Z(n26286) );
  IV U39012 ( .A(n26061), .Z(n26062) );
  NOR U39013 ( .A(n26063), .B(n26062), .Z(n32737) );
  IV U39014 ( .A(n26064), .Z(n26065) );
  NOR U39015 ( .A(n26066), .B(n26065), .Z(n32732) );
  NOR U39016 ( .A(n32737), .B(n32732), .Z(n29326) );
  IV U39017 ( .A(n26067), .Z(n26068) );
  NOR U39018 ( .A(n26069), .B(n26068), .Z(n32744) );
  IV U39019 ( .A(n26070), .Z(n26071) );
  NOR U39020 ( .A(n26072), .B(n26071), .Z(n32740) );
  NOR U39021 ( .A(n32744), .B(n32740), .Z(n29167) );
  IV U39022 ( .A(n26073), .Z(n26075) );
  NOR U39023 ( .A(n26075), .B(n26074), .Z(n29172) );
  IV U39024 ( .A(n26076), .Z(n26077) );
  NOR U39025 ( .A(n26078), .B(n26077), .Z(n29168) );
  NOR U39026 ( .A(n29172), .B(n29168), .Z(n26257) );
  IV U39027 ( .A(n26079), .Z(n26081) );
  NOR U39028 ( .A(n26081), .B(n26080), .Z(n32948) );
  IV U39029 ( .A(n26082), .Z(n26083) );
  NOR U39030 ( .A(n26084), .B(n26083), .Z(n32760) );
  NOR U39031 ( .A(n32948), .B(n32760), .Z(n29176) );
  IV U39032 ( .A(n26085), .Z(n26087) );
  NOR U39033 ( .A(n26087), .B(n26086), .Z(n32936) );
  IV U39034 ( .A(n26088), .Z(n26089) );
  NOR U39035 ( .A(n26090), .B(n26089), .Z(n32766) );
  NOR U39036 ( .A(n32936), .B(n32766), .Z(n29181) );
  IV U39037 ( .A(n26091), .Z(n26092) );
  NOR U39038 ( .A(n26093), .B(n26092), .Z(n29199) );
  IV U39039 ( .A(n26094), .Z(n26095) );
  NOR U39040 ( .A(n26096), .B(n26095), .Z(n29193) );
  IV U39041 ( .A(n26097), .Z(n26098) );
  NOR U39042 ( .A(n26099), .B(n26098), .Z(n29195) );
  NOR U39043 ( .A(n29193), .B(n29195), .Z(n26229) );
  IV U39044 ( .A(n26100), .Z(n26102) );
  NOR U39045 ( .A(n26102), .B(n26101), .Z(n29215) );
  IV U39046 ( .A(n26103), .Z(n26104) );
  NOR U39047 ( .A(n26105), .B(n26104), .Z(n32860) );
  IV U39048 ( .A(n26106), .Z(n26108) );
  NOR U39049 ( .A(n26108), .B(n26107), .Z(n29294) );
  IV U39050 ( .A(n26109), .Z(n26110) );
  NOR U39051 ( .A(n26111), .B(n26110), .Z(n29247) );
  NOR U39052 ( .A(n29294), .B(n29247), .Z(n26158) );
  IV U39053 ( .A(n26112), .Z(n26114) );
  NOR U39054 ( .A(n26114), .B(n26113), .Z(n29291) );
  IV U39055 ( .A(n26115), .Z(n26117) );
  NOR U39056 ( .A(n26117), .B(n26116), .Z(n29250) );
  IV U39057 ( .A(n26118), .Z(n26120) );
  NOR U39058 ( .A(n26120), .B(n26119), .Z(n29288) );
  NOR U39059 ( .A(n29250), .B(n29288), .Z(n26156) );
  IV U39060 ( .A(n26121), .Z(n26122) );
  NOR U39061 ( .A(n26123), .B(n26122), .Z(n29283) );
  IV U39062 ( .A(n26124), .Z(n26126) );
  NOR U39063 ( .A(n26126), .B(n26125), .Z(n29253) );
  NOR U39064 ( .A(n29283), .B(n29253), .Z(n26155) );
  IV U39065 ( .A(n26127), .Z(n26128) );
  NOR U39066 ( .A(n26129), .B(n26128), .Z(n29263) );
  IV U39067 ( .A(n26130), .Z(n26131) );
  NOR U39068 ( .A(n26132), .B(n26131), .Z(n29273) );
  IV U39069 ( .A(n26133), .Z(n26135) );
  NOR U39070 ( .A(n26135), .B(n26134), .Z(n26136) );
  IV U39071 ( .A(n26136), .Z(n29257) );
  IV U39072 ( .A(n26137), .Z(n26139) );
  NOR U39073 ( .A(n26139), .B(n26138), .Z(n29271) );
  XOR U39074 ( .A(n29257), .B(n29271), .Z(n26140) );
  NOR U39075 ( .A(n29273), .B(n26140), .Z(n26147) );
  IV U39076 ( .A(n29273), .Z(n26144) );
  IV U39077 ( .A(n26141), .Z(n26143) );
  NOR U39078 ( .A(n26143), .B(n26142), .Z(n29270) );
  XOR U39079 ( .A(n26144), .B(n29270), .Z(n26145) );
  NOR U39080 ( .A(n29271), .B(n26145), .Z(n26146) );
  NOR U39081 ( .A(n26147), .B(n26146), .Z(n29264) );
  XOR U39082 ( .A(n29263), .B(n29264), .Z(n29284) );
  IV U39083 ( .A(n26148), .Z(n26150) );
  NOR U39084 ( .A(n26150), .B(n26149), .Z(n29285) );
  IV U39085 ( .A(n26151), .Z(n26153) );
  NOR U39086 ( .A(n26153), .B(n26152), .Z(n29259) );
  NOR U39087 ( .A(n29285), .B(n29259), .Z(n26154) );
  XOR U39088 ( .A(n29284), .B(n26154), .Z(n29254) );
  XOR U39089 ( .A(n26155), .B(n29254), .Z(n29290) );
  XOR U39090 ( .A(n26156), .B(n29290), .Z(n26157) );
  IV U39091 ( .A(n26157), .Z(n29295) );
  XOR U39092 ( .A(n29291), .B(n29295), .Z(n29248) );
  XOR U39093 ( .A(n26158), .B(n29248), .Z(n26159) );
  IV U39094 ( .A(n26159), .Z(n29246) );
  IV U39095 ( .A(n26160), .Z(n26161) );
  NOR U39096 ( .A(n26162), .B(n26161), .Z(n29244) );
  IV U39097 ( .A(n26163), .Z(n26164) );
  NOR U39098 ( .A(n26165), .B(n26164), .Z(n29242) );
  NOR U39099 ( .A(n29244), .B(n29242), .Z(n26166) );
  XOR U39100 ( .A(n29246), .B(n26166), .Z(n29237) );
  IV U39101 ( .A(n26167), .Z(n26168) );
  NOR U39102 ( .A(n26169), .B(n26168), .Z(n29239) );
  IV U39103 ( .A(n26170), .Z(n26171) );
  NOR U39104 ( .A(n26172), .B(n26171), .Z(n29236) );
  NOR U39105 ( .A(n29239), .B(n29236), .Z(n26173) );
  XOR U39106 ( .A(n29237), .B(n26173), .Z(n32848) );
  XOR U39107 ( .A(n32860), .B(n32848), .Z(n29234) );
  IV U39108 ( .A(n26174), .Z(n26176) );
  NOR U39109 ( .A(n26176), .B(n26175), .Z(n29297) );
  IV U39110 ( .A(n26177), .Z(n26178) );
  NOR U39111 ( .A(n26179), .B(n26178), .Z(n29233) );
  NOR U39112 ( .A(n29297), .B(n29233), .Z(n26180) );
  XOR U39113 ( .A(n29234), .B(n26180), .Z(n29225) );
  IV U39114 ( .A(n26181), .Z(n26182) );
  NOR U39115 ( .A(n26183), .B(n26182), .Z(n29226) );
  IV U39116 ( .A(n26184), .Z(n26185) );
  NOR U39117 ( .A(n26186), .B(n26185), .Z(n29228) );
  NOR U39118 ( .A(n29226), .B(n29228), .Z(n26187) );
  XOR U39119 ( .A(n29225), .B(n26187), .Z(n29223) );
  IV U39120 ( .A(n26188), .Z(n26190) );
  NOR U39121 ( .A(n26190), .B(n26189), .Z(n29222) );
  IV U39122 ( .A(n26191), .Z(n26193) );
  NOR U39123 ( .A(n26193), .B(n26192), .Z(n29220) );
  NOR U39124 ( .A(n29222), .B(n29220), .Z(n26194) );
  XOR U39125 ( .A(n29223), .B(n26194), .Z(n29217) );
  IV U39126 ( .A(n26195), .Z(n26196) );
  NOR U39127 ( .A(n26197), .B(n26196), .Z(n29218) );
  IV U39128 ( .A(n26198), .Z(n26199) );
  NOR U39129 ( .A(n26200), .B(n26199), .Z(n29300) );
  NOR U39130 ( .A(n29218), .B(n29300), .Z(n26201) );
  XOR U39131 ( .A(n29217), .B(n26201), .Z(n29304) );
  XOR U39132 ( .A(n29215), .B(n29304), .Z(n29310) );
  IV U39133 ( .A(n26202), .Z(n26204) );
  NOR U39134 ( .A(n26204), .B(n26203), .Z(n29303) );
  IV U39135 ( .A(n26205), .Z(n26206) );
  NOR U39136 ( .A(n26207), .B(n26206), .Z(n29309) );
  NOR U39137 ( .A(n29303), .B(n29309), .Z(n26208) );
  XOR U39138 ( .A(n29310), .B(n26208), .Z(n29307) );
  IV U39139 ( .A(n26209), .Z(n26210) );
  NOR U39140 ( .A(n26211), .B(n26210), .Z(n32785) );
  IV U39141 ( .A(n26212), .Z(n26214) );
  NOR U39142 ( .A(n26214), .B(n26213), .Z(n32780) );
  NOR U39143 ( .A(n32785), .B(n32780), .Z(n29308) );
  XOR U39144 ( .A(n29307), .B(n29308), .Z(n29213) );
  IV U39145 ( .A(n26215), .Z(n26217) );
  NOR U39146 ( .A(n26217), .B(n26216), .Z(n29212) );
  IV U39147 ( .A(n26218), .Z(n26219) );
  NOR U39148 ( .A(n26220), .B(n26219), .Z(n29210) );
  NOR U39149 ( .A(n29212), .B(n29210), .Z(n26221) );
  XOR U39150 ( .A(n29213), .B(n26221), .Z(n29205) );
  IV U39151 ( .A(n26222), .Z(n26223) );
  NOR U39152 ( .A(n26224), .B(n26223), .Z(n29207) );
  IV U39153 ( .A(n26225), .Z(n26226) );
  NOR U39154 ( .A(n26227), .B(n26226), .Z(n29204) );
  NOR U39155 ( .A(n29207), .B(n29204), .Z(n26228) );
  XOR U39156 ( .A(n29205), .B(n26228), .Z(n29197) );
  XOR U39157 ( .A(n26229), .B(n29197), .Z(n26230) );
  IV U39158 ( .A(n26230), .Z(n29200) );
  XOR U39159 ( .A(n29199), .B(n29200), .Z(n29189) );
  IV U39160 ( .A(n26231), .Z(n26233) );
  NOR U39161 ( .A(n26233), .B(n26232), .Z(n29191) );
  IV U39162 ( .A(n26234), .Z(n26236) );
  NOR U39163 ( .A(n26236), .B(n26235), .Z(n29188) );
  NOR U39164 ( .A(n29191), .B(n29188), .Z(n26237) );
  XOR U39165 ( .A(n29189), .B(n26237), .Z(n29186) );
  IV U39166 ( .A(n26238), .Z(n26239) );
  NOR U39167 ( .A(n26240), .B(n26239), .Z(n32928) );
  IV U39168 ( .A(n26241), .Z(n26243) );
  NOR U39169 ( .A(n26243), .B(n26242), .Z(n32920) );
  NOR U39170 ( .A(n32928), .B(n32920), .Z(n29187) );
  XOR U39171 ( .A(n29186), .B(n29187), .Z(n32767) );
  XOR U39172 ( .A(n29181), .B(n32767), .Z(n29178) );
  IV U39173 ( .A(n26244), .Z(n26245) );
  NOR U39174 ( .A(n26246), .B(n26245), .Z(n29182) );
  IV U39175 ( .A(n26247), .Z(n26248) );
  NOR U39176 ( .A(n26249), .B(n26248), .Z(n29177) );
  NOR U39177 ( .A(n29182), .B(n29177), .Z(n26250) );
  XOR U39178 ( .A(n29178), .B(n26250), .Z(n32763) );
  XOR U39179 ( .A(n29176), .B(n32763), .Z(n29170) );
  IV U39180 ( .A(n26251), .Z(n26253) );
  NOR U39181 ( .A(n26253), .B(n26252), .Z(n32757) );
  IV U39182 ( .A(n26254), .Z(n26255) );
  NOR U39183 ( .A(n26256), .B(n26255), .Z(n32752) );
  NOR U39184 ( .A(n32757), .B(n32752), .Z(n29171) );
  XOR U39185 ( .A(n29170), .B(n29171), .Z(n29173) );
  XOR U39186 ( .A(n26257), .B(n29173), .Z(n29166) );
  XOR U39187 ( .A(n29167), .B(n29166), .Z(n32734) );
  XOR U39188 ( .A(n29326), .B(n32734), .Z(n29161) );
  IV U39189 ( .A(n26258), .Z(n26259) );
  NOR U39190 ( .A(n26260), .B(n26259), .Z(n29322) );
  IV U39191 ( .A(n26261), .Z(n26262) );
  NOR U39192 ( .A(n26263), .B(n26262), .Z(n29164) );
  NOR U39193 ( .A(n29322), .B(n29164), .Z(n26264) );
  XOR U39194 ( .A(n29161), .B(n26264), .Z(n29158) );
  IV U39195 ( .A(n26265), .Z(n26266) );
  NOR U39196 ( .A(n26267), .B(n26266), .Z(n29160) );
  IV U39197 ( .A(n26268), .Z(n26269) );
  NOR U39198 ( .A(n26270), .B(n26269), .Z(n29157) );
  NOR U39199 ( .A(n29160), .B(n29157), .Z(n26271) );
  XOR U39200 ( .A(n29158), .B(n26271), .Z(n29150) );
  IV U39201 ( .A(n26272), .Z(n26273) );
  NOR U39202 ( .A(n26274), .B(n26273), .Z(n29151) );
  IV U39203 ( .A(n26275), .Z(n26276) );
  NOR U39204 ( .A(n26277), .B(n26276), .Z(n29153) );
  NOR U39205 ( .A(n29151), .B(n29153), .Z(n26278) );
  XOR U39206 ( .A(n29150), .B(n26278), .Z(n29148) );
  NOR U39207 ( .A(n26286), .B(n29148), .Z(n29336) );
  IV U39208 ( .A(n26279), .Z(n26280) );
  NOR U39209 ( .A(n26281), .B(n26280), .Z(n29144) );
  IV U39210 ( .A(n26282), .Z(n26284) );
  NOR U39211 ( .A(n26284), .B(n26283), .Z(n26285) );
  IV U39212 ( .A(n26285), .Z(n29149) );
  XOR U39213 ( .A(n29149), .B(n29148), .Z(n29145) );
  XOR U39214 ( .A(n29144), .B(n29145), .Z(n26288) );
  NOR U39215 ( .A(n29145), .B(n26286), .Z(n26287) );
  NOR U39216 ( .A(n26288), .B(n26287), .Z(n26289) );
  NOR U39217 ( .A(n29336), .B(n26289), .Z(n29142) );
  IV U39218 ( .A(n26290), .Z(n26291) );
  NOR U39219 ( .A(n26292), .B(n26291), .Z(n36075) );
  IV U39220 ( .A(n26293), .Z(n26295) );
  NOR U39221 ( .A(n26295), .B(n26294), .Z(n29347) );
  NOR U39222 ( .A(n36075), .B(n29347), .Z(n26296) );
  XOR U39223 ( .A(n29142), .B(n26296), .Z(n29140) );
  XOR U39224 ( .A(n29141), .B(n29140), .Z(n29138) );
  IV U39225 ( .A(n26297), .Z(n26299) );
  NOR U39226 ( .A(n26299), .B(n26298), .Z(n32718) );
  IV U39227 ( .A(n26300), .Z(n26302) );
  NOR U39228 ( .A(n26302), .B(n26301), .Z(n32713) );
  NOR U39229 ( .A(n32718), .B(n32713), .Z(n29139) );
  XOR U39230 ( .A(n29138), .B(n29139), .Z(n29136) );
  XOR U39231 ( .A(n29133), .B(n29136), .Z(n29369) );
  XOR U39232 ( .A(n26303), .B(n29369), .Z(n29363) );
  XOR U39233 ( .A(n26304), .B(n29363), .Z(n29385) );
  XOR U39234 ( .A(n29382), .B(n29385), .Z(n29131) );
  XOR U39235 ( .A(n26305), .B(n29131), .Z(n29127) );
  IV U39236 ( .A(n26306), .Z(n26308) );
  NOR U39237 ( .A(n26308), .B(n26307), .Z(n29128) );
  IV U39238 ( .A(n26309), .Z(n26310) );
  NOR U39239 ( .A(n26311), .B(n26310), .Z(n29390) );
  NOR U39240 ( .A(n29128), .B(n29390), .Z(n26312) );
  XOR U39241 ( .A(n29127), .B(n26312), .Z(n32694) );
  XOR U39242 ( .A(n29122), .B(n32694), .Z(n29123) );
  IV U39243 ( .A(n26313), .Z(n26314) );
  NOR U39244 ( .A(n26315), .B(n26314), .Z(n32687) );
  IV U39245 ( .A(n26316), .Z(n26317) );
  NOR U39246 ( .A(n26318), .B(n26317), .Z(n32986) );
  NOR U39247 ( .A(n32687), .B(n32986), .Z(n29124) );
  XOR U39248 ( .A(n29123), .B(n29124), .Z(n29398) );
  XOR U39249 ( .A(n26319), .B(n29398), .Z(n26329) );
  NOR U39250 ( .A(n26328), .B(n26329), .Z(n26320) );
  IV U39251 ( .A(n26320), .Z(n26324) );
  IV U39252 ( .A(n26321), .Z(n26322) );
  NOR U39253 ( .A(n26323), .B(n26322), .Z(n26325) );
  NOR U39254 ( .A(n26324), .B(n26325), .Z(n26334) );
  IV U39255 ( .A(n26325), .Z(n26327) );
  XOR U39256 ( .A(n29120), .B(n29398), .Z(n26326) );
  NOR U39257 ( .A(n26327), .B(n26326), .Z(n32683) );
  IV U39258 ( .A(n26328), .Z(n26331) );
  IV U39259 ( .A(n26329), .Z(n26330) );
  NOR U39260 ( .A(n26331), .B(n26330), .Z(n29119) );
  NOR U39261 ( .A(n32683), .B(n29119), .Z(n26332) );
  IV U39262 ( .A(n26332), .Z(n26333) );
  NOR U39263 ( .A(n26334), .B(n26333), .Z(n26335) );
  IV U39264 ( .A(n26335), .Z(n36037) );
  XOR U39265 ( .A(n29115), .B(n36037), .Z(n29116) );
  IV U39266 ( .A(n26336), .Z(n26337) );
  NOR U39267 ( .A(n26338), .B(n26337), .Z(n29411) );
  IV U39268 ( .A(n26339), .Z(n26340) );
  NOR U39269 ( .A(n26341), .B(n26340), .Z(n29415) );
  NOR U39270 ( .A(n29411), .B(n29415), .Z(n26342) );
  XOR U39271 ( .A(n29116), .B(n26342), .Z(n29406) );
  IV U39272 ( .A(n26343), .Z(n26344) );
  NOR U39273 ( .A(n26345), .B(n26344), .Z(n29410) );
  IV U39274 ( .A(n26346), .Z(n26348) );
  NOR U39275 ( .A(n26348), .B(n26347), .Z(n29405) );
  NOR U39276 ( .A(n29410), .B(n29405), .Z(n26349) );
  XOR U39277 ( .A(n29406), .B(n26349), .Z(n29111) );
  NOR U39278 ( .A(n29112), .B(n29111), .Z(n26354) );
  IV U39279 ( .A(n26350), .Z(n26351) );
  NOR U39280 ( .A(n26352), .B(n26351), .Z(n26355) );
  IV U39281 ( .A(n26355), .Z(n26353) );
  NOR U39282 ( .A(n26354), .B(n26353), .Z(n32670) );
  XOR U39283 ( .A(n29112), .B(n29111), .Z(n29108) );
  NOR U39284 ( .A(n26355), .B(n29108), .Z(n26356) );
  NOR U39285 ( .A(n32670), .B(n26356), .Z(n29104) );
  IV U39286 ( .A(n26357), .Z(n26359) );
  NOR U39287 ( .A(n26359), .B(n26358), .Z(n29107) );
  IV U39288 ( .A(n26360), .Z(n26362) );
  NOR U39289 ( .A(n26362), .B(n26361), .Z(n29103) );
  NOR U39290 ( .A(n29107), .B(n29103), .Z(n26363) );
  XOR U39291 ( .A(n29104), .B(n26363), .Z(n32664) );
  XOR U39292 ( .A(n29098), .B(n32664), .Z(n26364) );
  IV U39293 ( .A(n26364), .Z(n36013) );
  XOR U39294 ( .A(n29099), .B(n36013), .Z(n29432) );
  XOR U39295 ( .A(n29096), .B(n29432), .Z(n29094) );
  XOR U39296 ( .A(n26365), .B(n29094), .Z(n32647) );
  XOR U39297 ( .A(n29434), .B(n32647), .Z(n33008) );
  XOR U39298 ( .A(n29436), .B(n33008), .Z(n29091) );
  XOR U39299 ( .A(n29092), .B(n29091), .Z(n33019) );
  XOR U39300 ( .A(n33022), .B(n33019), .Z(n29088) );
  IV U39301 ( .A(n26366), .Z(n26367) );
  NOR U39302 ( .A(n26368), .B(n26367), .Z(n29087) );
  IV U39303 ( .A(n26369), .Z(n26370) );
  NOR U39304 ( .A(n26371), .B(n26370), .Z(n29442) );
  NOR U39305 ( .A(n29087), .B(n29442), .Z(n26372) );
  XOR U39306 ( .A(n29088), .B(n26372), .Z(n29086) );
  IV U39307 ( .A(n26373), .Z(n26374) );
  NOR U39308 ( .A(n26375), .B(n26374), .Z(n29084) );
  IV U39309 ( .A(n26376), .Z(n26377) );
  NOR U39310 ( .A(n26378), .B(n26377), .Z(n29082) );
  NOR U39311 ( .A(n29084), .B(n29082), .Z(n26379) );
  XOR U39312 ( .A(n29086), .B(n26379), .Z(n29077) );
  IV U39313 ( .A(n26380), .Z(n26382) );
  NOR U39314 ( .A(n26382), .B(n26381), .Z(n29079) );
  IV U39315 ( .A(n26383), .Z(n26385) );
  NOR U39316 ( .A(n26385), .B(n26384), .Z(n29076) );
  NOR U39317 ( .A(n29079), .B(n29076), .Z(n26386) );
  XOR U39318 ( .A(n29077), .B(n26386), .Z(n29455) );
  XOR U39319 ( .A(n29452), .B(n29455), .Z(n29449) );
  XOR U39320 ( .A(n26387), .B(n29449), .Z(n29459) );
  IV U39321 ( .A(n26388), .Z(n26389) );
  NOR U39322 ( .A(n26390), .B(n26389), .Z(n29460) );
  IV U39323 ( .A(n26391), .Z(n26392) );
  NOR U39324 ( .A(n26393), .B(n26392), .Z(n29468) );
  NOR U39325 ( .A(n29460), .B(n29468), .Z(n26394) );
  XOR U39326 ( .A(n29459), .B(n26394), .Z(n29474) );
  XOR U39327 ( .A(n29471), .B(n29474), .Z(n29479) );
  XOR U39328 ( .A(n26395), .B(n29479), .Z(n29477) );
  XOR U39329 ( .A(n35958), .B(n29477), .Z(n29074) );
  XOR U39330 ( .A(n26396), .B(n29074), .Z(n26407) );
  NOR U39331 ( .A(n26397), .B(n26407), .Z(n26400) );
  IV U39332 ( .A(n26397), .Z(n26399) );
  XOR U39333 ( .A(n29073), .B(n29074), .Z(n26398) );
  NOR U39334 ( .A(n26399), .B(n26398), .Z(n33043) );
  NOR U39335 ( .A(n26400), .B(n33043), .Z(n26401) );
  NOR U39336 ( .A(n26406), .B(n26401), .Z(n26410) );
  IV U39337 ( .A(n26402), .Z(n26404) );
  NOR U39338 ( .A(n26404), .B(n26403), .Z(n26411) );
  IV U39339 ( .A(n26411), .Z(n26405) );
  NOR U39340 ( .A(n26410), .B(n26405), .Z(n33050) );
  IV U39341 ( .A(n26406), .Z(n26409) );
  IV U39342 ( .A(n26407), .Z(n26408) );
  NOR U39343 ( .A(n26409), .B(n26408), .Z(n33047) );
  NOR U39344 ( .A(n26410), .B(n33047), .Z(n26418) );
  NOR U39345 ( .A(n26411), .B(n26418), .Z(n26412) );
  NOR U39346 ( .A(n33050), .B(n26412), .Z(n26421) );
  IV U39347 ( .A(n26421), .Z(n26413) );
  NOR U39348 ( .A(n26414), .B(n26413), .Z(n33057) );
  IV U39349 ( .A(n26415), .Z(n26417) );
  NOR U39350 ( .A(n26417), .B(n26416), .Z(n26422) );
  IV U39351 ( .A(n26422), .Z(n26420) );
  IV U39352 ( .A(n26418), .Z(n26419) );
  NOR U39353 ( .A(n26420), .B(n26419), .Z(n33054) );
  NOR U39354 ( .A(n26422), .B(n26421), .Z(n26423) );
  NOR U39355 ( .A(n33054), .B(n26423), .Z(n29482) );
  NOR U39356 ( .A(n26424), .B(n29482), .Z(n26425) );
  NOR U39357 ( .A(n33057), .B(n26425), .Z(n26426) );
  IV U39358 ( .A(n26426), .Z(n32608) );
  XOR U39359 ( .A(n32610), .B(n32608), .Z(n29068) );
  IV U39360 ( .A(n26427), .Z(n26428) );
  NOR U39361 ( .A(n26429), .B(n26428), .Z(n29491) );
  IV U39362 ( .A(n26430), .Z(n26431) );
  NOR U39363 ( .A(n26432), .B(n26431), .Z(n29069) );
  NOR U39364 ( .A(n29491), .B(n29069), .Z(n26433) );
  XOR U39365 ( .A(n29068), .B(n26433), .Z(n29064) );
  XOR U39366 ( .A(n29063), .B(n29064), .Z(n32602) );
  XOR U39367 ( .A(n29066), .B(n32602), .Z(n29058) );
  IV U39368 ( .A(n26434), .Z(n26435) );
  NOR U39369 ( .A(n26436), .B(n26435), .Z(n32598) );
  IV U39370 ( .A(n26437), .Z(n26438) );
  NOR U39371 ( .A(n26439), .B(n26438), .Z(n32593) );
  NOR U39372 ( .A(n32598), .B(n32593), .Z(n29059) );
  XOR U39373 ( .A(n29058), .B(n29059), .Z(n32587) );
  XOR U39374 ( .A(n29060), .B(n32587), .Z(n29052) );
  IV U39375 ( .A(n26440), .Z(n26441) );
  NOR U39376 ( .A(n26442), .B(n26441), .Z(n29055) );
  IV U39377 ( .A(n26443), .Z(n26444) );
  NOR U39378 ( .A(n26445), .B(n26444), .Z(n29051) );
  NOR U39379 ( .A(n29055), .B(n29051), .Z(n26446) );
  XOR U39380 ( .A(n29052), .B(n26446), .Z(n29050) );
  IV U39381 ( .A(n26447), .Z(n26449) );
  NOR U39382 ( .A(n26449), .B(n26448), .Z(n29048) );
  IV U39383 ( .A(n26450), .Z(n26451) );
  NOR U39384 ( .A(n26452), .B(n26451), .Z(n29046) );
  NOR U39385 ( .A(n29048), .B(n29046), .Z(n26453) );
  XOR U39386 ( .A(n29050), .B(n26453), .Z(n32567) );
  XOR U39387 ( .A(n32572), .B(n32567), .Z(n32561) );
  IV U39388 ( .A(n26454), .Z(n26456) );
  NOR U39389 ( .A(n26456), .B(n26455), .Z(n32566) );
  IV U39390 ( .A(n26457), .Z(n26459) );
  NOR U39391 ( .A(n26459), .B(n26458), .Z(n32559) );
  NOR U39392 ( .A(n32566), .B(n32559), .Z(n26460) );
  IV U39393 ( .A(n26460), .Z(n29498) );
  XOR U39394 ( .A(n32561), .B(n29498), .Z(n29508) );
  IV U39395 ( .A(n26461), .Z(n26462) );
  NOR U39396 ( .A(n26463), .B(n26462), .Z(n29506) );
  IV U39397 ( .A(n26464), .Z(n26466) );
  NOR U39398 ( .A(n26466), .B(n26465), .Z(n29504) );
  NOR U39399 ( .A(n29506), .B(n29504), .Z(n26467) );
  XOR U39400 ( .A(n29508), .B(n26467), .Z(n29502) );
  XOR U39401 ( .A(n29503), .B(n29502), .Z(n29043) );
  IV U39402 ( .A(n26468), .Z(n26469) );
  NOR U39403 ( .A(n26470), .B(n26469), .Z(n29513) );
  IV U39404 ( .A(n26471), .Z(n26472) );
  NOR U39405 ( .A(n26473), .B(n26472), .Z(n29042) );
  NOR U39406 ( .A(n29513), .B(n29042), .Z(n26474) );
  XOR U39407 ( .A(n29043), .B(n26474), .Z(n29035) );
  IV U39408 ( .A(n26475), .Z(n26477) );
  NOR U39409 ( .A(n26477), .B(n26476), .Z(n29039) );
  IV U39410 ( .A(n26478), .Z(n26479) );
  NOR U39411 ( .A(n26480), .B(n26479), .Z(n29036) );
  NOR U39412 ( .A(n29039), .B(n29036), .Z(n26481) );
  XOR U39413 ( .A(n29035), .B(n26481), .Z(n29519) );
  IV U39414 ( .A(n26482), .Z(n26484) );
  NOR U39415 ( .A(n26484), .B(n26483), .Z(n29518) );
  IV U39416 ( .A(n26485), .Z(n26486) );
  NOR U39417 ( .A(n26487), .B(n26486), .Z(n29522) );
  NOR U39418 ( .A(n29518), .B(n29522), .Z(n29034) );
  XOR U39419 ( .A(n29519), .B(n29034), .Z(n26488) );
  IV U39420 ( .A(n26488), .Z(n29536) );
  XOR U39421 ( .A(n29533), .B(n29536), .Z(n29529) );
  XOR U39422 ( .A(n26489), .B(n29529), .Z(n33097) );
  XOR U39423 ( .A(n29030), .B(n33097), .Z(n29032) );
  XOR U39424 ( .A(n29033), .B(n29032), .Z(n26490) );
  IV U39425 ( .A(n26490), .Z(n32538) );
  XOR U39426 ( .A(n29548), .B(n32538), .Z(n29561) );
  XOR U39427 ( .A(n29559), .B(n29561), .Z(n29554) );
  XOR U39428 ( .A(n29555), .B(n29554), .Z(n29551) );
  IV U39429 ( .A(n26491), .Z(n26492) );
  NOR U39430 ( .A(n26493), .B(n26492), .Z(n29550) );
  IV U39431 ( .A(n26494), .Z(n26495) );
  NOR U39432 ( .A(n26496), .B(n26495), .Z(n29577) );
  NOR U39433 ( .A(n29550), .B(n29577), .Z(n26497) );
  XOR U39434 ( .A(n29551), .B(n26497), .Z(n32518) );
  XOR U39435 ( .A(n29029), .B(n32518), .Z(n26498) );
  IV U39436 ( .A(n26498), .Z(n29592) );
  IV U39437 ( .A(n26499), .Z(n26500) );
  NOR U39438 ( .A(n26501), .B(n26500), .Z(n29591) );
  IV U39439 ( .A(n26502), .Z(n26503) );
  NOR U39440 ( .A(n26504), .B(n26503), .Z(n29589) );
  NOR U39441 ( .A(n29591), .B(n29589), .Z(n26505) );
  XOR U39442 ( .A(n29592), .B(n26505), .Z(n29027) );
  IV U39443 ( .A(n26506), .Z(n26508) );
  NOR U39444 ( .A(n26508), .B(n26507), .Z(n29585) );
  IV U39445 ( .A(n26509), .Z(n26510) );
  NOR U39446 ( .A(n26511), .B(n26510), .Z(n29026) );
  NOR U39447 ( .A(n29585), .B(n29026), .Z(n26512) );
  XOR U39448 ( .A(n29027), .B(n26512), .Z(n29025) );
  XOR U39449 ( .A(n29024), .B(n29025), .Z(n29018) );
  IV U39450 ( .A(n26513), .Z(n26515) );
  NOR U39451 ( .A(n26515), .B(n26514), .Z(n29021) );
  IV U39452 ( .A(n26516), .Z(n26517) );
  NOR U39453 ( .A(n26518), .B(n26517), .Z(n29017) );
  NOR U39454 ( .A(n29021), .B(n29017), .Z(n26519) );
  XOR U39455 ( .A(n29018), .B(n26519), .Z(n29617) );
  XOR U39456 ( .A(n29015), .B(n29617), .Z(n26520) );
  NOR U39457 ( .A(n26521), .B(n26520), .Z(n29620) );
  IV U39458 ( .A(n26522), .Z(n26523) );
  NOR U39459 ( .A(n26524), .B(n26523), .Z(n29615) );
  NOR U39460 ( .A(n29015), .B(n29615), .Z(n26525) );
  XOR U39461 ( .A(n29617), .B(n26525), .Z(n29610) );
  NOR U39462 ( .A(n26526), .B(n29610), .Z(n26527) );
  NOR U39463 ( .A(n29620), .B(n26527), .Z(n29626) );
  IV U39464 ( .A(n26528), .Z(n26530) );
  NOR U39465 ( .A(n26530), .B(n26529), .Z(n29609) );
  IV U39466 ( .A(n26531), .Z(n26532) );
  NOR U39467 ( .A(n26533), .B(n26532), .Z(n29625) );
  NOR U39468 ( .A(n29609), .B(n29625), .Z(n26534) );
  XOR U39469 ( .A(n29626), .B(n26534), .Z(n33158) );
  XOR U39470 ( .A(n29624), .B(n33158), .Z(n29631) );
  IV U39471 ( .A(n26535), .Z(n26536) );
  NOR U39472 ( .A(n26537), .B(n26536), .Z(n32502) );
  IV U39473 ( .A(n26538), .Z(n26539) );
  NOR U39474 ( .A(n26540), .B(n26539), .Z(n33169) );
  NOR U39475 ( .A(n32502), .B(n33169), .Z(n29632) );
  XOR U39476 ( .A(n29631), .B(n29632), .Z(n29638) );
  XOR U39477 ( .A(n26541), .B(n29638), .Z(n29640) );
  IV U39478 ( .A(n26542), .Z(n26544) );
  NOR U39479 ( .A(n26544), .B(n26543), .Z(n32499) );
  IV U39480 ( .A(n26545), .Z(n26547) );
  NOR U39481 ( .A(n26547), .B(n26546), .Z(n32494) );
  NOR U39482 ( .A(n32499), .B(n32494), .Z(n29641) );
  XOR U39483 ( .A(n29640), .B(n29641), .Z(n35834) );
  XOR U39484 ( .A(n29644), .B(n35834), .Z(n29645) );
  IV U39485 ( .A(n26548), .Z(n26550) );
  NOR U39486 ( .A(n26550), .B(n26549), .Z(n29652) );
  IV U39487 ( .A(n26551), .Z(n26553) );
  NOR U39488 ( .A(n26553), .B(n26552), .Z(n29648) );
  NOR U39489 ( .A(n29652), .B(n29648), .Z(n26554) );
  XOR U39490 ( .A(n29645), .B(n26554), .Z(n29660) );
  IV U39491 ( .A(n26555), .Z(n26556) );
  NOR U39492 ( .A(n26557), .B(n26556), .Z(n29650) );
  IV U39493 ( .A(n26558), .Z(n26559) );
  NOR U39494 ( .A(n26560), .B(n26559), .Z(n29659) );
  NOR U39495 ( .A(n29650), .B(n29659), .Z(n26561) );
  XOR U39496 ( .A(n29660), .B(n26561), .Z(n29657) );
  XOR U39497 ( .A(n29658), .B(n29657), .Z(n29013) );
  XOR U39498 ( .A(n29010), .B(n29013), .Z(n29008) );
  XOR U39499 ( .A(n26562), .B(n29008), .Z(n29005) );
  XOR U39500 ( .A(n29003), .B(n29005), .Z(n29000) );
  IV U39501 ( .A(n26563), .Z(n26564) );
  NOR U39502 ( .A(n26565), .B(n26564), .Z(n28999) );
  IV U39503 ( .A(n26566), .Z(n26567) );
  NOR U39504 ( .A(n26568), .B(n26567), .Z(n28997) );
  NOR U39505 ( .A(n28999), .B(n28997), .Z(n26569) );
  XOR U39506 ( .A(n29000), .B(n26569), .Z(n28990) );
  XOR U39507 ( .A(n26570), .B(n28990), .Z(n28988) );
  XOR U39508 ( .A(n28985), .B(n28988), .Z(n28980) );
  IV U39509 ( .A(n26571), .Z(n26572) );
  NOR U39510 ( .A(n26573), .B(n26572), .Z(n28986) );
  IV U39511 ( .A(n26574), .Z(n26576) );
  NOR U39512 ( .A(n26576), .B(n26575), .Z(n28979) );
  NOR U39513 ( .A(n28986), .B(n28979), .Z(n26577) );
  XOR U39514 ( .A(n28980), .B(n26577), .Z(n28978) );
  XOR U39515 ( .A(n28976), .B(n28978), .Z(n26578) );
  NOR U39516 ( .A(n26579), .B(n26578), .Z(n33199) );
  IV U39517 ( .A(n26580), .Z(n26581) );
  NOR U39518 ( .A(n26582), .B(n26581), .Z(n28974) );
  NOR U39519 ( .A(n28976), .B(n28974), .Z(n26583) );
  XOR U39520 ( .A(n28978), .B(n26583), .Z(n29668) );
  NOR U39521 ( .A(n26584), .B(n29668), .Z(n26585) );
  NOR U39522 ( .A(n33199), .B(n26585), .Z(n28971) );
  IV U39523 ( .A(n26586), .Z(n26588) );
  NOR U39524 ( .A(n26588), .B(n26587), .Z(n29667) );
  IV U39525 ( .A(n26589), .Z(n26590) );
  NOR U39526 ( .A(n26591), .B(n26590), .Z(n28970) );
  NOR U39527 ( .A(n29667), .B(n28970), .Z(n26592) );
  XOR U39528 ( .A(n28971), .B(n26592), .Z(n32451) );
  XOR U39529 ( .A(n29671), .B(n32451), .Z(n29673) );
  XOR U39530 ( .A(n26593), .B(n29673), .Z(n29678) );
  XOR U39531 ( .A(n29677), .B(n29678), .Z(n28964) );
  IV U39532 ( .A(n26594), .Z(n26596) );
  NOR U39533 ( .A(n26596), .B(n26595), .Z(n28967) );
  IV U39534 ( .A(n26597), .Z(n26599) );
  NOR U39535 ( .A(n26599), .B(n26598), .Z(n28963) );
  NOR U39536 ( .A(n28967), .B(n28963), .Z(n26600) );
  XOR U39537 ( .A(n28964), .B(n26600), .Z(n36564) );
  IV U39538 ( .A(n26601), .Z(n26603) );
  NOR U39539 ( .A(n26603), .B(n26602), .Z(n36559) );
  IV U39540 ( .A(n26604), .Z(n26605) );
  NOR U39541 ( .A(n26606), .B(n26605), .Z(n36574) );
  NOR U39542 ( .A(n36559), .B(n36574), .Z(n29685) );
  XOR U39543 ( .A(n36564), .B(n29685), .Z(n33223) );
  XOR U39544 ( .A(n28962), .B(n33223), .Z(n29694) );
  XOR U39545 ( .A(n29695), .B(n29694), .Z(n29691) );
  XOR U39546 ( .A(n29692), .B(n29691), .Z(n28959) );
  IV U39547 ( .A(n26607), .Z(n26609) );
  NOR U39548 ( .A(n26609), .B(n26608), .Z(n28958) );
  IV U39549 ( .A(n26610), .Z(n26612) );
  NOR U39550 ( .A(n26612), .B(n26611), .Z(n28956) );
  NOR U39551 ( .A(n28958), .B(n28956), .Z(n26613) );
  XOR U39552 ( .A(n28959), .B(n26613), .Z(n28952) );
  XOR U39553 ( .A(n33242), .B(n28952), .Z(n32433) );
  IV U39554 ( .A(n26614), .Z(n26616) );
  NOR U39555 ( .A(n26616), .B(n26615), .Z(n33244) );
  IV U39556 ( .A(n26617), .Z(n26618) );
  NOR U39557 ( .A(n26619), .B(n26618), .Z(n32431) );
  NOR U39558 ( .A(n33244), .B(n32431), .Z(n28953) );
  XOR U39559 ( .A(n32433), .B(n28953), .Z(n28949) );
  XOR U39560 ( .A(n28950), .B(n28949), .Z(n35758) );
  XOR U39561 ( .A(n28951), .B(n35758), .Z(n26620) );
  IV U39562 ( .A(n26620), .Z(n29712) );
  XOR U39563 ( .A(n29709), .B(n29712), .Z(n28947) );
  XOR U39564 ( .A(n26621), .B(n28947), .Z(n29723) );
  XOR U39565 ( .A(n29724), .B(n29723), .Z(n28944) );
  XOR U39566 ( .A(n28943), .B(n28944), .Z(n33256) );
  XOR U39567 ( .A(n29730), .B(n33256), .Z(n28941) );
  IV U39568 ( .A(n26622), .Z(n26623) );
  NOR U39569 ( .A(n26624), .B(n26623), .Z(n28940) );
  IV U39570 ( .A(n26625), .Z(n26627) );
  NOR U39571 ( .A(n26627), .B(n26626), .Z(n29739) );
  NOR U39572 ( .A(n28940), .B(n29739), .Z(n26628) );
  XOR U39573 ( .A(n28941), .B(n26628), .Z(n32423) );
  XOR U39574 ( .A(n33278), .B(n32423), .Z(n29747) );
  IV U39575 ( .A(n26629), .Z(n26631) );
  NOR U39576 ( .A(n26631), .B(n26630), .Z(n29746) );
  IV U39577 ( .A(n26632), .Z(n26633) );
  NOR U39578 ( .A(n26634), .B(n26633), .Z(n29749) );
  NOR U39579 ( .A(n29746), .B(n29749), .Z(n26635) );
  XOR U39580 ( .A(n29747), .B(n26635), .Z(n29753) );
  XOR U39581 ( .A(n26636), .B(n29753), .Z(n26647) );
  IV U39582 ( .A(n26647), .Z(n26637) );
  NOR U39583 ( .A(n26646), .B(n26637), .Z(n32416) );
  IV U39584 ( .A(n26638), .Z(n26639) );
  NOR U39585 ( .A(n26640), .B(n26639), .Z(n26643) );
  IV U39586 ( .A(n26643), .Z(n26642) );
  XOR U39587 ( .A(n29752), .B(n29753), .Z(n26641) );
  NOR U39588 ( .A(n26642), .B(n26641), .Z(n33288) );
  NOR U39589 ( .A(n32416), .B(n33288), .Z(n29758) );
  IV U39590 ( .A(n29758), .Z(n26645) );
  NOR U39591 ( .A(n26643), .B(n26647), .Z(n26644) );
  NOR U39592 ( .A(n26645), .B(n26644), .Z(n26649) );
  NOR U39593 ( .A(n26647), .B(n26646), .Z(n26648) );
  NOR U39594 ( .A(n26649), .B(n26648), .Z(n29761) );
  IV U39595 ( .A(n26650), .Z(n26651) );
  NOR U39596 ( .A(n26652), .B(n26651), .Z(n29759) );
  IV U39597 ( .A(n26653), .Z(n26654) );
  NOR U39598 ( .A(n26655), .B(n26654), .Z(n28935) );
  NOR U39599 ( .A(n29759), .B(n28935), .Z(n26656) );
  XOR U39600 ( .A(n29761), .B(n26656), .Z(n28933) );
  IV U39601 ( .A(n26657), .Z(n26659) );
  NOR U39602 ( .A(n26659), .B(n26658), .Z(n28937) );
  IV U39603 ( .A(n26660), .Z(n26661) );
  NOR U39604 ( .A(n26662), .B(n26661), .Z(n28932) );
  NOR U39605 ( .A(n28937), .B(n28932), .Z(n26663) );
  XOR U39606 ( .A(n28933), .B(n26663), .Z(n28931) );
  IV U39607 ( .A(n26664), .Z(n26666) );
  NOR U39608 ( .A(n26666), .B(n26665), .Z(n28929) );
  IV U39609 ( .A(n26667), .Z(n26669) );
  NOR U39610 ( .A(n26669), .B(n26668), .Z(n28927) );
  NOR U39611 ( .A(n28929), .B(n28927), .Z(n26670) );
  XOR U39612 ( .A(n28931), .B(n26670), .Z(n29766) );
  NOR U39613 ( .A(n26671), .B(n29766), .Z(n26674) );
  IV U39614 ( .A(n26671), .Z(n26673) );
  XOR U39615 ( .A(n28929), .B(n28931), .Z(n26672) );
  NOR U39616 ( .A(n26673), .B(n26672), .Z(n29774) );
  NOR U39617 ( .A(n26674), .B(n29774), .Z(n28924) );
  IV U39618 ( .A(n26675), .Z(n26677) );
  NOR U39619 ( .A(n26677), .B(n26676), .Z(n29765) );
  IV U39620 ( .A(n26678), .Z(n26680) );
  NOR U39621 ( .A(n26680), .B(n26679), .Z(n28923) );
  NOR U39622 ( .A(n29765), .B(n28923), .Z(n26681) );
  XOR U39623 ( .A(n28924), .B(n26681), .Z(n33300) );
  XOR U39624 ( .A(n28922), .B(n33300), .Z(n26682) );
  IV U39625 ( .A(n26682), .Z(n29791) );
  XOR U39626 ( .A(n29790), .B(n29791), .Z(n29780) );
  XOR U39627 ( .A(n26683), .B(n29780), .Z(n29786) );
  XOR U39628 ( .A(n26684), .B(n29786), .Z(n32380) );
  IV U39629 ( .A(n32380), .Z(n32394) );
  XOR U39630 ( .A(n32378), .B(n32394), .Z(n28913) );
  IV U39631 ( .A(n26685), .Z(n26687) );
  NOR U39632 ( .A(n26687), .B(n26686), .Z(n32389) );
  IV U39633 ( .A(n26688), .Z(n26689) );
  NOR U39634 ( .A(n26690), .B(n26689), .Z(n32377) );
  NOR U39635 ( .A(n32389), .B(n32377), .Z(n28915) );
  XOR U39636 ( .A(n28913), .B(n28915), .Z(n28917) );
  XOR U39637 ( .A(n26691), .B(n28917), .Z(n29807) );
  XOR U39638 ( .A(n29806), .B(n29807), .Z(n29815) );
  XOR U39639 ( .A(n26692), .B(n29815), .Z(n29825) );
  XOR U39640 ( .A(n29803), .B(n29825), .Z(n29829) );
  IV U39641 ( .A(n26693), .Z(n26695) );
  NOR U39642 ( .A(n26695), .B(n26694), .Z(n29824) );
  IV U39643 ( .A(n26696), .Z(n26698) );
  NOR U39644 ( .A(n26698), .B(n26697), .Z(n29828) );
  NOR U39645 ( .A(n29824), .B(n29828), .Z(n26699) );
  XOR U39646 ( .A(n29829), .B(n26699), .Z(n29833) );
  IV U39647 ( .A(n26700), .Z(n26702) );
  NOR U39648 ( .A(n26702), .B(n26701), .Z(n29834) );
  IV U39649 ( .A(n26703), .Z(n26704) );
  NOR U39650 ( .A(n26705), .B(n26704), .Z(n32352) );
  NOR U39651 ( .A(n29834), .B(n32352), .Z(n26706) );
  XOR U39652 ( .A(n29833), .B(n26706), .Z(n32347) );
  IV U39653 ( .A(n26707), .Z(n26708) );
  NOR U39654 ( .A(n26709), .B(n26708), .Z(n33324) );
  IV U39655 ( .A(n26710), .Z(n26712) );
  NOR U39656 ( .A(n26712), .B(n26711), .Z(n32346) );
  NOR U39657 ( .A(n33324), .B(n32346), .Z(n26713) );
  IV U39658 ( .A(n26713), .Z(n29836) );
  XOR U39659 ( .A(n32347), .B(n29836), .Z(n28910) );
  XOR U39660 ( .A(n28908), .B(n28910), .Z(n28904) );
  XOR U39661 ( .A(n26714), .B(n28904), .Z(n28896) );
  XOR U39662 ( .A(n26715), .B(n28896), .Z(n29843) );
  XOR U39663 ( .A(n28894), .B(n29843), .Z(n28891) );
  XOR U39664 ( .A(n26716), .B(n28891), .Z(n29845) );
  XOR U39665 ( .A(n29846), .B(n29845), .Z(n29852) );
  XOR U39666 ( .A(n29847), .B(n29852), .Z(n28888) );
  XOR U39667 ( .A(n26717), .B(n28888), .Z(n29856) );
  XOR U39668 ( .A(n26718), .B(n29856), .Z(n28885) );
  XOR U39669 ( .A(n26719), .B(n28885), .Z(n26731) );
  NOR U39670 ( .A(n26720), .B(n26731), .Z(n26723) );
  IV U39671 ( .A(n26720), .Z(n26722) );
  XOR U39672 ( .A(n28884), .B(n28885), .Z(n26721) );
  NOR U39673 ( .A(n26722), .B(n26721), .Z(n28880) );
  NOR U39674 ( .A(n26723), .B(n28880), .Z(n26734) );
  IV U39675 ( .A(n26734), .Z(n26724) );
  NOR U39676 ( .A(n26737), .B(n26724), .Z(n33376) );
  IV U39677 ( .A(n26725), .Z(n26726) );
  NOR U39678 ( .A(n26727), .B(n26726), .Z(n28876) );
  IV U39679 ( .A(n26728), .Z(n26729) );
  NOR U39680 ( .A(n26730), .B(n26729), .Z(n26735) );
  IV U39681 ( .A(n26735), .Z(n26733) );
  IV U39682 ( .A(n26731), .Z(n26732) );
  NOR U39683 ( .A(n26733), .B(n26732), .Z(n32329) );
  NOR U39684 ( .A(n26735), .B(n26734), .Z(n26736) );
  NOR U39685 ( .A(n32329), .B(n26736), .Z(n28877) );
  XOR U39686 ( .A(n28876), .B(n28877), .Z(n26739) );
  NOR U39687 ( .A(n28877), .B(n26737), .Z(n26738) );
  NOR U39688 ( .A(n26739), .B(n26738), .Z(n26740) );
  NOR U39689 ( .A(n33376), .B(n26740), .Z(n26741) );
  IV U39690 ( .A(n26741), .Z(n28874) );
  XOR U39691 ( .A(n26742), .B(n28874), .Z(n33387) );
  XOR U39692 ( .A(n28866), .B(n33387), .Z(n33396) );
  XOR U39693 ( .A(n28868), .B(n33396), .Z(n29878) );
  XOR U39694 ( .A(n26743), .B(n29878), .Z(n29871) );
  XOR U39695 ( .A(n26744), .B(n29871), .Z(n32321) );
  XOR U39696 ( .A(n29887), .B(n32321), .Z(n29888) );
  XOR U39697 ( .A(n29889), .B(n29888), .Z(n28864) );
  XOR U39698 ( .A(n28863), .B(n28864), .Z(n29896) );
  IV U39699 ( .A(n26745), .Z(n26747) );
  NOR U39700 ( .A(n26747), .B(n26746), .Z(n28861) );
  IV U39701 ( .A(n26748), .Z(n26749) );
  NOR U39702 ( .A(n26750), .B(n26749), .Z(n29895) );
  NOR U39703 ( .A(n28861), .B(n29895), .Z(n26751) );
  XOR U39704 ( .A(n29896), .B(n26751), .Z(n28858) );
  IV U39705 ( .A(n26752), .Z(n26753) );
  NOR U39706 ( .A(n26754), .B(n26753), .Z(n29892) );
  IV U39707 ( .A(n26755), .Z(n26757) );
  NOR U39708 ( .A(n26757), .B(n26756), .Z(n28859) );
  NOR U39709 ( .A(n29892), .B(n28859), .Z(n26758) );
  XOR U39710 ( .A(n28858), .B(n26758), .Z(n36747) );
  IV U39711 ( .A(n26759), .Z(n26760) );
  NOR U39712 ( .A(n26761), .B(n26760), .Z(n36742) );
  IV U39713 ( .A(n26762), .Z(n26764) );
  NOR U39714 ( .A(n26764), .B(n26763), .Z(n36754) );
  NOR U39715 ( .A(n36742), .B(n36754), .Z(n28856) );
  XOR U39716 ( .A(n36747), .B(n28856), .Z(n26765) );
  IV U39717 ( .A(n26765), .Z(n28853) );
  XOR U39718 ( .A(n28850), .B(n28853), .Z(n28847) );
  XOR U39719 ( .A(n26766), .B(n28847), .Z(n29904) );
  XOR U39720 ( .A(n29905), .B(n29904), .Z(n29918) );
  XOR U39721 ( .A(n26767), .B(n29918), .Z(n29910) );
  IV U39722 ( .A(n26768), .Z(n26769) );
  NOR U39723 ( .A(n26770), .B(n26769), .Z(n29914) );
  IV U39724 ( .A(n26771), .Z(n26773) );
  NOR U39725 ( .A(n26773), .B(n26772), .Z(n29911) );
  NOR U39726 ( .A(n29914), .B(n29911), .Z(n26774) );
  XOR U39727 ( .A(n29910), .B(n26774), .Z(n33440) );
  XOR U39728 ( .A(n29925), .B(n33440), .Z(n28843) );
  IV U39729 ( .A(n26775), .Z(n26776) );
  NOR U39730 ( .A(n26777), .B(n26776), .Z(n36784) );
  IV U39731 ( .A(n26778), .Z(n26780) );
  NOR U39732 ( .A(n26780), .B(n26779), .Z(n36798) );
  NOR U39733 ( .A(n36784), .B(n36798), .Z(n28844) );
  XOR U39734 ( .A(n28843), .B(n28844), .Z(n29936) );
  XOR U39735 ( .A(n26781), .B(n29936), .Z(n26791) );
  IV U39736 ( .A(n26782), .Z(n26783) );
  NOR U39737 ( .A(n26784), .B(n26783), .Z(n26794) );
  IV U39738 ( .A(n26785), .Z(n26786) );
  NOR U39739 ( .A(n26787), .B(n26786), .Z(n26790) );
  NOR U39740 ( .A(n26794), .B(n26790), .Z(n26788) );
  IV U39741 ( .A(n26788), .Z(n26789) );
  NOR U39742 ( .A(n26791), .B(n26789), .Z(n26798) );
  IV U39743 ( .A(n26790), .Z(n26793) );
  IV U39744 ( .A(n26791), .Z(n26792) );
  NOR U39745 ( .A(n26793), .B(n26792), .Z(n33454) );
  IV U39746 ( .A(n26794), .Z(n26796) );
  XOR U39747 ( .A(n29923), .B(n29936), .Z(n26795) );
  NOR U39748 ( .A(n26796), .B(n26795), .Z(n32286) );
  NOR U39749 ( .A(n33454), .B(n32286), .Z(n26797) );
  IV U39750 ( .A(n26797), .Z(n29938) );
  NOR U39751 ( .A(n26798), .B(n29938), .Z(n28836) );
  IV U39752 ( .A(n26799), .Z(n26801) );
  NOR U39753 ( .A(n26801), .B(n26800), .Z(n28835) );
  IV U39754 ( .A(n26802), .Z(n26804) );
  NOR U39755 ( .A(n26804), .B(n26803), .Z(n28838) );
  NOR U39756 ( .A(n28835), .B(n28838), .Z(n26805) );
  XOR U39757 ( .A(n28836), .B(n26805), .Z(n29942) );
  XOR U39758 ( .A(n28833), .B(n29942), .Z(n28831) );
  IV U39759 ( .A(n26806), .Z(n26807) );
  NOR U39760 ( .A(n26808), .B(n26807), .Z(n29941) );
  IV U39761 ( .A(n26809), .Z(n26811) );
  NOR U39762 ( .A(n26811), .B(n26810), .Z(n28830) );
  NOR U39763 ( .A(n29941), .B(n28830), .Z(n26812) );
  XOR U39764 ( .A(n28831), .B(n26812), .Z(n28824) );
  XOR U39765 ( .A(n28825), .B(n28824), .Z(n28822) );
  XOR U39766 ( .A(n28821), .B(n28822), .Z(n28816) );
  XOR U39767 ( .A(n26813), .B(n28816), .Z(n32267) );
  XOR U39768 ( .A(n29945), .B(n32267), .Z(n29951) );
  IV U39769 ( .A(n26814), .Z(n26815) );
  NOR U39770 ( .A(n26816), .B(n26815), .Z(n29946) );
  IV U39771 ( .A(n26817), .Z(n26818) );
  NOR U39772 ( .A(n26819), .B(n26818), .Z(n29950) );
  NOR U39773 ( .A(n29946), .B(n29950), .Z(n26820) );
  XOR U39774 ( .A(n29951), .B(n26820), .Z(n28813) );
  IV U39775 ( .A(n26821), .Z(n26822) );
  NOR U39776 ( .A(n26823), .B(n26822), .Z(n32260) );
  IV U39777 ( .A(n26824), .Z(n26825) );
  NOR U39778 ( .A(n26826), .B(n26825), .Z(n32252) );
  NOR U39779 ( .A(n32260), .B(n32252), .Z(n28814) );
  XOR U39780 ( .A(n28813), .B(n28814), .Z(n32246) );
  IV U39781 ( .A(n26827), .Z(n26829) );
  NOR U39782 ( .A(n26829), .B(n26828), .Z(n32249) );
  IV U39783 ( .A(n26830), .Z(n26831) );
  NOR U39784 ( .A(n26832), .B(n26831), .Z(n32245) );
  NOR U39785 ( .A(n32249), .B(n32245), .Z(n29958) );
  XOR U39786 ( .A(n32246), .B(n29958), .Z(n28811) );
  XOR U39787 ( .A(n26833), .B(n28811), .Z(n29973) );
  XOR U39788 ( .A(n29970), .B(n29973), .Z(n28808) );
  IV U39789 ( .A(n26834), .Z(n26835) );
  NOR U39790 ( .A(n26836), .B(n26835), .Z(n29972) );
  IV U39791 ( .A(n26837), .Z(n26838) );
  NOR U39792 ( .A(n26839), .B(n26838), .Z(n28807) );
  NOR U39793 ( .A(n29972), .B(n28807), .Z(n26840) );
  XOR U39794 ( .A(n28808), .B(n26840), .Z(n28799) );
  IV U39795 ( .A(n26841), .Z(n26843) );
  NOR U39796 ( .A(n26843), .B(n26842), .Z(n28804) );
  IV U39797 ( .A(n26844), .Z(n26846) );
  NOR U39798 ( .A(n26846), .B(n26845), .Z(n28800) );
  NOR U39799 ( .A(n28804), .B(n28800), .Z(n26847) );
  XOR U39800 ( .A(n28799), .B(n26847), .Z(n29979) );
  XOR U39801 ( .A(n28802), .B(n29979), .Z(n29984) );
  IV U39802 ( .A(n26848), .Z(n26849) );
  NOR U39803 ( .A(n26850), .B(n26849), .Z(n29978) );
  IV U39804 ( .A(n26851), .Z(n26853) );
  NOR U39805 ( .A(n26853), .B(n26852), .Z(n29983) );
  NOR U39806 ( .A(n29978), .B(n29983), .Z(n26854) );
  XOR U39807 ( .A(n29984), .B(n26854), .Z(n29981) );
  IV U39808 ( .A(n26855), .Z(n26857) );
  NOR U39809 ( .A(n26857), .B(n26856), .Z(n32231) );
  IV U39810 ( .A(n26858), .Z(n26860) );
  NOR U39811 ( .A(n26860), .B(n26859), .Z(n32226) );
  NOR U39812 ( .A(n32231), .B(n32226), .Z(n29982) );
  XOR U39813 ( .A(n29981), .B(n29982), .Z(n29991) );
  IV U39814 ( .A(n26861), .Z(n26862) );
  NOR U39815 ( .A(n26863), .B(n26862), .Z(n29990) );
  IV U39816 ( .A(n26864), .Z(n26865) );
  NOR U39817 ( .A(n26866), .B(n26865), .Z(n29988) );
  NOR U39818 ( .A(n29990), .B(n29988), .Z(n26867) );
  XOR U39819 ( .A(n29991), .B(n26867), .Z(n28793) );
  IV U39820 ( .A(n26868), .Z(n26870) );
  NOR U39821 ( .A(n26870), .B(n26869), .Z(n28796) );
  IV U39822 ( .A(n26871), .Z(n26872) );
  NOR U39823 ( .A(n26873), .B(n26872), .Z(n28792) );
  NOR U39824 ( .A(n28796), .B(n28792), .Z(n26874) );
  XOR U39825 ( .A(n28793), .B(n26874), .Z(n32207) );
  XOR U39826 ( .A(n29994), .B(n32207), .Z(n29995) );
  XOR U39827 ( .A(n29996), .B(n29995), .Z(n33511) );
  IV U39828 ( .A(n33511), .Z(n26881) );
  IV U39829 ( .A(n26875), .Z(n26877) );
  NOR U39830 ( .A(n26877), .B(n26876), .Z(n33509) );
  IV U39831 ( .A(n26878), .Z(n26879) );
  NOR U39832 ( .A(n26880), .B(n26879), .Z(n33520) );
  NOR U39833 ( .A(n33509), .B(n33520), .Z(n30002) );
  XOR U39834 ( .A(n26881), .B(n30002), .Z(n30004) );
  XOR U39835 ( .A(n30003), .B(n30004), .Z(n28790) );
  XOR U39836 ( .A(n26882), .B(n28790), .Z(n28787) );
  XOR U39837 ( .A(n28788), .B(n28787), .Z(n30016) );
  XOR U39838 ( .A(n30015), .B(n30016), .Z(n30013) );
  XOR U39839 ( .A(n30012), .B(n30013), .Z(n26889) );
  NOR U39840 ( .A(n26883), .B(n26889), .Z(n33536) );
  IV U39841 ( .A(n26884), .Z(n26886) );
  NOR U39842 ( .A(n26886), .B(n26885), .Z(n26890) );
  IV U39843 ( .A(n26890), .Z(n26887) );
  NOR U39844 ( .A(n26887), .B(n30013), .Z(n30010) );
  NOR U39845 ( .A(n33536), .B(n30010), .Z(n26888) );
  IV U39846 ( .A(n26888), .Z(n26896) );
  IV U39847 ( .A(n26889), .Z(n26894) );
  NOR U39848 ( .A(n26891), .B(n26890), .Z(n26892) );
  IV U39849 ( .A(n26892), .Z(n26893) );
  NOR U39850 ( .A(n26894), .B(n26893), .Z(n26895) );
  NOR U39851 ( .A(n26896), .B(n26895), .Z(n26897) );
  IV U39852 ( .A(n26897), .Z(n30033) );
  XOR U39853 ( .A(n30030), .B(n30033), .Z(n28785) );
  IV U39854 ( .A(n26898), .Z(n26899) );
  NOR U39855 ( .A(n26900), .B(n26899), .Z(n30032) );
  IV U39856 ( .A(n26901), .Z(n26902) );
  NOR U39857 ( .A(n26903), .B(n26902), .Z(n28784) );
  NOR U39858 ( .A(n30032), .B(n28784), .Z(n26904) );
  XOR U39859 ( .A(n28785), .B(n26904), .Z(n26910) );
  XOR U39860 ( .A(n26905), .B(n26910), .Z(n26913) );
  NOR U39861 ( .A(n26906), .B(n26913), .Z(n33545) );
  IV U39862 ( .A(n26907), .Z(n26908) );
  NOR U39863 ( .A(n26909), .B(n26908), .Z(n26915) );
  IV U39864 ( .A(n26915), .Z(n26912) );
  IV U39865 ( .A(n26910), .Z(n28782) );
  XOR U39866 ( .A(n28778), .B(n28782), .Z(n26911) );
  NOR U39867 ( .A(n26912), .B(n26911), .Z(n32183) );
  IV U39868 ( .A(n26913), .Z(n26914) );
  NOR U39869 ( .A(n26915), .B(n26914), .Z(n26916) );
  NOR U39870 ( .A(n32183), .B(n26916), .Z(n30038) );
  NOR U39871 ( .A(n26917), .B(n30038), .Z(n26918) );
  NOR U39872 ( .A(n33545), .B(n26918), .Z(n30042) );
  IV U39873 ( .A(n26919), .Z(n26921) );
  NOR U39874 ( .A(n26921), .B(n26920), .Z(n30037) );
  IV U39875 ( .A(n26922), .Z(n26924) );
  NOR U39876 ( .A(n26924), .B(n26923), .Z(n30041) );
  NOR U39877 ( .A(n30037), .B(n30041), .Z(n26925) );
  XOR U39878 ( .A(n30042), .B(n26925), .Z(n30049) );
  IV U39879 ( .A(n26926), .Z(n26927) );
  NOR U39880 ( .A(n26928), .B(n26927), .Z(n30045) );
  IV U39881 ( .A(n26929), .Z(n26930) );
  NOR U39882 ( .A(n26931), .B(n26930), .Z(n30047) );
  NOR U39883 ( .A(n30045), .B(n30047), .Z(n26932) );
  XOR U39884 ( .A(n30049), .B(n26932), .Z(n26933) );
  NOR U39885 ( .A(n26934), .B(n26933), .Z(n26937) );
  IV U39886 ( .A(n26934), .Z(n26936) );
  XOR U39887 ( .A(n30045), .B(n30049), .Z(n26935) );
  NOR U39888 ( .A(n26936), .B(n26935), .Z(n32176) );
  NOR U39889 ( .A(n26937), .B(n32176), .Z(n30053) );
  XOR U39890 ( .A(n26938), .B(n30053), .Z(n30065) );
  IV U39891 ( .A(n26939), .Z(n26941) );
  NOR U39892 ( .A(n26941), .B(n26940), .Z(n28776) );
  IV U39893 ( .A(n26942), .Z(n26944) );
  NOR U39894 ( .A(n26944), .B(n26943), .Z(n30064) );
  NOR U39895 ( .A(n28776), .B(n30064), .Z(n26945) );
  XOR U39896 ( .A(n30065), .B(n26945), .Z(n28774) );
  XOR U39897 ( .A(n28775), .B(n28774), .Z(n30072) );
  IV U39898 ( .A(n30072), .Z(n26952) );
  IV U39899 ( .A(n26946), .Z(n26947) );
  NOR U39900 ( .A(n26948), .B(n26947), .Z(n30075) );
  IV U39901 ( .A(n26949), .Z(n26951) );
  NOR U39902 ( .A(n26951), .B(n26950), .Z(n30070) );
  NOR U39903 ( .A(n30075), .B(n30070), .Z(n28773) );
  XOR U39904 ( .A(n26952), .B(n28773), .Z(n30081) );
  NOR U39905 ( .A(n26960), .B(n30081), .Z(n32160) );
  IV U39906 ( .A(n26953), .Z(n26954) );
  NOR U39907 ( .A(n26955), .B(n26954), .Z(n28767) );
  IV U39908 ( .A(n26956), .Z(n26957) );
  NOR U39909 ( .A(n26958), .B(n26957), .Z(n26959) );
  IV U39910 ( .A(n26959), .Z(n30082) );
  XOR U39911 ( .A(n30082), .B(n30081), .Z(n28768) );
  XOR U39912 ( .A(n28767), .B(n28768), .Z(n26962) );
  NOR U39913 ( .A(n28768), .B(n26960), .Z(n26961) );
  NOR U39914 ( .A(n26962), .B(n26961), .Z(n26963) );
  NOR U39915 ( .A(n32160), .B(n26963), .Z(n26964) );
  IV U39916 ( .A(n26964), .Z(n28765) );
  XOR U39917 ( .A(n28764), .B(n28765), .Z(n28760) );
  IV U39918 ( .A(n26965), .Z(n26967) );
  NOR U39919 ( .A(n26967), .B(n26966), .Z(n28762) );
  IV U39920 ( .A(n26968), .Z(n26969) );
  NOR U39921 ( .A(n26970), .B(n26969), .Z(n28759) );
  NOR U39922 ( .A(n28762), .B(n28759), .Z(n26971) );
  XOR U39923 ( .A(n28760), .B(n26971), .Z(n28752) );
  IV U39924 ( .A(n26972), .Z(n26974) );
  NOR U39925 ( .A(n26974), .B(n26973), .Z(n28753) );
  IV U39926 ( .A(n26975), .Z(n26977) );
  NOR U39927 ( .A(n26977), .B(n26976), .Z(n28755) );
  NOR U39928 ( .A(n28753), .B(n28755), .Z(n26978) );
  XOR U39929 ( .A(n28752), .B(n26978), .Z(n28750) );
  IV U39930 ( .A(n26979), .Z(n26981) );
  NOR U39931 ( .A(n26981), .B(n26980), .Z(n28749) );
  IV U39932 ( .A(n26982), .Z(n26983) );
  NOR U39933 ( .A(n26984), .B(n26983), .Z(n28746) );
  NOR U39934 ( .A(n28749), .B(n28746), .Z(n26985) );
  XOR U39935 ( .A(n28750), .B(n26985), .Z(n28742) );
  XOR U39936 ( .A(n28743), .B(n28742), .Z(n30090) );
  XOR U39937 ( .A(n26986), .B(n30090), .Z(n26998) );
  IV U39938 ( .A(n26987), .Z(n26988) );
  NOR U39939 ( .A(n26989), .B(n26988), .Z(n30092) );
  IV U39940 ( .A(n26990), .Z(n26992) );
  NOR U39941 ( .A(n26992), .B(n26991), .Z(n28740) );
  NOR U39942 ( .A(n30092), .B(n28740), .Z(n26993) );
  XOR U39943 ( .A(n26998), .B(n26993), .Z(n27001) );
  NOR U39944 ( .A(n26994), .B(n27001), .Z(n32134) );
  IV U39945 ( .A(n26995), .Z(n26996) );
  NOR U39946 ( .A(n26997), .B(n26996), .Z(n27003) );
  IV U39947 ( .A(n27003), .Z(n27000) );
  IV U39948 ( .A(n26998), .Z(n30093) );
  XOR U39949 ( .A(n30092), .B(n30093), .Z(n26999) );
  NOR U39950 ( .A(n27000), .B(n26999), .Z(n32132) );
  IV U39951 ( .A(n27001), .Z(n27002) );
  NOR U39952 ( .A(n27003), .B(n27002), .Z(n27004) );
  NOR U39953 ( .A(n32132), .B(n27004), .Z(n27012) );
  NOR U39954 ( .A(n27005), .B(n27012), .Z(n27006) );
  NOR U39955 ( .A(n32134), .B(n27006), .Z(n27020) );
  IV U39956 ( .A(n27020), .Z(n27007) );
  NOR U39957 ( .A(n27008), .B(n27007), .Z(n32129) );
  IV U39958 ( .A(n27009), .Z(n27010) );
  NOR U39959 ( .A(n27011), .B(n27010), .Z(n27016) );
  IV U39960 ( .A(n27016), .Z(n27014) );
  IV U39961 ( .A(n27012), .Z(n27013) );
  NOR U39962 ( .A(n27014), .B(n27013), .Z(n33596) );
  NOR U39963 ( .A(n32129), .B(n33596), .Z(n27015) );
  IV U39964 ( .A(n27015), .Z(n28739) );
  NOR U39965 ( .A(n27017), .B(n27016), .Z(n27018) );
  IV U39966 ( .A(n27018), .Z(n27019) );
  NOR U39967 ( .A(n27020), .B(n27019), .Z(n27021) );
  NOR U39968 ( .A(n28739), .B(n27021), .Z(n28734) );
  XOR U39969 ( .A(n27022), .B(n28734), .Z(n30105) );
  IV U39970 ( .A(n27023), .Z(n27025) );
  NOR U39971 ( .A(n27025), .B(n27024), .Z(n30104) );
  IV U39972 ( .A(n27026), .Z(n27028) );
  NOR U39973 ( .A(n27028), .B(n27027), .Z(n30101) );
  NOR U39974 ( .A(n30104), .B(n30101), .Z(n27029) );
  XOR U39975 ( .A(n30105), .B(n27029), .Z(n28730) );
  IV U39976 ( .A(n27030), .Z(n27032) );
  NOR U39977 ( .A(n27032), .B(n27031), .Z(n28731) );
  IV U39978 ( .A(n27033), .Z(n27034) );
  NOR U39979 ( .A(n27035), .B(n27034), .Z(n30115) );
  NOR U39980 ( .A(n28731), .B(n30115), .Z(n27036) );
  XOR U39981 ( .A(n28730), .B(n27036), .Z(n28728) );
  IV U39982 ( .A(n27037), .Z(n27038) );
  NOR U39983 ( .A(n27039), .B(n27038), .Z(n28727) );
  IV U39984 ( .A(n27040), .Z(n27042) );
  NOR U39985 ( .A(n27042), .B(n27041), .Z(n28725) );
  NOR U39986 ( .A(n28727), .B(n28725), .Z(n27043) );
  XOR U39987 ( .A(n28728), .B(n27043), .Z(n30122) );
  XOR U39988 ( .A(n27044), .B(n30122), .Z(n35398) );
  XOR U39989 ( .A(n30120), .B(n35398), .Z(n32107) );
  XOR U39990 ( .A(n27045), .B(n32107), .Z(n33626) );
  IV U39991 ( .A(n33626), .Z(n27052) );
  IV U39992 ( .A(n27046), .Z(n27048) );
  NOR U39993 ( .A(n27048), .B(n27047), .Z(n32106) );
  IV U39994 ( .A(n27049), .Z(n27051) );
  NOR U39995 ( .A(n27051), .B(n27050), .Z(n33624) );
  NOR U39996 ( .A(n32106), .B(n33624), .Z(n28718) );
  XOR U39997 ( .A(n27052), .B(n28718), .Z(n28714) );
  XOR U39998 ( .A(n28711), .B(n28714), .Z(n27053) );
  NOR U39999 ( .A(n27054), .B(n27053), .Z(n32094) );
  IV U40000 ( .A(n27055), .Z(n27056) );
  NOR U40001 ( .A(n27057), .B(n27056), .Z(n28713) );
  NOR U40002 ( .A(n28711), .B(n28713), .Z(n27058) );
  XOR U40003 ( .A(n27058), .B(n28714), .Z(n28708) );
  NOR U40004 ( .A(n27059), .B(n28708), .Z(n27060) );
  NOR U40005 ( .A(n32094), .B(n27060), .Z(n28702) );
  XOR U40006 ( .A(n27061), .B(n28702), .Z(n32088) );
  XOR U40007 ( .A(n28700), .B(n32088), .Z(n27062) );
  IV U40008 ( .A(n27062), .Z(n28697) );
  XOR U40009 ( .A(n28696), .B(n28697), .Z(n27069) );
  NOR U40010 ( .A(n27063), .B(n27069), .Z(n33644) );
  IV U40011 ( .A(n27064), .Z(n27065) );
  NOR U40012 ( .A(n27066), .B(n27065), .Z(n27070) );
  IV U40013 ( .A(n27070), .Z(n27067) );
  NOR U40014 ( .A(n27067), .B(n28697), .Z(n33637) );
  NOR U40015 ( .A(n33644), .B(n33637), .Z(n27068) );
  IV U40016 ( .A(n27068), .Z(n30137) );
  IV U40017 ( .A(n27069), .Z(n27074) );
  NOR U40018 ( .A(n27071), .B(n27070), .Z(n27072) );
  IV U40019 ( .A(n27072), .Z(n27073) );
  NOR U40020 ( .A(n27074), .B(n27073), .Z(n27075) );
  NOR U40021 ( .A(n30137), .B(n27075), .Z(n27076) );
  IV U40022 ( .A(n27076), .Z(n30140) );
  XOR U40023 ( .A(n30135), .B(n30140), .Z(n28694) );
  XOR U40024 ( .A(n27077), .B(n28694), .Z(n27078) );
  IV U40025 ( .A(n27078), .Z(n28692) );
  IV U40026 ( .A(n27079), .Z(n27080) );
  NOR U40027 ( .A(n27081), .B(n27080), .Z(n28690) );
  IV U40028 ( .A(n27082), .Z(n27083) );
  NOR U40029 ( .A(n27084), .B(n27083), .Z(n28688) );
  NOR U40030 ( .A(n28690), .B(n28688), .Z(n27085) );
  XOR U40031 ( .A(n28692), .B(n27085), .Z(n30143) );
  IV U40032 ( .A(n27086), .Z(n27087) );
  NOR U40033 ( .A(n27088), .B(n27087), .Z(n30142) );
  IV U40034 ( .A(n27089), .Z(n27091) );
  NOR U40035 ( .A(n27091), .B(n27090), .Z(n30145) );
  NOR U40036 ( .A(n30142), .B(n30145), .Z(n27092) );
  XOR U40037 ( .A(n30143), .B(n27092), .Z(n28686) );
  XOR U40038 ( .A(n28685), .B(n28686), .Z(n27096) );
  NOR U40039 ( .A(n27095), .B(n27096), .Z(n27093) );
  IV U40040 ( .A(n27093), .Z(n27094) );
  NOR U40041 ( .A(n27099), .B(n27094), .Z(n35343) );
  IV U40042 ( .A(n27095), .Z(n27098) );
  IV U40043 ( .A(n27096), .Z(n27097) );
  NOR U40044 ( .A(n27098), .B(n27097), .Z(n33668) );
  IV U40045 ( .A(n27099), .Z(n27100) );
  NOR U40046 ( .A(n28686), .B(n27100), .Z(n33671) );
  NOR U40047 ( .A(n33668), .B(n33671), .Z(n30153) );
  IV U40048 ( .A(n30153), .Z(n35337) );
  NOR U40049 ( .A(n35343), .B(n35337), .Z(n30159) );
  IV U40050 ( .A(n27101), .Z(n27102) );
  NOR U40051 ( .A(n27103), .B(n27102), .Z(n36986) );
  IV U40052 ( .A(n27104), .Z(n27105) );
  NOR U40053 ( .A(n27106), .B(n27105), .Z(n35334) );
  NOR U40054 ( .A(n36986), .B(n35334), .Z(n30161) );
  XOR U40055 ( .A(n30159), .B(n30161), .Z(n30166) );
  XOR U40056 ( .A(n27107), .B(n30166), .Z(n28679) );
  IV U40057 ( .A(n27108), .Z(n27109) );
  NOR U40058 ( .A(n27110), .B(n27109), .Z(n28678) );
  IV U40059 ( .A(n27111), .Z(n27112) );
  NOR U40060 ( .A(n27113), .B(n27112), .Z(n28681) );
  NOR U40061 ( .A(n28678), .B(n28681), .Z(n27114) );
  XOR U40062 ( .A(n28679), .B(n27114), .Z(n28676) );
  XOR U40063 ( .A(n27115), .B(n28676), .Z(n30172) );
  IV U40064 ( .A(n27116), .Z(n27117) );
  NOR U40065 ( .A(n27118), .B(n27117), .Z(n35314) );
  IV U40066 ( .A(n27119), .Z(n27120) );
  NOR U40067 ( .A(n27121), .B(n27120), .Z(n27122) );
  NOR U40068 ( .A(n35314), .B(n27122), .Z(n30173) );
  XOR U40069 ( .A(n30172), .B(n30173), .Z(n28671) );
  XOR U40070 ( .A(n27123), .B(n28671), .Z(n28666) );
  IV U40071 ( .A(n27124), .Z(n27126) );
  NOR U40072 ( .A(n27126), .B(n27125), .Z(n28665) );
  IV U40073 ( .A(n27127), .Z(n27129) );
  NOR U40074 ( .A(n27129), .B(n27128), .Z(n30185) );
  NOR U40075 ( .A(n28665), .B(n30185), .Z(n27130) );
  XOR U40076 ( .A(n28666), .B(n27130), .Z(n32070) );
  IV U40077 ( .A(n27131), .Z(n27132) );
  NOR U40078 ( .A(n27133), .B(n27132), .Z(n33708) );
  IV U40079 ( .A(n27134), .Z(n27135) );
  NOR U40080 ( .A(n27136), .B(n27135), .Z(n27137) );
  NOR U40081 ( .A(n33708), .B(n27137), .Z(n30184) );
  XOR U40082 ( .A(n32070), .B(n30184), .Z(n30190) );
  IV U40083 ( .A(n27138), .Z(n27139) );
  NOR U40084 ( .A(n27140), .B(n27139), .Z(n30194) );
  IV U40085 ( .A(n27141), .Z(n27142) );
  NOR U40086 ( .A(n27143), .B(n27142), .Z(n30196) );
  NOR U40087 ( .A(n30194), .B(n30196), .Z(n27144) );
  XOR U40088 ( .A(n30190), .B(n27144), .Z(n30209) );
  IV U40089 ( .A(n27145), .Z(n27147) );
  NOR U40090 ( .A(n27147), .B(n27146), .Z(n30189) );
  IV U40091 ( .A(n27148), .Z(n27150) );
  NOR U40092 ( .A(n27150), .B(n27149), .Z(n30208) );
  NOR U40093 ( .A(n30189), .B(n30208), .Z(n27151) );
  XOR U40094 ( .A(n30209), .B(n27151), .Z(n30211) );
  XOR U40095 ( .A(n30212), .B(n30211), .Z(n30213) );
  NOR U40096 ( .A(n27159), .B(n30213), .Z(n33722) );
  IV U40097 ( .A(n27152), .Z(n27153) );
  NOR U40098 ( .A(n27154), .B(n27153), .Z(n28661) );
  IV U40099 ( .A(n27155), .Z(n27156) );
  NOR U40100 ( .A(n27157), .B(n27156), .Z(n27158) );
  IV U40101 ( .A(n27158), .Z(n30214) );
  XOR U40102 ( .A(n30214), .B(n30213), .Z(n28662) );
  XOR U40103 ( .A(n28661), .B(n28662), .Z(n27161) );
  NOR U40104 ( .A(n28662), .B(n27159), .Z(n27160) );
  NOR U40105 ( .A(n27161), .B(n27160), .Z(n27162) );
  NOR U40106 ( .A(n33722), .B(n27162), .Z(n27163) );
  IV U40107 ( .A(n27163), .Z(n33725) );
  XOR U40108 ( .A(n28656), .B(n33725), .Z(n28650) );
  IV U40109 ( .A(n27164), .Z(n27166) );
  NOR U40110 ( .A(n27166), .B(n27165), .Z(n28657) );
  IV U40111 ( .A(n27167), .Z(n27169) );
  NOR U40112 ( .A(n27169), .B(n27168), .Z(n28649) );
  NOR U40113 ( .A(n28657), .B(n28649), .Z(n27170) );
  XOR U40114 ( .A(n28650), .B(n27170), .Z(n28654) );
  XOR U40115 ( .A(n28647), .B(n28654), .Z(n28645) );
  XOR U40116 ( .A(n27171), .B(n28645), .Z(n28642) );
  XOR U40117 ( .A(n28638), .B(n28642), .Z(n28636) );
  IV U40118 ( .A(n27172), .Z(n27173) );
  NOR U40119 ( .A(n27174), .B(n27173), .Z(n28640) );
  IV U40120 ( .A(n27175), .Z(n27176) );
  NOR U40121 ( .A(n27177), .B(n27176), .Z(n28635) );
  NOR U40122 ( .A(n28640), .B(n28635), .Z(n27178) );
  XOR U40123 ( .A(n28636), .B(n27178), .Z(n28632) );
  IV U40124 ( .A(n27179), .Z(n27181) );
  NOR U40125 ( .A(n27181), .B(n27180), .Z(n30219) );
  IV U40126 ( .A(n27182), .Z(n27184) );
  NOR U40127 ( .A(n27184), .B(n27183), .Z(n28633) );
  NOR U40128 ( .A(n30219), .B(n28633), .Z(n27185) );
  XOR U40129 ( .A(n28632), .B(n27185), .Z(n28630) );
  XOR U40130 ( .A(n28629), .B(n28630), .Z(n28625) );
  IV U40131 ( .A(n27186), .Z(n27188) );
  NOR U40132 ( .A(n27188), .B(n27187), .Z(n28627) );
  IV U40133 ( .A(n27189), .Z(n27191) );
  NOR U40134 ( .A(n27191), .B(n27190), .Z(n28624) );
  NOR U40135 ( .A(n28627), .B(n28624), .Z(n27192) );
  XOR U40136 ( .A(n28625), .B(n27192), .Z(n28622) );
  IV U40137 ( .A(n27193), .Z(n27195) );
  NOR U40138 ( .A(n27195), .B(n27194), .Z(n33765) );
  IV U40139 ( .A(n27196), .Z(n27197) );
  NOR U40140 ( .A(n27198), .B(n27197), .Z(n27199) );
  NOR U40141 ( .A(n33765), .B(n27199), .Z(n28623) );
  XOR U40142 ( .A(n28622), .B(n28623), .Z(n30232) );
  XOR U40143 ( .A(n30227), .B(n30232), .Z(n30224) );
  IV U40144 ( .A(n27200), .Z(n27202) );
  NOR U40145 ( .A(n27202), .B(n27201), .Z(n30223) );
  IV U40146 ( .A(n27203), .Z(n27204) );
  NOR U40147 ( .A(n27205), .B(n27204), .Z(n30245) );
  NOR U40148 ( .A(n30223), .B(n30245), .Z(n27206) );
  XOR U40149 ( .A(n30224), .B(n27206), .Z(n28621) );
  XOR U40150 ( .A(n27207), .B(n28621), .Z(n28612) );
  XOR U40151 ( .A(n28613), .B(n28612), .Z(n30249) );
  IV U40152 ( .A(n30249), .Z(n27215) );
  IV U40153 ( .A(n27208), .Z(n27210) );
  NOR U40154 ( .A(n27210), .B(n27209), .Z(n28614) );
  IV U40155 ( .A(n27211), .Z(n27213) );
  NOR U40156 ( .A(n27213), .B(n27212), .Z(n30248) );
  NOR U40157 ( .A(n28614), .B(n30248), .Z(n27214) );
  XOR U40158 ( .A(n27215), .B(n27214), .Z(n28611) );
  XOR U40159 ( .A(n28609), .B(n28611), .Z(n27216) );
  NOR U40160 ( .A(n27224), .B(n27216), .Z(n32013) );
  IV U40161 ( .A(n27217), .Z(n27219) );
  NOR U40162 ( .A(n27219), .B(n27218), .Z(n28596) );
  IV U40163 ( .A(n27220), .Z(n27221) );
  NOR U40164 ( .A(n27222), .B(n27221), .Z(n28607) );
  NOR U40165 ( .A(n28609), .B(n28607), .Z(n27223) );
  XOR U40166 ( .A(n28611), .B(n27223), .Z(n28597) );
  XOR U40167 ( .A(n28596), .B(n28597), .Z(n27226) );
  NOR U40168 ( .A(n28597), .B(n27224), .Z(n27225) );
  NOR U40169 ( .A(n27226), .B(n27225), .Z(n27227) );
  NOR U40170 ( .A(n32013), .B(n27227), .Z(n27228) );
  IV U40171 ( .A(n27228), .Z(n28603) );
  XOR U40172 ( .A(n28600), .B(n28603), .Z(n30258) );
  IV U40173 ( .A(n27229), .Z(n27230) );
  NOR U40174 ( .A(n27231), .B(n27230), .Z(n28602) );
  IV U40175 ( .A(n27232), .Z(n27233) );
  NOR U40176 ( .A(n27234), .B(n27233), .Z(n30257) );
  NOR U40177 ( .A(n28602), .B(n30257), .Z(n27235) );
  XOR U40178 ( .A(n30258), .B(n27235), .Z(n28593) );
  IV U40179 ( .A(n27236), .Z(n27238) );
  NOR U40180 ( .A(n27238), .B(n27237), .Z(n30254) );
  IV U40181 ( .A(n27239), .Z(n27241) );
  NOR U40182 ( .A(n27241), .B(n27240), .Z(n28594) );
  NOR U40183 ( .A(n30254), .B(n28594), .Z(n27242) );
  XOR U40184 ( .A(n28593), .B(n27242), .Z(n32000) );
  XOR U40185 ( .A(n28592), .B(n32000), .Z(n28590) );
  IV U40186 ( .A(n27243), .Z(n27245) );
  NOR U40187 ( .A(n27245), .B(n27244), .Z(n31993) );
  IV U40188 ( .A(n27246), .Z(n27247) );
  NOR U40189 ( .A(n27248), .B(n27247), .Z(n27249) );
  NOR U40190 ( .A(n31993), .B(n27249), .Z(n28591) );
  XOR U40191 ( .A(n28590), .B(n28591), .Z(n31986) );
  XOR U40192 ( .A(n27250), .B(n31986), .Z(n30270) );
  XOR U40193 ( .A(n28588), .B(n30270), .Z(n28586) );
  IV U40194 ( .A(n27251), .Z(n27253) );
  NOR U40195 ( .A(n27253), .B(n27252), .Z(n30269) );
  IV U40196 ( .A(n27254), .Z(n27255) );
  NOR U40197 ( .A(n27256), .B(n27255), .Z(n28585) );
  NOR U40198 ( .A(n30269), .B(n28585), .Z(n27257) );
  XOR U40199 ( .A(n28586), .B(n27257), .Z(n30273) );
  IV U40200 ( .A(n27258), .Z(n27259) );
  NOR U40201 ( .A(n27260), .B(n27259), .Z(n30278) );
  IV U40202 ( .A(n27261), .Z(n27263) );
  NOR U40203 ( .A(n27263), .B(n27262), .Z(n30274) );
  NOR U40204 ( .A(n30278), .B(n30274), .Z(n27264) );
  XOR U40205 ( .A(n30273), .B(n27264), .Z(n30286) );
  IV U40206 ( .A(n27265), .Z(n27266) );
  NOR U40207 ( .A(n27267), .B(n27266), .Z(n30287) );
  IV U40208 ( .A(n27268), .Z(n27269) );
  NOR U40209 ( .A(n27270), .B(n27269), .Z(n28581) );
  NOR U40210 ( .A(n30287), .B(n28581), .Z(n27271) );
  XOR U40211 ( .A(n30286), .B(n27271), .Z(n28577) );
  IV U40212 ( .A(n27272), .Z(n27274) );
  NOR U40213 ( .A(n27274), .B(n27273), .Z(n30285) );
  IV U40214 ( .A(n27275), .Z(n27277) );
  NOR U40215 ( .A(n27277), .B(n27276), .Z(n28576) );
  NOR U40216 ( .A(n30285), .B(n28576), .Z(n27278) );
  XOR U40217 ( .A(n28577), .B(n27278), .Z(n31966) );
  XOR U40218 ( .A(n30292), .B(n31966), .Z(n27279) );
  IV U40219 ( .A(n27279), .Z(n30294) );
  XOR U40220 ( .A(n30293), .B(n30294), .Z(n30304) );
  XOR U40221 ( .A(n27280), .B(n30304), .Z(n28573) );
  XOR U40222 ( .A(n27281), .B(n28573), .Z(n31950) );
  XOR U40223 ( .A(n30311), .B(n31950), .Z(n30313) );
  IV U40224 ( .A(n27282), .Z(n27283) );
  NOR U40225 ( .A(n27284), .B(n27283), .Z(n30312) );
  IV U40226 ( .A(n27285), .Z(n27286) );
  NOR U40227 ( .A(n27287), .B(n27286), .Z(n30317) );
  NOR U40228 ( .A(n30312), .B(n30317), .Z(n27288) );
  XOR U40229 ( .A(n30313), .B(n27288), .Z(n28572) );
  XOR U40230 ( .A(n28568), .B(n28572), .Z(n27289) );
  NOR U40231 ( .A(n27290), .B(n27289), .Z(n33803) );
  IV U40232 ( .A(n27291), .Z(n27292) );
  NOR U40233 ( .A(n27293), .B(n27292), .Z(n28570) );
  NOR U40234 ( .A(n28568), .B(n28570), .Z(n27294) );
  XOR U40235 ( .A(n28572), .B(n27294), .Z(n30321) );
  NOR U40236 ( .A(n27295), .B(n30321), .Z(n27296) );
  NOR U40237 ( .A(n33803), .B(n27296), .Z(n27297) );
  IV U40238 ( .A(n27297), .Z(n28566) );
  IV U40239 ( .A(n27298), .Z(n27300) );
  NOR U40240 ( .A(n27300), .B(n27299), .Z(n30320) );
  IV U40241 ( .A(n27301), .Z(n27303) );
  NOR U40242 ( .A(n27303), .B(n27302), .Z(n28565) );
  NOR U40243 ( .A(n30320), .B(n28565), .Z(n27304) );
  XOR U40244 ( .A(n28566), .B(n27304), .Z(n30327) );
  NOR U40245 ( .A(n30328), .B(n30327), .Z(n27309) );
  IV U40246 ( .A(n27305), .Z(n27306) );
  NOR U40247 ( .A(n27307), .B(n27306), .Z(n27310) );
  IV U40248 ( .A(n27310), .Z(n27308) );
  NOR U40249 ( .A(n27309), .B(n27308), .Z(n30333) );
  XOR U40250 ( .A(n30328), .B(n30327), .Z(n27313) );
  NOR U40251 ( .A(n27310), .B(n27313), .Z(n27311) );
  NOR U40252 ( .A(n30333), .B(n27311), .Z(n28562) );
  NOR U40253 ( .A(n27312), .B(n28562), .Z(n27316) );
  IV U40254 ( .A(n27312), .Z(n27315) );
  IV U40255 ( .A(n27313), .Z(n27314) );
  NOR U40256 ( .A(n27315), .B(n27314), .Z(n30335) );
  NOR U40257 ( .A(n27316), .B(n30335), .Z(n28558) );
  IV U40258 ( .A(n27317), .Z(n27319) );
  NOR U40259 ( .A(n27319), .B(n27318), .Z(n28561) );
  IV U40260 ( .A(n27320), .Z(n27322) );
  NOR U40261 ( .A(n27322), .B(n27321), .Z(n28557) );
  NOR U40262 ( .A(n28561), .B(n28557), .Z(n27323) );
  XOR U40263 ( .A(n28558), .B(n27323), .Z(n33826) );
  XOR U40264 ( .A(n33828), .B(n33826), .Z(n27324) );
  IV U40265 ( .A(n27324), .Z(n28553) );
  XOR U40266 ( .A(n28552), .B(n28553), .Z(n30341) );
  XOR U40267 ( .A(n27325), .B(n30341), .Z(n28539) );
  IV U40268 ( .A(n27326), .Z(n27328) );
  NOR U40269 ( .A(n27328), .B(n27327), .Z(n30337) );
  IV U40270 ( .A(n27329), .Z(n27331) );
  NOR U40271 ( .A(n27331), .B(n27330), .Z(n28540) );
  NOR U40272 ( .A(n30337), .B(n28540), .Z(n27332) );
  XOR U40273 ( .A(n28539), .B(n27332), .Z(n28545) );
  XOR U40274 ( .A(n28542), .B(n28545), .Z(n30347) );
  XOR U40275 ( .A(n27333), .B(n30347), .Z(n28537) );
  XOR U40276 ( .A(n27334), .B(n28537), .Z(n30357) );
  IV U40277 ( .A(n27335), .Z(n27336) );
  NOR U40278 ( .A(n27337), .B(n27336), .Z(n30361) );
  IV U40279 ( .A(n27338), .Z(n27339) );
  NOR U40280 ( .A(n27340), .B(n27339), .Z(n30356) );
  NOR U40281 ( .A(n30361), .B(n30356), .Z(n27341) );
  XOR U40282 ( .A(n30357), .B(n27341), .Z(n28532) );
  XOR U40283 ( .A(n28533), .B(n28532), .Z(n28535) );
  XOR U40284 ( .A(n27342), .B(n28535), .Z(n30377) );
  IV U40285 ( .A(n27343), .Z(n27345) );
  NOR U40286 ( .A(n27345), .B(n27344), .Z(n31916) );
  IV U40287 ( .A(n27346), .Z(n27347) );
  NOR U40288 ( .A(n27348), .B(n27347), .Z(n31909) );
  NOR U40289 ( .A(n31916), .B(n31909), .Z(n30378) );
  XOR U40290 ( .A(n30377), .B(n30378), .Z(n31904) );
  XOR U40291 ( .A(n31905), .B(n31904), .Z(n30383) );
  IV U40292 ( .A(n27349), .Z(n27351) );
  NOR U40293 ( .A(n27351), .B(n27350), .Z(n35135) );
  IV U40294 ( .A(n27352), .Z(n27353) );
  NOR U40295 ( .A(n27354), .B(n27353), .Z(n35130) );
  NOR U40296 ( .A(n35135), .B(n35130), .Z(n31903) );
  XOR U40297 ( .A(n30383), .B(n31903), .Z(n30388) );
  NOR U40298 ( .A(n27362), .B(n30388), .Z(n31895) );
  IV U40299 ( .A(n27355), .Z(n27357) );
  NOR U40300 ( .A(n27357), .B(n27356), .Z(n30391) );
  IV U40301 ( .A(n27358), .Z(n27359) );
  NOR U40302 ( .A(n27360), .B(n27359), .Z(n27361) );
  IV U40303 ( .A(n27361), .Z(n30389) );
  XOR U40304 ( .A(n30389), .B(n30388), .Z(n30392) );
  XOR U40305 ( .A(n30391), .B(n30392), .Z(n27364) );
  NOR U40306 ( .A(n30392), .B(n27362), .Z(n27363) );
  NOR U40307 ( .A(n27364), .B(n27363), .Z(n27365) );
  NOR U40308 ( .A(n31895), .B(n27365), .Z(n30395) );
  IV U40309 ( .A(n27366), .Z(n27368) );
  NOR U40310 ( .A(n27368), .B(n27367), .Z(n31889) );
  IV U40311 ( .A(n27369), .Z(n27370) );
  NOR U40312 ( .A(n27371), .B(n27370), .Z(n31884) );
  NOR U40313 ( .A(n31889), .B(n31884), .Z(n30396) );
  XOR U40314 ( .A(n30395), .B(n30396), .Z(n30399) );
  NOR U40315 ( .A(n27379), .B(n30399), .Z(n31878) );
  IV U40316 ( .A(n27372), .Z(n27373) );
  NOR U40317 ( .A(n27374), .B(n27373), .Z(n28525) );
  IV U40318 ( .A(n27375), .Z(n27376) );
  NOR U40319 ( .A(n27377), .B(n27376), .Z(n27378) );
  IV U40320 ( .A(n27378), .Z(n30400) );
  XOR U40321 ( .A(n30400), .B(n30399), .Z(n28526) );
  XOR U40322 ( .A(n28525), .B(n28526), .Z(n27381) );
  NOR U40323 ( .A(n28526), .B(n27379), .Z(n27380) );
  NOR U40324 ( .A(n27381), .B(n27380), .Z(n27382) );
  NOR U40325 ( .A(n31878), .B(n27382), .Z(n30403) );
  XOR U40326 ( .A(n30404), .B(n30403), .Z(n30409) );
  XOR U40327 ( .A(n27383), .B(n30409), .Z(n30412) );
  IV U40328 ( .A(n27384), .Z(n27386) );
  NOR U40329 ( .A(n27386), .B(n27385), .Z(n30411) );
  IV U40330 ( .A(n27387), .Z(n27388) );
  NOR U40331 ( .A(n27389), .B(n27388), .Z(n30415) );
  NOR U40332 ( .A(n30411), .B(n30415), .Z(n27390) );
  XOR U40333 ( .A(n30412), .B(n27390), .Z(n30422) );
  IV U40334 ( .A(n27391), .Z(n27393) );
  NOR U40335 ( .A(n27393), .B(n27392), .Z(n30418) );
  IV U40336 ( .A(n27394), .Z(n27395) );
  NOR U40337 ( .A(n27396), .B(n27395), .Z(n30421) );
  NOR U40338 ( .A(n30418), .B(n30421), .Z(n27397) );
  XOR U40339 ( .A(n30422), .B(n27397), .Z(n28520) );
  XOR U40340 ( .A(n27398), .B(n28520), .Z(n30435) );
  IV U40341 ( .A(n27399), .Z(n27401) );
  NOR U40342 ( .A(n27401), .B(n27400), .Z(n28519) );
  IV U40343 ( .A(n27402), .Z(n27404) );
  NOR U40344 ( .A(n27404), .B(n27403), .Z(n30434) );
  NOR U40345 ( .A(n28519), .B(n30434), .Z(n27405) );
  XOR U40346 ( .A(n30435), .B(n27405), .Z(n28518) );
  XOR U40347 ( .A(n35094), .B(n28518), .Z(n35085) );
  XOR U40348 ( .A(n30440), .B(n35085), .Z(n28511) );
  IV U40349 ( .A(n27406), .Z(n27407) );
  NOR U40350 ( .A(n27408), .B(n27407), .Z(n30443) );
  IV U40351 ( .A(n27409), .Z(n27411) );
  NOR U40352 ( .A(n27411), .B(n27410), .Z(n28510) );
  NOR U40353 ( .A(n30443), .B(n28510), .Z(n27412) );
  XOR U40354 ( .A(n28511), .B(n27412), .Z(n28516) );
  IV U40355 ( .A(n27413), .Z(n27415) );
  NOR U40356 ( .A(n27415), .B(n27414), .Z(n28508) );
  IV U40357 ( .A(n27416), .Z(n27418) );
  NOR U40358 ( .A(n27418), .B(n27417), .Z(n28514) );
  NOR U40359 ( .A(n28508), .B(n28514), .Z(n27419) );
  XOR U40360 ( .A(n28516), .B(n27419), .Z(n27420) );
  NOR U40361 ( .A(n27421), .B(n27420), .Z(n28506) );
  IV U40362 ( .A(n27421), .Z(n27423) );
  XOR U40363 ( .A(n28508), .B(n28516), .Z(n27422) );
  NOR U40364 ( .A(n27423), .B(n27422), .Z(n31840) );
  NOR U40365 ( .A(n28506), .B(n31840), .Z(n31834) );
  IV U40366 ( .A(n27424), .Z(n27425) );
  NOR U40367 ( .A(n27426), .B(n27425), .Z(n28505) );
  IV U40368 ( .A(n28505), .Z(n37239) );
  XOR U40369 ( .A(n31834), .B(n37239), .Z(n28503) );
  XOR U40370 ( .A(n27427), .B(n28503), .Z(n28496) );
  XOR U40371 ( .A(n28497), .B(n28496), .Z(n28499) );
  XOR U40372 ( .A(n27428), .B(n28499), .Z(n27429) );
  IV U40373 ( .A(n27429), .Z(n28488) );
  IV U40374 ( .A(n27430), .Z(n27432) );
  NOR U40375 ( .A(n27432), .B(n27431), .Z(n28493) );
  IV U40376 ( .A(n27433), .Z(n27434) );
  NOR U40377 ( .A(n27435), .B(n27434), .Z(n28487) );
  NOR U40378 ( .A(n28493), .B(n28487), .Z(n27436) );
  XOR U40379 ( .A(n28488), .B(n27436), .Z(n28480) );
  IV U40380 ( .A(n27437), .Z(n27439) );
  NOR U40381 ( .A(n27439), .B(n27438), .Z(n28484) );
  IV U40382 ( .A(n27440), .Z(n27442) );
  NOR U40383 ( .A(n27442), .B(n27441), .Z(n28481) );
  NOR U40384 ( .A(n28484), .B(n28481), .Z(n27443) );
  XOR U40385 ( .A(n28480), .B(n27443), .Z(n30456) );
  IV U40386 ( .A(n27444), .Z(n27445) );
  NOR U40387 ( .A(n27446), .B(n27445), .Z(n30459) );
  IV U40388 ( .A(n27447), .Z(n27448) );
  NOR U40389 ( .A(n27449), .B(n27448), .Z(n30454) );
  NOR U40390 ( .A(n30459), .B(n30454), .Z(n28479) );
  XOR U40391 ( .A(n30456), .B(n28479), .Z(n30466) );
  XOR U40392 ( .A(n27450), .B(n30466), .Z(n28471) );
  IV U40393 ( .A(n27451), .Z(n27452) );
  NOR U40394 ( .A(n27453), .B(n27452), .Z(n28476) );
  IV U40395 ( .A(n27454), .Z(n27456) );
  NOR U40396 ( .A(n27456), .B(n27455), .Z(n28470) );
  NOR U40397 ( .A(n28476), .B(n28470), .Z(n27457) );
  XOR U40398 ( .A(n28471), .B(n27457), .Z(n28464) );
  IV U40399 ( .A(n27458), .Z(n27460) );
  NOR U40400 ( .A(n27460), .B(n27459), .Z(n28467) );
  IV U40401 ( .A(n27461), .Z(n27462) );
  NOR U40402 ( .A(n27463), .B(n27462), .Z(n28465) );
  NOR U40403 ( .A(n28467), .B(n28465), .Z(n27464) );
  XOR U40404 ( .A(n28464), .B(n27464), .Z(n30474) );
  IV U40405 ( .A(n27465), .Z(n27466) );
  NOR U40406 ( .A(n27467), .B(n27466), .Z(n30473) );
  IV U40407 ( .A(n27468), .Z(n27469) );
  NOR U40408 ( .A(n27470), .B(n27469), .Z(n28462) );
  NOR U40409 ( .A(n30473), .B(n28462), .Z(n27471) );
  XOR U40410 ( .A(n30474), .B(n27471), .Z(n30479) );
  IV U40411 ( .A(n27472), .Z(n27474) );
  NOR U40412 ( .A(n27474), .B(n27473), .Z(n28459) );
  IV U40413 ( .A(n27475), .Z(n27477) );
  NOR U40414 ( .A(n27477), .B(n27476), .Z(n30478) );
  NOR U40415 ( .A(n28459), .B(n30478), .Z(n27478) );
  XOR U40416 ( .A(n30479), .B(n27478), .Z(n30491) );
  IV U40417 ( .A(n27479), .Z(n27480) );
  NOR U40418 ( .A(n27481), .B(n27480), .Z(n28457) );
  IV U40419 ( .A(n27482), .Z(n27483) );
  NOR U40420 ( .A(n27484), .B(n27483), .Z(n30489) );
  NOR U40421 ( .A(n28457), .B(n30489), .Z(n27485) );
  XOR U40422 ( .A(n30491), .B(n27485), .Z(n30487) );
  IV U40423 ( .A(n27486), .Z(n27488) );
  NOR U40424 ( .A(n27488), .B(n27487), .Z(n30486) );
  IV U40425 ( .A(n27489), .Z(n27490) );
  NOR U40426 ( .A(n27491), .B(n27490), .Z(n30498) );
  NOR U40427 ( .A(n30486), .B(n30498), .Z(n27492) );
  XOR U40428 ( .A(n30487), .B(n27492), .Z(n30503) );
  XOR U40429 ( .A(n30493), .B(n30503), .Z(n28451) );
  XOR U40430 ( .A(n28452), .B(n28451), .Z(n28454) );
  IV U40431 ( .A(n27493), .Z(n27494) );
  NOR U40432 ( .A(n27495), .B(n27494), .Z(n28453) );
  IV U40433 ( .A(n27496), .Z(n27497) );
  NOR U40434 ( .A(n27498), .B(n27497), .Z(n28449) );
  NOR U40435 ( .A(n28453), .B(n28449), .Z(n27499) );
  XOR U40436 ( .A(n28454), .B(n27499), .Z(n30511) );
  IV U40437 ( .A(n27500), .Z(n27501) );
  NOR U40438 ( .A(n27502), .B(n27501), .Z(n33911) );
  IV U40439 ( .A(n27503), .Z(n27504) );
  NOR U40440 ( .A(n27505), .B(n27504), .Z(n31775) );
  NOR U40441 ( .A(n33911), .B(n31775), .Z(n30512) );
  XOR U40442 ( .A(n30511), .B(n30512), .Z(n30516) );
  XOR U40443 ( .A(n30513), .B(n30516), .Z(n30524) );
  IV U40444 ( .A(n27506), .Z(n27507) );
  NOR U40445 ( .A(n27508), .B(n27507), .Z(n30515) );
  IV U40446 ( .A(n27509), .Z(n27511) );
  NOR U40447 ( .A(n27511), .B(n27510), .Z(n30523) );
  NOR U40448 ( .A(n30515), .B(n30523), .Z(n27512) );
  XOR U40449 ( .A(n30524), .B(n27512), .Z(n30521) );
  IV U40450 ( .A(n27513), .Z(n27514) );
  NOR U40451 ( .A(n27515), .B(n27514), .Z(n31768) );
  IV U40452 ( .A(n27516), .Z(n27517) );
  NOR U40453 ( .A(n27518), .B(n27517), .Z(n31763) );
  NOR U40454 ( .A(n31768), .B(n31763), .Z(n30522) );
  XOR U40455 ( .A(n30521), .B(n30522), .Z(n28447) );
  XOR U40456 ( .A(n28446), .B(n28447), .Z(n30531) );
  IV U40457 ( .A(n27519), .Z(n27520) );
  NOR U40458 ( .A(n27521), .B(n27520), .Z(n28444) );
  IV U40459 ( .A(n27522), .Z(n27523) );
  NOR U40460 ( .A(n27524), .B(n27523), .Z(n30530) );
  NOR U40461 ( .A(n28444), .B(n30530), .Z(n27525) );
  XOR U40462 ( .A(n30531), .B(n27525), .Z(n30528) );
  IV U40463 ( .A(n27526), .Z(n27527) );
  NOR U40464 ( .A(n27528), .B(n27527), .Z(n34996) );
  IV U40465 ( .A(n27529), .Z(n27530) );
  NOR U40466 ( .A(n27531), .B(n27530), .Z(n34988) );
  NOR U40467 ( .A(n34996), .B(n34988), .Z(n30529) );
  XOR U40468 ( .A(n30528), .B(n30529), .Z(n30547) );
  XOR U40469 ( .A(n30539), .B(n30547), .Z(n30535) );
  IV U40470 ( .A(n27532), .Z(n27534) );
  NOR U40471 ( .A(n27534), .B(n27533), .Z(n30546) );
  IV U40472 ( .A(n27535), .Z(n27536) );
  NOR U40473 ( .A(n27537), .B(n27536), .Z(n30534) );
  NOR U40474 ( .A(n30546), .B(n30534), .Z(n27538) );
  XOR U40475 ( .A(n30535), .B(n27538), .Z(n28437) );
  IV U40476 ( .A(n27539), .Z(n27540) );
  NOR U40477 ( .A(n27541), .B(n27540), .Z(n37308) );
  IV U40478 ( .A(n27542), .Z(n27544) );
  NOR U40479 ( .A(n27544), .B(n27543), .Z(n34974) );
  NOR U40480 ( .A(n37308), .B(n34974), .Z(n28438) );
  XOR U40481 ( .A(n28437), .B(n28438), .Z(n28442) );
  XOR U40482 ( .A(n28439), .B(n28442), .Z(n28435) );
  IV U40483 ( .A(n27545), .Z(n27546) );
  NOR U40484 ( .A(n27547), .B(n27546), .Z(n28441) );
  IV U40485 ( .A(n27548), .Z(n27549) );
  NOR U40486 ( .A(n27550), .B(n27549), .Z(n28434) );
  NOR U40487 ( .A(n28441), .B(n28434), .Z(n27551) );
  XOR U40488 ( .A(n28435), .B(n27551), .Z(n30553) );
  IV U40489 ( .A(n27552), .Z(n27554) );
  NOR U40490 ( .A(n27554), .B(n27553), .Z(n37323) );
  IV U40491 ( .A(n27555), .Z(n27557) );
  NOR U40492 ( .A(n27557), .B(n27556), .Z(n34966) );
  NOR U40493 ( .A(n37323), .B(n34966), .Z(n30554) );
  XOR U40494 ( .A(n30553), .B(n30554), .Z(n28432) );
  IV U40495 ( .A(n27558), .Z(n27559) );
  NOR U40496 ( .A(n27560), .B(n27559), .Z(n28431) );
  IV U40497 ( .A(n27561), .Z(n27562) );
  NOR U40498 ( .A(n27563), .B(n27562), .Z(n28429) );
  NOR U40499 ( .A(n28431), .B(n28429), .Z(n27564) );
  XOR U40500 ( .A(n28432), .B(n27564), .Z(n27577) );
  IV U40501 ( .A(n27577), .Z(n27565) );
  NOR U40502 ( .A(n27566), .B(n27565), .Z(n31740) );
  IV U40503 ( .A(n27567), .Z(n27569) );
  NOR U40504 ( .A(n27569), .B(n27568), .Z(n27573) );
  IV U40505 ( .A(n27573), .Z(n27571) );
  XOR U40506 ( .A(n28431), .B(n28432), .Z(n27570) );
  NOR U40507 ( .A(n27571), .B(n27570), .Z(n33934) );
  NOR U40508 ( .A(n31740), .B(n33934), .Z(n27572) );
  IV U40509 ( .A(n27572), .Z(n30564) );
  NOR U40510 ( .A(n27574), .B(n27573), .Z(n27575) );
  IV U40511 ( .A(n27575), .Z(n27576) );
  NOR U40512 ( .A(n27577), .B(n27576), .Z(n27578) );
  NOR U40513 ( .A(n30564), .B(n27578), .Z(n30562) );
  IV U40514 ( .A(n27579), .Z(n27580) );
  NOR U40515 ( .A(n27581), .B(n27580), .Z(n33936) );
  IV U40516 ( .A(n27582), .Z(n27584) );
  NOR U40517 ( .A(n27584), .B(n27583), .Z(n33944) );
  NOR U40518 ( .A(n33936), .B(n33944), .Z(n30563) );
  XOR U40519 ( .A(n30562), .B(n30563), .Z(n30567) );
  NOR U40520 ( .A(n27592), .B(n30567), .Z(n33951) );
  IV U40521 ( .A(n27585), .Z(n27586) );
  NOR U40522 ( .A(n27587), .B(n27586), .Z(n28425) );
  IV U40523 ( .A(n27588), .Z(n27590) );
  NOR U40524 ( .A(n27590), .B(n27589), .Z(n27591) );
  IV U40525 ( .A(n27591), .Z(n30568) );
  XOR U40526 ( .A(n30568), .B(n30567), .Z(n28426) );
  XOR U40527 ( .A(n28425), .B(n28426), .Z(n27594) );
  NOR U40528 ( .A(n28426), .B(n27592), .Z(n27593) );
  NOR U40529 ( .A(n27594), .B(n27593), .Z(n27595) );
  NOR U40530 ( .A(n33951), .B(n27595), .Z(n30571) );
  XOR U40531 ( .A(n30572), .B(n30571), .Z(n30583) );
  XOR U40532 ( .A(n27596), .B(n30583), .Z(n30579) );
  IV U40533 ( .A(n27597), .Z(n27598) );
  NOR U40534 ( .A(n27599), .B(n27598), .Z(n30578) );
  IV U40535 ( .A(n27600), .Z(n27602) );
  NOR U40536 ( .A(n27602), .B(n27601), .Z(n30594) );
  NOR U40537 ( .A(n30578), .B(n30594), .Z(n27603) );
  XOR U40538 ( .A(n30579), .B(n27603), .Z(n30601) );
  XOR U40539 ( .A(n30592), .B(n30601), .Z(n27604) );
  NOR U40540 ( .A(n27605), .B(n27604), .Z(n31727) );
  IV U40541 ( .A(n27606), .Z(n27607) );
  NOR U40542 ( .A(n27608), .B(n27607), .Z(n30599) );
  NOR U40543 ( .A(n30592), .B(n30599), .Z(n27609) );
  XOR U40544 ( .A(n30601), .B(n27609), .Z(n27613) );
  NOR U40545 ( .A(n27610), .B(n27613), .Z(n27611) );
  NOR U40546 ( .A(n31727), .B(n27611), .Z(n30603) );
  NOR U40547 ( .A(n27612), .B(n30603), .Z(n27616) );
  IV U40548 ( .A(n27612), .Z(n27615) );
  IV U40549 ( .A(n27613), .Z(n27614) );
  NOR U40550 ( .A(n27615), .B(n27614), .Z(n31730) );
  NOR U40551 ( .A(n27616), .B(n31730), .Z(n28420) );
  IV U40552 ( .A(n27617), .Z(n27619) );
  NOR U40553 ( .A(n27619), .B(n27618), .Z(n30602) );
  IV U40554 ( .A(n27620), .Z(n27621) );
  NOR U40555 ( .A(n27622), .B(n27621), .Z(n28419) );
  NOR U40556 ( .A(n30602), .B(n28419), .Z(n27623) );
  XOR U40557 ( .A(n28420), .B(n27623), .Z(n30610) );
  XOR U40558 ( .A(n30606), .B(n30610), .Z(n30616) );
  IV U40559 ( .A(n27624), .Z(n27626) );
  NOR U40560 ( .A(n27626), .B(n27625), .Z(n30608) );
  IV U40561 ( .A(n27627), .Z(n27628) );
  NOR U40562 ( .A(n27629), .B(n27628), .Z(n30615) );
  NOR U40563 ( .A(n30608), .B(n30615), .Z(n27630) );
  XOR U40564 ( .A(n30616), .B(n27630), .Z(n30612) );
  IV U40565 ( .A(n27631), .Z(n27632) );
  NOR U40566 ( .A(n27633), .B(n27632), .Z(n30613) );
  IV U40567 ( .A(n27634), .Z(n27635) );
  NOR U40568 ( .A(n27636), .B(n27635), .Z(n30620) );
  NOR U40569 ( .A(n30613), .B(n30620), .Z(n27637) );
  XOR U40570 ( .A(n30612), .B(n27637), .Z(n31716) );
  XOR U40571 ( .A(n30619), .B(n31716), .Z(n28417) );
  IV U40572 ( .A(n27638), .Z(n27639) );
  NOR U40573 ( .A(n27640), .B(n27639), .Z(n28416) );
  IV U40574 ( .A(n27641), .Z(n27642) );
  NOR U40575 ( .A(n27643), .B(n27642), .Z(n30626) );
  NOR U40576 ( .A(n28416), .B(n30626), .Z(n27644) );
  XOR U40577 ( .A(n28417), .B(n27644), .Z(n30630) );
  XOR U40578 ( .A(n27645), .B(n30630), .Z(n27646) );
  NOR U40579 ( .A(n27647), .B(n27646), .Z(n27650) );
  IV U40580 ( .A(n27647), .Z(n27649) );
  XOR U40581 ( .A(n30629), .B(n30630), .Z(n27648) );
  NOR U40582 ( .A(n27649), .B(n27648), .Z(n31703) );
  NOR U40583 ( .A(n27650), .B(n31703), .Z(n27651) );
  IV U40584 ( .A(n27651), .Z(n28411) );
  XOR U40585 ( .A(n28410), .B(n28411), .Z(n27652) );
  NOR U40586 ( .A(n27653), .B(n27652), .Z(n31698) );
  IV U40587 ( .A(n27654), .Z(n27656) );
  NOR U40588 ( .A(n27656), .B(n27655), .Z(n28408) );
  NOR U40589 ( .A(n28410), .B(n28408), .Z(n27657) );
  XOR U40590 ( .A(n27657), .B(n28411), .Z(n27667) );
  NOR U40591 ( .A(n27658), .B(n27667), .Z(n27659) );
  NOR U40592 ( .A(n31698), .B(n27659), .Z(n27665) );
  IV U40593 ( .A(n27665), .Z(n27660) );
  NOR U40594 ( .A(n27661), .B(n27660), .Z(n31693) );
  IV U40595 ( .A(n27662), .Z(n27663) );
  NOR U40596 ( .A(n27664), .B(n27663), .Z(n27666) );
  NOR U40597 ( .A(n27666), .B(n27665), .Z(n27670) );
  IV U40598 ( .A(n27666), .Z(n27669) );
  IV U40599 ( .A(n27667), .Z(n27668) );
  NOR U40600 ( .A(n27669), .B(n27668), .Z(n31695) );
  NOR U40601 ( .A(n27670), .B(n31695), .Z(n27671) );
  NOR U40602 ( .A(n27672), .B(n27671), .Z(n27673) );
  NOR U40603 ( .A(n31693), .B(n27673), .Z(n28404) );
  XOR U40604 ( .A(n27674), .B(n28404), .Z(n30640) );
  XOR U40605 ( .A(n27675), .B(n30640), .Z(n28401) );
  XOR U40606 ( .A(n28402), .B(n28401), .Z(n30667) );
  IV U40607 ( .A(n30667), .Z(n27682) );
  IV U40608 ( .A(n27676), .Z(n27677) );
  NOR U40609 ( .A(n27678), .B(n27677), .Z(n30670) );
  IV U40610 ( .A(n27679), .Z(n27680) );
  NOR U40611 ( .A(n27681), .B(n27680), .Z(n30664) );
  NOR U40612 ( .A(n30670), .B(n30664), .Z(n30661) );
  XOR U40613 ( .A(n27682), .B(n30661), .Z(n37370) );
  XOR U40614 ( .A(n28399), .B(n37370), .Z(n34860) );
  XOR U40615 ( .A(n30679), .B(n34860), .Z(n28397) );
  IV U40616 ( .A(n27683), .Z(n27684) );
  NOR U40617 ( .A(n27685), .B(n27684), .Z(n34009) );
  IV U40618 ( .A(n27686), .Z(n27688) );
  NOR U40619 ( .A(n27688), .B(n27687), .Z(n34001) );
  NOR U40620 ( .A(n34009), .B(n34001), .Z(n28398) );
  XOR U40621 ( .A(n28397), .B(n28398), .Z(n30690) );
  XOR U40622 ( .A(n30687), .B(n30690), .Z(n30695) );
  XOR U40623 ( .A(n27689), .B(n30695), .Z(n30702) );
  XOR U40624 ( .A(n30698), .B(n30702), .Z(n28395) );
  IV U40625 ( .A(n27690), .Z(n27692) );
  NOR U40626 ( .A(n27692), .B(n27691), .Z(n30700) );
  IV U40627 ( .A(n27693), .Z(n27694) );
  NOR U40628 ( .A(n27695), .B(n27694), .Z(n28394) );
  NOR U40629 ( .A(n30700), .B(n28394), .Z(n27696) );
  XOR U40630 ( .A(n28395), .B(n27696), .Z(n30707) );
  XOR U40631 ( .A(n30708), .B(n30707), .Z(n30710) );
  IV U40632 ( .A(n27697), .Z(n27698) );
  NOR U40633 ( .A(n27699), .B(n27698), .Z(n30709) );
  IV U40634 ( .A(n27700), .Z(n27701) );
  NOR U40635 ( .A(n27702), .B(n27701), .Z(n30704) );
  NOR U40636 ( .A(n30709), .B(n30704), .Z(n27703) );
  XOR U40637 ( .A(n30710), .B(n27703), .Z(n27704) );
  IV U40638 ( .A(n27704), .Z(n30728) );
  XOR U40639 ( .A(n30719), .B(n30728), .Z(n28392) );
  XOR U40640 ( .A(n27705), .B(n28392), .Z(n28385) );
  IV U40641 ( .A(n27706), .Z(n27707) );
  NOR U40642 ( .A(n27708), .B(n27707), .Z(n28388) );
  IV U40643 ( .A(n27709), .Z(n27710) );
  NOR U40644 ( .A(n27711), .B(n27710), .Z(n28386) );
  NOR U40645 ( .A(n28388), .B(n28386), .Z(n27712) );
  XOR U40646 ( .A(n28385), .B(n27712), .Z(n31640) );
  XOR U40647 ( .A(n30733), .B(n31640), .Z(n27713) );
  IV U40648 ( .A(n27713), .Z(n30735) );
  IV U40649 ( .A(n27714), .Z(n27715) );
  NOR U40650 ( .A(n27716), .B(n27715), .Z(n30734) );
  IV U40651 ( .A(n27717), .Z(n27718) );
  NOR U40652 ( .A(n27719), .B(n27718), .Z(n28383) );
  NOR U40653 ( .A(n30734), .B(n28383), .Z(n27720) );
  XOR U40654 ( .A(n30735), .B(n27720), .Z(n30741) );
  IV U40655 ( .A(n27721), .Z(n27723) );
  NOR U40656 ( .A(n27723), .B(n27722), .Z(n30740) );
  IV U40657 ( .A(n27724), .Z(n27726) );
  NOR U40658 ( .A(n27726), .B(n27725), .Z(n30748) );
  NOR U40659 ( .A(n30740), .B(n30748), .Z(n27727) );
  XOR U40660 ( .A(n30741), .B(n27727), .Z(n30755) );
  XOR U40661 ( .A(n30751), .B(n30755), .Z(n30758) );
  IV U40662 ( .A(n27728), .Z(n27729) );
  NOR U40663 ( .A(n27730), .B(n27729), .Z(n30753) );
  IV U40664 ( .A(n27731), .Z(n27733) );
  NOR U40665 ( .A(n27733), .B(n27732), .Z(n30757) );
  NOR U40666 ( .A(n30753), .B(n30757), .Z(n27734) );
  XOR U40667 ( .A(n30758), .B(n27734), .Z(n28381) );
  XOR U40668 ( .A(n28382), .B(n28381), .Z(n31615) );
  XOR U40669 ( .A(n28376), .B(n31615), .Z(n28374) );
  XOR U40670 ( .A(n27735), .B(n28374), .Z(n30770) );
  XOR U40671 ( .A(n27736), .B(n30770), .Z(n28368) );
  IV U40672 ( .A(n27737), .Z(n27738) );
  NOR U40673 ( .A(n27739), .B(n27738), .Z(n30762) );
  IV U40674 ( .A(n27740), .Z(n27741) );
  NOR U40675 ( .A(n27742), .B(n27741), .Z(n34826) );
  NOR U40676 ( .A(n30762), .B(n34826), .Z(n27743) );
  XOR U40677 ( .A(n28368), .B(n27743), .Z(n34048) );
  XOR U40678 ( .A(n28366), .B(n34048), .Z(n34054) );
  XOR U40679 ( .A(n30777), .B(n34054), .Z(n30778) );
  XOR U40680 ( .A(n34061), .B(n30778), .Z(n30783) );
  IV U40681 ( .A(n27744), .Z(n27746) );
  NOR U40682 ( .A(n27746), .B(n27745), .Z(n30782) );
  IV U40683 ( .A(n27747), .Z(n27748) );
  NOR U40684 ( .A(n27749), .B(n27748), .Z(n28364) );
  NOR U40685 ( .A(n30782), .B(n28364), .Z(n27750) );
  XOR U40686 ( .A(n30783), .B(n27750), .Z(n30786) );
  IV U40687 ( .A(n27751), .Z(n27752) );
  NOR U40688 ( .A(n27753), .B(n27752), .Z(n30787) );
  IV U40689 ( .A(n27754), .Z(n27756) );
  NOR U40690 ( .A(n27756), .B(n27755), .Z(n30789) );
  NOR U40691 ( .A(n30787), .B(n30789), .Z(n27757) );
  XOR U40692 ( .A(n30786), .B(n27757), .Z(n28362) );
  XOR U40693 ( .A(n28361), .B(n28362), .Z(n28357) );
  IV U40694 ( .A(n27758), .Z(n27760) );
  NOR U40695 ( .A(n27760), .B(n27759), .Z(n28359) );
  IV U40696 ( .A(n27761), .Z(n27762) );
  NOR U40697 ( .A(n27763), .B(n27762), .Z(n28356) );
  NOR U40698 ( .A(n28359), .B(n28356), .Z(n27764) );
  XOR U40699 ( .A(n28357), .B(n27764), .Z(n30801) );
  XOR U40700 ( .A(n30802), .B(n30801), .Z(n34789) );
  IV U40701 ( .A(n27765), .Z(n27766) );
  NOR U40702 ( .A(n27767), .B(n27766), .Z(n34784) );
  IV U40703 ( .A(n27768), .Z(n27769) );
  NOR U40704 ( .A(n27770), .B(n27769), .Z(n37482) );
  NOR U40705 ( .A(n34784), .B(n37482), .Z(n30803) );
  XOR U40706 ( .A(n34789), .B(n30803), .Z(n28353) );
  XOR U40707 ( .A(n27771), .B(n28353), .Z(n28351) );
  XOR U40708 ( .A(n27772), .B(n28351), .Z(n27773) );
  IV U40709 ( .A(n27773), .Z(n30814) );
  XOR U40710 ( .A(n30811), .B(n30814), .Z(n30821) );
  XOR U40711 ( .A(n27774), .B(n30821), .Z(n28341) );
  XOR U40712 ( .A(n27775), .B(n28341), .Z(n34774) );
  IV U40713 ( .A(n27776), .Z(n27778) );
  NOR U40714 ( .A(n27778), .B(n27777), .Z(n28344) );
  IV U40715 ( .A(n27779), .Z(n27781) );
  NOR U40716 ( .A(n27781), .B(n27780), .Z(n28336) );
  NOR U40717 ( .A(n28344), .B(n28336), .Z(n27782) );
  XOR U40718 ( .A(n34774), .B(n27782), .Z(n28338) );
  IV U40719 ( .A(n27783), .Z(n27784) );
  NOR U40720 ( .A(n27785), .B(n27784), .Z(n28339) );
  IV U40721 ( .A(n27786), .Z(n27787) );
  NOR U40722 ( .A(n27788), .B(n27787), .Z(n30824) );
  NOR U40723 ( .A(n28339), .B(n30824), .Z(n27789) );
  XOR U40724 ( .A(n28338), .B(n27789), .Z(n31578) );
  XOR U40725 ( .A(n30827), .B(n31578), .Z(n30828) );
  IV U40726 ( .A(n27790), .Z(n27792) );
  NOR U40727 ( .A(n27792), .B(n27791), .Z(n30838) );
  IV U40728 ( .A(n27793), .Z(n27794) );
  NOR U40729 ( .A(n27795), .B(n27794), .Z(n30841) );
  NOR U40730 ( .A(n30838), .B(n30841), .Z(n27796) );
  XOR U40731 ( .A(n30828), .B(n27796), .Z(n30833) );
  XOR U40732 ( .A(n27797), .B(n30833), .Z(n28333) );
  IV U40733 ( .A(n27798), .Z(n27799) );
  NOR U40734 ( .A(n27800), .B(n27799), .Z(n30851) );
  IV U40735 ( .A(n27801), .Z(n27802) );
  NOR U40736 ( .A(n27803), .B(n27802), .Z(n28334) );
  NOR U40737 ( .A(n30851), .B(n28334), .Z(n27804) );
  XOR U40738 ( .A(n28333), .B(n27804), .Z(n34742) );
  XOR U40739 ( .A(n30858), .B(n34742), .Z(n28331) );
  IV U40740 ( .A(n27805), .Z(n27806) );
  NOR U40741 ( .A(n27807), .B(n27806), .Z(n30859) );
  IV U40742 ( .A(n27808), .Z(n27810) );
  NOR U40743 ( .A(n27810), .B(n27809), .Z(n28330) );
  NOR U40744 ( .A(n30859), .B(n28330), .Z(n27811) );
  XOR U40745 ( .A(n28331), .B(n27811), .Z(n30865) );
  IV U40746 ( .A(n27812), .Z(n27814) );
  NOR U40747 ( .A(n27814), .B(n27813), .Z(n30864) );
  IV U40748 ( .A(n27815), .Z(n27817) );
  NOR U40749 ( .A(n27817), .B(n27816), .Z(n28328) );
  NOR U40750 ( .A(n30864), .B(n28328), .Z(n27818) );
  XOR U40751 ( .A(n30865), .B(n27818), .Z(n28322) );
  IV U40752 ( .A(n27819), .Z(n27820) );
  NOR U40753 ( .A(n27821), .B(n27820), .Z(n28325) );
  IV U40754 ( .A(n27822), .Z(n27823) );
  NOR U40755 ( .A(n27824), .B(n27823), .Z(n28323) );
  NOR U40756 ( .A(n28325), .B(n28323), .Z(n27825) );
  XOR U40757 ( .A(n28322), .B(n27825), .Z(n30880) );
  XOR U40758 ( .A(n27826), .B(n30880), .Z(n30874) );
  IV U40759 ( .A(n27827), .Z(n27828) );
  NOR U40760 ( .A(n27829), .B(n27828), .Z(n30883) );
  IV U40761 ( .A(n27830), .Z(n27832) );
  NOR U40762 ( .A(n27832), .B(n27831), .Z(n30873) );
  NOR U40763 ( .A(n30883), .B(n30873), .Z(n27833) );
  XOR U40764 ( .A(n30874), .B(n27833), .Z(n31543) );
  IV U40765 ( .A(n27834), .Z(n27836) );
  NOR U40766 ( .A(n27836), .B(n27835), .Z(n31546) );
  IV U40767 ( .A(n27837), .Z(n27839) );
  NOR U40768 ( .A(n27839), .B(n27838), .Z(n31540) );
  NOR U40769 ( .A(n31546), .B(n31540), .Z(n28318) );
  XOR U40770 ( .A(n31543), .B(n28318), .Z(n28320) );
  IV U40771 ( .A(n27840), .Z(n27841) );
  NOR U40772 ( .A(n27842), .B(n27841), .Z(n28319) );
  IV U40773 ( .A(n27843), .Z(n27845) );
  NOR U40774 ( .A(n27845), .B(n27844), .Z(n30893) );
  NOR U40775 ( .A(n28319), .B(n30893), .Z(n27846) );
  XOR U40776 ( .A(n28320), .B(n27846), .Z(n34115) );
  XOR U40777 ( .A(n27847), .B(n34115), .Z(n28316) );
  XOR U40778 ( .A(n28315), .B(n28316), .Z(n28311) );
  IV U40779 ( .A(n27848), .Z(n27849) );
  NOR U40780 ( .A(n27850), .B(n27849), .Z(n28313) );
  IV U40781 ( .A(n27851), .Z(n27853) );
  NOR U40782 ( .A(n27853), .B(n27852), .Z(n28310) );
  NOR U40783 ( .A(n28313), .B(n28310), .Z(n27854) );
  XOR U40784 ( .A(n28311), .B(n27854), .Z(n28304) );
  IV U40785 ( .A(n27855), .Z(n27857) );
  NOR U40786 ( .A(n27857), .B(n27856), .Z(n28307) );
  IV U40787 ( .A(n27858), .Z(n27859) );
  NOR U40788 ( .A(n27860), .B(n27859), .Z(n28305) );
  NOR U40789 ( .A(n28307), .B(n28305), .Z(n27861) );
  XOR U40790 ( .A(n28304), .B(n27861), .Z(n30907) );
  IV U40791 ( .A(n27862), .Z(n27863) );
  NOR U40792 ( .A(n27864), .B(n27863), .Z(n28302) );
  IV U40793 ( .A(n27865), .Z(n27867) );
  NOR U40794 ( .A(n27867), .B(n27866), .Z(n30906) );
  NOR U40795 ( .A(n28302), .B(n30906), .Z(n27868) );
  XOR U40796 ( .A(n30907), .B(n27868), .Z(n30899) );
  IV U40797 ( .A(n27869), .Z(n27871) );
  NOR U40798 ( .A(n27871), .B(n27870), .Z(n30903) );
  IV U40799 ( .A(n27872), .Z(n27873) );
  NOR U40800 ( .A(n27874), .B(n27873), .Z(n30898) );
  NOR U40801 ( .A(n30903), .B(n30898), .Z(n27875) );
  XOR U40802 ( .A(n30899), .B(n27875), .Z(n30919) );
  IV U40803 ( .A(n27876), .Z(n27877) );
  NOR U40804 ( .A(n27878), .B(n27877), .Z(n30915) );
  IV U40805 ( .A(n27879), .Z(n27881) );
  NOR U40806 ( .A(n27881), .B(n27880), .Z(n30917) );
  NOR U40807 ( .A(n30915), .B(n30917), .Z(n27882) );
  XOR U40808 ( .A(n30919), .B(n27882), .Z(n30921) );
  IV U40809 ( .A(n27883), .Z(n27885) );
  NOR U40810 ( .A(n27885), .B(n27884), .Z(n30920) );
  IV U40811 ( .A(n27886), .Z(n27887) );
  NOR U40812 ( .A(n27888), .B(n27887), .Z(n30924) );
  NOR U40813 ( .A(n30920), .B(n30924), .Z(n27889) );
  XOR U40814 ( .A(n30921), .B(n27889), .Z(n31518) );
  XOR U40815 ( .A(n28296), .B(n31518), .Z(n28294) );
  XOR U40816 ( .A(n27890), .B(n28294), .Z(n30930) );
  IV U40817 ( .A(n30930), .Z(n27898) );
  IV U40818 ( .A(n27891), .Z(n27893) );
  NOR U40819 ( .A(n27893), .B(n27892), .Z(n28291) );
  IV U40820 ( .A(n27894), .Z(n27896) );
  NOR U40821 ( .A(n27896), .B(n27895), .Z(n30928) );
  NOR U40822 ( .A(n28291), .B(n30928), .Z(n27897) );
  XOR U40823 ( .A(n27898), .B(n27897), .Z(n28289) );
  XOR U40824 ( .A(n28288), .B(n28289), .Z(n27899) );
  NOR U40825 ( .A(n27900), .B(n27899), .Z(n31500) );
  IV U40826 ( .A(n27901), .Z(n27902) );
  NOR U40827 ( .A(n27903), .B(n27902), .Z(n28285) );
  NOR U40828 ( .A(n28288), .B(n28285), .Z(n27904) );
  XOR U40829 ( .A(n27904), .B(n28289), .Z(n28281) );
  NOR U40830 ( .A(n27905), .B(n28281), .Z(n27906) );
  NOR U40831 ( .A(n31500), .B(n27906), .Z(n30940) );
  IV U40832 ( .A(n27907), .Z(n27909) );
  NOR U40833 ( .A(n27909), .B(n27908), .Z(n28280) );
  IV U40834 ( .A(n27910), .Z(n27911) );
  NOR U40835 ( .A(n27912), .B(n27911), .Z(n30939) );
  NOR U40836 ( .A(n28280), .B(n30939), .Z(n27913) );
  XOR U40837 ( .A(n30940), .B(n27913), .Z(n30938) );
  XOR U40838 ( .A(n27914), .B(n30938), .Z(n30945) );
  XOR U40839 ( .A(n30946), .B(n30945), .Z(n34670) );
  XOR U40840 ( .A(n28277), .B(n34670), .Z(n30951) );
  XOR U40841 ( .A(n30952), .B(n30951), .Z(n30963) );
  IV U40842 ( .A(n27915), .Z(n27916) );
  NOR U40843 ( .A(n27917), .B(n27916), .Z(n30964) );
  IV U40844 ( .A(n27918), .Z(n27919) );
  NOR U40845 ( .A(n27920), .B(n27919), .Z(n30960) );
  NOR U40846 ( .A(n30964), .B(n30960), .Z(n27921) );
  XOR U40847 ( .A(n30963), .B(n27921), .Z(n28272) );
  XOR U40848 ( .A(n27922), .B(n28272), .Z(n30977) );
  XOR U40849 ( .A(n30976), .B(n30977), .Z(n27923) );
  IV U40850 ( .A(n27923), .Z(n30972) );
  XOR U40851 ( .A(n30969), .B(n30972), .Z(n28269) );
  XOR U40852 ( .A(n27924), .B(n28269), .Z(n28262) );
  XOR U40853 ( .A(n28263), .B(n28262), .Z(n28265) );
  XOR U40854 ( .A(n28264), .B(n28265), .Z(n28258) );
  XOR U40855 ( .A(n27925), .B(n28258), .Z(n28254) );
  XOR U40856 ( .A(n27926), .B(n28254), .Z(n31006) );
  XOR U40857 ( .A(n31005), .B(n31006), .Z(n27927) );
  NOR U40858 ( .A(n27928), .B(n27927), .Z(n31009) );
  IV U40859 ( .A(n27929), .Z(n27930) );
  NOR U40860 ( .A(n27931), .B(n27930), .Z(n31003) );
  NOR U40861 ( .A(n31005), .B(n31003), .Z(n27932) );
  XOR U40862 ( .A(n27932), .B(n31006), .Z(n27933) );
  NOR U40863 ( .A(n27934), .B(n27933), .Z(n27935) );
  NOR U40864 ( .A(n31009), .B(n27935), .Z(n31011) );
  IV U40865 ( .A(n27936), .Z(n27938) );
  NOR U40866 ( .A(n27938), .B(n27937), .Z(n34165) );
  IV U40867 ( .A(n27939), .Z(n27940) );
  NOR U40868 ( .A(n27941), .B(n27940), .Z(n34172) );
  NOR U40869 ( .A(n34165), .B(n34172), .Z(n31012) );
  XOR U40870 ( .A(n31011), .B(n31012), .Z(n34177) );
  XOR U40871 ( .A(n34179), .B(n34177), .Z(n28249) );
  IV U40872 ( .A(n27942), .Z(n27943) );
  NOR U40873 ( .A(n27944), .B(n27943), .Z(n31451) );
  IV U40874 ( .A(n27945), .Z(n27947) );
  NOR U40875 ( .A(n27947), .B(n27946), .Z(n31445) );
  NOR U40876 ( .A(n31451), .B(n31445), .Z(n28250) );
  XOR U40877 ( .A(n28249), .B(n28250), .Z(n28252) );
  XOR U40878 ( .A(n27948), .B(n28252), .Z(n28245) );
  IV U40879 ( .A(n27949), .Z(n27951) );
  NOR U40880 ( .A(n27951), .B(n27950), .Z(n34182) );
  IV U40881 ( .A(n27952), .Z(n27953) );
  NOR U40882 ( .A(n27954), .B(n27953), .Z(n31434) );
  NOR U40883 ( .A(n34182), .B(n31434), .Z(n28246) );
  XOR U40884 ( .A(n28245), .B(n28246), .Z(n31025) );
  XOR U40885 ( .A(n28243), .B(n31025), .Z(n31031) );
  XOR U40886 ( .A(n31032), .B(n31031), .Z(n28241) );
  IV U40887 ( .A(n27955), .Z(n27956) );
  NOR U40888 ( .A(n27957), .B(n27956), .Z(n28240) );
  IV U40889 ( .A(n27958), .Z(n27959) );
  NOR U40890 ( .A(n27960), .B(n27959), .Z(n31043) );
  NOR U40891 ( .A(n28240), .B(n31043), .Z(n27961) );
  XOR U40892 ( .A(n28241), .B(n27961), .Z(n28238) );
  XOR U40893 ( .A(n28237), .B(n28238), .Z(n28233) );
  IV U40894 ( .A(n27962), .Z(n27964) );
  NOR U40895 ( .A(n27964), .B(n27963), .Z(n28235) );
  IV U40896 ( .A(n27965), .Z(n27966) );
  NOR U40897 ( .A(n27967), .B(n27966), .Z(n28232) );
  NOR U40898 ( .A(n28235), .B(n28232), .Z(n27968) );
  XOR U40899 ( .A(n28233), .B(n27968), .Z(n28226) );
  XOR U40900 ( .A(n27969), .B(n28226), .Z(n31415) );
  XOR U40901 ( .A(n28221), .B(n31415), .Z(n28223) );
  IV U40902 ( .A(n27970), .Z(n27971) );
  NOR U40903 ( .A(n27972), .B(n27971), .Z(n28222) );
  IV U40904 ( .A(n27973), .Z(n27975) );
  NOR U40905 ( .A(n27975), .B(n27974), .Z(n31062) );
  NOR U40906 ( .A(n28222), .B(n31062), .Z(n27976) );
  XOR U40907 ( .A(n28223), .B(n27976), .Z(n28219) );
  XOR U40908 ( .A(n28218), .B(n28219), .Z(n31076) );
  XOR U40909 ( .A(n27977), .B(n31076), .Z(n31072) );
  IV U40910 ( .A(n27978), .Z(n27980) );
  NOR U40911 ( .A(n27980), .B(n27979), .Z(n31073) );
  IV U40912 ( .A(n27981), .Z(n27983) );
  NOR U40913 ( .A(n27983), .B(n27982), .Z(n31081) );
  NOR U40914 ( .A(n31073), .B(n31081), .Z(n27984) );
  XOR U40915 ( .A(n31072), .B(n27984), .Z(n31086) );
  XOR U40916 ( .A(n31079), .B(n31086), .Z(n31089) );
  XOR U40917 ( .A(n27985), .B(n31089), .Z(n31092) );
  XOR U40918 ( .A(n31093), .B(n31092), .Z(n31095) );
  XOR U40919 ( .A(n31094), .B(n31095), .Z(n31389) );
  XOR U40920 ( .A(n31102), .B(n31389), .Z(n31099) );
  IV U40921 ( .A(n27986), .Z(n27987) );
  NOR U40922 ( .A(n27988), .B(n27987), .Z(n31103) );
  IV U40923 ( .A(n27989), .Z(n27990) );
  NOR U40924 ( .A(n27991), .B(n27990), .Z(n31098) );
  NOR U40925 ( .A(n31103), .B(n31098), .Z(n27992) );
  XOR U40926 ( .A(n31099), .B(n27992), .Z(n37699) );
  XOR U40927 ( .A(n31115), .B(n37699), .Z(n28007) );
  IV U40928 ( .A(n27993), .Z(n27994) );
  NOR U40929 ( .A(n27995), .B(n27994), .Z(n31111) );
  IV U40930 ( .A(n27996), .Z(n27997) );
  NOR U40931 ( .A(n27998), .B(n27997), .Z(n31109) );
  NOR U40932 ( .A(n31111), .B(n31109), .Z(n27999) );
  XOR U40933 ( .A(n28007), .B(n27999), .Z(n28010) );
  NOR U40934 ( .A(n28000), .B(n28010), .Z(n34221) );
  IV U40935 ( .A(n28001), .Z(n28002) );
  NOR U40936 ( .A(n28003), .B(n28002), .Z(n28018) );
  IV U40937 ( .A(n28018), .Z(n28015) );
  IV U40938 ( .A(n28004), .Z(n28006) );
  NOR U40939 ( .A(n28006), .B(n28005), .Z(n28012) );
  IV U40940 ( .A(n28012), .Z(n28009) );
  IV U40941 ( .A(n28007), .Z(n31112) );
  XOR U40942 ( .A(n31111), .B(n31112), .Z(n28008) );
  NOR U40943 ( .A(n28009), .B(n28008), .Z(n31380) );
  IV U40944 ( .A(n28010), .Z(n28011) );
  NOR U40945 ( .A(n28012), .B(n28011), .Z(n28013) );
  NOR U40946 ( .A(n31380), .B(n28013), .Z(n28021) );
  IV U40947 ( .A(n28021), .Z(n28014) );
  NOR U40948 ( .A(n28015), .B(n28014), .Z(n34230) );
  NOR U40949 ( .A(n34221), .B(n34230), .Z(n28016) );
  IV U40950 ( .A(n28016), .Z(n31125) );
  NOR U40951 ( .A(n28018), .B(n28017), .Z(n28019) );
  IV U40952 ( .A(n28019), .Z(n28020) );
  NOR U40953 ( .A(n28021), .B(n28020), .Z(n28022) );
  NOR U40954 ( .A(n31125), .B(n28022), .Z(n31128) );
  XOR U40955 ( .A(n31131), .B(n31128), .Z(n37725) );
  XOR U40956 ( .A(n31126), .B(n37725), .Z(n31137) );
  XOR U40957 ( .A(n31138), .B(n31137), .Z(n31374) );
  XOR U40958 ( .A(n31139), .B(n31374), .Z(n28207) );
  IV U40959 ( .A(n28023), .Z(n28024) );
  NOR U40960 ( .A(n28025), .B(n28024), .Z(n28212) );
  IV U40961 ( .A(n28026), .Z(n28028) );
  NOR U40962 ( .A(n28028), .B(n28027), .Z(n28206) );
  NOR U40963 ( .A(n28212), .B(n28206), .Z(n28029) );
  XOR U40964 ( .A(n28207), .B(n28029), .Z(n31148) );
  IV U40965 ( .A(n28030), .Z(n28032) );
  NOR U40966 ( .A(n28032), .B(n28031), .Z(n28209) );
  IV U40967 ( .A(n28033), .Z(n28034) );
  NOR U40968 ( .A(n28035), .B(n28034), .Z(n31147) );
  NOR U40969 ( .A(n28209), .B(n31147), .Z(n28036) );
  XOR U40970 ( .A(n31148), .B(n28036), .Z(n31144) );
  IV U40971 ( .A(n28037), .Z(n28038) );
  NOR U40972 ( .A(n28039), .B(n28038), .Z(n31145) );
  IV U40973 ( .A(n28040), .Z(n28042) );
  NOR U40974 ( .A(n28042), .B(n28041), .Z(n31151) );
  NOR U40975 ( .A(n31145), .B(n31151), .Z(n28043) );
  XOR U40976 ( .A(n31144), .B(n28043), .Z(n28204) );
  XOR U40977 ( .A(n28201), .B(n28204), .Z(n28198) );
  XOR U40978 ( .A(n28044), .B(n28198), .Z(n28195) );
  XOR U40979 ( .A(n28196), .B(n28195), .Z(n28193) );
  XOR U40980 ( .A(n28190), .B(n28193), .Z(n28188) );
  XOR U40981 ( .A(n28045), .B(n28188), .Z(n31156) );
  XOR U40982 ( .A(n31157), .B(n31156), .Z(n31159) );
  XOR U40983 ( .A(n31158), .B(n31159), .Z(n28185) );
  XOR U40984 ( .A(n28046), .B(n28185), .Z(n31170) );
  IV U40985 ( .A(n28047), .Z(n28048) );
  NOR U40986 ( .A(n28049), .B(n28048), .Z(n34277) );
  IV U40987 ( .A(n28050), .Z(n28051) );
  NOR U40988 ( .A(n28052), .B(n28051), .Z(n28053) );
  NOR U40989 ( .A(n34277), .B(n28053), .Z(n31171) );
  XOR U40990 ( .A(n31170), .B(n31171), .Z(n34282) );
  XOR U40991 ( .A(n28181), .B(n34282), .Z(n31175) );
  IV U40992 ( .A(n28054), .Z(n28055) );
  NOR U40993 ( .A(n28056), .B(n28055), .Z(n31340) );
  IV U40994 ( .A(n28057), .Z(n28058) );
  NOR U40995 ( .A(n28059), .B(n28058), .Z(n31333) );
  NOR U40996 ( .A(n31340), .B(n31333), .Z(n31176) );
  XOR U40997 ( .A(n31175), .B(n31176), .Z(n31186) );
  XOR U40998 ( .A(n28060), .B(n31186), .Z(n31181) );
  XOR U40999 ( .A(n28061), .B(n31181), .Z(n31197) );
  XOR U41000 ( .A(n31196), .B(n31197), .Z(n28179) );
  XOR U41001 ( .A(n28062), .B(n28179), .Z(n31213) );
  XOR U41002 ( .A(n31214), .B(n31213), .Z(n34304) );
  XOR U41003 ( .A(n28063), .B(n34304), .Z(n31318) );
  XOR U41004 ( .A(n28170), .B(n31318), .Z(n28166) );
  IV U41005 ( .A(n28166), .Z(n28172) );
  XOR U41006 ( .A(n28171), .B(n28172), .Z(n31222) );
  XOR U41007 ( .A(n28064), .B(n31222), .Z(n28156) );
  IV U41008 ( .A(n28065), .Z(n28067) );
  NOR U41009 ( .A(n28067), .B(n28066), .Z(n31218) );
  IV U41010 ( .A(n28068), .Z(n28070) );
  NOR U41011 ( .A(n28070), .B(n28069), .Z(n28157) );
  NOR U41012 ( .A(n31218), .B(n28157), .Z(n28071) );
  XOR U41013 ( .A(n28156), .B(n28071), .Z(n28162) );
  XOR U41014 ( .A(n28072), .B(n28162), .Z(n31298) );
  XOR U41015 ( .A(n28151), .B(n31298), .Z(n34332) );
  XOR U41016 ( .A(n28153), .B(n34332), .Z(n28150) );
  XOR U41017 ( .A(n28148), .B(n28150), .Z(n28144) );
  IV U41018 ( .A(n28073), .Z(n28075) );
  NOR U41019 ( .A(n28075), .B(n28074), .Z(n28146) );
  IV U41020 ( .A(n28076), .Z(n28077) );
  NOR U41021 ( .A(n28078), .B(n28077), .Z(n28143) );
  NOR U41022 ( .A(n28146), .B(n28143), .Z(n28079) );
  XOR U41023 ( .A(n28144), .B(n28079), .Z(n28136) );
  IV U41024 ( .A(n28080), .Z(n28081) );
  NOR U41025 ( .A(n28082), .B(n28081), .Z(n34343) );
  IV U41026 ( .A(n28083), .Z(n28085) );
  NOR U41027 ( .A(n28085), .B(n28084), .Z(n31288) );
  NOR U41028 ( .A(n34343), .B(n31288), .Z(n28137) );
  XOR U41029 ( .A(n28136), .B(n28137), .Z(n28139) );
  XOR U41030 ( .A(n28138), .B(n28139), .Z(n28128) );
  IV U41031 ( .A(n28086), .Z(n28087) );
  NOR U41032 ( .A(n28088), .B(n28087), .Z(n28134) );
  IV U41033 ( .A(n28089), .Z(n28091) );
  NOR U41034 ( .A(n28091), .B(n28090), .Z(n28127) );
  NOR U41035 ( .A(n28134), .B(n28127), .Z(n28092) );
  XOR U41036 ( .A(n28128), .B(n28092), .Z(n28130) );
  IV U41037 ( .A(n28093), .Z(n28095) );
  NOR U41038 ( .A(n28095), .B(n28094), .Z(n28131) );
  IV U41039 ( .A(n28096), .Z(n28098) );
  NOR U41040 ( .A(n28098), .B(n28097), .Z(n31232) );
  NOR U41041 ( .A(n28131), .B(n31232), .Z(n28099) );
  XOR U41042 ( .A(n28130), .B(n28099), .Z(n31230) );
  XOR U41043 ( .A(n31229), .B(n31230), .Z(n28123) );
  IV U41044 ( .A(n28100), .Z(n28101) );
  NOR U41045 ( .A(n28102), .B(n28101), .Z(n28125) );
  IV U41046 ( .A(n28103), .Z(n28105) );
  NOR U41047 ( .A(n28105), .B(n28104), .Z(n28122) );
  NOR U41048 ( .A(n28125), .B(n28122), .Z(n28106) );
  XOR U41049 ( .A(n28123), .B(n28106), .Z(n28119) );
  IV U41050 ( .A(n28107), .Z(n28109) );
  NOR U41051 ( .A(n28109), .B(n28108), .Z(n31238) );
  IV U41052 ( .A(n28110), .Z(n28111) );
  NOR U41053 ( .A(n28112), .B(n28111), .Z(n28120) );
  NOR U41054 ( .A(n31238), .B(n28120), .Z(n28113) );
  XOR U41055 ( .A(n28119), .B(n28113), .Z(n31247) );
  NOR U41056 ( .A(n28114), .B(n31247), .Z(n34441) );
  IV U41057 ( .A(n28115), .Z(n28117) );
  NOR U41058 ( .A(n28117), .B(n28116), .Z(n31254) );
  IV U41059 ( .A(n31254), .Z(n28118) );
  NOR U41060 ( .A(n28118), .B(n31247), .Z(n37881) );
  NOR U41061 ( .A(n34441), .B(n37881), .Z(n31272) );
  IV U41062 ( .A(n28119), .Z(n31240) );
  IV U41063 ( .A(n28120), .Z(n28121) );
  NOR U41064 ( .A(n31240), .B(n28121), .Z(n31242) );
  IV U41065 ( .A(n31242), .Z(n31237) );
  IV U41066 ( .A(n28122), .Z(n28124) );
  NOR U41067 ( .A(n28124), .B(n28123), .Z(n34358) );
  IV U41068 ( .A(n28125), .Z(n28126) );
  NOR U41069 ( .A(n28126), .B(n31230), .Z(n34355) );
  IV U41070 ( .A(n28127), .Z(n28129) );
  NOR U41071 ( .A(n28129), .B(n28128), .Z(n31281) );
  IV U41072 ( .A(n28130), .Z(n31234) );
  IV U41073 ( .A(n28131), .Z(n28132) );
  NOR U41074 ( .A(n31234), .B(n28132), .Z(n28133) );
  IV U41075 ( .A(n28133), .Z(n34347) );
  IV U41076 ( .A(n28134), .Z(n28135) );
  NOR U41077 ( .A(n28135), .B(n28139), .Z(n31279) );
  IV U41078 ( .A(n28136), .Z(n31289) );
  NOR U41079 ( .A(n31289), .B(n28137), .Z(n28141) );
  IV U41080 ( .A(n28138), .Z(n28140) );
  NOR U41081 ( .A(n28140), .B(n28139), .Z(n31285) );
  NOR U41082 ( .A(n28141), .B(n31285), .Z(n28142) );
  IV U41083 ( .A(n28142), .Z(n31227) );
  IV U41084 ( .A(n28143), .Z(n28145) );
  NOR U41085 ( .A(n28145), .B(n28144), .Z(n34339) );
  IV U41086 ( .A(n28146), .Z(n28147) );
  NOR U41087 ( .A(n28150), .B(n28147), .Z(n34336) );
  IV U41088 ( .A(n28148), .Z(n28149) );
  NOR U41089 ( .A(n28150), .B(n28149), .Z(n31292) );
  IV U41090 ( .A(n28151), .Z(n28152) );
  NOR U41091 ( .A(n31298), .B(n28152), .Z(n28155) );
  NOR U41092 ( .A(n28153), .B(n34332), .Z(n28154) );
  NOR U41093 ( .A(n28155), .B(n28154), .Z(n31226) );
  IV U41094 ( .A(n28156), .Z(n31220) );
  IV U41095 ( .A(n28157), .Z(n28158) );
  NOR U41096 ( .A(n31220), .B(n28158), .Z(n34325) );
  IV U41097 ( .A(n28159), .Z(n28160) );
  NOR U41098 ( .A(n28160), .B(n28162), .Z(n31306) );
  IV U41099 ( .A(n28161), .Z(n28163) );
  NOR U41100 ( .A(n28163), .B(n28162), .Z(n34328) );
  NOR U41101 ( .A(n31306), .B(n34328), .Z(n28164) );
  IV U41102 ( .A(n28164), .Z(n28165) );
  NOR U41103 ( .A(n34325), .B(n28165), .Z(n31225) );
  NOR U41104 ( .A(n28171), .B(n28166), .Z(n28169) );
  IV U41105 ( .A(n28167), .Z(n28168) );
  NOR U41106 ( .A(n28169), .B(n28168), .Z(n34318) );
  NOR U41107 ( .A(n28170), .B(n31318), .Z(n28174) );
  IV U41108 ( .A(n28171), .Z(n28173) );
  NOR U41109 ( .A(n28173), .B(n28172), .Z(n31311) );
  NOR U41110 ( .A(n28174), .B(n31311), .Z(n28175) );
  IV U41111 ( .A(n28175), .Z(n31217) );
  IV U41112 ( .A(n28176), .Z(n28177) );
  NOR U41113 ( .A(n28177), .B(n31197), .Z(n31209) );
  IV U41114 ( .A(n28178), .Z(n28180) );
  NOR U41115 ( .A(n28180), .B(n28179), .Z(n31206) );
  IV U41116 ( .A(n31206), .Z(n31195) );
  NOR U41117 ( .A(n28181), .B(n34282), .Z(n31173) );
  IV U41118 ( .A(n31173), .Z(n31169) );
  IV U41119 ( .A(n28182), .Z(n28183) );
  NOR U41120 ( .A(n28183), .B(n28185), .Z(n34261) );
  IV U41121 ( .A(n28184), .Z(n28186) );
  NOR U41122 ( .A(n28186), .B(n28185), .Z(n31163) );
  IV U41123 ( .A(n28187), .Z(n28189) );
  NOR U41124 ( .A(n28189), .B(n28188), .Z(n34253) );
  IV U41125 ( .A(n28190), .Z(n28191) );
  NOR U41126 ( .A(n28191), .B(n28193), .Z(n37782) );
  IV U41127 ( .A(n28192), .Z(n28194) );
  NOR U41128 ( .A(n28194), .B(n28193), .Z(n34511) );
  NOR U41129 ( .A(n37782), .B(n34511), .Z(n31350) );
  IV U41130 ( .A(n28195), .Z(n31353) );
  NOR U41131 ( .A(n31353), .B(n28196), .Z(n28200) );
  IV U41132 ( .A(n28197), .Z(n28199) );
  NOR U41133 ( .A(n28199), .B(n28198), .Z(n31357) );
  NOR U41134 ( .A(n28200), .B(n31357), .Z(n31154) );
  IV U41135 ( .A(n28201), .Z(n28202) );
  NOR U41136 ( .A(n28202), .B(n28204), .Z(n37994) );
  IV U41137 ( .A(n28203), .Z(n28205) );
  NOR U41138 ( .A(n28205), .B(n28204), .Z(n40921) );
  NOR U41139 ( .A(n37994), .B(n40921), .Z(n31356) );
  IV U41140 ( .A(n28206), .Z(n28208) );
  IV U41141 ( .A(n28207), .Z(n28213) );
  NOR U41142 ( .A(n28208), .B(n28213), .Z(n31366) );
  IV U41143 ( .A(n28209), .Z(n28211) );
  XOR U41144 ( .A(n28212), .B(n28213), .Z(n28210) );
  NOR U41145 ( .A(n28211), .B(n28210), .Z(n31364) );
  NOR U41146 ( .A(n31366), .B(n31364), .Z(n31143) );
  IV U41147 ( .A(n28212), .Z(n28214) );
  NOR U41148 ( .A(n28214), .B(n28213), .Z(n31368) );
  IV U41149 ( .A(n28215), .Z(n28216) );
  NOR U41150 ( .A(n28216), .B(n28219), .Z(n28217) );
  IV U41151 ( .A(n28217), .Z(n31411) );
  IV U41152 ( .A(n28218), .Z(n28220) );
  NOR U41153 ( .A(n28220), .B(n28219), .Z(n31070) );
  IV U41154 ( .A(n31070), .Z(n31061) );
  NOR U41155 ( .A(n28221), .B(n31415), .Z(n31065) );
  IV U41156 ( .A(n28222), .Z(n28224) );
  IV U41157 ( .A(n28223), .Z(n31063) );
  NOR U41158 ( .A(n28224), .B(n31063), .Z(n34569) );
  NOR U41159 ( .A(n31065), .B(n34569), .Z(n28225) );
  IV U41160 ( .A(n28225), .Z(n31059) );
  IV U41161 ( .A(n28226), .Z(n28231) );
  IV U41162 ( .A(n28227), .Z(n28228) );
  NOR U41163 ( .A(n28231), .B(n28228), .Z(n31422) );
  IV U41164 ( .A(n28229), .Z(n28230) );
  NOR U41165 ( .A(n28231), .B(n28230), .Z(n31425) );
  IV U41166 ( .A(n28232), .Z(n28234) );
  NOR U41167 ( .A(n28234), .B(n28233), .Z(n31428) );
  NOR U41168 ( .A(n31425), .B(n31428), .Z(n31058) );
  IV U41169 ( .A(n28235), .Z(n28236) );
  NOR U41170 ( .A(n28236), .B(n28238), .Z(n31055) );
  IV U41171 ( .A(n28237), .Z(n28239) );
  NOR U41172 ( .A(n28239), .B(n28238), .Z(n31051) );
  IV U41173 ( .A(n31051), .Z(n31042) );
  IV U41174 ( .A(n28240), .Z(n28242) );
  IV U41175 ( .A(n28241), .Z(n31044) );
  NOR U41176 ( .A(n28242), .B(n31044), .Z(n31039) );
  IV U41177 ( .A(n31039), .Z(n31030) );
  IV U41178 ( .A(n28243), .Z(n31026) );
  IV U41179 ( .A(n28246), .Z(n28244) );
  NOR U41180 ( .A(n28245), .B(n28244), .Z(n31020) );
  IV U41181 ( .A(n28245), .Z(n31436) );
  NOR U41182 ( .A(n28246), .B(n31436), .Z(n31022) );
  IV U41183 ( .A(n28247), .Z(n28248) );
  NOR U41184 ( .A(n28248), .B(n28252), .Z(n31023) );
  IV U41185 ( .A(n31023), .Z(n31442) );
  IV U41186 ( .A(n28249), .Z(n31446) );
  NOR U41187 ( .A(n28250), .B(n31446), .Z(n31435) );
  IV U41188 ( .A(n28251), .Z(n28253) );
  NOR U41189 ( .A(n28253), .B(n28252), .Z(n31443) );
  NOR U41190 ( .A(n31435), .B(n31443), .Z(n31016) );
  IV U41191 ( .A(n31009), .Z(n31002) );
  IV U41192 ( .A(n28254), .Z(n30990) );
  IV U41193 ( .A(n28255), .Z(n28256) );
  NOR U41194 ( .A(n30990), .B(n28256), .Z(n30999) );
  IV U41195 ( .A(n30999), .Z(n30987) );
  IV U41196 ( .A(n28257), .Z(n28259) );
  NOR U41197 ( .A(n28259), .B(n28258), .Z(n31460) );
  IV U41198 ( .A(n28260), .Z(n28261) );
  NOR U41199 ( .A(n28261), .B(n28265), .Z(n31462) );
  NOR U41200 ( .A(n31460), .B(n31462), .Z(n30986) );
  IV U41201 ( .A(n28262), .Z(n31469) );
  NOR U41202 ( .A(n31469), .B(n28263), .Z(n28267) );
  IV U41203 ( .A(n28264), .Z(n28266) );
  NOR U41204 ( .A(n28266), .B(n28265), .Z(n31465) );
  NOR U41205 ( .A(n28267), .B(n31465), .Z(n30985) );
  IV U41206 ( .A(n28268), .Z(n28270) );
  NOR U41207 ( .A(n28270), .B(n28269), .Z(n31475) );
  IV U41208 ( .A(n28271), .Z(n28274) );
  IV U41209 ( .A(n28272), .Z(n28273) );
  NOR U41210 ( .A(n28274), .B(n28273), .Z(n28275) );
  IV U41211 ( .A(n28275), .Z(n31484) );
  IV U41212 ( .A(n30964), .Z(n28276) );
  NOR U41213 ( .A(n28276), .B(n30963), .Z(n30958) );
  IV U41214 ( .A(n30958), .Z(n30950) );
  NOR U41215 ( .A(n28277), .B(n34670), .Z(n30948) );
  IV U41216 ( .A(n30948), .Z(n30944) );
  IV U41217 ( .A(n28278), .Z(n28279) );
  NOR U41218 ( .A(n30938), .B(n28279), .Z(n34157) );
  IV U41219 ( .A(n28280), .Z(n28283) );
  IV U41220 ( .A(n28281), .Z(n28282) );
  NOR U41221 ( .A(n28283), .B(n28282), .Z(n28284) );
  IV U41222 ( .A(n28284), .Z(n31498) );
  IV U41223 ( .A(n28285), .Z(n28286) );
  NOR U41224 ( .A(n28286), .B(n28289), .Z(n31503) );
  NOR U41225 ( .A(n31503), .B(n31500), .Z(n28287) );
  IV U41226 ( .A(n28287), .Z(n30935) );
  IV U41227 ( .A(n28288), .Z(n28290) );
  NOR U41228 ( .A(n28290), .B(n28289), .Z(n31505) );
  IV U41229 ( .A(n28291), .Z(n28292) );
  NOR U41230 ( .A(n30930), .B(n28292), .Z(n31509) );
  IV U41231 ( .A(n28293), .Z(n28295) );
  IV U41232 ( .A(n28294), .Z(n28298) );
  NOR U41233 ( .A(n28295), .B(n28298), .Z(n31511) );
  NOR U41234 ( .A(n31509), .B(n31511), .Z(n30933) );
  NOR U41235 ( .A(n31518), .B(n28296), .Z(n28300) );
  IV U41236 ( .A(n28297), .Z(n28299) );
  NOR U41237 ( .A(n28299), .B(n28298), .Z(n31514) );
  NOR U41238 ( .A(n28300), .B(n31514), .Z(n28301) );
  IV U41239 ( .A(n28301), .Z(n30927) );
  IV U41240 ( .A(n28302), .Z(n28303) );
  NOR U41241 ( .A(n28303), .B(n30907), .Z(n31532) );
  IV U41242 ( .A(n28304), .Z(n28309) );
  IV U41243 ( .A(n28305), .Z(n28306) );
  NOR U41244 ( .A(n28309), .B(n28306), .Z(n34135) );
  IV U41245 ( .A(n28307), .Z(n28308) );
  NOR U41246 ( .A(n28309), .B(n28308), .Z(n34132) );
  IV U41247 ( .A(n28310), .Z(n28312) );
  NOR U41248 ( .A(n28312), .B(n28311), .Z(n34128) );
  IV U41249 ( .A(n28313), .Z(n28314) );
  NOR U41250 ( .A(n28314), .B(n28316), .Z(n34125) );
  IV U41251 ( .A(n28315), .Z(n28317) );
  NOR U41252 ( .A(n28317), .B(n28316), .Z(n34118) );
  NOR U41253 ( .A(n31543), .B(n28318), .Z(n50782) );
  IV U41254 ( .A(n28319), .Z(n28321) );
  IV U41255 ( .A(n28320), .Z(n30894) );
  NOR U41256 ( .A(n28321), .B(n30894), .Z(n31535) );
  NOR U41257 ( .A(n50782), .B(n31535), .Z(n30891) );
  IV U41258 ( .A(n28322), .Z(n28327) );
  IV U41259 ( .A(n28323), .Z(n28324) );
  NOR U41260 ( .A(n28327), .B(n28324), .Z(n31555) );
  IV U41261 ( .A(n28325), .Z(n28326) );
  NOR U41262 ( .A(n28327), .B(n28326), .Z(n31552) );
  IV U41263 ( .A(n28328), .Z(n28329) );
  NOR U41264 ( .A(n28329), .B(n30865), .Z(n31560) );
  IV U41265 ( .A(n28330), .Z(n28332) );
  IV U41266 ( .A(n28331), .Z(n30860) );
  NOR U41267 ( .A(n28332), .B(n30860), .Z(n34101) );
  IV U41268 ( .A(n34101), .Z(n30867) );
  IV U41269 ( .A(n28333), .Z(n30853) );
  IV U41270 ( .A(n28334), .Z(n28335) );
  NOR U41271 ( .A(n30853), .B(n28335), .Z(n30855) );
  IV U41272 ( .A(n28336), .Z(n28337) );
  NOR U41273 ( .A(n28337), .B(n34774), .Z(n34767) );
  IV U41274 ( .A(n28338), .Z(n30826) );
  IV U41275 ( .A(n28339), .Z(n28340) );
  NOR U41276 ( .A(n30826), .B(n28340), .Z(n34763) );
  NOR U41277 ( .A(n34767), .B(n34763), .Z(n34088) );
  IV U41278 ( .A(n28341), .Z(n30819) );
  IV U41279 ( .A(n28342), .Z(n28343) );
  NOR U41280 ( .A(n30819), .B(n28343), .Z(n37498) );
  IV U41281 ( .A(n28344), .Z(n28345) );
  NOR U41282 ( .A(n28345), .B(n34774), .Z(n28346) );
  NOR U41283 ( .A(n37498), .B(n28346), .Z(n31582) );
  IV U41284 ( .A(n28347), .Z(n28348) );
  NOR U41285 ( .A(n28351), .B(n28348), .Z(n34072) );
  IV U41286 ( .A(n28349), .Z(n28350) );
  NOR U41287 ( .A(n28351), .B(n28350), .Z(n34069) );
  IV U41288 ( .A(n28352), .Z(n28354) );
  IV U41289 ( .A(n28353), .Z(n30807) );
  NOR U41290 ( .A(n28354), .B(n30807), .Z(n31584) );
  NOR U41291 ( .A(n34069), .B(n31584), .Z(n28355) );
  IV U41292 ( .A(n28355), .Z(n30810) );
  IV U41293 ( .A(n28356), .Z(n28358) );
  NOR U41294 ( .A(n28358), .B(n28357), .Z(n30797) );
  IV U41295 ( .A(n28359), .Z(n28360) );
  NOR U41296 ( .A(n28360), .B(n28362), .Z(n31597) );
  IV U41297 ( .A(n28361), .Z(n28363) );
  NOR U41298 ( .A(n28363), .B(n28362), .Z(n30793) );
  IV U41299 ( .A(n30793), .Z(n30785) );
  IV U41300 ( .A(n28364), .Z(n28365) );
  NOR U41301 ( .A(n28365), .B(n30783), .Z(n31609) );
  IV U41302 ( .A(n28366), .Z(n28367) );
  NOR U41303 ( .A(n34048), .B(n28367), .Z(n28370) );
  IV U41304 ( .A(n34826), .Z(n28369) );
  IV U41305 ( .A(n28368), .Z(n30763) );
  NOR U41306 ( .A(n28369), .B(n30763), .Z(n37461) );
  NOR U41307 ( .A(n28370), .B(n37461), .Z(n34045) );
  IV U41308 ( .A(n28371), .Z(n28372) );
  NOR U41309 ( .A(n30770), .B(n28372), .Z(n31612) );
  IV U41310 ( .A(n28373), .Z(n28375) );
  IV U41311 ( .A(n28374), .Z(n28378) );
  NOR U41312 ( .A(n28375), .B(n28378), .Z(n34030) );
  NOR U41313 ( .A(n31612), .B(n34030), .Z(n30761) );
  NOR U41314 ( .A(n28376), .B(n31615), .Z(n28380) );
  IV U41315 ( .A(n28377), .Z(n28379) );
  NOR U41316 ( .A(n28379), .B(n28378), .Z(n34032) );
  NOR U41317 ( .A(n28380), .B(n34032), .Z(n30760) );
  IV U41318 ( .A(n28381), .Z(n31629) );
  NOR U41319 ( .A(n28382), .B(n31629), .Z(n31619) );
  IV U41320 ( .A(n28383), .Z(n28384) );
  NOR U41321 ( .A(n28384), .B(n30735), .Z(n31638) );
  IV U41322 ( .A(n31638), .Z(n41469) );
  IV U41323 ( .A(n28385), .Z(n28390) );
  IV U41324 ( .A(n28386), .Z(n28387) );
  NOR U41325 ( .A(n28390), .B(n28387), .Z(n31643) );
  IV U41326 ( .A(n28388), .Z(n28389) );
  NOR U41327 ( .A(n28390), .B(n28389), .Z(n31650) );
  IV U41328 ( .A(n28391), .Z(n28393) );
  NOR U41329 ( .A(n28393), .B(n28392), .Z(n30730) );
  IV U41330 ( .A(n30730), .Z(n30717) );
  IV U41331 ( .A(n28394), .Z(n28396) );
  NOR U41332 ( .A(n28396), .B(n28395), .Z(n31666) );
  IV U41333 ( .A(n28397), .Z(n34006) );
  NOR U41334 ( .A(n28398), .B(n34006), .Z(n30685) );
  IV U41335 ( .A(n30685), .Z(n30678) );
  IV U41336 ( .A(n28399), .Z(n28400) );
  NOR U41337 ( .A(n28400), .B(n37370), .Z(n30676) );
  IV U41338 ( .A(n30676), .Z(n30660) );
  IV U41339 ( .A(n28401), .Z(n30650) );
  NOR U41340 ( .A(n28402), .B(n30650), .Z(n30647) );
  IV U41341 ( .A(n28403), .Z(n28405) );
  IV U41342 ( .A(n28404), .Z(n30642) );
  NOR U41343 ( .A(n28405), .B(n30642), .Z(n31687) );
  XOR U41344 ( .A(n31693), .B(n31695), .Z(n28406) );
  NOR U41345 ( .A(n31687), .B(n28406), .Z(n28407) );
  IV U41346 ( .A(n28407), .Z(n30634) );
  IV U41347 ( .A(n28408), .Z(n28409) );
  NOR U41348 ( .A(n28409), .B(n28411), .Z(n33989) );
  IV U41349 ( .A(n28410), .Z(n28412) );
  NOR U41350 ( .A(n28412), .B(n28411), .Z(n33986) );
  IV U41351 ( .A(n28413), .Z(n28414) );
  NOR U41352 ( .A(n28414), .B(n30630), .Z(n31704) );
  XOR U41353 ( .A(n31703), .B(n31704), .Z(n28415) );
  NOR U41354 ( .A(n33986), .B(n28415), .Z(n30633) );
  IV U41355 ( .A(n28416), .Z(n28418) );
  IV U41356 ( .A(n28417), .Z(n30627) );
  NOR U41357 ( .A(n28418), .B(n30627), .Z(n31712) );
  IV U41358 ( .A(n28419), .Z(n28422) );
  IV U41359 ( .A(n28420), .Z(n28421) );
  NOR U41360 ( .A(n28422), .B(n28421), .Z(n33970) );
  IV U41361 ( .A(n28423), .Z(n28424) );
  NOR U41362 ( .A(n28424), .B(n30583), .Z(n30576) );
  IV U41363 ( .A(n30576), .Z(n30570) );
  IV U41364 ( .A(n28425), .Z(n28428) );
  IV U41365 ( .A(n28426), .Z(n28427) );
  NOR U41366 ( .A(n28428), .B(n28427), .Z(n33948) );
  IV U41367 ( .A(n28429), .Z(n28430) );
  NOR U41368 ( .A(n28430), .B(n28432), .Z(n30558) );
  IV U41369 ( .A(n28431), .Z(n28433) );
  NOR U41370 ( .A(n28433), .B(n28432), .Z(n30556) );
  IV U41371 ( .A(n30556), .Z(n30552) );
  IV U41372 ( .A(n28434), .Z(n28436) );
  NOR U41373 ( .A(n28436), .B(n28435), .Z(n31744) );
  IV U41374 ( .A(n28437), .Z(n34979) );
  NOR U41375 ( .A(n34979), .B(n28438), .Z(n33926) );
  IV U41376 ( .A(n28439), .Z(n28440) );
  NOR U41377 ( .A(n28440), .B(n28442), .Z(n37311) );
  IV U41378 ( .A(n28441), .Z(n28443) );
  NOR U41379 ( .A(n28443), .B(n28442), .Z(n37316) );
  NOR U41380 ( .A(n37311), .B(n37316), .Z(n31747) );
  IV U41381 ( .A(n28444), .Z(n28445) );
  NOR U41382 ( .A(n28445), .B(n28447), .Z(n31755) );
  IV U41383 ( .A(n28446), .Z(n28448) );
  NOR U41384 ( .A(n28448), .B(n28447), .Z(n31760) );
  IV U41385 ( .A(n28449), .Z(n28450) );
  NOR U41386 ( .A(n28450), .B(n28454), .Z(n33908) );
  IV U41387 ( .A(n28451), .Z(n33902) );
  NOR U41388 ( .A(n28452), .B(n33902), .Z(n28456) );
  IV U41389 ( .A(n28453), .Z(n28455) );
  NOR U41390 ( .A(n28455), .B(n28454), .Z(n31779) );
  NOR U41391 ( .A(n28456), .B(n31779), .Z(n30510) );
  IV U41392 ( .A(n28457), .Z(n28458) );
  NOR U41393 ( .A(n30491), .B(n28458), .Z(n30484) );
  IV U41394 ( .A(n30484), .Z(n30477) );
  IV U41395 ( .A(n28459), .Z(n28461) );
  XOR U41396 ( .A(n30473), .B(n30474), .Z(n28460) );
  NOR U41397 ( .A(n28461), .B(n28460), .Z(n33891) );
  IV U41398 ( .A(n28462), .Z(n28463) );
  NOR U41399 ( .A(n28463), .B(n30474), .Z(n31794) );
  IV U41400 ( .A(n28464), .Z(n28469) );
  IV U41401 ( .A(n28465), .Z(n28466) );
  NOR U41402 ( .A(n28469), .B(n28466), .Z(n31797) );
  IV U41403 ( .A(n28467), .Z(n28468) );
  NOR U41404 ( .A(n28469), .B(n28468), .Z(n31800) );
  IV U41405 ( .A(n28470), .Z(n28472) );
  NOR U41406 ( .A(n28472), .B(n28471), .Z(n31806) );
  XOR U41407 ( .A(n31800), .B(n31806), .Z(n28473) );
  NOR U41408 ( .A(n31797), .B(n28473), .Z(n28474) );
  IV U41409 ( .A(n28474), .Z(n30472) );
  XOR U41410 ( .A(n30465), .B(n30466), .Z(n28475) );
  NOR U41411 ( .A(n30468), .B(n28475), .Z(n28478) );
  IV U41412 ( .A(n28476), .Z(n28477) );
  NOR U41413 ( .A(n28478), .B(n28477), .Z(n31803) );
  NOR U41414 ( .A(n28479), .B(n30456), .Z(n30453) );
  IV U41415 ( .A(n28480), .Z(n28486) );
  IV U41416 ( .A(n28481), .Z(n28482) );
  NOR U41417 ( .A(n28486), .B(n28482), .Z(n28483) );
  IV U41418 ( .A(n28483), .Z(n31815) );
  IV U41419 ( .A(n28484), .Z(n28485) );
  NOR U41420 ( .A(n28486), .B(n28485), .Z(n31818) );
  IV U41421 ( .A(n28487), .Z(n28489) );
  NOR U41422 ( .A(n28489), .B(n28488), .Z(n31816) );
  NOR U41423 ( .A(n31818), .B(n31816), .Z(n28490) );
  IV U41424 ( .A(n28490), .Z(n30451) );
  IV U41425 ( .A(n28491), .Z(n28492) );
  NOR U41426 ( .A(n28492), .B(n28499), .Z(n33876) );
  IV U41427 ( .A(n28493), .Z(n28495) );
  XOR U41428 ( .A(n28498), .B(n28499), .Z(n28494) );
  NOR U41429 ( .A(n28495), .B(n28494), .Z(n31823) );
  NOR U41430 ( .A(n33876), .B(n31823), .Z(n30450) );
  IV U41431 ( .A(n28496), .Z(n31829) );
  NOR U41432 ( .A(n31829), .B(n28497), .Z(n28501) );
  IV U41433 ( .A(n28498), .Z(n28500) );
  NOR U41434 ( .A(n28500), .B(n28499), .Z(n33879) );
  NOR U41435 ( .A(n28501), .B(n33879), .Z(n30449) );
  IV U41436 ( .A(n28502), .Z(n28504) );
  NOR U41437 ( .A(n28504), .B(n28503), .Z(n31825) );
  NOR U41438 ( .A(n28505), .B(n35064), .Z(n31837) );
  NOR U41439 ( .A(n28506), .B(n31837), .Z(n28507) );
  NOR U41440 ( .A(n28507), .B(n31840), .Z(n30448) );
  IV U41441 ( .A(n28508), .Z(n28509) );
  NOR U41442 ( .A(n28516), .B(n28509), .Z(n37235) );
  IV U41443 ( .A(n28510), .Z(n28513) );
  IV U41444 ( .A(n28511), .Z(n28512) );
  NOR U41445 ( .A(n28513), .B(n28512), .Z(n35073) );
  NOR U41446 ( .A(n37235), .B(n35073), .Z(n31843) );
  IV U41447 ( .A(n31843), .Z(n28517) );
  IV U41448 ( .A(n28514), .Z(n28515) );
  NOR U41449 ( .A(n28516), .B(n28515), .Z(n31838) );
  NOR U41450 ( .A(n28517), .B(n31838), .Z(n30447) );
  IV U41451 ( .A(n28518), .Z(n30433) );
  IV U41452 ( .A(n28519), .Z(n28522) );
  IV U41453 ( .A(n28520), .Z(n30429) );
  XOR U41454 ( .A(n30427), .B(n30429), .Z(n28521) );
  NOR U41455 ( .A(n28522), .B(n28521), .Z(n33862) );
  IV U41456 ( .A(n28523), .Z(n28524) );
  NOR U41457 ( .A(n28524), .B(n30409), .Z(n30406) );
  IV U41458 ( .A(n30406), .Z(n30402) );
  IV U41459 ( .A(n28525), .Z(n28528) );
  IV U41460 ( .A(n28526), .Z(n28527) );
  NOR U41461 ( .A(n28528), .B(n28527), .Z(n31876) );
  IV U41462 ( .A(n28529), .Z(n28530) );
  NOR U41463 ( .A(n28530), .B(n28535), .Z(n28531) );
  IV U41464 ( .A(n28531), .Z(n31920) );
  IV U41465 ( .A(n28532), .Z(n31922) );
  NOR U41466 ( .A(n31922), .B(n28533), .Z(n31911) );
  IV U41467 ( .A(n28534), .Z(n28536) );
  NOR U41468 ( .A(n28536), .B(n28535), .Z(n33847) );
  NOR U41469 ( .A(n31911), .B(n33847), .Z(n30376) );
  IV U41470 ( .A(n28537), .Z(n30367) );
  IV U41471 ( .A(n30362), .Z(n28538) );
  NOR U41472 ( .A(n30367), .B(n28538), .Z(n30354) );
  IV U41473 ( .A(n30354), .Z(n30345) );
  IV U41474 ( .A(n28539), .Z(n30339) );
  IV U41475 ( .A(n28540), .Z(n28541) );
  NOR U41476 ( .A(n30339), .B(n28541), .Z(n31932) );
  IV U41477 ( .A(n28542), .Z(n28543) );
  NOR U41478 ( .A(n28543), .B(n28545), .Z(n31928) );
  IV U41479 ( .A(n28544), .Z(n28546) );
  NOR U41480 ( .A(n28546), .B(n28545), .Z(n31926) );
  NOR U41481 ( .A(n31928), .B(n31926), .Z(n28547) );
  IV U41482 ( .A(n28547), .Z(n28548) );
  NOR U41483 ( .A(n31932), .B(n28548), .Z(n30344) );
  IV U41484 ( .A(n28549), .Z(n28550) );
  NOR U41485 ( .A(n28550), .B(n28553), .Z(n28551) );
  IV U41486 ( .A(n28551), .Z(n33830) );
  NOR U41487 ( .A(n33826), .B(n33828), .Z(n28555) );
  IV U41488 ( .A(n28552), .Z(n28554) );
  NOR U41489 ( .A(n28554), .B(n28553), .Z(n33832) );
  NOR U41490 ( .A(n28555), .B(n33832), .Z(n28556) );
  IV U41491 ( .A(n28556), .Z(n30336) );
  IV U41492 ( .A(n28557), .Z(n28560) );
  IV U41493 ( .A(n28558), .Z(n28559) );
  NOR U41494 ( .A(n28560), .B(n28559), .Z(n33822) );
  IV U41495 ( .A(n28561), .Z(n28564) );
  IV U41496 ( .A(n28562), .Z(n28563) );
  NOR U41497 ( .A(n28564), .B(n28563), .Z(n33819) );
  IV U41498 ( .A(n30333), .Z(n30326) );
  IV U41499 ( .A(n28565), .Z(n28567) );
  NOR U41500 ( .A(n28567), .B(n28566), .Z(n33811) );
  IV U41501 ( .A(n28568), .Z(n28569) );
  NOR U41502 ( .A(n28572), .B(n28569), .Z(n35191) );
  IV U41503 ( .A(n28570), .Z(n28571) );
  NOR U41504 ( .A(n28572), .B(n28571), .Z(n35184) );
  NOR U41505 ( .A(n35191), .B(n35184), .Z(n33802) );
  IV U41506 ( .A(n28573), .Z(n30302) );
  IV U41507 ( .A(n28574), .Z(n28575) );
  NOR U41508 ( .A(n30302), .B(n28575), .Z(n30308) );
  IV U41509 ( .A(n28576), .Z(n28579) );
  IV U41510 ( .A(n28577), .Z(n28578) );
  NOR U41511 ( .A(n28579), .B(n28578), .Z(n28580) );
  IV U41512 ( .A(n28580), .Z(n33796) );
  IV U41513 ( .A(n28581), .Z(n28582) );
  NOR U41514 ( .A(n28582), .B(n30286), .Z(n31975) );
  IV U41515 ( .A(n30287), .Z(n28583) );
  NOR U41516 ( .A(n28583), .B(n30286), .Z(n28584) );
  IV U41517 ( .A(n28584), .Z(n31974) );
  IV U41518 ( .A(n28585), .Z(n28587) );
  NOR U41519 ( .A(n28587), .B(n28586), .Z(n31983) );
  IV U41520 ( .A(n28588), .Z(n28589) );
  NOR U41521 ( .A(n28589), .B(n30270), .Z(n30267) );
  IV U41522 ( .A(n30267), .Z(n30263) );
  IV U41523 ( .A(n28590), .Z(n31995) );
  NOR U41524 ( .A(n28591), .B(n31995), .Z(n31988) );
  NOR U41525 ( .A(n28592), .B(n32000), .Z(n30261) );
  IV U41526 ( .A(n28593), .Z(n30256) );
  IV U41527 ( .A(n28594), .Z(n28595) );
  NOR U41528 ( .A(n30256), .B(n28595), .Z(n33781) );
  IV U41529 ( .A(n28596), .Z(n28599) );
  IV U41530 ( .A(n28597), .Z(n28598) );
  NOR U41531 ( .A(n28599), .B(n28598), .Z(n35253) );
  IV U41532 ( .A(n28600), .Z(n28601) );
  NOR U41533 ( .A(n28601), .B(n28603), .Z(n35248) );
  IV U41534 ( .A(n28602), .Z(n28604) );
  NOR U41535 ( .A(n28604), .B(n28603), .Z(n35243) );
  NOR U41536 ( .A(n35248), .B(n35243), .Z(n28605) );
  IV U41537 ( .A(n28605), .Z(n28606) );
  NOR U41538 ( .A(n35253), .B(n28606), .Z(n32007) );
  IV U41539 ( .A(n28607), .Z(n28608) );
  NOR U41540 ( .A(n28611), .B(n28608), .Z(n33777) );
  IV U41541 ( .A(n28609), .Z(n28610) );
  NOR U41542 ( .A(n28611), .B(n28610), .Z(n33774) );
  IV U41543 ( .A(n28612), .Z(n32021) );
  NOR U41544 ( .A(n28613), .B(n32021), .Z(n28616) );
  IV U41545 ( .A(n28614), .Z(n28615) );
  NOR U41546 ( .A(n28615), .B(n30249), .Z(n32017) );
  NOR U41547 ( .A(n28616), .B(n32017), .Z(n30253) );
  IV U41548 ( .A(n28617), .Z(n28618) );
  NOR U41549 ( .A(n28621), .B(n28618), .Z(n32027) );
  IV U41550 ( .A(n28619), .Z(n28620) );
  NOR U41551 ( .A(n28621), .B(n28620), .Z(n32024) );
  IV U41552 ( .A(n28622), .Z(n33750) );
  NOR U41553 ( .A(n33750), .B(n28623), .Z(n33760) );
  IV U41554 ( .A(n28624), .Z(n28626) );
  NOR U41555 ( .A(n28626), .B(n28625), .Z(n32030) );
  IV U41556 ( .A(n28627), .Z(n28628) );
  NOR U41557 ( .A(n28628), .B(n28630), .Z(n33744) );
  IV U41558 ( .A(n28629), .Z(n28631) );
  NOR U41559 ( .A(n28631), .B(n28630), .Z(n35279) );
  IV U41560 ( .A(n28632), .Z(n30221) );
  IV U41561 ( .A(n28633), .Z(n28634) );
  NOR U41562 ( .A(n30221), .B(n28634), .Z(n37038) );
  NOR U41563 ( .A(n35279), .B(n37038), .Z(n32034) );
  IV U41564 ( .A(n28635), .Z(n28637) );
  NOR U41565 ( .A(n28637), .B(n28636), .Z(n32035) );
  IV U41566 ( .A(n28638), .Z(n28639) );
  NOR U41567 ( .A(n28642), .B(n28639), .Z(n32043) );
  IV U41568 ( .A(n28640), .Z(n28641) );
  NOR U41569 ( .A(n28642), .B(n28641), .Z(n32041) );
  NOR U41570 ( .A(n32043), .B(n32041), .Z(n28643) );
  IV U41571 ( .A(n28643), .Z(n30218) );
  IV U41572 ( .A(n28644), .Z(n28646) );
  NOR U41573 ( .A(n28646), .B(n28645), .Z(n32046) );
  IV U41574 ( .A(n28647), .Z(n28648) );
  NOR U41575 ( .A(n28654), .B(n28648), .Z(n38588) );
  IV U41576 ( .A(n28649), .Z(n28651) );
  IV U41577 ( .A(n28650), .Z(n28658) );
  NOR U41578 ( .A(n28651), .B(n28658), .Z(n38598) );
  NOR U41579 ( .A(n38588), .B(n38598), .Z(n33741) );
  IV U41580 ( .A(n33741), .Z(n28655) );
  IV U41581 ( .A(n28652), .Z(n28653) );
  NOR U41582 ( .A(n28654), .B(n28653), .Z(n32050) );
  NOR U41583 ( .A(n28655), .B(n32050), .Z(n30217) );
  NOR U41584 ( .A(n28656), .B(n33725), .Z(n28660) );
  IV U41585 ( .A(n28657), .Z(n28659) );
  NOR U41586 ( .A(n28659), .B(n28658), .Z(n33734) );
  NOR U41587 ( .A(n28660), .B(n33734), .Z(n30216) );
  IV U41588 ( .A(n28661), .Z(n28664) );
  IV U41589 ( .A(n28662), .Z(n28663) );
  NOR U41590 ( .A(n28664), .B(n28663), .Z(n32053) );
  IV U41591 ( .A(n28665), .Z(n28667) );
  IV U41592 ( .A(n28666), .Z(n30186) );
  NOR U41593 ( .A(n28667), .B(n30186), .Z(n30180) );
  IV U41594 ( .A(n28668), .Z(n28669) );
  NOR U41595 ( .A(n28669), .B(n28671), .Z(n33695) );
  IV U41596 ( .A(n28670), .Z(n28672) );
  NOR U41597 ( .A(n28672), .B(n28671), .Z(n30177) );
  IV U41598 ( .A(n30177), .Z(n30171) );
  IV U41599 ( .A(n28673), .Z(n28674) );
  NOR U41600 ( .A(n28674), .B(n28676), .Z(n30174) );
  IV U41601 ( .A(n30174), .Z(n32079) );
  IV U41602 ( .A(n28675), .Z(n28677) );
  NOR U41603 ( .A(n28677), .B(n28676), .Z(n32077) );
  IV U41604 ( .A(n28678), .Z(n28680) );
  IV U41605 ( .A(n28679), .Z(n28682) );
  NOR U41606 ( .A(n28680), .B(n28682), .Z(n32082) );
  IV U41607 ( .A(n28681), .Z(n28683) );
  NOR U41608 ( .A(n28683), .B(n28682), .Z(n32080) );
  XOR U41609 ( .A(n32082), .B(n32080), .Z(n28684) );
  NOR U41610 ( .A(n32077), .B(n28684), .Z(n30169) );
  NOR U41611 ( .A(n28686), .B(n28685), .Z(n28687) );
  IV U41612 ( .A(n28687), .Z(n30148) );
  IV U41613 ( .A(n28688), .Z(n28689) );
  NOR U41614 ( .A(n28692), .B(n28689), .Z(n33658) );
  IV U41615 ( .A(n28690), .Z(n28691) );
  NOR U41616 ( .A(n28692), .B(n28691), .Z(n33655) );
  IV U41617 ( .A(n28693), .Z(n28695) );
  NOR U41618 ( .A(n28695), .B(n28694), .Z(n33651) );
  IV U41619 ( .A(n28696), .Z(n28698) );
  NOR U41620 ( .A(n28698), .B(n28697), .Z(n28699) );
  IV U41621 ( .A(n28699), .Z(n33636) );
  NOR U41622 ( .A(n32088), .B(n28700), .Z(n28705) );
  IV U41623 ( .A(n28701), .Z(n28704) );
  IV U41624 ( .A(n28702), .Z(n28703) );
  NOR U41625 ( .A(n28704), .B(n28703), .Z(n32091) );
  NOR U41626 ( .A(n28705), .B(n32091), .Z(n28706) );
  IV U41627 ( .A(n28706), .Z(n30134) );
  IV U41628 ( .A(n28707), .Z(n28710) );
  IV U41629 ( .A(n28708), .Z(n28709) );
  NOR U41630 ( .A(n28710), .B(n28709), .Z(n32097) );
  IV U41631 ( .A(n28711), .Z(n28712) );
  NOR U41632 ( .A(n28712), .B(n28714), .Z(n32103) );
  IV U41633 ( .A(n28713), .Z(n28715) );
  NOR U41634 ( .A(n28715), .B(n28714), .Z(n32101) );
  NOR U41635 ( .A(n32103), .B(n32101), .Z(n30132) );
  IV U41636 ( .A(n28716), .Z(n28717) );
  IV U41637 ( .A(n32107), .Z(n28721) );
  NOR U41638 ( .A(n28717), .B(n28721), .Z(n33616) );
  NOR U41639 ( .A(n28718), .B(n33626), .Z(n28719) );
  NOR U41640 ( .A(n33616), .B(n28719), .Z(n30131) );
  IV U41641 ( .A(n28720), .Z(n32108) );
  NOR U41642 ( .A(n32108), .B(n28721), .Z(n30127) );
  IV U41643 ( .A(n28722), .Z(n28724) );
  XOR U41644 ( .A(n28727), .B(n28728), .Z(n28723) );
  NOR U41645 ( .A(n28724), .B(n28723), .Z(n33609) );
  IV U41646 ( .A(n28725), .Z(n28726) );
  NOR U41647 ( .A(n28726), .B(n28728), .Z(n32120) );
  IV U41648 ( .A(n28727), .Z(n28729) );
  NOR U41649 ( .A(n28729), .B(n28728), .Z(n32117) );
  IV U41650 ( .A(n28730), .Z(n30117) );
  IV U41651 ( .A(n28731), .Z(n28732) );
  NOR U41652 ( .A(n30117), .B(n28732), .Z(n30113) );
  IV U41653 ( .A(n30113), .Z(n30100) );
  IV U41654 ( .A(n28733), .Z(n28735) );
  IV U41655 ( .A(n28734), .Z(n28737) );
  NOR U41656 ( .A(n28735), .B(n28737), .Z(n30097) );
  IV U41657 ( .A(n28736), .Z(n28738) );
  NOR U41658 ( .A(n28738), .B(n28737), .Z(n32126) );
  NOR U41659 ( .A(n28739), .B(n32126), .Z(n30096) );
  IV U41660 ( .A(n28740), .Z(n28741) );
  NOR U41661 ( .A(n28741), .B(n30093), .Z(n33586) );
  IV U41662 ( .A(n28742), .Z(n32145) );
  NOR U41663 ( .A(n32145), .B(n28743), .Z(n33591) );
  IV U41664 ( .A(n28744), .Z(n28745) );
  NOR U41665 ( .A(n28745), .B(n30090), .Z(n32137) );
  NOR U41666 ( .A(n33591), .B(n32137), .Z(n30088) );
  IV U41667 ( .A(n28746), .Z(n28747) );
  NOR U41668 ( .A(n28747), .B(n28750), .Z(n28748) );
  IV U41669 ( .A(n28748), .Z(n33582) );
  IV U41670 ( .A(n28749), .Z(n28751) );
  NOR U41671 ( .A(n28751), .B(n28750), .Z(n33579) );
  IV U41672 ( .A(n28752), .Z(n28757) );
  IV U41673 ( .A(n28753), .Z(n28754) );
  NOR U41674 ( .A(n28757), .B(n28754), .Z(n33567) );
  IV U41675 ( .A(n28755), .Z(n28756) );
  NOR U41676 ( .A(n28757), .B(n28756), .Z(n33568) );
  XOR U41677 ( .A(n33567), .B(n33568), .Z(n28758) );
  NOR U41678 ( .A(n33579), .B(n28758), .Z(n30087) );
  IV U41679 ( .A(n28759), .Z(n28761) );
  NOR U41680 ( .A(n28761), .B(n28760), .Z(n33571) );
  IV U41681 ( .A(n28762), .Z(n28763) );
  NOR U41682 ( .A(n28763), .B(n28765), .Z(n32153) );
  IV U41683 ( .A(n28764), .Z(n28766) );
  NOR U41684 ( .A(n28766), .B(n28765), .Z(n32155) );
  IV U41685 ( .A(n28767), .Z(n28770) );
  IV U41686 ( .A(n28768), .Z(n28769) );
  NOR U41687 ( .A(n28770), .B(n28769), .Z(n32157) );
  NOR U41688 ( .A(n32155), .B(n32157), .Z(n28771) );
  IV U41689 ( .A(n28771), .Z(n28772) );
  NOR U41690 ( .A(n32153), .B(n28772), .Z(n30085) );
  NOR U41691 ( .A(n28773), .B(n30072), .Z(n30069) );
  IV U41692 ( .A(n28774), .Z(n32168) );
  NOR U41693 ( .A(n28775), .B(n32168), .Z(n30067) );
  IV U41694 ( .A(n28776), .Z(n28777) );
  NOR U41695 ( .A(n28777), .B(n30065), .Z(n30061) );
  IV U41696 ( .A(n30061), .Z(n30051) );
  IV U41697 ( .A(n28778), .Z(n28779) );
  NOR U41698 ( .A(n28782), .B(n28779), .Z(n32192) );
  IV U41699 ( .A(n28780), .Z(n28781) );
  NOR U41700 ( .A(n28782), .B(n28781), .Z(n32187) );
  NOR U41701 ( .A(n32192), .B(n32187), .Z(n28783) );
  IV U41702 ( .A(n28783), .Z(n30036) );
  IV U41703 ( .A(n28784), .Z(n28786) );
  NOR U41704 ( .A(n28786), .B(n28785), .Z(n32189) );
  IV U41705 ( .A(n28787), .Z(n32203) );
  NOR U41706 ( .A(n32203), .B(n28788), .Z(n30021) );
  IV U41707 ( .A(n28789), .Z(n28791) );
  NOR U41708 ( .A(n28791), .B(n28790), .Z(n33524) );
  IV U41709 ( .A(n28792), .Z(n28795) );
  IV U41710 ( .A(n28793), .Z(n28794) );
  NOR U41711 ( .A(n28795), .B(n28794), .Z(n32210) );
  IV U41712 ( .A(n28796), .Z(n28798) );
  XOR U41713 ( .A(n29990), .B(n29991), .Z(n28797) );
  NOR U41714 ( .A(n28798), .B(n28797), .Z(n32217) );
  IV U41715 ( .A(n28799), .Z(n28806) );
  IV U41716 ( .A(n28800), .Z(n28801) );
  NOR U41717 ( .A(n28806), .B(n28801), .Z(n33491) );
  IV U41718 ( .A(n28802), .Z(n28803) );
  NOR U41719 ( .A(n28803), .B(n29979), .Z(n32237) );
  NOR U41720 ( .A(n33491), .B(n32237), .Z(n29976) );
  IV U41721 ( .A(n28804), .Z(n28805) );
  NOR U41722 ( .A(n28806), .B(n28805), .Z(n33480) );
  IV U41723 ( .A(n28807), .Z(n28809) );
  NOR U41724 ( .A(n28809), .B(n28808), .Z(n32239) );
  IV U41725 ( .A(n28810), .Z(n28812) );
  IV U41726 ( .A(n28811), .Z(n29954) );
  NOR U41727 ( .A(n28812), .B(n29954), .Z(n29965) );
  IV U41728 ( .A(n28813), .Z(n32254) );
  NOR U41729 ( .A(n32254), .B(n28814), .Z(n29960) );
  IV U41730 ( .A(n28815), .Z(n28817) );
  NOR U41731 ( .A(n28817), .B(n28816), .Z(n28818) );
  IV U41732 ( .A(n28818), .Z(n32270) );
  IV U41733 ( .A(n28819), .Z(n28820) );
  NOR U41734 ( .A(n28820), .B(n28822), .Z(n32272) );
  IV U41735 ( .A(n28821), .Z(n28823) );
  NOR U41736 ( .A(n28823), .B(n28822), .Z(n32274) );
  IV U41737 ( .A(n28824), .Z(n32278) );
  NOR U41738 ( .A(n32278), .B(n28825), .Z(n28826) );
  NOR U41739 ( .A(n32274), .B(n28826), .Z(n28827) );
  IV U41740 ( .A(n28827), .Z(n28828) );
  NOR U41741 ( .A(n32272), .B(n28828), .Z(n28829) );
  IV U41742 ( .A(n28829), .Z(n29944) );
  IV U41743 ( .A(n28830), .Z(n28832) );
  NOR U41744 ( .A(n28832), .B(n28831), .Z(n33462) );
  IV U41745 ( .A(n28833), .Z(n28834) );
  NOR U41746 ( .A(n28834), .B(n29942), .Z(n33465) );
  IV U41747 ( .A(n28835), .Z(n28837) );
  IV U41748 ( .A(n28836), .Z(n28839) );
  NOR U41749 ( .A(n28837), .B(n28839), .Z(n32284) );
  IV U41750 ( .A(n28838), .Z(n28840) );
  NOR U41751 ( .A(n28840), .B(n28839), .Z(n32281) );
  XOR U41752 ( .A(n32284), .B(n32281), .Z(n28841) );
  NOR U41753 ( .A(n33465), .B(n28841), .Z(n28842) );
  IV U41754 ( .A(n28842), .Z(n29940) );
  IV U41755 ( .A(n28843), .Z(n36789) );
  NOR U41756 ( .A(n28844), .B(n36789), .Z(n28845) );
  IV U41757 ( .A(n28845), .Z(n29931) );
  IV U41758 ( .A(n28846), .Z(n28848) );
  NOR U41759 ( .A(n28848), .B(n28847), .Z(n28849) );
  IV U41760 ( .A(n28849), .Z(n32300) );
  IV U41761 ( .A(n28850), .Z(n28851) );
  NOR U41762 ( .A(n28851), .B(n28853), .Z(n32305) );
  IV U41763 ( .A(n28852), .Z(n28854) );
  NOR U41764 ( .A(n28854), .B(n28853), .Z(n32303) );
  NOR U41765 ( .A(n32305), .B(n32303), .Z(n28855) );
  IV U41766 ( .A(n28855), .Z(n28857) );
  NOR U41767 ( .A(n28856), .B(n36747), .Z(n33421) );
  NOR U41768 ( .A(n28857), .B(n33421), .Z(n29903) );
  IV U41769 ( .A(n28858), .Z(n29894) );
  IV U41770 ( .A(n28859), .Z(n28860) );
  NOR U41771 ( .A(n29894), .B(n28860), .Z(n29900) );
  IV U41772 ( .A(n28861), .Z(n28862) );
  NOR U41773 ( .A(n28862), .B(n28864), .Z(n33414) );
  IV U41774 ( .A(n28863), .Z(n28865) );
  NOR U41775 ( .A(n28865), .B(n28864), .Z(n33407) );
  IV U41776 ( .A(n28866), .Z(n28867) );
  NOR U41777 ( .A(n33387), .B(n28867), .Z(n28870) );
  NOR U41778 ( .A(n28868), .B(n33396), .Z(n28869) );
  NOR U41779 ( .A(n28870), .B(n28869), .Z(n29869) );
  IV U41780 ( .A(n28871), .Z(n28872) );
  NOR U41781 ( .A(n28872), .B(n28874), .Z(n33382) );
  IV U41782 ( .A(n28873), .Z(n28875) );
  NOR U41783 ( .A(n28875), .B(n28874), .Z(n33380) );
  IV U41784 ( .A(n28876), .Z(n28879) );
  IV U41785 ( .A(n28877), .Z(n28878) );
  NOR U41786 ( .A(n28879), .B(n28878), .Z(n33373) );
  IV U41787 ( .A(n28880), .Z(n32328) );
  IV U41788 ( .A(n28881), .Z(n28882) );
  NOR U41789 ( .A(n28882), .B(n28885), .Z(n28883) );
  IV U41790 ( .A(n28883), .Z(n33371) );
  IV U41791 ( .A(n28884), .Z(n28886) );
  NOR U41792 ( .A(n28886), .B(n28885), .Z(n29866) );
  IV U41793 ( .A(n29866), .Z(n29855) );
  IV U41794 ( .A(n28887), .Z(n28889) );
  NOR U41795 ( .A(n28889), .B(n28888), .Z(n33360) );
  IV U41796 ( .A(n28890), .Z(n28892) );
  NOR U41797 ( .A(n28892), .B(n28891), .Z(n28893) );
  IV U41798 ( .A(n28893), .Z(n32338) );
  IV U41799 ( .A(n28894), .Z(n28895) );
  NOR U41800 ( .A(n28895), .B(n29843), .Z(n33345) );
  IV U41801 ( .A(n28896), .Z(n28901) );
  IV U41802 ( .A(n28897), .Z(n28898) );
  NOR U41803 ( .A(n28901), .B(n28898), .Z(n33337) );
  IV U41804 ( .A(n28899), .Z(n28900) );
  NOR U41805 ( .A(n28901), .B(n28900), .Z(n32343) );
  XOR U41806 ( .A(n33337), .B(n32343), .Z(n28902) );
  NOR U41807 ( .A(n33345), .B(n28902), .Z(n29840) );
  IV U41808 ( .A(n28903), .Z(n28905) );
  NOR U41809 ( .A(n28905), .B(n28904), .Z(n33334) );
  IV U41810 ( .A(n28906), .Z(n28907) );
  NOR U41811 ( .A(n28910), .B(n28907), .Z(n33330) );
  IV U41812 ( .A(n28908), .Z(n28909) );
  NOR U41813 ( .A(n28910), .B(n28909), .Z(n33327) );
  IV U41814 ( .A(n29807), .Z(n32365) );
  NOR U41815 ( .A(n29806), .B(n32365), .Z(n29810) );
  IV U41816 ( .A(n28911), .Z(n28912) );
  NOR U41817 ( .A(n28912), .B(n28917), .Z(n32371) );
  IV U41818 ( .A(n28913), .Z(n28914) );
  NOR U41819 ( .A(n28915), .B(n28914), .Z(n28919) );
  IV U41820 ( .A(n28916), .Z(n28918) );
  NOR U41821 ( .A(n28918), .B(n28917), .Z(n32374) );
  NOR U41822 ( .A(n28919), .B(n32374), .Z(n29801) );
  IV U41823 ( .A(n28920), .Z(n28921) );
  NOR U41824 ( .A(n29786), .B(n28921), .Z(n32381) );
  NOR U41825 ( .A(n32378), .B(n32394), .Z(n32383) );
  NOR U41826 ( .A(n32381), .B(n32383), .Z(n29800) );
  NOR U41827 ( .A(n33300), .B(n28922), .Z(n29793) );
  IV U41828 ( .A(n28923), .Z(n28926) );
  IV U41829 ( .A(n28924), .Z(n28925) );
  NOR U41830 ( .A(n28926), .B(n28925), .Z(n29777) );
  IV U41831 ( .A(n29777), .Z(n29764) );
  IV U41832 ( .A(n28927), .Z(n28928) );
  NOR U41833 ( .A(n28931), .B(n28928), .Z(n32403) );
  IV U41834 ( .A(n28929), .Z(n28930) );
  NOR U41835 ( .A(n28931), .B(n28930), .Z(n33294) );
  IV U41836 ( .A(n28932), .Z(n28934) );
  IV U41837 ( .A(n28933), .Z(n28938) );
  NOR U41838 ( .A(n28934), .B(n28938), .Z(n33292) );
  NOR U41839 ( .A(n33294), .B(n33292), .Z(n29763) );
  IV U41840 ( .A(n28935), .Z(n28936) );
  NOR U41841 ( .A(n29761), .B(n28936), .Z(n32412) );
  IV U41842 ( .A(n28937), .Z(n28939) );
  NOR U41843 ( .A(n28939), .B(n28938), .Z(n32406) );
  NOR U41844 ( .A(n32412), .B(n32406), .Z(n29762) );
  IV U41845 ( .A(n28940), .Z(n28942) );
  IV U41846 ( .A(n28941), .Z(n29740) );
  NOR U41847 ( .A(n28942), .B(n29740), .Z(n32425) );
  IV U41848 ( .A(n32425), .Z(n29729) );
  IV U41849 ( .A(n28943), .Z(n28945) );
  NOR U41850 ( .A(n28945), .B(n28944), .Z(n29727) );
  IV U41851 ( .A(n29727), .Z(n29722) );
  IV U41852 ( .A(n28946), .Z(n28948) );
  NOR U41853 ( .A(n28948), .B(n28947), .Z(n29720) );
  IV U41854 ( .A(n29720), .Z(n29707) );
  IV U41855 ( .A(n28949), .Z(n38946) );
  NOR U41856 ( .A(n28950), .B(n38946), .Z(n33247) );
  NOR U41857 ( .A(n28951), .B(n35758), .Z(n33249) );
  NOR U41858 ( .A(n33247), .B(n33249), .Z(n29706) );
  IV U41859 ( .A(n28952), .Z(n33240) );
  NOR U41860 ( .A(n33242), .B(n33240), .Z(n28955) );
  NOR U41861 ( .A(n28953), .B(n32433), .Z(n28954) );
  NOR U41862 ( .A(n28955), .B(n28954), .Z(n29705) );
  IV U41863 ( .A(n28956), .Z(n28957) );
  NOR U41864 ( .A(n28957), .B(n28959), .Z(n33235) );
  IV U41865 ( .A(n28958), .Z(n28960) );
  NOR U41866 ( .A(n28960), .B(n28959), .Z(n33233) );
  IV U41867 ( .A(n33223), .Z(n28961) );
  NOR U41868 ( .A(n28962), .B(n28961), .Z(n29689) );
  IV U41869 ( .A(n29689), .Z(n29684) );
  IV U41870 ( .A(n28963), .Z(n28966) );
  IV U41871 ( .A(n28964), .Z(n28965) );
  NOR U41872 ( .A(n28966), .B(n28965), .Z(n32448) );
  IV U41873 ( .A(n28967), .Z(n28968) );
  NOR U41874 ( .A(n29678), .B(n28968), .Z(n28969) );
  IV U41875 ( .A(n28969), .Z(n33220) );
  IV U41876 ( .A(n28970), .Z(n28973) );
  IV U41877 ( .A(n28971), .Z(n28972) );
  NOR U41878 ( .A(n28973), .B(n28972), .Z(n33206) );
  IV U41879 ( .A(n28974), .Z(n28975) );
  NOR U41880 ( .A(n28978), .B(n28975), .Z(n33196) );
  IV U41881 ( .A(n28976), .Z(n28977) );
  NOR U41882 ( .A(n28978), .B(n28977), .Z(n33186) );
  IV U41883 ( .A(n28979), .Z(n28982) );
  IV U41884 ( .A(n28980), .Z(n28981) );
  NOR U41885 ( .A(n28982), .B(n28981), .Z(n33187) );
  XOR U41886 ( .A(n33186), .B(n33187), .Z(n28983) );
  NOR U41887 ( .A(n33196), .B(n28983), .Z(n28984) );
  IV U41888 ( .A(n28984), .Z(n29666) );
  NOR U41889 ( .A(n28988), .B(n28985), .Z(n42375) );
  IV U41890 ( .A(n28986), .Z(n28987) );
  NOR U41891 ( .A(n28988), .B(n28987), .Z(n43048) );
  NOR U41892 ( .A(n42375), .B(n43048), .Z(n33190) );
  IV U41893 ( .A(n33190), .Z(n28996) );
  IV U41894 ( .A(n28989), .Z(n28991) );
  IV U41895 ( .A(n28990), .Z(n28993) );
  NOR U41896 ( .A(n28991), .B(n28993), .Z(n32463) );
  IV U41897 ( .A(n28992), .Z(n28994) );
  NOR U41898 ( .A(n28994), .B(n28993), .Z(n32462) );
  XOR U41899 ( .A(n32463), .B(n32462), .Z(n28995) );
  NOR U41900 ( .A(n28996), .B(n28995), .Z(n29665) );
  IV U41901 ( .A(n28997), .Z(n28998) );
  NOR U41902 ( .A(n28998), .B(n29000), .Z(n32466) );
  IV U41903 ( .A(n28999), .Z(n29001) );
  NOR U41904 ( .A(n29001), .B(n29000), .Z(n33182) );
  NOR U41905 ( .A(n32466), .B(n33182), .Z(n29002) );
  IV U41906 ( .A(n29002), .Z(n29006) );
  IV U41907 ( .A(n29003), .Z(n29004) );
  NOR U41908 ( .A(n29005), .B(n29004), .Z(n32471) );
  NOR U41909 ( .A(n29006), .B(n32471), .Z(n29664) );
  IV U41910 ( .A(n29007), .Z(n29009) );
  NOR U41911 ( .A(n29009), .B(n29008), .Z(n32468) );
  IV U41912 ( .A(n29010), .Z(n29011) );
  NOR U41913 ( .A(n29011), .B(n29013), .Z(n35813) );
  IV U41914 ( .A(n29012), .Z(n29014) );
  NOR U41915 ( .A(n29014), .B(n29013), .Z(n35809) );
  NOR U41916 ( .A(n35813), .B(n35809), .Z(n32474) );
  IV U41917 ( .A(n29015), .Z(n29016) );
  NOR U41918 ( .A(n29617), .B(n29016), .Z(n33143) );
  IV U41919 ( .A(n29017), .Z(n29020) );
  IV U41920 ( .A(n29018), .Z(n29019) );
  NOR U41921 ( .A(n29020), .B(n29019), .Z(n29605) );
  IV U41922 ( .A(n29021), .Z(n29022) );
  NOR U41923 ( .A(n29025), .B(n29022), .Z(n29023) );
  IV U41924 ( .A(n29023), .Z(n32511) );
  NOR U41925 ( .A(n29025), .B(n29024), .Z(n33129) );
  IV U41926 ( .A(n29026), .Z(n29028) );
  IV U41927 ( .A(n29027), .Z(n29586) );
  NOR U41928 ( .A(n29028), .B(n29586), .Z(n29604) );
  NOR U41929 ( .A(n33129), .B(n29604), .Z(n29602) );
  NOR U41930 ( .A(n29029), .B(n32518), .Z(n29581) );
  IV U41931 ( .A(n29030), .Z(n29031) );
  NOR U41932 ( .A(n33097), .B(n29031), .Z(n33095) );
  NOR U41933 ( .A(n29033), .B(n29032), .Z(n33111) );
  NOR U41934 ( .A(n33095), .B(n33111), .Z(n29547) );
  NOR U41935 ( .A(n29034), .B(n29519), .Z(n29517) );
  IV U41936 ( .A(n29035), .Z(n29041) );
  IV U41937 ( .A(n29036), .Z(n29037) );
  NOR U41938 ( .A(n29041), .B(n29037), .Z(n29038) );
  IV U41939 ( .A(n29038), .Z(n35901) );
  IV U41940 ( .A(n29039), .Z(n29040) );
  NOR U41941 ( .A(n29041), .B(n29040), .Z(n33090) );
  IV U41942 ( .A(n29042), .Z(n29044) );
  NOR U41943 ( .A(n29044), .B(n29043), .Z(n33087) );
  NOR U41944 ( .A(n33090), .B(n33087), .Z(n29045) );
  IV U41945 ( .A(n29045), .Z(n29516) );
  IV U41946 ( .A(n29046), .Z(n29047) );
  NOR U41947 ( .A(n29050), .B(n29047), .Z(n33079) );
  IV U41948 ( .A(n29048), .Z(n29049) );
  NOR U41949 ( .A(n29050), .B(n29049), .Z(n32575) );
  IV U41950 ( .A(n29051), .Z(n29053) );
  IV U41951 ( .A(n29052), .Z(n29056) );
  NOR U41952 ( .A(n29053), .B(n29056), .Z(n32580) );
  NOR U41953 ( .A(n32575), .B(n32580), .Z(n29054) );
  IV U41954 ( .A(n29054), .Z(n29496) );
  IV U41955 ( .A(n29055), .Z(n29057) );
  NOR U41956 ( .A(n29057), .B(n29056), .Z(n32577) );
  IV U41957 ( .A(n29058), .Z(n32594) );
  NOR U41958 ( .A(n29059), .B(n32594), .Z(n29062) );
  NOR U41959 ( .A(n29060), .B(n32587), .Z(n29061) );
  NOR U41960 ( .A(n29062), .B(n29061), .Z(n29495) );
  IV U41961 ( .A(n29063), .Z(n29065) );
  NOR U41962 ( .A(n29065), .B(n29064), .Z(n32605) );
  NOR U41963 ( .A(n29066), .B(n32602), .Z(n29067) );
  NOR U41964 ( .A(n32605), .B(n29067), .Z(n29494) );
  IV U41965 ( .A(n29068), .Z(n29493) );
  IV U41966 ( .A(n29069), .Z(n29070) );
  NOR U41967 ( .A(n29493), .B(n29070), .Z(n33065) );
  IV U41968 ( .A(n29071), .Z(n29072) );
  NOR U41969 ( .A(n29072), .B(n29074), .Z(n33040) );
  IV U41970 ( .A(n29073), .Z(n29075) );
  NOR U41971 ( .A(n29075), .B(n29074), .Z(n32611) );
  IV U41972 ( .A(n29076), .Z(n29078) );
  IV U41973 ( .A(n29077), .Z(n29080) );
  NOR U41974 ( .A(n29078), .B(n29080), .Z(n33027) );
  IV U41975 ( .A(n29079), .Z(n29081) );
  NOR U41976 ( .A(n29081), .B(n29080), .Z(n33024) );
  IV U41977 ( .A(n29082), .Z(n29083) );
  NOR U41978 ( .A(n29086), .B(n29083), .Z(n32635) );
  IV U41979 ( .A(n29084), .Z(n29085) );
  NOR U41980 ( .A(n29086), .B(n29085), .Z(n32632) );
  NOR U41981 ( .A(n33022), .B(n33019), .Z(n29090) );
  IV U41982 ( .A(n29087), .Z(n29089) );
  IV U41983 ( .A(n29088), .Z(n29443) );
  NOR U41984 ( .A(n29089), .B(n29443), .Z(n32639) );
  NOR U41985 ( .A(n29090), .B(n32639), .Z(n29447) );
  IV U41986 ( .A(n29091), .Z(n32643) );
  NOR U41987 ( .A(n29092), .B(n32643), .Z(n29441) );
  IV U41988 ( .A(n29093), .Z(n29095) );
  NOR U41989 ( .A(n29095), .B(n29094), .Z(n32654) );
  IV U41990 ( .A(n29096), .Z(n29097) );
  NOR U41991 ( .A(n29097), .B(n29432), .Z(n32658) );
  NOR U41992 ( .A(n32664), .B(n29098), .Z(n29101) );
  IV U41993 ( .A(n29099), .Z(n29100) );
  NOR U41994 ( .A(n29100), .B(n36013), .Z(n32661) );
  NOR U41995 ( .A(n29101), .B(n32661), .Z(n29102) );
  IV U41996 ( .A(n29102), .Z(n29430) );
  IV U41997 ( .A(n29103), .Z(n29106) );
  IV U41998 ( .A(n29104), .Z(n29105) );
  NOR U41999 ( .A(n29106), .B(n29105), .Z(n32997) );
  IV U42000 ( .A(n29107), .Z(n29110) );
  IV U42001 ( .A(n29108), .Z(n29109) );
  NOR U42002 ( .A(n29110), .B(n29109), .Z(n32994) );
  IV U42003 ( .A(n29111), .Z(n29114) );
  IV U42004 ( .A(n29112), .Z(n29113) );
  NOR U42005 ( .A(n29114), .B(n29113), .Z(n29427) );
  IV U42006 ( .A(n29427), .Z(n29425) );
  NOR U42007 ( .A(n29115), .B(n36037), .Z(n29118) );
  IV U42008 ( .A(n29411), .Z(n29117) );
  IV U42009 ( .A(n29116), .Z(n29416) );
  NOR U42010 ( .A(n29117), .B(n29416), .Z(n36337) );
  NOR U42011 ( .A(n29118), .B(n36337), .Z(n32681) );
  IV U42012 ( .A(n29119), .Z(n29401) );
  IV U42013 ( .A(n29120), .Z(n29121) );
  NOR U42014 ( .A(n29121), .B(n29398), .Z(n32983) );
  NOR U42015 ( .A(n29122), .B(n32694), .Z(n29126) );
  IV U42016 ( .A(n29123), .Z(n32689) );
  NOR U42017 ( .A(n29124), .B(n32689), .Z(n29125) );
  NOR U42018 ( .A(n29126), .B(n29125), .Z(n29395) );
  IV U42019 ( .A(n29127), .Z(n29392) );
  IV U42020 ( .A(n29128), .Z(n29129) );
  NOR U42021 ( .A(n29392), .B(n29129), .Z(n32700) );
  IV U42022 ( .A(n29130), .Z(n29132) );
  NOR U42023 ( .A(n29132), .B(n29131), .Z(n32975) );
  NOR U42024 ( .A(n32700), .B(n32975), .Z(n29394) );
  IV U42025 ( .A(n29133), .Z(n29134) );
  NOR U42026 ( .A(n29134), .B(n29136), .Z(n32710) );
  IV U42027 ( .A(n29135), .Z(n29137) );
  NOR U42028 ( .A(n29137), .B(n29136), .Z(n32708) );
  NOR U42029 ( .A(n32710), .B(n32708), .Z(n29362) );
  IV U42030 ( .A(n29138), .Z(n32715) );
  NOR U42031 ( .A(n29139), .B(n32715), .Z(n29358) );
  NOR U42032 ( .A(n29141), .B(n29140), .Z(n29355) );
  IV U42033 ( .A(n29355), .Z(n29345) );
  IV U42034 ( .A(n36075), .Z(n29143) );
  IV U42035 ( .A(n29142), .Z(n36074) );
  NOR U42036 ( .A(n29143), .B(n36074), .Z(n29339) );
  IV U42037 ( .A(n29144), .Z(n29147) );
  IV U42038 ( .A(n29145), .Z(n29146) );
  NOR U42039 ( .A(n29147), .B(n29146), .Z(n32960) );
  NOR U42040 ( .A(n29149), .B(n29148), .Z(n32721) );
  IV U42041 ( .A(n29150), .Z(n29155) );
  IV U42042 ( .A(n29151), .Z(n29152) );
  NOR U42043 ( .A(n29155), .B(n29152), .Z(n32726) );
  IV U42044 ( .A(n29153), .Z(n29154) );
  NOR U42045 ( .A(n29155), .B(n29154), .Z(n32727) );
  XOR U42046 ( .A(n32726), .B(n32727), .Z(n29156) );
  NOR U42047 ( .A(n32721), .B(n29156), .Z(n29335) );
  IV U42048 ( .A(n29157), .Z(n29159) );
  NOR U42049 ( .A(n29159), .B(n29158), .Z(n32955) );
  IV U42050 ( .A(n29160), .Z(n29163) );
  IV U42051 ( .A(n29161), .Z(n29323) );
  XOR U42052 ( .A(n29322), .B(n29323), .Z(n29162) );
  NOR U42053 ( .A(n29163), .B(n29162), .Z(n32952) );
  IV U42054 ( .A(n29164), .Z(n29165) );
  NOR U42055 ( .A(n29165), .B(n29323), .Z(n29332) );
  IV U42056 ( .A(n29332), .Z(n29321) );
  IV U42057 ( .A(n29166), .Z(n32741) );
  NOR U42058 ( .A(n29167), .B(n32741), .Z(n29328) );
  IV U42059 ( .A(n29168), .Z(n29169) );
  NOR U42060 ( .A(n29169), .B(n29173), .Z(n32747) );
  IV U42061 ( .A(n29170), .Z(n32753) );
  NOR U42062 ( .A(n29171), .B(n32753), .Z(n29175) );
  IV U42063 ( .A(n29172), .Z(n29174) );
  NOR U42064 ( .A(n29174), .B(n29173), .Z(n32750) );
  NOR U42065 ( .A(n29175), .B(n32750), .Z(n29318) );
  NOR U42066 ( .A(n29176), .B(n32763), .Z(n29180) );
  IV U42067 ( .A(n29177), .Z(n29179) );
  IV U42068 ( .A(n29178), .Z(n29183) );
  NOR U42069 ( .A(n29179), .B(n29183), .Z(n32944) );
  NOR U42070 ( .A(n29180), .B(n32944), .Z(n29317) );
  NOR U42071 ( .A(n29181), .B(n32767), .Z(n29185) );
  IV U42072 ( .A(n29182), .Z(n29184) );
  NOR U42073 ( .A(n29184), .B(n29183), .Z(n32942) );
  NOR U42074 ( .A(n29185), .B(n32942), .Z(n29316) );
  IV U42075 ( .A(n29186), .Z(n32922) );
  NOR U42076 ( .A(n32922), .B(n29187), .Z(n29315) );
  IV U42077 ( .A(n29188), .Z(n29190) );
  NOR U42078 ( .A(n29190), .B(n29189), .Z(n32770) );
  IV U42079 ( .A(n29191), .Z(n29192) );
  NOR U42080 ( .A(n29192), .B(n29200), .Z(n32914) );
  IV U42081 ( .A(n29193), .Z(n29194) );
  NOR U42082 ( .A(n29197), .B(n29194), .Z(n32906) );
  IV U42083 ( .A(n29195), .Z(n29196) );
  NOR U42084 ( .A(n29197), .B(n29196), .Z(n32909) );
  NOR U42085 ( .A(n32906), .B(n32909), .Z(n29198) );
  IV U42086 ( .A(n29198), .Z(n29202) );
  IV U42087 ( .A(n29199), .Z(n29201) );
  NOR U42088 ( .A(n29201), .B(n29200), .Z(n32773) );
  NOR U42089 ( .A(n29202), .B(n32773), .Z(n29203) );
  IV U42090 ( .A(n29203), .Z(n29314) );
  IV U42091 ( .A(n29204), .Z(n29206) );
  IV U42092 ( .A(n29205), .Z(n29208) );
  NOR U42093 ( .A(n29206), .B(n29208), .Z(n32904) );
  IV U42094 ( .A(n29207), .Z(n29209) );
  NOR U42095 ( .A(n29209), .B(n29208), .Z(n32893) );
  IV U42096 ( .A(n29210), .Z(n29211) );
  NOR U42097 ( .A(n29211), .B(n29213), .Z(n32776) );
  IV U42098 ( .A(n29212), .Z(n29214) );
  NOR U42099 ( .A(n29214), .B(n29213), .Z(n32896) );
  IV U42100 ( .A(n29215), .Z(n29216) );
  NOR U42101 ( .A(n29216), .B(n29304), .Z(n32882) );
  IV U42102 ( .A(n29217), .Z(n29302) );
  IV U42103 ( .A(n29218), .Z(n29219) );
  NOR U42104 ( .A(n29302), .B(n29219), .Z(n32875) );
  IV U42105 ( .A(n29220), .Z(n29221) );
  NOR U42106 ( .A(n29221), .B(n29223), .Z(n32872) );
  IV U42107 ( .A(n29222), .Z(n29224) );
  NOR U42108 ( .A(n29224), .B(n29223), .Z(n32788) );
  IV U42109 ( .A(n29225), .Z(n29230) );
  IV U42110 ( .A(n29226), .Z(n29227) );
  NOR U42111 ( .A(n29230), .B(n29227), .Z(n32866) );
  IV U42112 ( .A(n29228), .Z(n29229) );
  NOR U42113 ( .A(n29230), .B(n29229), .Z(n32790) );
  XOR U42114 ( .A(n32866), .B(n32790), .Z(n29231) );
  NOR U42115 ( .A(n32788), .B(n29231), .Z(n29232) );
  IV U42116 ( .A(n29232), .Z(n29299) );
  IV U42117 ( .A(n29233), .Z(n29235) );
  NOR U42118 ( .A(n29235), .B(n29234), .Z(n32863) );
  IV U42119 ( .A(n29236), .Z(n29238) );
  IV U42120 ( .A(n29237), .Z(n29240) );
  NOR U42121 ( .A(n29238), .B(n29240), .Z(n32849) );
  IV U42122 ( .A(n29239), .Z(n29241) );
  NOR U42123 ( .A(n29241), .B(n29240), .Z(n32841) );
  IV U42124 ( .A(n29242), .Z(n29243) );
  NOR U42125 ( .A(n29246), .B(n29243), .Z(n32838) );
  IV U42126 ( .A(n29244), .Z(n29245) );
  NOR U42127 ( .A(n29246), .B(n29245), .Z(n32796) );
  IV U42128 ( .A(n29247), .Z(n29249) );
  NOR U42129 ( .A(n29249), .B(n29248), .Z(n32793) );
  IV U42130 ( .A(n29250), .Z(n29251) );
  NOR U42131 ( .A(n29290), .B(n29251), .Z(n29252) );
  IV U42132 ( .A(n29252), .Z(n32812) );
  IV U42133 ( .A(n29253), .Z(n29256) );
  IV U42134 ( .A(n29254), .Z(n29255) );
  NOR U42135 ( .A(n29256), .B(n29255), .Z(n32813) );
  IV U42136 ( .A(n29271), .Z(n29258) );
  NOR U42137 ( .A(n29258), .B(n29257), .Z(n29272) );
  IV U42138 ( .A(n29272), .Z(n29262) );
  IV U42139 ( .A(n29259), .Z(n29260) );
  NOR U42140 ( .A(n29260), .B(n29284), .Z(n29276) );
  IV U42141 ( .A(n29276), .Z(n29261) );
  NOR U42142 ( .A(n29262), .B(n29261), .Z(n32810) );
  IV U42143 ( .A(n29263), .Z(n29265) );
  NOR U42144 ( .A(n29265), .B(n29264), .Z(n29268) );
  IV U42145 ( .A(n29285), .Z(n29266) );
  NOR U42146 ( .A(n29266), .B(n29284), .Z(n29267) );
  NOR U42147 ( .A(n29268), .B(n29267), .Z(n29269) );
  IV U42148 ( .A(n29269), .Z(n29280) );
  NOR U42149 ( .A(n29271), .B(n29270), .Z(n29275) );
  NOR U42150 ( .A(n29273), .B(n29272), .Z(n29274) );
  NOR U42151 ( .A(n29275), .B(n29274), .Z(n29277) );
  NOR U42152 ( .A(n29277), .B(n29276), .Z(n29278) );
  IV U42153 ( .A(n29278), .Z(n29279) );
  NOR U42154 ( .A(n29280), .B(n29279), .Z(n29281) );
  NOR U42155 ( .A(n32810), .B(n29281), .Z(n29282) );
  IV U42156 ( .A(n29282), .Z(n32808) );
  IV U42157 ( .A(n29283), .Z(n29287) );
  XOR U42158 ( .A(n29285), .B(n29284), .Z(n29286) );
  NOR U42159 ( .A(n29287), .B(n29286), .Z(n32806) );
  XOR U42160 ( .A(n32808), .B(n32806), .Z(n32814) );
  XOR U42161 ( .A(n32813), .B(n32814), .Z(n32811) );
  XOR U42162 ( .A(n32812), .B(n32811), .Z(n32800) );
  IV U42163 ( .A(n29288), .Z(n29289) );
  NOR U42164 ( .A(n29290), .B(n29289), .Z(n32803) );
  IV U42165 ( .A(n29291), .Z(n29292) );
  NOR U42166 ( .A(n29292), .B(n29295), .Z(n32799) );
  NOR U42167 ( .A(n32803), .B(n32799), .Z(n29293) );
  XOR U42168 ( .A(n32800), .B(n29293), .Z(n32824) );
  IV U42169 ( .A(n29294), .Z(n29296) );
  NOR U42170 ( .A(n29296), .B(n29295), .Z(n32822) );
  XOR U42171 ( .A(n32824), .B(n32822), .Z(n32795) );
  XOR U42172 ( .A(n32793), .B(n32795), .Z(n32798) );
  XOR U42173 ( .A(n32796), .B(n32798), .Z(n32840) );
  XOR U42174 ( .A(n32838), .B(n32840), .Z(n32842) );
  XOR U42175 ( .A(n32841), .B(n32842), .Z(n32851) );
  XOR U42176 ( .A(n32849), .B(n32851), .Z(n32857) );
  NOR U42177 ( .A(n32860), .B(n29297), .Z(n29298) );
  NOR U42178 ( .A(n32848), .B(n29298), .Z(n32856) );
  XOR U42179 ( .A(n32857), .B(n32856), .Z(n32864) );
  XOR U42180 ( .A(n32863), .B(n32864), .Z(n32867) );
  XOR U42181 ( .A(n29299), .B(n32867), .Z(n32873) );
  XOR U42182 ( .A(n32872), .B(n32873), .Z(n32876) );
  XOR U42183 ( .A(n32875), .B(n32876), .Z(n32881) );
  IV U42184 ( .A(n29300), .Z(n29301) );
  NOR U42185 ( .A(n29302), .B(n29301), .Z(n32879) );
  XOR U42186 ( .A(n32881), .B(n32879), .Z(n32883) );
  XOR U42187 ( .A(n32882), .B(n32883), .Z(n32887) );
  IV U42188 ( .A(n29303), .Z(n29305) );
  NOR U42189 ( .A(n29305), .B(n29304), .Z(n29306) );
  IV U42190 ( .A(n29306), .Z(n32886) );
  XOR U42191 ( .A(n32887), .B(n32886), .Z(n32781) );
  IV U42192 ( .A(n29307), .Z(n32782) );
  NOR U42193 ( .A(n32782), .B(n29308), .Z(n29312) );
  IV U42194 ( .A(n29309), .Z(n29311) );
  NOR U42195 ( .A(n29311), .B(n29310), .Z(n32888) );
  NOR U42196 ( .A(n29312), .B(n32888), .Z(n29313) );
  XOR U42197 ( .A(n32781), .B(n29313), .Z(n32898) );
  XOR U42198 ( .A(n32896), .B(n32898), .Z(n32777) );
  XOR U42199 ( .A(n32776), .B(n32777), .Z(n32895) );
  XOR U42200 ( .A(n32893), .B(n32895), .Z(n32910) );
  XOR U42201 ( .A(n32904), .B(n32910), .Z(n32774) );
  XOR U42202 ( .A(n29314), .B(n32774), .Z(n32916) );
  XOR U42203 ( .A(n32914), .B(n32916), .Z(n32771) );
  XOR U42204 ( .A(n32770), .B(n32771), .Z(n32921) );
  XOR U42205 ( .A(n29315), .B(n32921), .Z(n32946) );
  XOR U42206 ( .A(n29316), .B(n32946), .Z(n32761) );
  XOR U42207 ( .A(n29317), .B(n32761), .Z(n32754) );
  XOR U42208 ( .A(n29318), .B(n32754), .Z(n29319) );
  IV U42209 ( .A(n29319), .Z(n32749) );
  XOR U42210 ( .A(n32747), .B(n32749), .Z(n32733) );
  XOR U42211 ( .A(n29328), .B(n32733), .Z(n29320) );
  NOR U42212 ( .A(n29321), .B(n29320), .Z(n36253) );
  IV U42213 ( .A(n29322), .Z(n29324) );
  NOR U42214 ( .A(n29324), .B(n29323), .Z(n29325) );
  IV U42215 ( .A(n29325), .Z(n32731) );
  NOR U42216 ( .A(n29326), .B(n32734), .Z(n29327) );
  NOR U42217 ( .A(n29328), .B(n29327), .Z(n29329) );
  IV U42218 ( .A(n29329), .Z(n29330) );
  XOR U42219 ( .A(n29330), .B(n32733), .Z(n32730) );
  XOR U42220 ( .A(n32731), .B(n32730), .Z(n29331) );
  NOR U42221 ( .A(n29332), .B(n29331), .Z(n29333) );
  NOR U42222 ( .A(n36253), .B(n29333), .Z(n29334) );
  IV U42223 ( .A(n29334), .Z(n32953) );
  XOR U42224 ( .A(n32952), .B(n32953), .Z(n32957) );
  XOR U42225 ( .A(n32955), .B(n32957), .Z(n32725) );
  XOR U42226 ( .A(n29335), .B(n32725), .Z(n29340) );
  NOR U42227 ( .A(n29336), .B(n29340), .Z(n29338) );
  IV U42228 ( .A(n29336), .Z(n29337) );
  NOR U42229 ( .A(n29337), .B(n32725), .Z(n36264) );
  NOR U42230 ( .A(n29338), .B(n36264), .Z(n32961) );
  XOR U42231 ( .A(n32960), .B(n32961), .Z(n29351) );
  NOR U42232 ( .A(n29339), .B(n29351), .Z(n29343) );
  IV U42233 ( .A(n29339), .Z(n29342) );
  IV U42234 ( .A(n29340), .Z(n29341) );
  NOR U42235 ( .A(n29342), .B(n29341), .Z(n36082) );
  NOR U42236 ( .A(n29343), .B(n36082), .Z(n29349) );
  IV U42237 ( .A(n29349), .Z(n29344) );
  NOR U42238 ( .A(n29345), .B(n29344), .Z(n36283) );
  NOR U42239 ( .A(n29358), .B(n36283), .Z(n29346) );
  IV U42240 ( .A(n29346), .Z(n29357) );
  IV U42241 ( .A(n29347), .Z(n29348) );
  NOR U42242 ( .A(n29348), .B(n36074), .Z(n29350) );
  NOR U42243 ( .A(n29350), .B(n29349), .Z(n29354) );
  IV U42244 ( .A(n29350), .Z(n29353) );
  IV U42245 ( .A(n29351), .Z(n29352) );
  NOR U42246 ( .A(n29353), .B(n29352), .Z(n36272) );
  NOR U42247 ( .A(n29354), .B(n36272), .Z(n32714) );
  NOR U42248 ( .A(n29355), .B(n32714), .Z(n29356) );
  NOR U42249 ( .A(n29357), .B(n29356), .Z(n29361) );
  IV U42250 ( .A(n29358), .Z(n29359) );
  NOR U42251 ( .A(n32714), .B(n29359), .Z(n29360) );
  NOR U42252 ( .A(n29361), .B(n29360), .Z(n32712) );
  XOR U42253 ( .A(n29362), .B(n32712), .Z(n29373) );
  IV U42254 ( .A(n29373), .Z(n29367) );
  IV U42255 ( .A(n29363), .Z(n29381) );
  IV U42256 ( .A(n29364), .Z(n29365) );
  NOR U42257 ( .A(n29381), .B(n29365), .Z(n29372) );
  IV U42258 ( .A(n29372), .Z(n29366) );
  NOR U42259 ( .A(n29367), .B(n29366), .Z(n36065) );
  IV U42260 ( .A(n29368), .Z(n29370) );
  NOR U42261 ( .A(n29370), .B(n29369), .Z(n29376) );
  IV U42262 ( .A(n29376), .Z(n29371) );
  NOR U42263 ( .A(n32712), .B(n29371), .Z(n32969) );
  NOR U42264 ( .A(n29373), .B(n29372), .Z(n29374) );
  IV U42265 ( .A(n29374), .Z(n29375) );
  NOR U42266 ( .A(n29376), .B(n29375), .Z(n29377) );
  NOR U42267 ( .A(n32969), .B(n29377), .Z(n29378) );
  IV U42268 ( .A(n29378), .Z(n32967) );
  NOR U42269 ( .A(n36065), .B(n32967), .Z(n32702) );
  IV U42270 ( .A(n29379), .Z(n29380) );
  NOR U42271 ( .A(n29381), .B(n29380), .Z(n32965) );
  IV U42272 ( .A(n29382), .Z(n29383) );
  NOR U42273 ( .A(n29383), .B(n29385), .Z(n32705) );
  IV U42274 ( .A(n29384), .Z(n29386) );
  NOR U42275 ( .A(n29386), .B(n29385), .Z(n32703) );
  NOR U42276 ( .A(n32705), .B(n32703), .Z(n29387) );
  IV U42277 ( .A(n29387), .Z(n29388) );
  NOR U42278 ( .A(n32965), .B(n29388), .Z(n29389) );
  XOR U42279 ( .A(n32702), .B(n29389), .Z(n32977) );
  IV U42280 ( .A(n29390), .Z(n29391) );
  NOR U42281 ( .A(n29392), .B(n29391), .Z(n32698) );
  XOR U42282 ( .A(n32977), .B(n32698), .Z(n29393) );
  XOR U42283 ( .A(n29394), .B(n29393), .Z(n32688) );
  XOR U42284 ( .A(n29395), .B(n32688), .Z(n32984) );
  XOR U42285 ( .A(n32983), .B(n32984), .Z(n29396) );
  NOR U42286 ( .A(n29401), .B(n29396), .Z(n36044) );
  IV U42287 ( .A(n29397), .Z(n29399) );
  NOR U42288 ( .A(n29399), .B(n29398), .Z(n32981) );
  NOR U42289 ( .A(n32983), .B(n32981), .Z(n29400) );
  XOR U42290 ( .A(n29400), .B(n32984), .Z(n32684) );
  XOR U42291 ( .A(n32683), .B(n32684), .Z(n29403) );
  NOR U42292 ( .A(n32684), .B(n29401), .Z(n29402) );
  NOR U42293 ( .A(n29403), .B(n29402), .Z(n29404) );
  NOR U42294 ( .A(n36044), .B(n29404), .Z(n29414) );
  XOR U42295 ( .A(n32681), .B(n29414), .Z(n29409) );
  IV U42296 ( .A(n29405), .Z(n29407) );
  NOR U42297 ( .A(n29407), .B(n29406), .Z(n29408) );
  IV U42298 ( .A(n29408), .Z(n29420) );
  NOR U42299 ( .A(n29409), .B(n29420), .Z(n36031) );
  IV U42300 ( .A(n29410), .Z(n29413) );
  XOR U42301 ( .A(n29411), .B(n29416), .Z(n29412) );
  NOR U42302 ( .A(n29413), .B(n29412), .Z(n32677) );
  IV U42303 ( .A(n29414), .Z(n36035) );
  IV U42304 ( .A(n29415), .Z(n29417) );
  NOR U42305 ( .A(n29417), .B(n29416), .Z(n32675) );
  IV U42306 ( .A(n32681), .Z(n29418) );
  NOR U42307 ( .A(n32675), .B(n29418), .Z(n29419) );
  XOR U42308 ( .A(n36035), .B(n29419), .Z(n32678) );
  XOR U42309 ( .A(n32677), .B(n32678), .Z(n29422) );
  NOR U42310 ( .A(n32678), .B(n29420), .Z(n29421) );
  NOR U42311 ( .A(n29422), .B(n29421), .Z(n29423) );
  NOR U42312 ( .A(n36031), .B(n29423), .Z(n29426) );
  IV U42313 ( .A(n29426), .Z(n29424) );
  NOR U42314 ( .A(n29425), .B(n29424), .Z(n36029) );
  NOR U42315 ( .A(n29427), .B(n29426), .Z(n32672) );
  XOR U42316 ( .A(n32672), .B(n32670), .Z(n29428) );
  NOR U42317 ( .A(n36029), .B(n29428), .Z(n29429) );
  IV U42318 ( .A(n29429), .Z(n32995) );
  XOR U42319 ( .A(n32994), .B(n32995), .Z(n32998) );
  XOR U42320 ( .A(n32997), .B(n32998), .Z(n36010) );
  XOR U42321 ( .A(n29430), .B(n36010), .Z(n32660) );
  XOR U42322 ( .A(n32658), .B(n32660), .Z(n32653) );
  IV U42323 ( .A(n29431), .Z(n29433) );
  NOR U42324 ( .A(n29433), .B(n29432), .Z(n32651) );
  XOR U42325 ( .A(n32653), .B(n32651), .Z(n32655) );
  XOR U42326 ( .A(n32654), .B(n32655), .Z(n33007) );
  IV U42327 ( .A(n29434), .Z(n29435) );
  NOR U42328 ( .A(n32647), .B(n29435), .Z(n29439) );
  IV U42329 ( .A(n29436), .Z(n29437) );
  NOR U42330 ( .A(n33008), .B(n29437), .Z(n29438) );
  NOR U42331 ( .A(n29439), .B(n29438), .Z(n29440) );
  XOR U42332 ( .A(n33007), .B(n29440), .Z(n33020) );
  XOR U42333 ( .A(n29441), .B(n33020), .Z(n32641) );
  IV U42334 ( .A(n29442), .Z(n29444) );
  NOR U42335 ( .A(n29444), .B(n29443), .Z(n29445) );
  IV U42336 ( .A(n29445), .Z(n32638) );
  XOR U42337 ( .A(n32641), .B(n32638), .Z(n29446) );
  XOR U42338 ( .A(n29447), .B(n29446), .Z(n32634) );
  XOR U42339 ( .A(n32632), .B(n32634), .Z(n32636) );
  XOR U42340 ( .A(n32635), .B(n32636), .Z(n33025) );
  XOR U42341 ( .A(n33024), .B(n33025), .Z(n33028) );
  XOR U42342 ( .A(n33027), .B(n33028), .Z(n32630) );
  IV U42343 ( .A(n29448), .Z(n29450) );
  NOR U42344 ( .A(n29450), .B(n29449), .Z(n29451) );
  IV U42345 ( .A(n29451), .Z(n29462) );
  NOR U42346 ( .A(n32630), .B(n29462), .Z(n35969) );
  IV U42347 ( .A(n29452), .Z(n29453) );
  NOR U42348 ( .A(n29453), .B(n29455), .Z(n32629) );
  IV U42349 ( .A(n29454), .Z(n29456) );
  NOR U42350 ( .A(n29456), .B(n29455), .Z(n32627) );
  NOR U42351 ( .A(n32629), .B(n32627), .Z(n29457) );
  IV U42352 ( .A(n29457), .Z(n29458) );
  XOR U42353 ( .A(n29458), .B(n32630), .Z(n32626) );
  IV U42354 ( .A(n29459), .Z(n29470) );
  IV U42355 ( .A(n29460), .Z(n29461) );
  NOR U42356 ( .A(n29470), .B(n29461), .Z(n29463) );
  IV U42357 ( .A(n29463), .Z(n32625) );
  XOR U42358 ( .A(n32626), .B(n32625), .Z(n29465) );
  NOR U42359 ( .A(n29463), .B(n29462), .Z(n29464) );
  NOR U42360 ( .A(n29465), .B(n29464), .Z(n29466) );
  NOR U42361 ( .A(n35969), .B(n29466), .Z(n29467) );
  IV U42362 ( .A(n29467), .Z(n32621) );
  IV U42363 ( .A(n29468), .Z(n29469) );
  NOR U42364 ( .A(n29470), .B(n29469), .Z(n32619) );
  XOR U42365 ( .A(n32621), .B(n32619), .Z(n32623) );
  IV U42366 ( .A(n29471), .Z(n29472) );
  NOR U42367 ( .A(n29472), .B(n29474), .Z(n32622) );
  IV U42368 ( .A(n29473), .Z(n29475) );
  NOR U42369 ( .A(n29475), .B(n29474), .Z(n32614) );
  NOR U42370 ( .A(n32622), .B(n32614), .Z(n29476) );
  XOR U42371 ( .A(n32623), .B(n29476), .Z(n32617) );
  IV U42372 ( .A(n29477), .Z(n35956) );
  NOR U42373 ( .A(n35956), .B(n35958), .Z(n33034) );
  IV U42374 ( .A(n29478), .Z(n29480) );
  NOR U42375 ( .A(n29480), .B(n29479), .Z(n32616) );
  NOR U42376 ( .A(n33034), .B(n32616), .Z(n29481) );
  XOR U42377 ( .A(n32617), .B(n29481), .Z(n32613) );
  XOR U42378 ( .A(n32611), .B(n32613), .Z(n33041) );
  XOR U42379 ( .A(n33040), .B(n33041), .Z(n33044) );
  XOR U42380 ( .A(n33043), .B(n33044), .Z(n33048) );
  XOR U42381 ( .A(n33047), .B(n33048), .Z(n33051) );
  XOR U42382 ( .A(n33050), .B(n33051), .Z(n33055) );
  XOR U42383 ( .A(n33054), .B(n33055), .Z(n33058) );
  IV U42384 ( .A(n29482), .Z(n29484) );
  IV U42385 ( .A(n29483), .Z(n35947) );
  NOR U42386 ( .A(n29484), .B(n35947), .Z(n29485) );
  NOR U42387 ( .A(n33057), .B(n29485), .Z(n29486) );
  XOR U42388 ( .A(n33058), .B(n29486), .Z(n29487) );
  IV U42389 ( .A(n29487), .Z(n29490) );
  IV U42390 ( .A(n29488), .Z(n36435) );
  NOR U42391 ( .A(n32608), .B(n36435), .Z(n29489) );
  XOR U42392 ( .A(n29490), .B(n29489), .Z(n33064) );
  IV U42393 ( .A(n29491), .Z(n29492) );
  NOR U42394 ( .A(n29493), .B(n29492), .Z(n33062) );
  XOR U42395 ( .A(n33064), .B(n33062), .Z(n33066) );
  XOR U42396 ( .A(n33065), .B(n33066), .Z(n32606) );
  XOR U42397 ( .A(n29494), .B(n32606), .Z(n32586) );
  XOR U42398 ( .A(n29495), .B(n32586), .Z(n32579) );
  XOR U42399 ( .A(n32577), .B(n32579), .Z(n32581) );
  XOR U42400 ( .A(n29496), .B(n32581), .Z(n33080) );
  XOR U42401 ( .A(n33079), .B(n33080), .Z(n32560) );
  NOR U42402 ( .A(n29497), .B(n32567), .Z(n29500) );
  NOR U42403 ( .A(n32561), .B(n29498), .Z(n29499) );
  NOR U42404 ( .A(n29500), .B(n29499), .Z(n29501) );
  XOR U42405 ( .A(n32560), .B(n29501), .Z(n32557) );
  IV U42406 ( .A(n29502), .Z(n29514) );
  NOR U42407 ( .A(n29503), .B(n29514), .Z(n32551) );
  IV U42408 ( .A(n29504), .Z(n29505) );
  NOR U42409 ( .A(n29508), .B(n29505), .Z(n32554) );
  IV U42410 ( .A(n29506), .Z(n29507) );
  NOR U42411 ( .A(n29508), .B(n29507), .Z(n32556) );
  NOR U42412 ( .A(n32554), .B(n32556), .Z(n29509) );
  IV U42413 ( .A(n29509), .Z(n29510) );
  NOR U42414 ( .A(n32551), .B(n29510), .Z(n29511) );
  XOR U42415 ( .A(n32557), .B(n29511), .Z(n29512) );
  IV U42416 ( .A(n29512), .Z(n33086) );
  IV U42417 ( .A(n29513), .Z(n29515) );
  NOR U42418 ( .A(n29515), .B(n29514), .Z(n33084) );
  XOR U42419 ( .A(n33086), .B(n33084), .Z(n35904) );
  XOR U42420 ( .A(n29516), .B(n35904), .Z(n32548) );
  XOR U42421 ( .A(n35901), .B(n32548), .Z(n29540) );
  NOR U42422 ( .A(n29517), .B(n29540), .Z(n29527) );
  IV U42423 ( .A(n29518), .Z(n29521) );
  NOR U42424 ( .A(n32548), .B(n29519), .Z(n29520) );
  IV U42425 ( .A(n29520), .Z(n29523) );
  NOR U42426 ( .A(n29521), .B(n29523), .Z(n36473) );
  IV U42427 ( .A(n29522), .Z(n29524) );
  NOR U42428 ( .A(n29524), .B(n29523), .Z(n36476) );
  NOR U42429 ( .A(n36473), .B(n36476), .Z(n29525) );
  IV U42430 ( .A(n29525), .Z(n29526) );
  NOR U42431 ( .A(n29527), .B(n29526), .Z(n29539) );
  IV U42432 ( .A(n29539), .Z(n29532) );
  IV U42433 ( .A(n29528), .Z(n29530) );
  NOR U42434 ( .A(n29530), .B(n29529), .Z(n29545) );
  IV U42435 ( .A(n29545), .Z(n29531) );
  NOR U42436 ( .A(n29532), .B(n29531), .Z(n32542) );
  IV U42437 ( .A(n29533), .Z(n29534) );
  NOR U42438 ( .A(n29534), .B(n29536), .Z(n32545) );
  IV U42439 ( .A(n29535), .Z(n29537) );
  NOR U42440 ( .A(n29537), .B(n29536), .Z(n32543) );
  NOR U42441 ( .A(n32545), .B(n32543), .Z(n29541) );
  IV U42442 ( .A(n29541), .Z(n29538) );
  NOR U42443 ( .A(n29539), .B(n29538), .Z(n29543) );
  IV U42444 ( .A(n29540), .Z(n32546) );
  NOR U42445 ( .A(n29541), .B(n32546), .Z(n29542) );
  NOR U42446 ( .A(n29543), .B(n29542), .Z(n29544) );
  NOR U42447 ( .A(n29545), .B(n29544), .Z(n29546) );
  NOR U42448 ( .A(n32542), .B(n29546), .Z(n33093) );
  XOR U42449 ( .A(n29547), .B(n33093), .Z(n32537) );
  NOR U42450 ( .A(n29548), .B(n32538), .Z(n32532) );
  IV U42451 ( .A(n29561), .Z(n32526) );
  NOR U42452 ( .A(n29559), .B(n32526), .Z(n29563) );
  NOR U42453 ( .A(n32532), .B(n29563), .Z(n29549) );
  XOR U42454 ( .A(n32537), .B(n29549), .Z(n29557) );
  IV U42455 ( .A(n29557), .Z(n35889) );
  IV U42456 ( .A(n29550), .Z(n29552) );
  IV U42457 ( .A(n29551), .Z(n29578) );
  NOR U42458 ( .A(n29552), .B(n29578), .Z(n29575) );
  IV U42459 ( .A(n29575), .Z(n29553) );
  NOR U42460 ( .A(n35889), .B(n29553), .Z(n36504) );
  NOR U42461 ( .A(n29555), .B(n29554), .Z(n29556) );
  NOR U42462 ( .A(n29557), .B(n29556), .Z(n29574) );
  IV U42463 ( .A(n29558), .Z(n29568) );
  IV U42464 ( .A(n29559), .Z(n29560) );
  NOR U42465 ( .A(n29561), .B(n29560), .Z(n29566) );
  XOR U42466 ( .A(n32532), .B(n32537), .Z(n29562) );
  NOR U42467 ( .A(n29563), .B(n29562), .Z(n29564) );
  IV U42468 ( .A(n29564), .Z(n29565) );
  NOR U42469 ( .A(n29566), .B(n29565), .Z(n29567) );
  IV U42470 ( .A(n29567), .Z(n29570) );
  NOR U42471 ( .A(n29568), .B(n29570), .Z(n36497) );
  IV U42472 ( .A(n29569), .Z(n29571) );
  NOR U42473 ( .A(n29571), .B(n29570), .Z(n36501) );
  NOR U42474 ( .A(n36497), .B(n36501), .Z(n29572) );
  IV U42475 ( .A(n29572), .Z(n29573) );
  NOR U42476 ( .A(n29574), .B(n29573), .Z(n32516) );
  NOR U42477 ( .A(n29575), .B(n32516), .Z(n29576) );
  NOR U42478 ( .A(n36504), .B(n29576), .Z(n32521) );
  IV U42479 ( .A(n29577), .Z(n29579) );
  NOR U42480 ( .A(n29579), .B(n29578), .Z(n29580) );
  IV U42481 ( .A(n29580), .Z(n35892) );
  XOR U42482 ( .A(n32521), .B(n35892), .Z(n29594) );
  NOR U42483 ( .A(n29581), .B(n29594), .Z(n29584) );
  IV U42484 ( .A(n29581), .Z(n29582) );
  NOR U42485 ( .A(n32516), .B(n29582), .Z(n29583) );
  NOR U42486 ( .A(n29584), .B(n29583), .Z(n35873) );
  IV U42487 ( .A(n29585), .Z(n29587) );
  NOR U42488 ( .A(n29587), .B(n29586), .Z(n29600) );
  IV U42489 ( .A(n29600), .Z(n29588) );
  NOR U42490 ( .A(n35873), .B(n29588), .Z(n35875) );
  IV U42491 ( .A(n29589), .Z(n29590) );
  NOR U42492 ( .A(n29590), .B(n29592), .Z(n33123) );
  IV U42493 ( .A(n29591), .Z(n29593) );
  NOR U42494 ( .A(n29593), .B(n29592), .Z(n29597) );
  IV U42495 ( .A(n29597), .Z(n29595) );
  NOR U42496 ( .A(n29595), .B(n29594), .Z(n35880) );
  IV U42497 ( .A(n35873), .Z(n29596) );
  NOR U42498 ( .A(n29597), .B(n29596), .Z(n29598) );
  NOR U42499 ( .A(n35880), .B(n29598), .Z(n33124) );
  XOR U42500 ( .A(n33123), .B(n33124), .Z(n29599) );
  NOR U42501 ( .A(n29600), .B(n29599), .Z(n29601) );
  NOR U42502 ( .A(n35875), .B(n29601), .Z(n32514) );
  XOR U42503 ( .A(n29602), .B(n32514), .Z(n32512) );
  XOR U42504 ( .A(n32511), .B(n32512), .Z(n29603) );
  NOR U42505 ( .A(n29605), .B(n29603), .Z(n29608) );
  IV U42506 ( .A(n29604), .Z(n35870) );
  XOR U42507 ( .A(n32514), .B(n35870), .Z(n29607) );
  IV U42508 ( .A(n29605), .Z(n29606) );
  NOR U42509 ( .A(n29607), .B(n29606), .Z(n39549) );
  NOR U42510 ( .A(n29608), .B(n39549), .Z(n29618) );
  IV U42511 ( .A(n29618), .Z(n33144) );
  XOR U42512 ( .A(n33143), .B(n33144), .Z(n29614) );
  IV U42513 ( .A(n29609), .Z(n29612) );
  IV U42514 ( .A(n29610), .Z(n29611) );
  NOR U42515 ( .A(n29612), .B(n29611), .Z(n29622) );
  IV U42516 ( .A(n29622), .Z(n29613) );
  NOR U42517 ( .A(n29614), .B(n29613), .Z(n35863) );
  IV U42518 ( .A(n29615), .Z(n29616) );
  NOR U42519 ( .A(n29617), .B(n29616), .Z(n33141) );
  NOR U42520 ( .A(n33143), .B(n33141), .Z(n29619) );
  XOR U42521 ( .A(n29619), .B(n29618), .Z(n32509) );
  IV U42522 ( .A(n29620), .Z(n32510) );
  XOR U42523 ( .A(n32509), .B(n32510), .Z(n29621) );
  NOR U42524 ( .A(n29622), .B(n29621), .Z(n29623) );
  NOR U42525 ( .A(n35863), .B(n29623), .Z(n32506) );
  NOR U42526 ( .A(n29624), .B(n33158), .Z(n29629) );
  IV U42527 ( .A(n29625), .Z(n29628) );
  IV U42528 ( .A(n29626), .Z(n29627) );
  NOR U42529 ( .A(n29628), .B(n29627), .Z(n32507) );
  NOR U42530 ( .A(n29629), .B(n32507), .Z(n29630) );
  XOR U42531 ( .A(n32506), .B(n29630), .Z(n33177) );
  IV U42532 ( .A(n29631), .Z(n32503) );
  NOR U42533 ( .A(n29632), .B(n32503), .Z(n29635) );
  IV U42534 ( .A(n29633), .Z(n29634) );
  NOR U42535 ( .A(n29634), .B(n29638), .Z(n33175) );
  NOR U42536 ( .A(n29635), .B(n33175), .Z(n29636) );
  XOR U42537 ( .A(n33177), .B(n29636), .Z(n32495) );
  IV U42538 ( .A(n29637), .Z(n29639) );
  NOR U42539 ( .A(n29639), .B(n29638), .Z(n33172) );
  IV U42540 ( .A(n29640), .Z(n32496) );
  NOR U42541 ( .A(n29641), .B(n32496), .Z(n29642) );
  NOR U42542 ( .A(n33172), .B(n29642), .Z(n29643) );
  XOR U42543 ( .A(n32495), .B(n29643), .Z(n35831) );
  NOR U42544 ( .A(n29644), .B(n35834), .Z(n32492) );
  IV U42545 ( .A(n29652), .Z(n29646) );
  IV U42546 ( .A(n29645), .Z(n29651) );
  NOR U42547 ( .A(n29646), .B(n29651), .Z(n32490) );
  NOR U42548 ( .A(n32492), .B(n32490), .Z(n29647) );
  XOR U42549 ( .A(n35831), .B(n29647), .Z(n29656) );
  IV U42550 ( .A(n29648), .Z(n29649) );
  NOR U42551 ( .A(n29649), .B(n29651), .Z(n32488) );
  IV U42552 ( .A(n29650), .Z(n29654) );
  XOR U42553 ( .A(n29652), .B(n29651), .Z(n29653) );
  NOR U42554 ( .A(n29654), .B(n29653), .Z(n32485) );
  NOR U42555 ( .A(n32488), .B(n32485), .Z(n29655) );
  XOR U42556 ( .A(n29656), .B(n29655), .Z(n32484) );
  IV U42557 ( .A(n29657), .Z(n32476) );
  NOR U42558 ( .A(n32476), .B(n29658), .Z(n29662) );
  IV U42559 ( .A(n29659), .Z(n29661) );
  NOR U42560 ( .A(n29661), .B(n29660), .Z(n32482) );
  NOR U42561 ( .A(n29662), .B(n32482), .Z(n29663) );
  XOR U42562 ( .A(n32484), .B(n29663), .Z(n32473) );
  XOR U42563 ( .A(n32474), .B(n32473), .Z(n32469) );
  XOR U42564 ( .A(n32468), .B(n32469), .Z(n33183) );
  XOR U42565 ( .A(n29664), .B(n33183), .Z(n32460) );
  XOR U42566 ( .A(n29665), .B(n32460), .Z(n33197) );
  XOR U42567 ( .A(n29666), .B(n33197), .Z(n33200) );
  XOR U42568 ( .A(n33199), .B(n33200), .Z(n33205) );
  IV U42569 ( .A(n29667), .Z(n29670) );
  IV U42570 ( .A(n29668), .Z(n29669) );
  NOR U42571 ( .A(n29670), .B(n29669), .Z(n33203) );
  XOR U42572 ( .A(n33205), .B(n33203), .Z(n33207) );
  XOR U42573 ( .A(n33206), .B(n33207), .Z(n33214) );
  NOR U42574 ( .A(n32451), .B(n29671), .Z(n29675) );
  IV U42575 ( .A(n29672), .Z(n29674) );
  IV U42576 ( .A(n29673), .Z(n29680) );
  NOR U42577 ( .A(n29674), .B(n29680), .Z(n33212) );
  NOR U42578 ( .A(n29675), .B(n33212), .Z(n29676) );
  XOR U42579 ( .A(n33214), .B(n29676), .Z(n33209) );
  NOR U42580 ( .A(n29678), .B(n29677), .Z(n33216) );
  IV U42581 ( .A(n29679), .Z(n29681) );
  NOR U42582 ( .A(n29681), .B(n29680), .Z(n33210) );
  NOR U42583 ( .A(n33216), .B(n33210), .Z(n29682) );
  XOR U42584 ( .A(n33209), .B(n29682), .Z(n33219) );
  XOR U42585 ( .A(n33220), .B(n33219), .Z(n29687) );
  IV U42586 ( .A(n29687), .Z(n36561) );
  XOR U42587 ( .A(n32448), .B(n36561), .Z(n29683) );
  NOR U42588 ( .A(n29684), .B(n29683), .Z(n36572) );
  NOR U42589 ( .A(n36564), .B(n29685), .Z(n32446) );
  NOR U42590 ( .A(n32446), .B(n32448), .Z(n29686) );
  XOR U42591 ( .A(n29687), .B(n29686), .Z(n29696) );
  IV U42592 ( .A(n29696), .Z(n29688) );
  NOR U42593 ( .A(n29689), .B(n29688), .Z(n29690) );
  NOR U42594 ( .A(n36572), .B(n29690), .Z(n32437) );
  IV U42595 ( .A(n29691), .Z(n32438) );
  NOR U42596 ( .A(n29692), .B(n32438), .Z(n29702) );
  IV U42597 ( .A(n29702), .Z(n29693) );
  NOR U42598 ( .A(n32437), .B(n29693), .Z(n29704) );
  NOR U42599 ( .A(n29695), .B(n29694), .Z(n29698) );
  IV U42600 ( .A(n29698), .Z(n29697) );
  NOR U42601 ( .A(n29697), .B(n29696), .Z(n32444) );
  NOR U42602 ( .A(n32437), .B(n29698), .Z(n29699) );
  NOR U42603 ( .A(n32444), .B(n29699), .Z(n29700) );
  IV U42604 ( .A(n29700), .Z(n29701) );
  NOR U42605 ( .A(n29702), .B(n29701), .Z(n29703) );
  NOR U42606 ( .A(n29704), .B(n29703), .Z(n33239) );
  XOR U42607 ( .A(n33233), .B(n33239), .Z(n33236) );
  XOR U42608 ( .A(n33235), .B(n33236), .Z(n32432) );
  XOR U42609 ( .A(n29705), .B(n32432), .Z(n29716) );
  XOR U42610 ( .A(n29706), .B(n29716), .Z(n29708) );
  NOR U42611 ( .A(n29707), .B(n29708), .Z(n35742) );
  IV U42612 ( .A(n29708), .Z(n29715) );
  IV U42613 ( .A(n29709), .Z(n29710) );
  NOR U42614 ( .A(n29710), .B(n29712), .Z(n35752) );
  IV U42615 ( .A(n29711), .Z(n29713) );
  NOR U42616 ( .A(n29713), .B(n29712), .Z(n35747) );
  NOR U42617 ( .A(n35752), .B(n35747), .Z(n29717) );
  IV U42618 ( .A(n29717), .Z(n29714) );
  NOR U42619 ( .A(n29715), .B(n29714), .Z(n29718) );
  IV U42620 ( .A(n29716), .Z(n35756) );
  XOR U42621 ( .A(n33247), .B(n35756), .Z(n35749) );
  NOR U42622 ( .A(n29717), .B(n35749), .Z(n33253) );
  NOR U42623 ( .A(n29718), .B(n33253), .Z(n29719) );
  NOR U42624 ( .A(n29720), .B(n29719), .Z(n29721) );
  NOR U42625 ( .A(n35742), .B(n29721), .Z(n29725) );
  IV U42626 ( .A(n29725), .Z(n32427) );
  NOR U42627 ( .A(n29722), .B(n32427), .Z(n33261) );
  IV U42628 ( .A(n29723), .Z(n32428) );
  NOR U42629 ( .A(n32428), .B(n29724), .Z(n29726) );
  XOR U42630 ( .A(n29726), .B(n29725), .Z(n29733) );
  NOR U42631 ( .A(n29727), .B(n29733), .Z(n29728) );
  NOR U42632 ( .A(n33261), .B(n29728), .Z(n29731) );
  IV U42633 ( .A(n29731), .Z(n35736) );
  NOR U42634 ( .A(n29729), .B(n35736), .Z(n42324) );
  NOR U42635 ( .A(n29730), .B(n33256), .Z(n29732) );
  NOR U42636 ( .A(n29731), .B(n29732), .Z(n29736) );
  IV U42637 ( .A(n29732), .Z(n29734) );
  IV U42638 ( .A(n29733), .Z(n33255) );
  NOR U42639 ( .A(n29734), .B(n33255), .Z(n29735) );
  NOR U42640 ( .A(n29736), .B(n29735), .Z(n29737) );
  NOR U42641 ( .A(n32425), .B(n29737), .Z(n29738) );
  NOR U42642 ( .A(n42324), .B(n29738), .Z(n32421) );
  IV U42643 ( .A(n29739), .Z(n29741) );
  NOR U42644 ( .A(n29741), .B(n29740), .Z(n42328) );
  NOR U42645 ( .A(n33278), .B(n32423), .Z(n29742) );
  NOR U42646 ( .A(n42328), .B(n29742), .Z(n29743) );
  XOR U42647 ( .A(n32421), .B(n29743), .Z(n38922) );
  IV U42648 ( .A(n29744), .Z(n29745) );
  NOR U42649 ( .A(n29745), .B(n29753), .Z(n33286) );
  IV U42650 ( .A(n29746), .Z(n29748) );
  IV U42651 ( .A(n29747), .Z(n29750) );
  NOR U42652 ( .A(n29748), .B(n29750), .Z(n33281) );
  IV U42653 ( .A(n33281), .Z(n38924) );
  IV U42654 ( .A(n29749), .Z(n29751) );
  NOR U42655 ( .A(n29751), .B(n29750), .Z(n39657) );
  IV U42656 ( .A(n29752), .Z(n29754) );
  NOR U42657 ( .A(n29754), .B(n29753), .Z(n33282) );
  NOR U42658 ( .A(n39657), .B(n33282), .Z(n29755) );
  XOR U42659 ( .A(n38924), .B(n29755), .Z(n29756) );
  NOR U42660 ( .A(n33286), .B(n29756), .Z(n29757) );
  XOR U42661 ( .A(n38922), .B(n29757), .Z(n32417) );
  XOR U42662 ( .A(n29758), .B(n32417), .Z(n32411) );
  IV U42663 ( .A(n29759), .Z(n29760) );
  NOR U42664 ( .A(n29761), .B(n29760), .Z(n32409) );
  XOR U42665 ( .A(n32411), .B(n32409), .Z(n32414) );
  XOR U42666 ( .A(n29762), .B(n32414), .Z(n29769) );
  XOR U42667 ( .A(n29763), .B(n29769), .Z(n32404) );
  XOR U42668 ( .A(n32403), .B(n32404), .Z(n29772) );
  NOR U42669 ( .A(n29764), .B(n29772), .Z(n36636) );
  IV U42670 ( .A(n29765), .Z(n29768) );
  IV U42671 ( .A(n29766), .Z(n29767) );
  NOR U42672 ( .A(n29768), .B(n29767), .Z(n32399) );
  IV U42673 ( .A(n29774), .Z(n29771) );
  IV U42674 ( .A(n29769), .Z(n33296) );
  XOR U42675 ( .A(n33296), .B(n33292), .Z(n29770) );
  NOR U42676 ( .A(n29771), .B(n29770), .Z(n38902) );
  IV U42677 ( .A(n29772), .Z(n29773) );
  NOR U42678 ( .A(n29774), .B(n29773), .Z(n29775) );
  NOR U42679 ( .A(n38902), .B(n29775), .Z(n32400) );
  XOR U42680 ( .A(n32399), .B(n32400), .Z(n29776) );
  NOR U42681 ( .A(n29777), .B(n29776), .Z(n29778) );
  NOR U42682 ( .A(n36636), .B(n29778), .Z(n29794) );
  IV U42683 ( .A(n29794), .Z(n33299) );
  XOR U42684 ( .A(n29793), .B(n33299), .Z(n29783) );
  IV U42685 ( .A(n29779), .Z(n29781) );
  NOR U42686 ( .A(n29781), .B(n29780), .Z(n29782) );
  IV U42687 ( .A(n29782), .Z(n29796) );
  NOR U42688 ( .A(n29783), .B(n29796), .Z(n33311) );
  IV U42689 ( .A(n29784), .Z(n29785) );
  NOR U42690 ( .A(n29786), .B(n29785), .Z(n33313) );
  IV U42691 ( .A(n29787), .Z(n29788) );
  NOR U42692 ( .A(n29788), .B(n29791), .Z(n29789) );
  IV U42693 ( .A(n29789), .Z(n33309) );
  IV U42694 ( .A(n29790), .Z(n29792) );
  NOR U42695 ( .A(n29792), .B(n29791), .Z(n32397) );
  NOR U42696 ( .A(n29793), .B(n32397), .Z(n29795) );
  XOR U42697 ( .A(n29795), .B(n29794), .Z(n33308) );
  XOR U42698 ( .A(n33309), .B(n33308), .Z(n33314) );
  XOR U42699 ( .A(n33313), .B(n33314), .Z(n29798) );
  NOR U42700 ( .A(n33314), .B(n29796), .Z(n29797) );
  NOR U42701 ( .A(n29798), .B(n29797), .Z(n29799) );
  NOR U42702 ( .A(n33311), .B(n29799), .Z(n32393) );
  XOR U42703 ( .A(n29800), .B(n32393), .Z(n32376) );
  XOR U42704 ( .A(n29801), .B(n32376), .Z(n29802) );
  IV U42705 ( .A(n29802), .Z(n32373) );
  XOR U42706 ( .A(n32371), .B(n32373), .Z(n29809) );
  XOR U42707 ( .A(n29810), .B(n29809), .Z(n43186) );
  IV U42708 ( .A(n29803), .Z(n29804) );
  NOR U42709 ( .A(n29804), .B(n29825), .Z(n29821) );
  IV U42710 ( .A(n29821), .Z(n29805) );
  NOR U42711 ( .A(n43186), .B(n29805), .Z(n35673) );
  IV U42712 ( .A(n29806), .Z(n29808) );
  NOR U42713 ( .A(n29808), .B(n29807), .Z(n29813) );
  NOR U42714 ( .A(n29810), .B(n29809), .Z(n29811) );
  IV U42715 ( .A(n29811), .Z(n29812) );
  NOR U42716 ( .A(n29813), .B(n29812), .Z(n29814) );
  IV U42717 ( .A(n29814), .Z(n35677) );
  NOR U42718 ( .A(n29816), .B(n35677), .Z(n33322) );
  NOR U42719 ( .A(n29816), .B(n29815), .Z(n29818) );
  IV U42720 ( .A(n43186), .Z(n29817) );
  NOR U42721 ( .A(n29818), .B(n29817), .Z(n29819) );
  NOR U42722 ( .A(n33322), .B(n29819), .Z(n29820) );
  NOR U42723 ( .A(n29821), .B(n29820), .Z(n29822) );
  NOR U42724 ( .A(n35673), .B(n29822), .Z(n29823) );
  IV U42725 ( .A(n29823), .Z(n32360) );
  IV U42726 ( .A(n29824), .Z(n29826) );
  NOR U42727 ( .A(n29826), .B(n29825), .Z(n32359) );
  XOR U42728 ( .A(n32360), .B(n32359), .Z(n32363) );
  IV U42729 ( .A(n32363), .Z(n29832) );
  IV U42730 ( .A(n29833), .Z(n32354) );
  IV U42731 ( .A(n29834), .Z(n29827) );
  NOR U42732 ( .A(n32354), .B(n29827), .Z(n32357) );
  IV U42733 ( .A(n29828), .Z(n29830) );
  NOR U42734 ( .A(n29830), .B(n29829), .Z(n32361) );
  NOR U42735 ( .A(n32357), .B(n32361), .Z(n29831) );
  XOR U42736 ( .A(n29832), .B(n29831), .Z(n32348) );
  XOR U42737 ( .A(n29834), .B(n29833), .Z(n29835) );
  NOR U42738 ( .A(n32352), .B(n29835), .Z(n29838) );
  NOR U42739 ( .A(n32347), .B(n29836), .Z(n29837) );
  NOR U42740 ( .A(n29838), .B(n29837), .Z(n29839) );
  XOR U42741 ( .A(n32348), .B(n29839), .Z(n33329) );
  XOR U42742 ( .A(n33327), .B(n33329), .Z(n33331) );
  XOR U42743 ( .A(n33330), .B(n33331), .Z(n33335) );
  XOR U42744 ( .A(n33334), .B(n33335), .Z(n33346) );
  XOR U42745 ( .A(n29840), .B(n33346), .Z(n29841) );
  IV U42746 ( .A(n29841), .Z(n33350) );
  IV U42747 ( .A(n29842), .Z(n29844) );
  NOR U42748 ( .A(n29844), .B(n29843), .Z(n33348) );
  XOR U42749 ( .A(n33350), .B(n33348), .Z(n32337) );
  XOR U42750 ( .A(n32338), .B(n32337), .Z(n33354) );
  IV U42751 ( .A(n29845), .Z(n32334) );
  NOR U42752 ( .A(n32334), .B(n29846), .Z(n29849) );
  IV U42753 ( .A(n29847), .Z(n29848) );
  NOR U42754 ( .A(n29848), .B(n29852), .Z(n33353) );
  NOR U42755 ( .A(n29849), .B(n33353), .Z(n29850) );
  XOR U42756 ( .A(n33354), .B(n29850), .Z(n33359) );
  IV U42757 ( .A(n29851), .Z(n29853) );
  NOR U42758 ( .A(n29853), .B(n29852), .Z(n33357) );
  XOR U42759 ( .A(n33359), .B(n33357), .Z(n33365) );
  XOR U42760 ( .A(n33360), .B(n33365), .Z(n29854) );
  NOR U42761 ( .A(n29855), .B(n29854), .Z(n43228) );
  IV U42762 ( .A(n29856), .Z(n29863) );
  IV U42763 ( .A(n29857), .Z(n29858) );
  NOR U42764 ( .A(n29863), .B(n29858), .Z(n33363) );
  NOR U42765 ( .A(n33363), .B(n33360), .Z(n29859) );
  IV U42766 ( .A(n29859), .Z(n29860) );
  XOR U42767 ( .A(n29860), .B(n33365), .Z(n33367) );
  IV U42768 ( .A(n29861), .Z(n29862) );
  NOR U42769 ( .A(n29863), .B(n29862), .Z(n29864) );
  IV U42770 ( .A(n29864), .Z(n33366) );
  XOR U42771 ( .A(n33367), .B(n33366), .Z(n29865) );
  NOR U42772 ( .A(n29866), .B(n29865), .Z(n29867) );
  NOR U42773 ( .A(n43228), .B(n29867), .Z(n33369) );
  XOR U42774 ( .A(n33371), .B(n33369), .Z(n33377) );
  XOR U42775 ( .A(n32328), .B(n33377), .Z(n32330) );
  NOR U42776 ( .A(n32329), .B(n33376), .Z(n29868) );
  XOR U42777 ( .A(n32330), .B(n29868), .Z(n33375) );
  XOR U42778 ( .A(n33373), .B(n33375), .Z(n33388) );
  XOR U42779 ( .A(n33380), .B(n33388), .Z(n33384) );
  XOR U42780 ( .A(n33382), .B(n33384), .Z(n33395) );
  XOR U42781 ( .A(n29869), .B(n33395), .Z(n33402) );
  IV U42782 ( .A(n29870), .Z(n29872) );
  IV U42783 ( .A(n29871), .Z(n29885) );
  NOR U42784 ( .A(n29872), .B(n29885), .Z(n29873) );
  IV U42785 ( .A(n29873), .Z(n29879) );
  NOR U42786 ( .A(n33402), .B(n29879), .Z(n35601) );
  IV U42787 ( .A(n29874), .Z(n29875) );
  NOR U42788 ( .A(n29878), .B(n29875), .Z(n33400) );
  XOR U42789 ( .A(n33402), .B(n33400), .Z(n33404) );
  IV U42790 ( .A(n29876), .Z(n29877) );
  NOR U42791 ( .A(n29878), .B(n29877), .Z(n29880) );
  IV U42792 ( .A(n29880), .Z(n33403) );
  XOR U42793 ( .A(n33404), .B(n33403), .Z(n29882) );
  NOR U42794 ( .A(n29880), .B(n29879), .Z(n29881) );
  NOR U42795 ( .A(n29882), .B(n29881), .Z(n29883) );
  NOR U42796 ( .A(n35601), .B(n29883), .Z(n32320) );
  IV U42797 ( .A(n29884), .Z(n29886) );
  NOR U42798 ( .A(n29886), .B(n29885), .Z(n32325) );
  XOR U42799 ( .A(n32320), .B(n32325), .Z(n32310) );
  NOR U42800 ( .A(n32321), .B(n29887), .Z(n32314) );
  IV U42801 ( .A(n29888), .Z(n32311) );
  NOR U42802 ( .A(n29889), .B(n32311), .Z(n29890) );
  NOR U42803 ( .A(n32314), .B(n29890), .Z(n29891) );
  XOR U42804 ( .A(n32310), .B(n29891), .Z(n33409) );
  XOR U42805 ( .A(n33407), .B(n33409), .Z(n33415) );
  XOR U42806 ( .A(n33414), .B(n33415), .Z(n33419) );
  IV U42807 ( .A(n29892), .Z(n29893) );
  NOR U42808 ( .A(n29894), .B(n29893), .Z(n32307) );
  IV U42809 ( .A(n29895), .Z(n29897) );
  NOR U42810 ( .A(n29897), .B(n29896), .Z(n33417) );
  NOR U42811 ( .A(n32307), .B(n33417), .Z(n29898) );
  XOR U42812 ( .A(n33419), .B(n29898), .Z(n29899) );
  NOR U42813 ( .A(n29900), .B(n29899), .Z(n33423) );
  IV U42814 ( .A(n29900), .Z(n29902) );
  XOR U42815 ( .A(n33417), .B(n33419), .Z(n29901) );
  NOR U42816 ( .A(n29902), .B(n29901), .Z(n36740) );
  NOR U42817 ( .A(n33423), .B(n36740), .Z(n32302) );
  XOR U42818 ( .A(n29903), .B(n32302), .Z(n32301) );
  XOR U42819 ( .A(n32300), .B(n32301), .Z(n33433) );
  IV U42820 ( .A(n29904), .Z(n32296) );
  NOR U42821 ( .A(n32296), .B(n29905), .Z(n29908) );
  IV U42822 ( .A(n29906), .Z(n29907) );
  NOR U42823 ( .A(n29907), .B(n29918), .Z(n33434) );
  NOR U42824 ( .A(n29908), .B(n33434), .Z(n29909) );
  XOR U42825 ( .A(n33433), .B(n29909), .Z(n33432) );
  IV U42826 ( .A(n29910), .Z(n29916) );
  IV U42827 ( .A(n29911), .Z(n29912) );
  NOR U42828 ( .A(n29916), .B(n29912), .Z(n29921) );
  IV U42829 ( .A(n29921), .Z(n29913) );
  NOR U42830 ( .A(n33432), .B(n29913), .Z(n35583) );
  IV U42831 ( .A(n29914), .Z(n29915) );
  NOR U42832 ( .A(n29916), .B(n29915), .Z(n32293) );
  IV U42833 ( .A(n29917), .Z(n29919) );
  NOR U42834 ( .A(n29919), .B(n29918), .Z(n33430) );
  NOR U42835 ( .A(n32293), .B(n33430), .Z(n29920) );
  XOR U42836 ( .A(n33432), .B(n29920), .Z(n29926) );
  NOR U42837 ( .A(n29921), .B(n29926), .Z(n29922) );
  NOR U42838 ( .A(n35583), .B(n29922), .Z(n29928) );
  IV U42839 ( .A(n29928), .Z(n36786) );
  NOR U42840 ( .A(n29931), .B(n36786), .Z(n33445) );
  IV U42841 ( .A(n29923), .Z(n29924) );
  NOR U42842 ( .A(n29924), .B(n29936), .Z(n33446) );
  NOR U42843 ( .A(n29925), .B(n33440), .Z(n29929) );
  IV U42844 ( .A(n29929), .Z(n29927) );
  IV U42845 ( .A(n29926), .Z(n33439) );
  NOR U42846 ( .A(n29927), .B(n33439), .Z(n32290) );
  NOR U42847 ( .A(n29929), .B(n29928), .Z(n29930) );
  NOR U42848 ( .A(n32290), .B(n29930), .Z(n33447) );
  XOR U42849 ( .A(n33446), .B(n33447), .Z(n29933) );
  NOR U42850 ( .A(n33447), .B(n29931), .Z(n29932) );
  NOR U42851 ( .A(n29933), .B(n29932), .Z(n29934) );
  NOR U42852 ( .A(n33445), .B(n29934), .Z(n32287) );
  IV U42853 ( .A(n29935), .Z(n29937) );
  NOR U42854 ( .A(n29937), .B(n29936), .Z(n33450) );
  NOR U42855 ( .A(n33450), .B(n29938), .Z(n29939) );
  XOR U42856 ( .A(n32287), .B(n29939), .Z(n33466) );
  XOR U42857 ( .A(n29940), .B(n33466), .Z(n33470) );
  IV U42858 ( .A(n29941), .Z(n29943) );
  NOR U42859 ( .A(n29943), .B(n29942), .Z(n33468) );
  XOR U42860 ( .A(n33470), .B(n33468), .Z(n33463) );
  XOR U42861 ( .A(n33462), .B(n33463), .Z(n32275) );
  XOR U42862 ( .A(n29944), .B(n32275), .Z(n32271) );
  XOR U42863 ( .A(n32270), .B(n32271), .Z(n32263) );
  IV U42864 ( .A(n29945), .Z(n32269) );
  NOR U42865 ( .A(n32267), .B(n32269), .Z(n29948) );
  IV U42866 ( .A(n29946), .Z(n29947) );
  NOR U42867 ( .A(n29947), .B(n29951), .Z(n32264) );
  NOR U42868 ( .A(n29948), .B(n32264), .Z(n29949) );
  XOR U42869 ( .A(n32263), .B(n29949), .Z(n32259) );
  IV U42870 ( .A(n29950), .Z(n29952) );
  NOR U42871 ( .A(n29952), .B(n29951), .Z(n32257) );
  XOR U42872 ( .A(n32259), .B(n32257), .Z(n32253) );
  XOR U42873 ( .A(n29960), .B(n32253), .Z(n29957) );
  IV U42874 ( .A(n29953), .Z(n29955) );
  NOR U42875 ( .A(n29955), .B(n29954), .Z(n29962) );
  IV U42876 ( .A(n29962), .Z(n29956) );
  NOR U42877 ( .A(n29957), .B(n29956), .Z(n35553) );
  NOR U42878 ( .A(n29958), .B(n32246), .Z(n29959) );
  NOR U42879 ( .A(n29960), .B(n29959), .Z(n29961) );
  XOR U42880 ( .A(n29961), .B(n32253), .Z(n29966) );
  NOR U42881 ( .A(n29962), .B(n29966), .Z(n29963) );
  NOR U42882 ( .A(n35553), .B(n29963), .Z(n29964) );
  NOR U42883 ( .A(n29965), .B(n29964), .Z(n29969) );
  IV U42884 ( .A(n29965), .Z(n29968) );
  IV U42885 ( .A(n29966), .Z(n29967) );
  NOR U42886 ( .A(n29968), .B(n29967), .Z(n39834) );
  NOR U42887 ( .A(n29969), .B(n39834), .Z(n32243) );
  IV U42888 ( .A(n29970), .Z(n29971) );
  NOR U42889 ( .A(n29971), .B(n29973), .Z(n32242) );
  IV U42890 ( .A(n29972), .Z(n29974) );
  NOR U42891 ( .A(n29974), .B(n29973), .Z(n33483) );
  NOR U42892 ( .A(n32242), .B(n33483), .Z(n29975) );
  XOR U42893 ( .A(n32243), .B(n29975), .Z(n42096) );
  XOR U42894 ( .A(n32239), .B(n42096), .Z(n33481) );
  XOR U42895 ( .A(n33480), .B(n33481), .Z(n33492) );
  XOR U42896 ( .A(n29976), .B(n33492), .Z(n29977) );
  IV U42897 ( .A(n29977), .Z(n33498) );
  IV U42898 ( .A(n29978), .Z(n29980) );
  NOR U42899 ( .A(n29980), .B(n29979), .Z(n33496) );
  XOR U42900 ( .A(n33498), .B(n33496), .Z(n32227) );
  IV U42901 ( .A(n29981), .Z(n32228) );
  NOR U42902 ( .A(n32228), .B(n29982), .Z(n29986) );
  IV U42903 ( .A(n29983), .Z(n29985) );
  NOR U42904 ( .A(n29985), .B(n29984), .Z(n32234) );
  NOR U42905 ( .A(n29986), .B(n32234), .Z(n29987) );
  XOR U42906 ( .A(n32227), .B(n29987), .Z(n32220) );
  IV U42907 ( .A(n29988), .Z(n29989) );
  NOR U42908 ( .A(n29989), .B(n29991), .Z(n32221) );
  IV U42909 ( .A(n29990), .Z(n29992) );
  NOR U42910 ( .A(n29992), .B(n29991), .Z(n32223) );
  NOR U42911 ( .A(n32221), .B(n32223), .Z(n29993) );
  XOR U42912 ( .A(n32220), .B(n29993), .Z(n32218) );
  XOR U42913 ( .A(n32217), .B(n32218), .Z(n32211) );
  XOR U42914 ( .A(n32210), .B(n32211), .Z(n33505) );
  NOR U42915 ( .A(n32207), .B(n29994), .Z(n29998) );
  IV U42916 ( .A(n29995), .Z(n33506) );
  NOR U42917 ( .A(n29996), .B(n33506), .Z(n29997) );
  NOR U42918 ( .A(n29998), .B(n29997), .Z(n29999) );
  XOR U42919 ( .A(n33505), .B(n29999), .Z(n33510) );
  IV U42920 ( .A(n30000), .Z(n30001) );
  NOR U42921 ( .A(n30001), .B(n30004), .Z(n33527) );
  NOR U42922 ( .A(n30002), .B(n33511), .Z(n30006) );
  IV U42923 ( .A(n30003), .Z(n30005) );
  NOR U42924 ( .A(n30005), .B(n30004), .Z(n33518) );
  NOR U42925 ( .A(n30006), .B(n33518), .Z(n30007) );
  IV U42926 ( .A(n30007), .Z(n30008) );
  NOR U42927 ( .A(n33527), .B(n30008), .Z(n30009) );
  XOR U42928 ( .A(n33510), .B(n30009), .Z(n33526) );
  XOR U42929 ( .A(n33524), .B(n33526), .Z(n32200) );
  XOR U42930 ( .A(n30021), .B(n32200), .Z(n30011) );
  IV U42931 ( .A(n30010), .Z(n30026) );
  NOR U42932 ( .A(n30011), .B(n30026), .Z(n35522) );
  IV U42933 ( .A(n30012), .Z(n30014) );
  NOR U42934 ( .A(n30014), .B(n30013), .Z(n30020) );
  IV U42935 ( .A(n30015), .Z(n30017) );
  NOR U42936 ( .A(n30017), .B(n30016), .Z(n32199) );
  NOR U42937 ( .A(n30021), .B(n32199), .Z(n30018) );
  XOR U42938 ( .A(n32200), .B(n30018), .Z(n30019) );
  NOR U42939 ( .A(n30020), .B(n30019), .Z(n30025) );
  IV U42940 ( .A(n30020), .Z(n30024) );
  NOR U42941 ( .A(n30021), .B(n32200), .Z(n30022) );
  IV U42942 ( .A(n30022), .Z(n30023) );
  NOR U42943 ( .A(n30024), .B(n30023), .Z(n36893) );
  NOR U42944 ( .A(n30025), .B(n36893), .Z(n33537) );
  XOR U42945 ( .A(n33536), .B(n33537), .Z(n30028) );
  NOR U42946 ( .A(n33537), .B(n30026), .Z(n30027) );
  NOR U42947 ( .A(n30028), .B(n30027), .Z(n30029) );
  NOR U42948 ( .A(n35522), .B(n30029), .Z(n32196) );
  IV U42949 ( .A(n30030), .Z(n30031) );
  NOR U42950 ( .A(n30031), .B(n30033), .Z(n33540) );
  IV U42951 ( .A(n30032), .Z(n30034) );
  NOR U42952 ( .A(n30034), .B(n30033), .Z(n32197) );
  NOR U42953 ( .A(n33540), .B(n32197), .Z(n30035) );
  XOR U42954 ( .A(n32196), .B(n30035), .Z(n32190) );
  XOR U42955 ( .A(n32189), .B(n32190), .Z(n32193) );
  XOR U42956 ( .A(n30036), .B(n32193), .Z(n32184) );
  XOR U42957 ( .A(n32183), .B(n32184), .Z(n33546) );
  XOR U42958 ( .A(n33545), .B(n33546), .Z(n33550) );
  IV U42959 ( .A(n30037), .Z(n30040) );
  IV U42960 ( .A(n30038), .Z(n30039) );
  NOR U42961 ( .A(n30040), .B(n30039), .Z(n33548) );
  XOR U42962 ( .A(n33550), .B(n33548), .Z(n32182) );
  IV U42963 ( .A(n30041), .Z(n30044) );
  IV U42964 ( .A(n30042), .Z(n30043) );
  NOR U42965 ( .A(n30044), .B(n30043), .Z(n32180) );
  XOR U42966 ( .A(n32182), .B(n32180), .Z(n35496) );
  IV U42967 ( .A(n30045), .Z(n30046) );
  NOR U42968 ( .A(n30049), .B(n30046), .Z(n35499) );
  IV U42969 ( .A(n30047), .Z(n30048) );
  NOR U42970 ( .A(n30049), .B(n30048), .Z(n35495) );
  NOR U42971 ( .A(n35499), .B(n35495), .Z(n32175) );
  XOR U42972 ( .A(n35496), .B(n32175), .Z(n30059) );
  IV U42973 ( .A(n30059), .Z(n32177) );
  XOR U42974 ( .A(n32176), .B(n32177), .Z(n30050) );
  NOR U42975 ( .A(n30051), .B(n30050), .Z(n35481) );
  IV U42976 ( .A(n30052), .Z(n30054) );
  IV U42977 ( .A(n30053), .Z(n30057) );
  NOR U42978 ( .A(n30054), .B(n30057), .Z(n30055) );
  IV U42979 ( .A(n30055), .Z(n32174) );
  IV U42980 ( .A(n30056), .Z(n30058) );
  NOR U42981 ( .A(n30058), .B(n30057), .Z(n32171) );
  NOR U42982 ( .A(n32176), .B(n32171), .Z(n30060) );
  XOR U42983 ( .A(n30060), .B(n30059), .Z(n32173) );
  XOR U42984 ( .A(n32174), .B(n32173), .Z(n32166) );
  NOR U42985 ( .A(n30061), .B(n32166), .Z(n30062) );
  NOR U42986 ( .A(n35481), .B(n30062), .Z(n30063) );
  IV U42987 ( .A(n30063), .Z(n33555) );
  IV U42988 ( .A(n30064), .Z(n30066) );
  NOR U42989 ( .A(n30066), .B(n30065), .Z(n33554) );
  XOR U42990 ( .A(n33555), .B(n33554), .Z(n30071) );
  XOR U42991 ( .A(n30067), .B(n30071), .Z(n32163) );
  IV U42992 ( .A(n32163), .Z(n30068) );
  NOR U42993 ( .A(n30069), .B(n30068), .Z(n30080) );
  IV U42994 ( .A(n30070), .Z(n30074) );
  NOR U42995 ( .A(n30072), .B(n30071), .Z(n30073) );
  IV U42996 ( .A(n30073), .Z(n30076) );
  NOR U42997 ( .A(n30074), .B(n30076), .Z(n35478) );
  IV U42998 ( .A(n30075), .Z(n30077) );
  NOR U42999 ( .A(n30077), .B(n30076), .Z(n35475) );
  NOR U43000 ( .A(n35478), .B(n35475), .Z(n30078) );
  IV U43001 ( .A(n30078), .Z(n30079) );
  NOR U43002 ( .A(n30080), .B(n30079), .Z(n30084) );
  NOR U43003 ( .A(n30082), .B(n30081), .Z(n32162) );
  NOR U43004 ( .A(n32162), .B(n32160), .Z(n30083) );
  XOR U43005 ( .A(n30084), .B(n30083), .Z(n32159) );
  XOR U43006 ( .A(n30085), .B(n32159), .Z(n30086) );
  IV U43007 ( .A(n30086), .Z(n33573) );
  XOR U43008 ( .A(n33571), .B(n33573), .Z(n33580) );
  XOR U43009 ( .A(n30087), .B(n33580), .Z(n32144) );
  XOR U43010 ( .A(n33582), .B(n32144), .Z(n33590) );
  XOR U43011 ( .A(n30088), .B(n33590), .Z(n32140) );
  IV U43012 ( .A(n30089), .Z(n30091) );
  NOR U43013 ( .A(n30091), .B(n30090), .Z(n32139) );
  IV U43014 ( .A(n30092), .Z(n30094) );
  NOR U43015 ( .A(n30094), .B(n30093), .Z(n33589) );
  NOR U43016 ( .A(n32139), .B(n33589), .Z(n30095) );
  XOR U43017 ( .A(n32140), .B(n30095), .Z(n33588) );
  XOR U43018 ( .A(n33586), .B(n33588), .Z(n33597) );
  XOR U43019 ( .A(n32132), .B(n33597), .Z(n32135) );
  XOR U43020 ( .A(n32134), .B(n32135), .Z(n32127) );
  XOR U43021 ( .A(n30096), .B(n32127), .Z(n30103) );
  NOR U43022 ( .A(n30097), .B(n30103), .Z(n30099) );
  IV U43023 ( .A(n30097), .Z(n30098) );
  NOR U43024 ( .A(n30098), .B(n32127), .Z(n32125) );
  NOR U43025 ( .A(n30099), .B(n32125), .Z(n30109) );
  IV U43026 ( .A(n30109), .Z(n32123) );
  NOR U43027 ( .A(n30100), .B(n32123), .Z(n36947) );
  IV U43028 ( .A(n30101), .Z(n30102) );
  NOR U43029 ( .A(n30102), .B(n30105), .Z(n33603) );
  IV U43030 ( .A(n30103), .Z(n30108) );
  IV U43031 ( .A(n30104), .Z(n30106) );
  NOR U43032 ( .A(n30106), .B(n30105), .Z(n30110) );
  IV U43033 ( .A(n30110), .Z(n30107) );
  NOR U43034 ( .A(n30108), .B(n30107), .Z(n35422) );
  NOR U43035 ( .A(n30110), .B(n30109), .Z(n30111) );
  NOR U43036 ( .A(n35422), .B(n30111), .Z(n33604) );
  XOR U43037 ( .A(n33603), .B(n33604), .Z(n30112) );
  NOR U43038 ( .A(n30113), .B(n30112), .Z(n30114) );
  NOR U43039 ( .A(n36947), .B(n30114), .Z(n30119) );
  IV U43040 ( .A(n30115), .Z(n30116) );
  NOR U43041 ( .A(n30117), .B(n30116), .Z(n30118) );
  IV U43042 ( .A(n30118), .Z(n32124) );
  XOR U43043 ( .A(n30119), .B(n32124), .Z(n32118) );
  XOR U43044 ( .A(n32117), .B(n32118), .Z(n32121) );
  XOR U43045 ( .A(n32120), .B(n32121), .Z(n33611) );
  XOR U43046 ( .A(n33609), .B(n33611), .Z(n35394) );
  NOR U43047 ( .A(n35398), .B(n30120), .Z(n32115) );
  IV U43048 ( .A(n30121), .Z(n30124) );
  IV U43049 ( .A(n30122), .Z(n30123) );
  NOR U43050 ( .A(n30124), .B(n30123), .Z(n33612) );
  NOR U43051 ( .A(n32115), .B(n33612), .Z(n30125) );
  XOR U43052 ( .A(n35394), .B(n30125), .Z(n30126) );
  NOR U43053 ( .A(n30127), .B(n30126), .Z(n30130) );
  IV U43054 ( .A(n30127), .Z(n30129) );
  XOR U43055 ( .A(n33612), .B(n35394), .Z(n30128) );
  NOR U43056 ( .A(n30129), .B(n30128), .Z(n35388) );
  NOR U43057 ( .A(n30130), .B(n35388), .Z(n32109) );
  XOR U43058 ( .A(n30131), .B(n32109), .Z(n32105) );
  XOR U43059 ( .A(n30132), .B(n32105), .Z(n30133) );
  IV U43060 ( .A(n30133), .Z(n32095) );
  XOR U43061 ( .A(n32094), .B(n32095), .Z(n32099) );
  XOR U43062 ( .A(n32097), .B(n32099), .Z(n32093) );
  XOR U43063 ( .A(n30134), .B(n32093), .Z(n33646) );
  XOR U43064 ( .A(n33636), .B(n33646), .Z(n33641) );
  IV U43065 ( .A(n30135), .Z(n30136) );
  NOR U43066 ( .A(n30136), .B(n30140), .Z(n33640) );
  NOR U43067 ( .A(n33640), .B(n30137), .Z(n30138) );
  XOR U43068 ( .A(n33641), .B(n30138), .Z(n33650) );
  IV U43069 ( .A(n30139), .Z(n30141) );
  NOR U43070 ( .A(n30141), .B(n30140), .Z(n33648) );
  XOR U43071 ( .A(n33650), .B(n33648), .Z(n33653) );
  XOR U43072 ( .A(n33651), .B(n33653), .Z(n33657) );
  XOR U43073 ( .A(n33655), .B(n33657), .Z(n33659) );
  XOR U43074 ( .A(n33658), .B(n33659), .Z(n33664) );
  NOR U43075 ( .A(n30148), .B(n33664), .Z(n36982) );
  IV U43076 ( .A(n30142), .Z(n30144) );
  IV U43077 ( .A(n30143), .Z(n30146) );
  NOR U43078 ( .A(n30144), .B(n30146), .Z(n33662) );
  XOR U43079 ( .A(n33664), .B(n33662), .Z(n33666) );
  IV U43080 ( .A(n30145), .Z(n30147) );
  NOR U43081 ( .A(n30147), .B(n30146), .Z(n30149) );
  IV U43082 ( .A(n30149), .Z(n33665) );
  XOR U43083 ( .A(n33666), .B(n33665), .Z(n30151) );
  NOR U43084 ( .A(n30149), .B(n30148), .Z(n30150) );
  NOR U43085 ( .A(n30151), .B(n30150), .Z(n30152) );
  NOR U43086 ( .A(n36982), .B(n30152), .Z(n30158) );
  XOR U43087 ( .A(n30153), .B(n30158), .Z(n30157) );
  IV U43088 ( .A(n30154), .Z(n30155) );
  NOR U43089 ( .A(n30155), .B(n30166), .Z(n30163) );
  IV U43090 ( .A(n30163), .Z(n30156) );
  NOR U43091 ( .A(n30157), .B(n30156), .Z(n35331) );
  IV U43092 ( .A(n30158), .Z(n35336) );
  IV U43093 ( .A(n30159), .Z(n30160) );
  NOR U43094 ( .A(n30161), .B(n30160), .Z(n32085) );
  NOR U43095 ( .A(n32085), .B(n35337), .Z(n30162) );
  XOR U43096 ( .A(n35336), .B(n30162), .Z(n35324) );
  NOR U43097 ( .A(n30163), .B(n35324), .Z(n30164) );
  NOR U43098 ( .A(n35331), .B(n30164), .Z(n33679) );
  IV U43099 ( .A(n30165), .Z(n30167) );
  NOR U43100 ( .A(n30167), .B(n30166), .Z(n30168) );
  IV U43101 ( .A(n30168), .Z(n33681) );
  XOR U43102 ( .A(n33679), .B(n33681), .Z(n32083) );
  XOR U43103 ( .A(n30169), .B(n32083), .Z(n32075) );
  XOR U43104 ( .A(n32079), .B(n32075), .Z(n30170) );
  NOR U43105 ( .A(n30171), .B(n30170), .Z(n35313) );
  IV U43106 ( .A(n30172), .Z(n35316) );
  NOR U43107 ( .A(n30173), .B(n35316), .Z(n32074) );
  NOR U43108 ( .A(n30174), .B(n32074), .Z(n30175) );
  XOR U43109 ( .A(n30175), .B(n32075), .Z(n30181) );
  IV U43110 ( .A(n30181), .Z(n30176) );
  NOR U43111 ( .A(n30177), .B(n30176), .Z(n30178) );
  NOR U43112 ( .A(n35313), .B(n30178), .Z(n33696) );
  XOR U43113 ( .A(n33695), .B(n33696), .Z(n30179) );
  NOR U43114 ( .A(n30180), .B(n30179), .Z(n30183) );
  IV U43115 ( .A(n30180), .Z(n30182) );
  NOR U43116 ( .A(n30182), .B(n30181), .Z(n35304) );
  NOR U43117 ( .A(n30183), .B(n35304), .Z(n32068) );
  NOR U43118 ( .A(n32070), .B(n30184), .Z(n33703) );
  IV U43119 ( .A(n30185), .Z(n30187) );
  NOR U43120 ( .A(n30187), .B(n30186), .Z(n32067) );
  NOR U43121 ( .A(n33703), .B(n32067), .Z(n30188) );
  XOR U43122 ( .A(n32068), .B(n30188), .Z(n30200) );
  IV U43123 ( .A(n30189), .Z(n30192) );
  IV U43124 ( .A(n30190), .Z(n30197) );
  XOR U43125 ( .A(n30194), .B(n30197), .Z(n30191) );
  NOR U43126 ( .A(n30192), .B(n30191), .Z(n30206) );
  IV U43127 ( .A(n30206), .Z(n30193) );
  NOR U43128 ( .A(n30200), .B(n30193), .Z(n37006) );
  XOR U43129 ( .A(n32067), .B(n32068), .Z(n32065) );
  IV U43130 ( .A(n30194), .Z(n30195) );
  NOR U43131 ( .A(n30195), .B(n30197), .Z(n33700) );
  IV U43132 ( .A(n30196), .Z(n30198) );
  NOR U43133 ( .A(n30198), .B(n30197), .Z(n32064) );
  NOR U43134 ( .A(n33700), .B(n32064), .Z(n30199) );
  NOR U43135 ( .A(n32065), .B(n30199), .Z(n30203) );
  IV U43136 ( .A(n30199), .Z(n30201) );
  NOR U43137 ( .A(n30201), .B(n30200), .Z(n30202) );
  NOR U43138 ( .A(n30203), .B(n30202), .Z(n30204) );
  IV U43139 ( .A(n30204), .Z(n30205) );
  NOR U43140 ( .A(n30206), .B(n30205), .Z(n30207) );
  NOR U43141 ( .A(n37006), .B(n30207), .Z(n33710) );
  IV U43142 ( .A(n30208), .Z(n30210) );
  NOR U43143 ( .A(n30210), .B(n30209), .Z(n33711) );
  XOR U43144 ( .A(n33710), .B(n33711), .Z(n32058) );
  IV U43145 ( .A(n30211), .Z(n33716) );
  NOR U43146 ( .A(n33716), .B(n30212), .Z(n32060) );
  NOR U43147 ( .A(n30214), .B(n30213), .Z(n32057) );
  NOR U43148 ( .A(n32060), .B(n32057), .Z(n30215) );
  XOR U43149 ( .A(n32058), .B(n30215), .Z(n33726) );
  XOR U43150 ( .A(n33722), .B(n33726), .Z(n32054) );
  XOR U43151 ( .A(n32053), .B(n32054), .Z(n33736) );
  XOR U43152 ( .A(n30216), .B(n33736), .Z(n32049) );
  XOR U43153 ( .A(n30217), .B(n32049), .Z(n32048) );
  XOR U43154 ( .A(n32046), .B(n32048), .Z(n32044) );
  XOR U43155 ( .A(n30218), .B(n32044), .Z(n32037) );
  XOR U43156 ( .A(n32035), .B(n32037), .Z(n32040) );
  IV U43157 ( .A(n30219), .Z(n30220) );
  NOR U43158 ( .A(n30221), .B(n30220), .Z(n32038) );
  XOR U43159 ( .A(n32040), .B(n32038), .Z(n35280) );
  XOR U43160 ( .A(n32034), .B(n35280), .Z(n30222) );
  IV U43161 ( .A(n30222), .Z(n33745) );
  XOR U43162 ( .A(n33744), .B(n33745), .Z(n32031) );
  XOR U43163 ( .A(n32030), .B(n32031), .Z(n33761) );
  XOR U43164 ( .A(n33760), .B(n33761), .Z(n30228) );
  IV U43165 ( .A(n30223), .Z(n30225) );
  IV U43166 ( .A(n30224), .Z(n30246) );
  NOR U43167 ( .A(n30225), .B(n30246), .Z(n30242) );
  IV U43168 ( .A(n30242), .Z(n30226) );
  NOR U43169 ( .A(n30228), .B(n30226), .Z(n35273) );
  NOR U43170 ( .A(n30227), .B(n30232), .Z(n30230) );
  IV U43171 ( .A(n30228), .Z(n30229) );
  NOR U43172 ( .A(n30230), .B(n30229), .Z(n30240) );
  IV U43173 ( .A(n30231), .Z(n30234) );
  NOR U43174 ( .A(n30232), .B(n33761), .Z(n30233) );
  IV U43175 ( .A(n30233), .Z(n30236) );
  NOR U43176 ( .A(n30234), .B(n30236), .Z(n35270) );
  IV U43177 ( .A(n30235), .Z(n30237) );
  NOR U43178 ( .A(n30237), .B(n30236), .Z(n37052) );
  NOR U43179 ( .A(n35270), .B(n37052), .Z(n30238) );
  IV U43180 ( .A(n30238), .Z(n30239) );
  NOR U43181 ( .A(n30240), .B(n30239), .Z(n30241) );
  NOR U43182 ( .A(n30242), .B(n30241), .Z(n30243) );
  NOR U43183 ( .A(n35273), .B(n30243), .Z(n30244) );
  IV U43184 ( .A(n30244), .Z(n33768) );
  IV U43185 ( .A(n30245), .Z(n30247) );
  NOR U43186 ( .A(n30247), .B(n30246), .Z(n33766) );
  XOR U43187 ( .A(n33768), .B(n33766), .Z(n32025) );
  XOR U43188 ( .A(n32024), .B(n32025), .Z(n32028) );
  XOR U43189 ( .A(n32027), .B(n32028), .Z(n32018) );
  IV U43190 ( .A(n30248), .Z(n30250) );
  NOR U43191 ( .A(n30250), .B(n30249), .Z(n30251) );
  IV U43192 ( .A(n30251), .Z(n32015) );
  XOR U43193 ( .A(n32018), .B(n32015), .Z(n30252) );
  XOR U43194 ( .A(n30253), .B(n30252), .Z(n33776) );
  XOR U43195 ( .A(n33774), .B(n33776), .Z(n33778) );
  XOR U43196 ( .A(n33777), .B(n33778), .Z(n35245) );
  XOR U43197 ( .A(n32013), .B(n35245), .Z(n35255) );
  XOR U43198 ( .A(n32007), .B(n35255), .Z(n32004) );
  IV U43199 ( .A(n30254), .Z(n30255) );
  NOR U43200 ( .A(n30256), .B(n30255), .Z(n32003) );
  IV U43201 ( .A(n30257), .Z(n30259) );
  NOR U43202 ( .A(n30259), .B(n30258), .Z(n32008) );
  NOR U43203 ( .A(n32003), .B(n32008), .Z(n30260) );
  XOR U43204 ( .A(n32004), .B(n30260), .Z(n33782) );
  XOR U43205 ( .A(n33781), .B(n33782), .Z(n31994) );
  XOR U43206 ( .A(n30261), .B(n31994), .Z(n31989) );
  XOR U43207 ( .A(n31988), .B(n31989), .Z(n30262) );
  NOR U43208 ( .A(n30263), .B(n30262), .Z(n35221) );
  NOR U43209 ( .A(n31986), .B(n35227), .Z(n30264) );
  NOR U43210 ( .A(n31988), .B(n30264), .Z(n30265) );
  XOR U43211 ( .A(n31989), .B(n30265), .Z(n30266) );
  NOR U43212 ( .A(n30267), .B(n30266), .Z(n30268) );
  NOR U43213 ( .A(n35221), .B(n30268), .Z(n31980) );
  IV U43214 ( .A(n30269), .Z(n30271) );
  NOR U43215 ( .A(n30271), .B(n30270), .Z(n30272) );
  IV U43216 ( .A(n30272), .Z(n31981) );
  XOR U43217 ( .A(n31980), .B(n31981), .Z(n31985) );
  XOR U43218 ( .A(n31983), .B(n31985), .Z(n30277) );
  IV U43219 ( .A(n30273), .Z(n30280) );
  IV U43220 ( .A(n30274), .Z(n30275) );
  NOR U43221 ( .A(n30280), .B(n30275), .Z(n30283) );
  IV U43222 ( .A(n30283), .Z(n30276) );
  NOR U43223 ( .A(n30277), .B(n30276), .Z(n37083) );
  IV U43224 ( .A(n30278), .Z(n30279) );
  NOR U43225 ( .A(n30280), .B(n30279), .Z(n31978) );
  NOR U43226 ( .A(n31983), .B(n31978), .Z(n30281) );
  XOR U43227 ( .A(n31985), .B(n30281), .Z(n30282) );
  NOR U43228 ( .A(n30283), .B(n30282), .Z(n30284) );
  NOR U43229 ( .A(n37083), .B(n30284), .Z(n31972) );
  XOR U43230 ( .A(n31974), .B(n31972), .Z(n31976) );
  XOR U43231 ( .A(n31975), .B(n31976), .Z(n33794) );
  IV U43232 ( .A(n30285), .Z(n30289) );
  XOR U43233 ( .A(n30287), .B(n30286), .Z(n30288) );
  NOR U43234 ( .A(n30289), .B(n30288), .Z(n33792) );
  XOR U43235 ( .A(n33794), .B(n33792), .Z(n33795) );
  XOR U43236 ( .A(n33796), .B(n33795), .Z(n31959) );
  IV U43237 ( .A(n30290), .Z(n30291) );
  NOR U43238 ( .A(n30291), .B(n30294), .Z(n31960) );
  NOR U43239 ( .A(n31966), .B(n30292), .Z(n30296) );
  IV U43240 ( .A(n30293), .Z(n30295) );
  NOR U43241 ( .A(n30295), .B(n30294), .Z(n31962) );
  NOR U43242 ( .A(n30296), .B(n31962), .Z(n30297) );
  IV U43243 ( .A(n30297), .Z(n30298) );
  NOR U43244 ( .A(n31960), .B(n30298), .Z(n30299) );
  XOR U43245 ( .A(n31959), .B(n30299), .Z(n31957) );
  IV U43246 ( .A(n30300), .Z(n30301) );
  NOR U43247 ( .A(n30302), .B(n30301), .Z(n31955) );
  IV U43248 ( .A(n30303), .Z(n30305) );
  NOR U43249 ( .A(n30305), .B(n30304), .Z(n31953) );
  NOR U43250 ( .A(n31955), .B(n31953), .Z(n30306) );
  XOR U43251 ( .A(n31957), .B(n30306), .Z(n30307) );
  NOR U43252 ( .A(n30308), .B(n30307), .Z(n30310) );
  IV U43253 ( .A(n30308), .Z(n30309) );
  XOR U43254 ( .A(n31957), .B(n31953), .Z(n31949) );
  NOR U43255 ( .A(n30309), .B(n31949), .Z(n35194) );
  NOR U43256 ( .A(n30310), .B(n35194), .Z(n31944) );
  NOR U43257 ( .A(n30311), .B(n31950), .Z(n30315) );
  IV U43258 ( .A(n30312), .Z(n30314) );
  IV U43259 ( .A(n30313), .Z(n30318) );
  NOR U43260 ( .A(n30314), .B(n30318), .Z(n31945) );
  NOR U43261 ( .A(n30315), .B(n31945), .Z(n30316) );
  XOR U43262 ( .A(n31944), .B(n30316), .Z(n31943) );
  IV U43263 ( .A(n30317), .Z(n30319) );
  NOR U43264 ( .A(n30319), .B(n30318), .Z(n31941) );
  XOR U43265 ( .A(n31943), .B(n31941), .Z(n35185) );
  XOR U43266 ( .A(n33802), .B(n35185), .Z(n33804) );
  IV U43267 ( .A(n30320), .Z(n30323) );
  IV U43268 ( .A(n30321), .Z(n30322) );
  NOR U43269 ( .A(n30323), .B(n30322), .Z(n33808) );
  NOR U43270 ( .A(n33803), .B(n33808), .Z(n30324) );
  XOR U43271 ( .A(n33804), .B(n30324), .Z(n33812) );
  XOR U43272 ( .A(n33811), .B(n33812), .Z(n30325) );
  NOR U43273 ( .A(n30326), .B(n30325), .Z(n37131) );
  IV U43274 ( .A(n30327), .Z(n30330) );
  IV U43275 ( .A(n30328), .Z(n30329) );
  NOR U43276 ( .A(n30330), .B(n30329), .Z(n31939) );
  NOR U43277 ( .A(n31939), .B(n33811), .Z(n30331) );
  XOR U43278 ( .A(n30331), .B(n33812), .Z(n30332) );
  NOR U43279 ( .A(n30333), .B(n30332), .Z(n30334) );
  NOR U43280 ( .A(n37131), .B(n30334), .Z(n33815) );
  IV U43281 ( .A(n30335), .Z(n33817) );
  XOR U43282 ( .A(n33815), .B(n33817), .Z(n33820) );
  XOR U43283 ( .A(n33819), .B(n33820), .Z(n33825) );
  XOR U43284 ( .A(n33822), .B(n33825), .Z(n33833) );
  XOR U43285 ( .A(n30336), .B(n33833), .Z(n33831) );
  XOR U43286 ( .A(n33830), .B(n33831), .Z(n31931) );
  IV U43287 ( .A(n30337), .Z(n30338) );
  NOR U43288 ( .A(n30339), .B(n30338), .Z(n31934) );
  IV U43289 ( .A(n30340), .Z(n30342) );
  NOR U43290 ( .A(n30342), .B(n30341), .Z(n31936) );
  NOR U43291 ( .A(n31934), .B(n31936), .Z(n30343) );
  XOR U43292 ( .A(n31931), .B(n30343), .Z(n31929) );
  XOR U43293 ( .A(n30344), .B(n31929), .Z(n30352) );
  IV U43294 ( .A(n30352), .Z(n35151) );
  NOR U43295 ( .A(n30345), .B(n35151), .Z(n31925) );
  XOR U43296 ( .A(n31932), .B(n31929), .Z(n30350) );
  IV U43297 ( .A(n30346), .Z(n30348) );
  NOR U43298 ( .A(n30348), .B(n30347), .Z(n30351) );
  IV U43299 ( .A(n30351), .Z(n30349) );
  NOR U43300 ( .A(n30350), .B(n30349), .Z(n33837) );
  NOR U43301 ( .A(n30352), .B(n30351), .Z(n30353) );
  NOR U43302 ( .A(n33837), .B(n30353), .Z(n30368) );
  NOR U43303 ( .A(n30354), .B(n30368), .Z(n30355) );
  NOR U43304 ( .A(n31925), .B(n30355), .Z(n30370) );
  IV U43305 ( .A(n30370), .Z(n30360) );
  IV U43306 ( .A(n30356), .Z(n30358) );
  NOR U43307 ( .A(n30358), .B(n30357), .Z(n30374) );
  IV U43308 ( .A(n30374), .Z(n30359) );
  NOR U43309 ( .A(n30360), .B(n30359), .Z(n38437) );
  IV U43310 ( .A(n30361), .Z(n30364) );
  XOR U43311 ( .A(n30362), .B(n30367), .Z(n30363) );
  NOR U43312 ( .A(n30364), .B(n30363), .Z(n33842) );
  IV U43313 ( .A(n30365), .Z(n30366) );
  NOR U43314 ( .A(n30367), .B(n30366), .Z(n30371) );
  IV U43315 ( .A(n30371), .Z(n35154) );
  IV U43316 ( .A(n30368), .Z(n30369) );
  NOR U43317 ( .A(n35154), .B(n30369), .Z(n33845) );
  NOR U43318 ( .A(n30371), .B(n30370), .Z(n30372) );
  NOR U43319 ( .A(n33845), .B(n30372), .Z(n33841) );
  XOR U43320 ( .A(n33842), .B(n33841), .Z(n30373) );
  NOR U43321 ( .A(n30374), .B(n30373), .Z(n30375) );
  NOR U43322 ( .A(n38437), .B(n30375), .Z(n31910) );
  XOR U43323 ( .A(n30376), .B(n31910), .Z(n31919) );
  XOR U43324 ( .A(n31920), .B(n31919), .Z(n31907) );
  IV U43325 ( .A(n30377), .Z(n31913) );
  NOR U43326 ( .A(n30378), .B(n31913), .Z(n30381) );
  IV U43327 ( .A(n30379), .Z(n30380) );
  NOR U43328 ( .A(n30380), .B(n31904), .Z(n37191) );
  NOR U43329 ( .A(n30381), .B(n37191), .Z(n30382) );
  XOR U43330 ( .A(n31907), .B(n30382), .Z(n31901) );
  IV U43331 ( .A(n30383), .Z(n31900) );
  NOR U43332 ( .A(n31903), .B(n31900), .Z(n30386) );
  IV U43333 ( .A(n30384), .Z(n30385) );
  NOR U43334 ( .A(n30385), .B(n31904), .Z(n35138) );
  NOR U43335 ( .A(n30386), .B(n35138), .Z(n30387) );
  XOR U43336 ( .A(n31901), .B(n30387), .Z(n31893) );
  NOR U43337 ( .A(n30389), .B(n30388), .Z(n31897) );
  NOR U43338 ( .A(n31897), .B(n31895), .Z(n30390) );
  XOR U43339 ( .A(n31893), .B(n30390), .Z(n31886) );
  IV U43340 ( .A(n30391), .Z(n30394) );
  IV U43341 ( .A(n30392), .Z(n30393) );
  NOR U43342 ( .A(n30394), .B(n30393), .Z(n31892) );
  IV U43343 ( .A(n30395), .Z(n31885) );
  NOR U43344 ( .A(n30396), .B(n31885), .Z(n30397) );
  NOR U43345 ( .A(n31892), .B(n30397), .Z(n30398) );
  XOR U43346 ( .A(n31886), .B(n30398), .Z(n31879) );
  NOR U43347 ( .A(n30400), .B(n30399), .Z(n31881) );
  NOR U43348 ( .A(n31881), .B(n31878), .Z(n30401) );
  XOR U43349 ( .A(n31879), .B(n30401), .Z(n35117) );
  XOR U43350 ( .A(n31876), .B(n35117), .Z(n31872) );
  NOR U43351 ( .A(n30402), .B(n31872), .Z(n35109) );
  IV U43352 ( .A(n30403), .Z(n35120) );
  NOR U43353 ( .A(n30404), .B(n35120), .Z(n31874) );
  NOR U43354 ( .A(n31876), .B(n31874), .Z(n30405) );
  XOR U43355 ( .A(n35117), .B(n30405), .Z(n31868) );
  NOR U43356 ( .A(n30406), .B(n31868), .Z(n30407) );
  NOR U43357 ( .A(n35109), .B(n30407), .Z(n31864) );
  IV U43358 ( .A(n30408), .Z(n30410) );
  NOR U43359 ( .A(n30410), .B(n30409), .Z(n31871) );
  IV U43360 ( .A(n30411), .Z(n30413) );
  IV U43361 ( .A(n30412), .Z(n30416) );
  NOR U43362 ( .A(n30413), .B(n30416), .Z(n31867) );
  NOR U43363 ( .A(n31871), .B(n31867), .Z(n30414) );
  XOR U43364 ( .A(n31864), .B(n30414), .Z(n31862) );
  IV U43365 ( .A(n30415), .Z(n30417) );
  NOR U43366 ( .A(n30417), .B(n30416), .Z(n31863) );
  IV U43367 ( .A(n30418), .Z(n30419) );
  NOR U43368 ( .A(n30419), .B(n30422), .Z(n31860) );
  NOR U43369 ( .A(n31863), .B(n31860), .Z(n30420) );
  XOR U43370 ( .A(n31862), .B(n30420), .Z(n31855) );
  IV U43371 ( .A(n30421), .Z(n30423) );
  NOR U43372 ( .A(n30423), .B(n30422), .Z(n30424) );
  IV U43373 ( .A(n30424), .Z(n31856) );
  XOR U43374 ( .A(n31855), .B(n31856), .Z(n33860) );
  IV U43375 ( .A(n33860), .Z(n30431) );
  IV U43376 ( .A(n30425), .Z(n30426) );
  NOR U43377 ( .A(n30429), .B(n30426), .Z(n33859) );
  IV U43378 ( .A(n30427), .Z(n30428) );
  NOR U43379 ( .A(n30429), .B(n30428), .Z(n31858) );
  NOR U43380 ( .A(n33859), .B(n31858), .Z(n30430) );
  XOR U43381 ( .A(n30431), .B(n30430), .Z(n33863) );
  XOR U43382 ( .A(n33862), .B(n33863), .Z(n31853) );
  NOR U43383 ( .A(n30433), .B(n31853), .Z(n30432) );
  IV U43384 ( .A(n30432), .Z(n35092) );
  NOR U43385 ( .A(n35092), .B(n35094), .Z(n33866) );
  NOR U43386 ( .A(n30433), .B(n35094), .Z(n30438) );
  IV U43387 ( .A(n30434), .Z(n30436) );
  NOR U43388 ( .A(n30436), .B(n30435), .Z(n30437) );
  IV U43389 ( .A(n30437), .Z(n31854) );
  XOR U43390 ( .A(n31854), .B(n31853), .Z(n31851) );
  NOR U43391 ( .A(n30438), .B(n31851), .Z(n30439) );
  NOR U43392 ( .A(n33866), .B(n30439), .Z(n31844) );
  NOR U43393 ( .A(n30440), .B(n35085), .Z(n31850) );
  IV U43394 ( .A(n35085), .Z(n30442) );
  IV U43395 ( .A(n30440), .Z(n30441) );
  NOR U43396 ( .A(n30442), .B(n30441), .Z(n30445) );
  IV U43397 ( .A(n30443), .Z(n30444) );
  NOR U43398 ( .A(n30445), .B(n30444), .Z(n30446) );
  NOR U43399 ( .A(n31850), .B(n30446), .Z(n31846) );
  XOR U43400 ( .A(n31844), .B(n31846), .Z(n35075) );
  XOR U43401 ( .A(n30447), .B(n35075), .Z(n31833) );
  XOR U43402 ( .A(n30448), .B(n31833), .Z(n31828) );
  XOR U43403 ( .A(n31825), .B(n31828), .Z(n33880) );
  XOR U43404 ( .A(n30449), .B(n33880), .Z(n31822) );
  XOR U43405 ( .A(n30450), .B(n31822), .Z(n31819) );
  XOR U43406 ( .A(n30451), .B(n31819), .Z(n31814) );
  XOR U43407 ( .A(n31815), .B(n31814), .Z(n30452) );
  NOR U43408 ( .A(n30453), .B(n30452), .Z(n30464) );
  IV U43409 ( .A(n30454), .Z(n30458) );
  XOR U43410 ( .A(n31816), .B(n31819), .Z(n30455) );
  NOR U43411 ( .A(n30456), .B(n30455), .Z(n30457) );
  IV U43412 ( .A(n30457), .Z(n30460) );
  NOR U43413 ( .A(n30458), .B(n30460), .Z(n35040) );
  IV U43414 ( .A(n30459), .Z(n30461) );
  NOR U43415 ( .A(n30461), .B(n30460), .Z(n31813) );
  NOR U43416 ( .A(n35040), .B(n31813), .Z(n30462) );
  IV U43417 ( .A(n30462), .Z(n30463) );
  NOR U43418 ( .A(n30464), .B(n30463), .Z(n31811) );
  IV U43419 ( .A(n30465), .Z(n30467) );
  IV U43420 ( .A(n30466), .Z(n30469) );
  NOR U43421 ( .A(n30467), .B(n30469), .Z(n33884) );
  IV U43422 ( .A(n30468), .Z(n30470) );
  NOR U43423 ( .A(n30470), .B(n30469), .Z(n31810) );
  NOR U43424 ( .A(n33884), .B(n31810), .Z(n30471) );
  XOR U43425 ( .A(n31811), .B(n30471), .Z(n31804) );
  XOR U43426 ( .A(n31803), .B(n31804), .Z(n31808) );
  XOR U43427 ( .A(n30472), .B(n31808), .Z(n35027) );
  IV U43428 ( .A(n30473), .Z(n30475) );
  NOR U43429 ( .A(n30475), .B(n30474), .Z(n31793) );
  XOR U43430 ( .A(n35027), .B(n31793), .Z(n33896) );
  XOR U43431 ( .A(n31794), .B(n33896), .Z(n33893) );
  XOR U43432 ( .A(n33891), .B(n33893), .Z(n30476) );
  NOR U43433 ( .A(n30477), .B(n30476), .Z(n41627) );
  IV U43434 ( .A(n30478), .Z(n30481) );
  IV U43435 ( .A(n30479), .Z(n30480) );
  NOR U43436 ( .A(n30481), .B(n30480), .Z(n33894) );
  XOR U43437 ( .A(n31794), .B(n33891), .Z(n30482) );
  NOR U43438 ( .A(n33894), .B(n30482), .Z(n30483) );
  XOR U43439 ( .A(n30483), .B(n33896), .Z(n31789) );
  NOR U43440 ( .A(n30484), .B(n31789), .Z(n30485) );
  NOR U43441 ( .A(n41627), .B(n30485), .Z(n31785) );
  IV U43442 ( .A(n30486), .Z(n30488) );
  IV U43443 ( .A(n30487), .Z(n30499) );
  NOR U43444 ( .A(n30488), .B(n30499), .Z(n31786) );
  IV U43445 ( .A(n30489), .Z(n30490) );
  NOR U43446 ( .A(n30491), .B(n30490), .Z(n31790) );
  NOR U43447 ( .A(n31786), .B(n31790), .Z(n30492) );
  XOR U43448 ( .A(n31785), .B(n30492), .Z(n37282) );
  NOR U43449 ( .A(n30503), .B(n30493), .Z(n30494) );
  IV U43450 ( .A(n30494), .Z(n30495) );
  NOR U43451 ( .A(n37282), .B(n30495), .Z(n33899) );
  IV U43452 ( .A(n30496), .Z(n30497) );
  NOR U43453 ( .A(n30503), .B(n30497), .Z(n37285) );
  IV U43454 ( .A(n30498), .Z(n30500) );
  NOR U43455 ( .A(n30500), .B(n30499), .Z(n30505) );
  IV U43456 ( .A(n30505), .Z(n31784) );
  XOR U43457 ( .A(n37282), .B(n31784), .Z(n30507) );
  IV U43458 ( .A(n30501), .Z(n30502) );
  NOR U43459 ( .A(n30503), .B(n30502), .Z(n30504) );
  IV U43460 ( .A(n30504), .Z(n37284) );
  NOR U43461 ( .A(n30505), .B(n37284), .Z(n30506) );
  NOR U43462 ( .A(n30507), .B(n30506), .Z(n33901) );
  IV U43463 ( .A(n33901), .Z(n30508) );
  NOR U43464 ( .A(n37285), .B(n30508), .Z(n30509) );
  NOR U43465 ( .A(n33899), .B(n30509), .Z(n31780) );
  XOR U43466 ( .A(n30510), .B(n31780), .Z(n33910) );
  XOR U43467 ( .A(n33908), .B(n33910), .Z(n35016) );
  IV U43468 ( .A(n30511), .Z(n31776) );
  NOR U43469 ( .A(n31776), .B(n30512), .Z(n30519) );
  IV U43470 ( .A(n30513), .Z(n30514) );
  NOR U43471 ( .A(n30514), .B(n30516), .Z(n35014) );
  IV U43472 ( .A(n30515), .Z(n30517) );
  NOR U43473 ( .A(n30517), .B(n30516), .Z(n37298) );
  NOR U43474 ( .A(n35014), .B(n37298), .Z(n31774) );
  IV U43475 ( .A(n31774), .Z(n30518) );
  NOR U43476 ( .A(n30519), .B(n30518), .Z(n30520) );
  XOR U43477 ( .A(n35016), .B(n30520), .Z(n31764) );
  IV U43478 ( .A(n30521), .Z(n31765) );
  NOR U43479 ( .A(n31765), .B(n30522), .Z(n30526) );
  IV U43480 ( .A(n30523), .Z(n30525) );
  NOR U43481 ( .A(n30525), .B(n30524), .Z(n31771) );
  NOR U43482 ( .A(n30526), .B(n31771), .Z(n30527) );
  XOR U43483 ( .A(n31764), .B(n30527), .Z(n31761) );
  XOR U43484 ( .A(n31760), .B(n31761), .Z(n31756) );
  XOR U43485 ( .A(n31755), .B(n31756), .Z(n34990) );
  IV U43486 ( .A(n30528), .Z(n34993) );
  NOR U43487 ( .A(n34993), .B(n30529), .Z(n31753) );
  IV U43488 ( .A(n30530), .Z(n30532) );
  NOR U43489 ( .A(n30532), .B(n30531), .Z(n31758) );
  NOR U43490 ( .A(n31753), .B(n31758), .Z(n30533) );
  XOR U43491 ( .A(n34990), .B(n30533), .Z(n30543) );
  IV U43492 ( .A(n30543), .Z(n30538) );
  IV U43493 ( .A(n30534), .Z(n30536) );
  NOR U43494 ( .A(n30536), .B(n30535), .Z(n30549) );
  IV U43495 ( .A(n30549), .Z(n30537) );
  NOR U43496 ( .A(n30538), .B(n30537), .Z(n34982) );
  IV U43497 ( .A(n30539), .Z(n30540) );
  NOR U43498 ( .A(n30540), .B(n30547), .Z(n30544) );
  IV U43499 ( .A(n30544), .Z(n30542) );
  XOR U43500 ( .A(n31758), .B(n34990), .Z(n30541) );
  NOR U43501 ( .A(n30542), .B(n30541), .Z(n33919) );
  NOR U43502 ( .A(n30544), .B(n30543), .Z(n30545) );
  NOR U43503 ( .A(n33919), .B(n30545), .Z(n31748) );
  IV U43504 ( .A(n30546), .Z(n30548) );
  NOR U43505 ( .A(n30548), .B(n30547), .Z(n31749) );
  XOR U43506 ( .A(n31748), .B(n31749), .Z(n33925) );
  NOR U43507 ( .A(n33925), .B(n30549), .Z(n30550) );
  NOR U43508 ( .A(n34982), .B(n30550), .Z(n31746) );
  XOR U43509 ( .A(n31747), .B(n31746), .Z(n30551) );
  XOR U43510 ( .A(n33926), .B(n30551), .Z(n34968) );
  XOR U43511 ( .A(n31744), .B(n34968), .Z(n34959) );
  NOR U43512 ( .A(n30552), .B(n34959), .Z(n34963) );
  NOR U43513 ( .A(n30558), .B(n34963), .Z(n33931) );
  IV U43514 ( .A(n33931), .Z(n30557) );
  IV U43515 ( .A(n30553), .Z(n34971) );
  NOR U43516 ( .A(n34971), .B(n30554), .Z(n31742) );
  NOR U43517 ( .A(n31742), .B(n31744), .Z(n30555) );
  XOR U43518 ( .A(n30555), .B(n34968), .Z(n30559) );
  NOR U43519 ( .A(n30556), .B(n30559), .Z(n33932) );
  NOR U43520 ( .A(n30557), .B(n33932), .Z(n30561) );
  IV U43521 ( .A(n30558), .Z(n34962) );
  NOR U43522 ( .A(n30559), .B(n34962), .Z(n30560) );
  NOR U43523 ( .A(n30561), .B(n30560), .Z(n33938) );
  IV U43524 ( .A(n30562), .Z(n33937) );
  NOR U43525 ( .A(n30563), .B(n33937), .Z(n30565) );
  NOR U43526 ( .A(n30565), .B(n30564), .Z(n30566) );
  XOR U43527 ( .A(n33938), .B(n30566), .Z(n33942) );
  NOR U43528 ( .A(n30568), .B(n30567), .Z(n33941) );
  NOR U43529 ( .A(n33941), .B(n33951), .Z(n30569) );
  XOR U43530 ( .A(n33942), .B(n30569), .Z(n33950) );
  XOR U43531 ( .A(n33948), .B(n33950), .Z(n30585) );
  NOR U43532 ( .A(n30570), .B(n30585), .Z(n34941) );
  IV U43533 ( .A(n30571), .Z(n31737) );
  NOR U43534 ( .A(n31737), .B(n30572), .Z(n30573) );
  NOR U43535 ( .A(n33948), .B(n30573), .Z(n30574) );
  XOR U43536 ( .A(n33950), .B(n30574), .Z(n30575) );
  NOR U43537 ( .A(n30576), .B(n30575), .Z(n30577) );
  NOR U43538 ( .A(n34941), .B(n30577), .Z(n30587) );
  IV U43539 ( .A(n30587), .Z(n31735) );
  IV U43540 ( .A(n30578), .Z(n30580) );
  IV U43541 ( .A(n30579), .Z(n30595) );
  NOR U43542 ( .A(n30580), .B(n30595), .Z(n30590) );
  IV U43543 ( .A(n30590), .Z(n30581) );
  NOR U43544 ( .A(n31735), .B(n30581), .Z(n37338) );
  IV U43545 ( .A(n30582), .Z(n30584) );
  NOR U43546 ( .A(n30584), .B(n30583), .Z(n30588) );
  IV U43547 ( .A(n30588), .Z(n30586) );
  NOR U43548 ( .A(n30586), .B(n30585), .Z(n37335) );
  NOR U43549 ( .A(n30588), .B(n30587), .Z(n30589) );
  NOR U43550 ( .A(n37335), .B(n30589), .Z(n33962) );
  NOR U43551 ( .A(n30590), .B(n33962), .Z(n30591) );
  NOR U43552 ( .A(n37338), .B(n30591), .Z(n30598) );
  IV U43553 ( .A(n30592), .Z(n30593) );
  NOR U43554 ( .A(n30601), .B(n30593), .Z(n33961) );
  IV U43555 ( .A(n30594), .Z(n30596) );
  NOR U43556 ( .A(n30596), .B(n30595), .Z(n31733) );
  NOR U43557 ( .A(n33961), .B(n31733), .Z(n30597) );
  XOR U43558 ( .A(n30598), .B(n30597), .Z(n33960) );
  IV U43559 ( .A(n30599), .Z(n30600) );
  NOR U43560 ( .A(n30601), .B(n30600), .Z(n33958) );
  XOR U43561 ( .A(n33960), .B(n33958), .Z(n31728) );
  XOR U43562 ( .A(n31727), .B(n31728), .Z(n31731) );
  XOR U43563 ( .A(n31730), .B(n31731), .Z(n33969) );
  IV U43564 ( .A(n30602), .Z(n30605) );
  IV U43565 ( .A(n30603), .Z(n30604) );
  NOR U43566 ( .A(n30605), .B(n30604), .Z(n33967) );
  XOR U43567 ( .A(n33969), .B(n33967), .Z(n33971) );
  XOR U43568 ( .A(n33970), .B(n33971), .Z(n33976) );
  IV U43569 ( .A(n30606), .Z(n30607) );
  NOR U43570 ( .A(n30610), .B(n30607), .Z(n33975) );
  IV U43571 ( .A(n30608), .Z(n30609) );
  NOR U43572 ( .A(n30610), .B(n30609), .Z(n31722) );
  NOR U43573 ( .A(n33975), .B(n31722), .Z(n30611) );
  XOR U43574 ( .A(n33976), .B(n30611), .Z(n31724) );
  IV U43575 ( .A(n30612), .Z(n30622) );
  IV U43576 ( .A(n30613), .Z(n30614) );
  NOR U43577 ( .A(n30622), .B(n30614), .Z(n33981) );
  IV U43578 ( .A(n30615), .Z(n30617) );
  NOR U43579 ( .A(n30617), .B(n30616), .Z(n31725) );
  NOR U43580 ( .A(n33981), .B(n31725), .Z(n30618) );
  XOR U43581 ( .A(n31724), .B(n30618), .Z(n33979) );
  NOR U43582 ( .A(n30619), .B(n31716), .Z(n30623) );
  IV U43583 ( .A(n30620), .Z(n30621) );
  NOR U43584 ( .A(n30622), .B(n30621), .Z(n33978) );
  NOR U43585 ( .A(n30623), .B(n33978), .Z(n30624) );
  XOR U43586 ( .A(n33979), .B(n30624), .Z(n30625) );
  IV U43587 ( .A(n30625), .Z(n31714) );
  XOR U43588 ( .A(n31712), .B(n31714), .Z(n31708) );
  IV U43589 ( .A(n30626), .Z(n30628) );
  NOR U43590 ( .A(n30628), .B(n30627), .Z(n31710) );
  IV U43591 ( .A(n30629), .Z(n30631) );
  NOR U43592 ( .A(n30631), .B(n30630), .Z(n31707) );
  NOR U43593 ( .A(n31710), .B(n31707), .Z(n30632) );
  XOR U43594 ( .A(n31708), .B(n30632), .Z(n31701) );
  XOR U43595 ( .A(n30633), .B(n31701), .Z(n33990) );
  XOR U43596 ( .A(n33989), .B(n33990), .Z(n31699) );
  XOR U43597 ( .A(n31698), .B(n31699), .Z(n31694) );
  XOR U43598 ( .A(n30634), .B(n31694), .Z(n31691) );
  IV U43599 ( .A(n30635), .Z(n30636) );
  NOR U43600 ( .A(n30640), .B(n30636), .Z(n30645) );
  IV U43601 ( .A(n30645), .Z(n30637) );
  NOR U43602 ( .A(n31691), .B(n30637), .Z(n34874) );
  IV U43603 ( .A(n30638), .Z(n30639) );
  NOR U43604 ( .A(n30640), .B(n30639), .Z(n31685) );
  IV U43605 ( .A(n30641), .Z(n30643) );
  NOR U43606 ( .A(n30643), .B(n30642), .Z(n31689) );
  NOR U43607 ( .A(n31685), .B(n31689), .Z(n30644) );
  XOR U43608 ( .A(n31691), .B(n30644), .Z(n30649) );
  NOR U43609 ( .A(n30645), .B(n30649), .Z(n30646) );
  NOR U43610 ( .A(n34874), .B(n30646), .Z(n30665) );
  NOR U43611 ( .A(n30647), .B(n30665), .Z(n30659) );
  IV U43612 ( .A(n30648), .Z(n30653) );
  IV U43613 ( .A(n30649), .Z(n30651) );
  NOR U43614 ( .A(n30651), .B(n30650), .Z(n30652) );
  IV U43615 ( .A(n30652), .Z(n30655) );
  NOR U43616 ( .A(n30653), .B(n30655), .Z(n34870) );
  IV U43617 ( .A(n30654), .Z(n30656) );
  NOR U43618 ( .A(n30656), .B(n30655), .Z(n34867) );
  NOR U43619 ( .A(n34870), .B(n34867), .Z(n30657) );
  IV U43620 ( .A(n30657), .Z(n30658) );
  NOR U43621 ( .A(n30659), .B(n30658), .Z(n30662) );
  IV U43622 ( .A(n30662), .Z(n37373) );
  NOR U43623 ( .A(n30660), .B(n37373), .Z(n37368) );
  NOR U43624 ( .A(n30661), .B(n30667), .Z(n30663) );
  NOR U43625 ( .A(n30663), .B(n30662), .Z(n30675) );
  IV U43626 ( .A(n30664), .Z(n30669) );
  IV U43627 ( .A(n30665), .Z(n30666) );
  NOR U43628 ( .A(n30667), .B(n30666), .Z(n30668) );
  IV U43629 ( .A(n30668), .Z(n30671) );
  NOR U43630 ( .A(n30669), .B(n30671), .Z(n37365) );
  IV U43631 ( .A(n30670), .Z(n30672) );
  NOR U43632 ( .A(n30672), .B(n30671), .Z(n34865) );
  NOR U43633 ( .A(n37365), .B(n34865), .Z(n30673) );
  IV U43634 ( .A(n30673), .Z(n30674) );
  NOR U43635 ( .A(n30675), .B(n30674), .Z(n30680) );
  NOR U43636 ( .A(n30676), .B(n30680), .Z(n30677) );
  NOR U43637 ( .A(n37368), .B(n30677), .Z(n30682) );
  IV U43638 ( .A(n30682), .Z(n34003) );
  NOR U43639 ( .A(n30678), .B(n34003), .Z(n34000) );
  NOR U43640 ( .A(n30679), .B(n34860), .Z(n30683) );
  IV U43641 ( .A(n30683), .Z(n30681) );
  IV U43642 ( .A(n30680), .Z(n34857) );
  NOR U43643 ( .A(n30681), .B(n34857), .Z(n33997) );
  NOR U43644 ( .A(n30683), .B(n30682), .Z(n30684) );
  NOR U43645 ( .A(n33997), .B(n30684), .Z(n31679) );
  NOR U43646 ( .A(n30685), .B(n31679), .Z(n30686) );
  NOR U43647 ( .A(n34000), .B(n30686), .Z(n30693) );
  IV U43648 ( .A(n30687), .Z(n30688) );
  NOR U43649 ( .A(n30688), .B(n30690), .Z(n31682) );
  IV U43650 ( .A(n30689), .Z(n30691) );
  NOR U43651 ( .A(n30691), .B(n30690), .Z(n31680) );
  NOR U43652 ( .A(n31682), .B(n31680), .Z(n30692) );
  XOR U43653 ( .A(n30693), .B(n30692), .Z(n31678) );
  IV U43654 ( .A(n30694), .Z(n30696) );
  NOR U43655 ( .A(n30696), .B(n30695), .Z(n30697) );
  IV U43656 ( .A(n30697), .Z(n31677) );
  XOR U43657 ( .A(n31678), .B(n31677), .Z(n31661) );
  IV U43658 ( .A(n30698), .Z(n30699) );
  NOR U43659 ( .A(n30702), .B(n30699), .Z(n31674) );
  IV U43660 ( .A(n30700), .Z(n30701) );
  NOR U43661 ( .A(n30702), .B(n30701), .Z(n31672) );
  NOR U43662 ( .A(n31674), .B(n31672), .Z(n30703) );
  XOR U43663 ( .A(n31661), .B(n30703), .Z(n31667) );
  XOR U43664 ( .A(n31666), .B(n31667), .Z(n31659) );
  IV U43665 ( .A(n30704), .Z(n30705) );
  NOR U43666 ( .A(n30705), .B(n30710), .Z(n30714) );
  IV U43667 ( .A(n30714), .Z(n30706) );
  NOR U43668 ( .A(n31659), .B(n30706), .Z(n37399) );
  IV U43669 ( .A(n30707), .Z(n31663) );
  NOR U43670 ( .A(n30708), .B(n31663), .Z(n30712) );
  IV U43671 ( .A(n30709), .Z(n30711) );
  NOR U43672 ( .A(n30711), .B(n30710), .Z(n31657) );
  NOR U43673 ( .A(n30712), .B(n31657), .Z(n30713) );
  XOR U43674 ( .A(n30713), .B(n31659), .Z(n30718) );
  NOR U43675 ( .A(n30714), .B(n30718), .Z(n30715) );
  NOR U43676 ( .A(n37399), .B(n30715), .Z(n30723) );
  IV U43677 ( .A(n30723), .Z(n30716) );
  NOR U43678 ( .A(n30717), .B(n30716), .Z(n37408) );
  IV U43679 ( .A(n30718), .Z(n30722) );
  IV U43680 ( .A(n30719), .Z(n30720) );
  NOR U43681 ( .A(n30728), .B(n30720), .Z(n30724) );
  IV U43682 ( .A(n30724), .Z(n30721) );
  NOR U43683 ( .A(n30722), .B(n30721), .Z(n37402) );
  NOR U43684 ( .A(n30724), .B(n30723), .Z(n30725) );
  NOR U43685 ( .A(n37402), .B(n30725), .Z(n31653) );
  IV U43686 ( .A(n30726), .Z(n30727) );
  NOR U43687 ( .A(n30728), .B(n30727), .Z(n31654) );
  XOR U43688 ( .A(n31653), .B(n31654), .Z(n30729) );
  NOR U43689 ( .A(n30730), .B(n30729), .Z(n30731) );
  NOR U43690 ( .A(n37408), .B(n30731), .Z(n30732) );
  IV U43691 ( .A(n30732), .Z(n31651) );
  XOR U43692 ( .A(n31650), .B(n31651), .Z(n31645) );
  XOR U43693 ( .A(n31643), .B(n31645), .Z(n40506) );
  NOR U43694 ( .A(n41469), .B(n40506), .Z(n30747) );
  NOR U43695 ( .A(n30733), .B(n31640), .Z(n30737) );
  IV U43696 ( .A(n30734), .Z(n30736) );
  NOR U43697 ( .A(n30736), .B(n30735), .Z(n41470) );
  NOR U43698 ( .A(n30737), .B(n41470), .Z(n30738) );
  IV U43699 ( .A(n30738), .Z(n30739) );
  XOR U43700 ( .A(n30739), .B(n40506), .Z(n31636) );
  IV U43701 ( .A(n30740), .Z(n30742) );
  IV U43702 ( .A(n30741), .Z(n30749) );
  NOR U43703 ( .A(n30742), .B(n30749), .Z(n30743) );
  IV U43704 ( .A(n30743), .Z(n31635) );
  XOR U43705 ( .A(n31636), .B(n31635), .Z(n30745) );
  NOR U43706 ( .A(n30743), .B(n41469), .Z(n30744) );
  NOR U43707 ( .A(n30745), .B(n30744), .Z(n30746) );
  NOR U43708 ( .A(n30747), .B(n30746), .Z(n34022) );
  IV U43709 ( .A(n30748), .Z(n30750) );
  NOR U43710 ( .A(n30750), .B(n30749), .Z(n34023) );
  XOR U43711 ( .A(n34022), .B(n34023), .Z(n31632) );
  IV U43712 ( .A(n30751), .Z(n30752) );
  NOR U43713 ( .A(n30755), .B(n30752), .Z(n34026) );
  IV U43714 ( .A(n30753), .Z(n30754) );
  NOR U43715 ( .A(n30755), .B(n30754), .Z(n31633) );
  NOR U43716 ( .A(n34026), .B(n31633), .Z(n30756) );
  XOR U43717 ( .A(n31632), .B(n30756), .Z(n47246) );
  IV U43718 ( .A(n30757), .Z(n30759) );
  NOR U43719 ( .A(n30759), .B(n30758), .Z(n47244) );
  XOR U43720 ( .A(n47246), .B(n47244), .Z(n47236) );
  XOR U43721 ( .A(n31619), .B(n47236), .Z(n34033) );
  XOR U43722 ( .A(n30760), .B(n34033), .Z(n30767) );
  XOR U43723 ( .A(n30761), .B(n30767), .Z(n30766) );
  IV U43724 ( .A(n30762), .Z(n30764) );
  NOR U43725 ( .A(n30764), .B(n30763), .Z(n30774) );
  IV U43726 ( .A(n30774), .Z(n30765) );
  NOR U43727 ( .A(n30766), .B(n30765), .Z(n34042) );
  IV U43728 ( .A(n30767), .Z(n34039) );
  IV U43729 ( .A(n30768), .Z(n30769) );
  NOR U43730 ( .A(n30770), .B(n30769), .Z(n34037) );
  NOR U43731 ( .A(n34037), .B(n31612), .Z(n30771) );
  IV U43732 ( .A(n30771), .Z(n30772) );
  NOR U43733 ( .A(n34030), .B(n30772), .Z(n30773) );
  XOR U43734 ( .A(n34039), .B(n30773), .Z(n37462) );
  NOR U43735 ( .A(n30774), .B(n37462), .Z(n30775) );
  NOR U43736 ( .A(n34042), .B(n30775), .Z(n30776) );
  IV U43737 ( .A(n30776), .Z(n34044) );
  XOR U43738 ( .A(n34045), .B(n34044), .Z(n34047) );
  NOR U43739 ( .A(n30777), .B(n34054), .Z(n30780) );
  IV U43740 ( .A(n30778), .Z(n34059) );
  NOR U43741 ( .A(n34061), .B(n34059), .Z(n30779) );
  NOR U43742 ( .A(n30780), .B(n30779), .Z(n30781) );
  XOR U43743 ( .A(n34047), .B(n30781), .Z(n31608) );
  IV U43744 ( .A(n30782), .Z(n30784) );
  NOR U43745 ( .A(n30784), .B(n30783), .Z(n31606) );
  XOR U43746 ( .A(n31608), .B(n31606), .Z(n31610) );
  XOR U43747 ( .A(n31609), .B(n31610), .Z(n31602) );
  NOR U43748 ( .A(n30785), .B(n31602), .Z(n37475) );
  IV U43749 ( .A(n30786), .Z(n30791) );
  IV U43750 ( .A(n30787), .Z(n30788) );
  NOR U43751 ( .A(n30791), .B(n30788), .Z(n31601) );
  XOR U43752 ( .A(n31601), .B(n31602), .Z(n31605) );
  IV U43753 ( .A(n30789), .Z(n30790) );
  NOR U43754 ( .A(n30791), .B(n30790), .Z(n30792) );
  IV U43755 ( .A(n30792), .Z(n31604) );
  XOR U43756 ( .A(n31605), .B(n31604), .Z(n30796) );
  NOR U43757 ( .A(n30793), .B(n30796), .Z(n30794) );
  NOR U43758 ( .A(n37475), .B(n30794), .Z(n31596) );
  XOR U43759 ( .A(n31597), .B(n31596), .Z(n30795) );
  NOR U43760 ( .A(n30797), .B(n30795), .Z(n30800) );
  IV U43761 ( .A(n30796), .Z(n30799) );
  IV U43762 ( .A(n30797), .Z(n30798) );
  NOR U43763 ( .A(n30799), .B(n30798), .Z(n34799) );
  NOR U43764 ( .A(n30800), .B(n34799), .Z(n31589) );
  IV U43765 ( .A(n30801), .Z(n31590) );
  NOR U43766 ( .A(n30802), .B(n31590), .Z(n30804) );
  NOR U43767 ( .A(n30803), .B(n34789), .Z(n34066) );
  NOR U43768 ( .A(n30804), .B(n34066), .Z(n30805) );
  XOR U43769 ( .A(n31589), .B(n30805), .Z(n34071) );
  IV U43770 ( .A(n30806), .Z(n30808) );
  NOR U43771 ( .A(n30808), .B(n30807), .Z(n31586) );
  XOR U43772 ( .A(n34071), .B(n31586), .Z(n30809) );
  XOR U43773 ( .A(n30810), .B(n30809), .Z(n34074) );
  XOR U43774 ( .A(n34072), .B(n34074), .Z(n34080) );
  IV U43775 ( .A(n30811), .Z(n30812) );
  NOR U43776 ( .A(n30812), .B(n30814), .Z(n34075) );
  IV U43777 ( .A(n30813), .Z(n30815) );
  NOR U43778 ( .A(n30815), .B(n30814), .Z(n34081) );
  NOR U43779 ( .A(n34075), .B(n34081), .Z(n30816) );
  XOR U43780 ( .A(n34080), .B(n30816), .Z(n34085) );
  IV U43781 ( .A(n30817), .Z(n30818) );
  NOR U43782 ( .A(n30819), .B(n30818), .Z(n34084) );
  IV U43783 ( .A(n30820), .Z(n30822) );
  NOR U43784 ( .A(n30822), .B(n30821), .Z(n34079) );
  NOR U43785 ( .A(n34084), .B(n34079), .Z(n30823) );
  XOR U43786 ( .A(n34085), .B(n30823), .Z(n31581) );
  XOR U43787 ( .A(n31582), .B(n31581), .Z(n34087) );
  XOR U43788 ( .A(n34088), .B(n34087), .Z(n34091) );
  IV U43789 ( .A(n30824), .Z(n30825) );
  NOR U43790 ( .A(n30826), .B(n30825), .Z(n34089) );
  XOR U43791 ( .A(n34091), .B(n34089), .Z(n31575) );
  NOR U43792 ( .A(n30827), .B(n31578), .Z(n30830) );
  IV U43793 ( .A(n30838), .Z(n30829) );
  IV U43794 ( .A(n30828), .Z(n30842) );
  NOR U43795 ( .A(n30829), .B(n30842), .Z(n31574) );
  NOR U43796 ( .A(n30830), .B(n31574), .Z(n30831) );
  XOR U43797 ( .A(n31575), .B(n30831), .Z(n30845) );
  IV U43798 ( .A(n30845), .Z(n30836) );
  IV U43799 ( .A(n30832), .Z(n30834) );
  NOR U43800 ( .A(n30834), .B(n30833), .Z(n30849) );
  IV U43801 ( .A(n30849), .Z(n30835) );
  NOR U43802 ( .A(n30836), .B(n30835), .Z(n37519) );
  IV U43803 ( .A(n30837), .Z(n30840) );
  XOR U43804 ( .A(n30838), .B(n30842), .Z(n30839) );
  NOR U43805 ( .A(n30840), .B(n30839), .Z(n31570) );
  IV U43806 ( .A(n30841), .Z(n30843) );
  NOR U43807 ( .A(n30843), .B(n30842), .Z(n30846) );
  IV U43808 ( .A(n30846), .Z(n30844) );
  NOR U43809 ( .A(n30844), .B(n31575), .Z(n34754) );
  NOR U43810 ( .A(n30846), .B(n30845), .Z(n30847) );
  NOR U43811 ( .A(n34754), .B(n30847), .Z(n31571) );
  XOR U43812 ( .A(n31570), .B(n31571), .Z(n30848) );
  NOR U43813 ( .A(n30849), .B(n30848), .Z(n30850) );
  NOR U43814 ( .A(n37519), .B(n30850), .Z(n30856) );
  IV U43815 ( .A(n30851), .Z(n30852) );
  NOR U43816 ( .A(n30853), .B(n30852), .Z(n31566) );
  XOR U43817 ( .A(n30856), .B(n31566), .Z(n30854) );
  NOR U43818 ( .A(n30855), .B(n30854), .Z(n31564) );
  IV U43819 ( .A(n30855), .Z(n30857) );
  IV U43820 ( .A(n30856), .Z(n31568) );
  NOR U43821 ( .A(n30857), .B(n31568), .Z(n34748) );
  NOR U43822 ( .A(n31564), .B(n34748), .Z(n30862) );
  IV U43823 ( .A(n30862), .Z(n34736) );
  NOR U43824 ( .A(n30867), .B(n34736), .Z(n34732) );
  NOR U43825 ( .A(n30858), .B(n34742), .Z(n31563) );
  IV U43826 ( .A(n30859), .Z(n30861) );
  NOR U43827 ( .A(n30861), .B(n30860), .Z(n34735) );
  NOR U43828 ( .A(n31563), .B(n34735), .Z(n30863) );
  XOR U43829 ( .A(n30863), .B(n30862), .Z(n31559) );
  IV U43830 ( .A(n30864), .Z(n30866) );
  NOR U43831 ( .A(n30866), .B(n30865), .Z(n30868) );
  IV U43832 ( .A(n30868), .Z(n31558) );
  XOR U43833 ( .A(n31559), .B(n31558), .Z(n30870) );
  NOR U43834 ( .A(n30868), .B(n30867), .Z(n30869) );
  NOR U43835 ( .A(n30870), .B(n30869), .Z(n30871) );
  NOR U43836 ( .A(n34732), .B(n30871), .Z(n30872) );
  IV U43837 ( .A(n30872), .Z(n31561) );
  XOR U43838 ( .A(n31560), .B(n31561), .Z(n31553) );
  XOR U43839 ( .A(n31552), .B(n31553), .Z(n31557) );
  XOR U43840 ( .A(n31555), .B(n31557), .Z(n34109) );
  IV U43841 ( .A(n30873), .Z(n30875) );
  IV U43842 ( .A(n30874), .Z(n30884) );
  NOR U43843 ( .A(n30875), .B(n30884), .Z(n30888) );
  IV U43844 ( .A(n30888), .Z(n30876) );
  NOR U43845 ( .A(n34109), .B(n30876), .Z(n34721) );
  IV U43846 ( .A(n30877), .Z(n30878) );
  NOR U43847 ( .A(n30878), .B(n30880), .Z(n31550) );
  IV U43848 ( .A(n30879), .Z(n30881) );
  NOR U43849 ( .A(n30881), .B(n30880), .Z(n34108) );
  NOR U43850 ( .A(n31550), .B(n34108), .Z(n30882) );
  IV U43851 ( .A(n30882), .Z(n30886) );
  IV U43852 ( .A(n30883), .Z(n30885) );
  NOR U43853 ( .A(n30885), .B(n30884), .Z(n34106) );
  NOR U43854 ( .A(n30886), .B(n34106), .Z(n30887) );
  XOR U43855 ( .A(n30887), .B(n34109), .Z(n31541) );
  NOR U43856 ( .A(n30888), .B(n31541), .Z(n30889) );
  NOR U43857 ( .A(n34721), .B(n30889), .Z(n30890) );
  IV U43858 ( .A(n30890), .Z(n50781) );
  XOR U43859 ( .A(n30891), .B(n50781), .Z(n31537) );
  NOR U43860 ( .A(n30892), .B(n34115), .Z(n30896) );
  IV U43861 ( .A(n30893), .Z(n30895) );
  NOR U43862 ( .A(n30895), .B(n30894), .Z(n31538) );
  NOR U43863 ( .A(n30896), .B(n31538), .Z(n30897) );
  XOR U43864 ( .A(n31537), .B(n30897), .Z(n34120) );
  XOR U43865 ( .A(n34118), .B(n34120), .Z(n34126) );
  XOR U43866 ( .A(n34125), .B(n34126), .Z(n34129) );
  XOR U43867 ( .A(n34128), .B(n34129), .Z(n34133) );
  XOR U43868 ( .A(n34132), .B(n34133), .Z(n34137) );
  XOR U43869 ( .A(n34135), .B(n34137), .Z(n31533) );
  XOR U43870 ( .A(n31532), .B(n31533), .Z(n30902) );
  IV U43871 ( .A(n30898), .Z(n30900) );
  IV U43872 ( .A(n30899), .Z(n30904) );
  NOR U43873 ( .A(n30900), .B(n30904), .Z(n30913) );
  IV U43874 ( .A(n30913), .Z(n30901) );
  NOR U43875 ( .A(n30902), .B(n30901), .Z(n34699) );
  IV U43876 ( .A(n30903), .Z(n30905) );
  NOR U43877 ( .A(n30905), .B(n30904), .Z(n31528) );
  IV U43878 ( .A(n30906), .Z(n30908) );
  NOR U43879 ( .A(n30908), .B(n30907), .Z(n31530) );
  NOR U43880 ( .A(n31530), .B(n31532), .Z(n30909) );
  IV U43881 ( .A(n30909), .Z(n30910) );
  NOR U43882 ( .A(n31528), .B(n30910), .Z(n30911) );
  XOR U43883 ( .A(n30911), .B(n31533), .Z(n30912) );
  NOR U43884 ( .A(n30913), .B(n30912), .Z(n30914) );
  NOR U43885 ( .A(n34699), .B(n30914), .Z(n31524) );
  IV U43886 ( .A(n30915), .Z(n30916) );
  NOR U43887 ( .A(n30919), .B(n30916), .Z(n31525) );
  XOR U43888 ( .A(n31524), .B(n31525), .Z(n34141) );
  IV U43889 ( .A(n30917), .Z(n30918) );
  NOR U43890 ( .A(n30919), .B(n30918), .Z(n34142) );
  IV U43891 ( .A(n30920), .Z(n30922) );
  IV U43892 ( .A(n30921), .Z(n30925) );
  NOR U43893 ( .A(n30922), .B(n30925), .Z(n34149) );
  NOR U43894 ( .A(n34142), .B(n34149), .Z(n30923) );
  XOR U43895 ( .A(n34141), .B(n30923), .Z(n34148) );
  IV U43896 ( .A(n30924), .Z(n30926) );
  NOR U43897 ( .A(n30926), .B(n30925), .Z(n34146) );
  XOR U43898 ( .A(n34148), .B(n34146), .Z(n31516) );
  XOR U43899 ( .A(n30927), .B(n31516), .Z(n31513) );
  IV U43900 ( .A(n30928), .Z(n30929) );
  NOR U43901 ( .A(n30930), .B(n30929), .Z(n30931) );
  IV U43902 ( .A(n30931), .Z(n31508) );
  XOR U43903 ( .A(n31513), .B(n31508), .Z(n30932) );
  XOR U43904 ( .A(n30933), .B(n30932), .Z(n31507) );
  XOR U43905 ( .A(n31505), .B(n31507), .Z(n30934) );
  XOR U43906 ( .A(n30935), .B(n30934), .Z(n31499) );
  XOR U43907 ( .A(n31498), .B(n31499), .Z(n31495) );
  IV U43908 ( .A(n30936), .Z(n30937) );
  NOR U43909 ( .A(n30938), .B(n30937), .Z(n34154) );
  IV U43910 ( .A(n30939), .Z(n30942) );
  IV U43911 ( .A(n30940), .Z(n30941) );
  NOR U43912 ( .A(n30942), .B(n30941), .Z(n31496) );
  NOR U43913 ( .A(n34154), .B(n31496), .Z(n30943) );
  XOR U43914 ( .A(n31495), .B(n30943), .Z(n34678) );
  XOR U43915 ( .A(n34157), .B(n34678), .Z(n34667) );
  NOR U43916 ( .A(n30944), .B(n34667), .Z(n34161) );
  IV U43917 ( .A(n30945), .Z(n34681) );
  NOR U43918 ( .A(n30946), .B(n34681), .Z(n31493) );
  NOR U43919 ( .A(n34157), .B(n31493), .Z(n30947) );
  XOR U43920 ( .A(n30947), .B(n34678), .Z(n30953) );
  NOR U43921 ( .A(n30948), .B(n30953), .Z(n30949) );
  NOR U43922 ( .A(n34161), .B(n30949), .Z(n30955) );
  IV U43923 ( .A(n30955), .Z(n31491) );
  NOR U43924 ( .A(n30950), .B(n31491), .Z(n34648) );
  IV U43925 ( .A(n30951), .Z(n34659) );
  NOR U43926 ( .A(n30952), .B(n34659), .Z(n30956) );
  IV U43927 ( .A(n30956), .Z(n30954) );
  IV U43928 ( .A(n30953), .Z(n34656) );
  NOR U43929 ( .A(n30954), .B(n34656), .Z(n34162) );
  NOR U43930 ( .A(n30956), .B(n30955), .Z(n30957) );
  NOR U43931 ( .A(n34162), .B(n30957), .Z(n31486) );
  NOR U43932 ( .A(n30958), .B(n31486), .Z(n30959) );
  NOR U43933 ( .A(n34648), .B(n30959), .Z(n30968) );
  IV U43934 ( .A(n30960), .Z(n30961) );
  NOR U43935 ( .A(n30961), .B(n30963), .Z(n31490) );
  IV U43936 ( .A(n30962), .Z(n30966) );
  XOR U43937 ( .A(n30964), .B(n30963), .Z(n30965) );
  NOR U43938 ( .A(n30966), .B(n30965), .Z(n31487) );
  NOR U43939 ( .A(n31490), .B(n31487), .Z(n30967) );
  XOR U43940 ( .A(n30968), .B(n30967), .Z(n31485) );
  XOR U43941 ( .A(n31484), .B(n31485), .Z(n31478) );
  IV U43942 ( .A(n30969), .Z(n30970) );
  NOR U43943 ( .A(n30970), .B(n30972), .Z(n31481) );
  IV U43944 ( .A(n30971), .Z(n30973) );
  NOR U43945 ( .A(n30973), .B(n30972), .Z(n31479) );
  NOR U43946 ( .A(n31481), .B(n31479), .Z(n30974) );
  NOR U43947 ( .A(n31478), .B(n30974), .Z(n30984) );
  IV U43948 ( .A(n30974), .Z(n30982) );
  NOR U43949 ( .A(n30977), .B(n31485), .Z(n30975) );
  IV U43950 ( .A(n30975), .Z(n34636) );
  NOR U43951 ( .A(n30976), .B(n34636), .Z(n34163) );
  NOR U43952 ( .A(n30977), .B(n30976), .Z(n30978) );
  NOR U43953 ( .A(n30978), .B(n31478), .Z(n30979) );
  NOR U43954 ( .A(n34163), .B(n30979), .Z(n30980) );
  IV U43955 ( .A(n30980), .Z(n30981) );
  NOR U43956 ( .A(n30982), .B(n30981), .Z(n30983) );
  NOR U43957 ( .A(n30984), .B(n30983), .Z(n31477) );
  XOR U43958 ( .A(n31475), .B(n31477), .Z(n31466) );
  XOR U43959 ( .A(n30985), .B(n31466), .Z(n30991) );
  XOR U43960 ( .A(n30986), .B(n30991), .Z(n30994) );
  NOR U43961 ( .A(n30987), .B(n30994), .Z(n38049) );
  IV U43962 ( .A(n30988), .Z(n30989) );
  NOR U43963 ( .A(n30990), .B(n30989), .Z(n30996) );
  IV U43964 ( .A(n30996), .Z(n30993) );
  IV U43965 ( .A(n30991), .Z(n31464) );
  XOR U43966 ( .A(n31464), .B(n31462), .Z(n30992) );
  NOR U43967 ( .A(n30993), .B(n30992), .Z(n34622) );
  IV U43968 ( .A(n30994), .Z(n30995) );
  NOR U43969 ( .A(n30996), .B(n30995), .Z(n30997) );
  NOR U43970 ( .A(n34622), .B(n30997), .Z(n30998) );
  NOR U43971 ( .A(n30999), .B(n30998), .Z(n31000) );
  NOR U43972 ( .A(n38049), .B(n31000), .Z(n31001) );
  IV U43973 ( .A(n31001), .Z(n31458) );
  NOR U43974 ( .A(n31002), .B(n31458), .Z(n34617) );
  IV U43975 ( .A(n31003), .Z(n31004) );
  NOR U43976 ( .A(n31004), .B(n31006), .Z(n31454) );
  IV U43977 ( .A(n31005), .Z(n31007) );
  NOR U43978 ( .A(n31007), .B(n31006), .Z(n31457) );
  NOR U43979 ( .A(n31454), .B(n31457), .Z(n31008) );
  XOR U43980 ( .A(n31008), .B(n31458), .Z(n34166) );
  NOR U43981 ( .A(n31009), .B(n34166), .Z(n31010) );
  NOR U43982 ( .A(n34617), .B(n31010), .Z(n34175) );
  IV U43983 ( .A(n31011), .Z(n34167) );
  NOR U43984 ( .A(n31012), .B(n34167), .Z(n31014) );
  NOR U43985 ( .A(n34179), .B(n34177), .Z(n31013) );
  NOR U43986 ( .A(n31014), .B(n31013), .Z(n31015) );
  XOR U43987 ( .A(n34175), .B(n31015), .Z(n31447) );
  XOR U43988 ( .A(n31016), .B(n31447), .Z(n31440) );
  XOR U43989 ( .A(n31442), .B(n31440), .Z(n31017) );
  NOR U43990 ( .A(n31022), .B(n31017), .Z(n31018) );
  IV U43991 ( .A(n31018), .Z(n31019) );
  NOR U43992 ( .A(n31020), .B(n31019), .Z(n31021) );
  IV U43993 ( .A(n31021), .Z(n34188) );
  NOR U43994 ( .A(n31026), .B(n34188), .Z(n31433) );
  NOR U43995 ( .A(n31023), .B(n31022), .Z(n31024) );
  XOR U43996 ( .A(n31024), .B(n31440), .Z(n31034) );
  IV U43997 ( .A(n31034), .Z(n31028) );
  NOR U43998 ( .A(n31026), .B(n31025), .Z(n31027) );
  NOR U43999 ( .A(n31028), .B(n31027), .Z(n31029) );
  NOR U44000 ( .A(n31433), .B(n31029), .Z(n31035) );
  IV U44001 ( .A(n31035), .Z(n31046) );
  NOR U44002 ( .A(n31030), .B(n31046), .Z(n37659) );
  NOR U44003 ( .A(n31032), .B(n31031), .Z(n31036) );
  IV U44004 ( .A(n31036), .Z(n31033) );
  NOR U44005 ( .A(n31034), .B(n31033), .Z(n34185) );
  NOR U44006 ( .A(n31036), .B(n31035), .Z(n31037) );
  NOR U44007 ( .A(n34185), .B(n31037), .Z(n31038) );
  NOR U44008 ( .A(n31039), .B(n31038), .Z(n31040) );
  NOR U44009 ( .A(n37659), .B(n31040), .Z(n31048) );
  IV U44010 ( .A(n31048), .Z(n31041) );
  NOR U44011 ( .A(n31042), .B(n31041), .Z(n34584) );
  IV U44012 ( .A(n31043), .Z(n31045) );
  NOR U44013 ( .A(n31045), .B(n31044), .Z(n31049) );
  IV U44014 ( .A(n31049), .Z(n31047) );
  NOR U44015 ( .A(n31047), .B(n31046), .Z(n37662) );
  NOR U44016 ( .A(n31049), .B(n31048), .Z(n31050) );
  NOR U44017 ( .A(n37662), .B(n31050), .Z(n31054) );
  NOR U44018 ( .A(n31051), .B(n31054), .Z(n31052) );
  NOR U44019 ( .A(n34584), .B(n31052), .Z(n31053) );
  NOR U44020 ( .A(n31055), .B(n31053), .Z(n31057) );
  IV U44021 ( .A(n31054), .Z(n31430) );
  IV U44022 ( .A(n31055), .Z(n31056) );
  NOR U44023 ( .A(n31430), .B(n31056), .Z(n37665) );
  NOR U44024 ( .A(n31057), .B(n37665), .Z(n31423) );
  XOR U44025 ( .A(n31058), .B(n31423), .Z(n31416) );
  XOR U44026 ( .A(n31422), .B(n31416), .Z(n34571) );
  XOR U44027 ( .A(n31059), .B(n34571), .Z(n31060) );
  NOR U44028 ( .A(n31061), .B(n31060), .Z(n34563) );
  IV U44029 ( .A(n31062), .Z(n31064) );
  NOR U44030 ( .A(n31064), .B(n31063), .Z(n34559) );
  NOR U44031 ( .A(n31065), .B(n34559), .Z(n31066) );
  IV U44032 ( .A(n31066), .Z(n31067) );
  NOR U44033 ( .A(n34569), .B(n31067), .Z(n31068) );
  XOR U44034 ( .A(n34571), .B(n31068), .Z(n31069) );
  NOR U44035 ( .A(n31070), .B(n31069), .Z(n31071) );
  NOR U44036 ( .A(n34563), .B(n31071), .Z(n31409) );
  XOR U44037 ( .A(n31411), .B(n31409), .Z(n37681) );
  IV U44038 ( .A(n31072), .Z(n31083) );
  IV U44039 ( .A(n31073), .Z(n31074) );
  NOR U44040 ( .A(n31083), .B(n31074), .Z(n31405) );
  IV U44041 ( .A(n31075), .Z(n31077) );
  NOR U44042 ( .A(n31077), .B(n31076), .Z(n31407) );
  NOR U44043 ( .A(n31405), .B(n31407), .Z(n31078) );
  XOR U44044 ( .A(n37681), .B(n31078), .Z(n31400) );
  IV U44045 ( .A(n31079), .Z(n31080) );
  NOR U44046 ( .A(n31080), .B(n31086), .Z(n31401) );
  IV U44047 ( .A(n31081), .Z(n31082) );
  NOR U44048 ( .A(n31083), .B(n31082), .Z(n31403) );
  NOR U44049 ( .A(n31401), .B(n31403), .Z(n31084) );
  XOR U44050 ( .A(n31400), .B(n31084), .Z(n34197) );
  IV U44051 ( .A(n31085), .Z(n31087) );
  NOR U44052 ( .A(n31087), .B(n31086), .Z(n34195) );
  XOR U44053 ( .A(n34197), .B(n34195), .Z(n34211) );
  IV U44054 ( .A(n31088), .Z(n31090) );
  NOR U44055 ( .A(n31090), .B(n31089), .Z(n31091) );
  IV U44056 ( .A(n31091), .Z(n34198) );
  XOR U44057 ( .A(n34211), .B(n34198), .Z(n31396) );
  IV U44058 ( .A(n31092), .Z(n34203) );
  NOR U44059 ( .A(n34203), .B(n31093), .Z(n34210) );
  IV U44060 ( .A(n31094), .Z(n31096) );
  NOR U44061 ( .A(n31096), .B(n31095), .Z(n31395) );
  NOR U44062 ( .A(n34210), .B(n31395), .Z(n31097) );
  XOR U44063 ( .A(n31396), .B(n31097), .Z(n40873) );
  IV U44064 ( .A(n31098), .Z(n31100) );
  IV U44065 ( .A(n31099), .Z(n31104) );
  NOR U44066 ( .A(n31100), .B(n31104), .Z(n31386) );
  IV U44067 ( .A(n31386), .Z(n31101) );
  NOR U44068 ( .A(n40873), .B(n31101), .Z(n40877) );
  NOR U44069 ( .A(n31102), .B(n31389), .Z(n31106) );
  IV U44070 ( .A(n31103), .Z(n31105) );
  NOR U44071 ( .A(n31105), .B(n31104), .Z(n40870) );
  NOR U44072 ( .A(n31106), .B(n40870), .Z(n31107) );
  XOR U44073 ( .A(n40873), .B(n31107), .Z(n31116) );
  NOR U44074 ( .A(n31386), .B(n31116), .Z(n31108) );
  NOR U44075 ( .A(n40877), .B(n31108), .Z(n31384) );
  IV U44076 ( .A(n31109), .Z(n31110) );
  NOR U44077 ( .A(n31110), .B(n31112), .Z(n34218) );
  IV U44078 ( .A(n31111), .Z(n31113) );
  NOR U44079 ( .A(n31113), .B(n31112), .Z(n31383) );
  NOR U44080 ( .A(n34218), .B(n31383), .Z(n31114) );
  NOR U44081 ( .A(n31384), .B(n31114), .Z(n31124) );
  IV U44082 ( .A(n31114), .Z(n31122) );
  NOR U44083 ( .A(n31115), .B(n37699), .Z(n31118) );
  IV U44084 ( .A(n31118), .Z(n31117) );
  IV U44085 ( .A(n31116), .Z(n37700) );
  NOR U44086 ( .A(n31117), .B(n37700), .Z(n37707) );
  NOR U44087 ( .A(n31118), .B(n31384), .Z(n31119) );
  NOR U44088 ( .A(n37707), .B(n31119), .Z(n31120) );
  IV U44089 ( .A(n31120), .Z(n31121) );
  NOR U44090 ( .A(n31122), .B(n31121), .Z(n31123) );
  NOR U44091 ( .A(n31124), .B(n31123), .Z(n34231) );
  XOR U44092 ( .A(n31380), .B(n34231), .Z(n34222) );
  XOR U44093 ( .A(n31125), .B(n34222), .Z(n37722) );
  NOR U44094 ( .A(n31126), .B(n37725), .Z(n31135) );
  IV U44095 ( .A(n31135), .Z(n31127) );
  NOR U44096 ( .A(n37722), .B(n31127), .Z(n34233) );
  IV U44097 ( .A(n31128), .Z(n31130) );
  NOR U44098 ( .A(n31130), .B(n34222), .Z(n31129) );
  IV U44099 ( .A(n31129), .Z(n34536) );
  NOR U44100 ( .A(n31131), .B(n34536), .Z(n34234) );
  NOR U44101 ( .A(n31131), .B(n31130), .Z(n31133) );
  IV U44102 ( .A(n37722), .Z(n31132) );
  NOR U44103 ( .A(n31133), .B(n31132), .Z(n31134) );
  NOR U44104 ( .A(n34234), .B(n31134), .Z(n34237) );
  NOR U44105 ( .A(n31135), .B(n34237), .Z(n31136) );
  NOR U44106 ( .A(n34233), .B(n31136), .Z(n31372) );
  IV U44107 ( .A(n31137), .Z(n34532) );
  NOR U44108 ( .A(n31138), .B(n34532), .Z(n34238) );
  NOR U44109 ( .A(n31139), .B(n31374), .Z(n31140) );
  NOR U44110 ( .A(n34238), .B(n31140), .Z(n31141) );
  XOR U44111 ( .A(n31372), .B(n31141), .Z(n31370) );
  XOR U44112 ( .A(n31368), .B(n31370), .Z(n31142) );
  XOR U44113 ( .A(n31143), .B(n31142), .Z(n31361) );
  IV U44114 ( .A(n31144), .Z(n31153) );
  IV U44115 ( .A(n31145), .Z(n31146) );
  NOR U44116 ( .A(n31153), .B(n31146), .Z(n34245) );
  IV U44117 ( .A(n31147), .Z(n31149) );
  NOR U44118 ( .A(n31149), .B(n31148), .Z(n31362) );
  NOR U44119 ( .A(n34245), .B(n31362), .Z(n31150) );
  XOR U44120 ( .A(n31361), .B(n31150), .Z(n34244) );
  IV U44121 ( .A(n31151), .Z(n31152) );
  NOR U44122 ( .A(n31153), .B(n31152), .Z(n34242) );
  XOR U44123 ( .A(n34244), .B(n34242), .Z(n38000) );
  XOR U44124 ( .A(n31356), .B(n38000), .Z(n31352) );
  XOR U44125 ( .A(n31154), .B(n31352), .Z(n34513) );
  XOR U44126 ( .A(n31350), .B(n34513), .Z(n31155) );
  IV U44127 ( .A(n31155), .Z(n34254) );
  XOR U44128 ( .A(n34253), .B(n34254), .Z(n31344) );
  IV U44129 ( .A(n31156), .Z(n31347) );
  NOR U44130 ( .A(n31347), .B(n31157), .Z(n31164) );
  IV U44131 ( .A(n31158), .Z(n31160) );
  NOR U44132 ( .A(n31160), .B(n31159), .Z(n31343) );
  NOR U44133 ( .A(n31164), .B(n31343), .Z(n31161) );
  XOR U44134 ( .A(n31344), .B(n31161), .Z(n31162) );
  NOR U44135 ( .A(n31163), .B(n31162), .Z(n31167) );
  IV U44136 ( .A(n31163), .Z(n31166) );
  XOR U44137 ( .A(n31164), .B(n31344), .Z(n31165) );
  NOR U44138 ( .A(n31166), .B(n31165), .Z(n34500) );
  NOR U44139 ( .A(n31167), .B(n34500), .Z(n31168) );
  IV U44140 ( .A(n31168), .Z(n34273) );
  XOR U44141 ( .A(n34261), .B(n34273), .Z(n34281) );
  NOR U44142 ( .A(n31169), .B(n34281), .Z(n34269) );
  IV U44143 ( .A(n31170), .Z(n34263) );
  NOR U44144 ( .A(n31171), .B(n34263), .Z(n34272) );
  NOR U44145 ( .A(n34261), .B(n34272), .Z(n31172) );
  XOR U44146 ( .A(n31172), .B(n34273), .Z(n31334) );
  NOR U44147 ( .A(n31173), .B(n31334), .Z(n31174) );
  NOR U44148 ( .A(n34269), .B(n31174), .Z(n31329) );
  IV U44149 ( .A(n31175), .Z(n31336) );
  NOR U44150 ( .A(n31176), .B(n31336), .Z(n31179) );
  IV U44151 ( .A(n31177), .Z(n31178) );
  NOR U44152 ( .A(n31178), .B(n31186), .Z(n31328) );
  NOR U44153 ( .A(n31179), .B(n31328), .Z(n31180) );
  XOR U44154 ( .A(n31329), .B(n31180), .Z(n34296) );
  IV U44155 ( .A(n31181), .Z(n31193) );
  IV U44156 ( .A(n31182), .Z(n31183) );
  NOR U44157 ( .A(n31193), .B(n31183), .Z(n31189) );
  IV U44158 ( .A(n31189), .Z(n31184) );
  NOR U44159 ( .A(n34296), .B(n31184), .Z(n37801) );
  IV U44160 ( .A(n31185), .Z(n31187) );
  NOR U44161 ( .A(n31187), .B(n31186), .Z(n31188) );
  IV U44162 ( .A(n31188), .Z(n34295) );
  XOR U44163 ( .A(n34295), .B(n34296), .Z(n31199) );
  NOR U44164 ( .A(n31189), .B(n31199), .Z(n31190) );
  NOR U44165 ( .A(n37801), .B(n31190), .Z(n31325) );
  IV U44166 ( .A(n31191), .Z(n31192) );
  NOR U44167 ( .A(n31193), .B(n31192), .Z(n31194) );
  IV U44168 ( .A(n31194), .Z(n31327) );
  XOR U44169 ( .A(n31325), .B(n31327), .Z(n31201) );
  NOR U44170 ( .A(n31195), .B(n31201), .Z(n37812) );
  IV U44171 ( .A(n31196), .Z(n31198) );
  NOR U44172 ( .A(n31198), .B(n31197), .Z(n31203) );
  IV U44173 ( .A(n31203), .Z(n31200) );
  IV U44174 ( .A(n31199), .Z(n31210) );
  NOR U44175 ( .A(n31200), .B(n31210), .Z(n34489) );
  IV U44176 ( .A(n31201), .Z(n31202) );
  NOR U44177 ( .A(n31203), .B(n31202), .Z(n31204) );
  NOR U44178 ( .A(n34489), .B(n31204), .Z(n31205) );
  NOR U44179 ( .A(n31206), .B(n31205), .Z(n31207) );
  NOR U44180 ( .A(n37812), .B(n31207), .Z(n31208) );
  NOR U44181 ( .A(n31209), .B(n31208), .Z(n31212) );
  IV U44182 ( .A(n31209), .Z(n31211) );
  NOR U44183 ( .A(n31211), .B(n31210), .Z(n34487) );
  NOR U44184 ( .A(n31212), .B(n34487), .Z(n31315) );
  IV U44185 ( .A(n31213), .Z(n34300) );
  NOR U44186 ( .A(n34300), .B(n31214), .Z(n31316) );
  NOR U44187 ( .A(n31215), .B(n34304), .Z(n34312) );
  NOR U44188 ( .A(n31316), .B(n34312), .Z(n31216) );
  XOR U44189 ( .A(n31315), .B(n31216), .Z(n31312) );
  XOR U44190 ( .A(n31217), .B(n31312), .Z(n34320) );
  XOR U44191 ( .A(n34318), .B(n34320), .Z(n37825) );
  IV U44192 ( .A(n31218), .Z(n31219) );
  NOR U44193 ( .A(n31220), .B(n31219), .Z(n31309) );
  IV U44194 ( .A(n31221), .Z(n31223) );
  NOR U44195 ( .A(n31223), .B(n31222), .Z(n34321) );
  NOR U44196 ( .A(n31309), .B(n34321), .Z(n31224) );
  XOR U44197 ( .A(n37825), .B(n31224), .Z(n31307) );
  XOR U44198 ( .A(n31225), .B(n31307), .Z(n34331) );
  XOR U44199 ( .A(n31226), .B(n34331), .Z(n31293) );
  XOR U44200 ( .A(n31292), .B(n31293), .Z(n34338) );
  XOR U44201 ( .A(n34336), .B(n34338), .Z(n34341) );
  XOR U44202 ( .A(n34339), .B(n34341), .Z(n31286) );
  XOR U44203 ( .A(n31227), .B(n31286), .Z(n37870) );
  XOR U44204 ( .A(n31279), .B(n37870), .Z(n31283) );
  XOR U44205 ( .A(n34347), .B(n31283), .Z(n31228) );
  XOR U44206 ( .A(n31281), .B(n31228), .Z(n31276) );
  IV U44207 ( .A(n31229), .Z(n31231) );
  NOR U44208 ( .A(n31231), .B(n31230), .Z(n34351) );
  IV U44209 ( .A(n31232), .Z(n31233) );
  NOR U44210 ( .A(n31234), .B(n31233), .Z(n31277) );
  NOR U44211 ( .A(n34351), .B(n31277), .Z(n31235) );
  XOR U44212 ( .A(n31276), .B(n31235), .Z(n34357) );
  XOR U44213 ( .A(n34355), .B(n34357), .Z(n34360) );
  XOR U44214 ( .A(n34358), .B(n34360), .Z(n31236) );
  NOR U44215 ( .A(n31237), .B(n31236), .Z(n34450) );
  IV U44216 ( .A(n31238), .Z(n31239) );
  NOR U44217 ( .A(n31240), .B(n31239), .Z(n31274) );
  NOR U44218 ( .A(n31274), .B(n34358), .Z(n31241) );
  XOR U44219 ( .A(n31241), .B(n34360), .Z(n34442) );
  NOR U44220 ( .A(n31242), .B(n34442), .Z(n31243) );
  NOR U44221 ( .A(n34450), .B(n31243), .Z(n31270) );
  XOR U44222 ( .A(n31272), .B(n31270), .Z(n34366) );
  IV U44223 ( .A(n31244), .Z(n31245) );
  NOR U44224 ( .A(n31246), .B(n31245), .Z(n31253) );
  IV U44225 ( .A(n31253), .Z(n31249) );
  XOR U44226 ( .A(n31248), .B(n31247), .Z(n31256) );
  NOR U44227 ( .A(n31249), .B(n31256), .Z(n34364) );
  IV U44228 ( .A(n31250), .Z(n31252) );
  NOR U44229 ( .A(n31252), .B(n31251), .Z(n31262) );
  IV U44230 ( .A(n31262), .Z(n34368) );
  NOR U44231 ( .A(n31254), .B(n31253), .Z(n31255) );
  XOR U44232 ( .A(n31256), .B(n31255), .Z(n31264) );
  IV U44233 ( .A(n31264), .Z(n34370) );
  NOR U44234 ( .A(n34368), .B(n34370), .Z(n31257) );
  NOR U44235 ( .A(n34364), .B(n31257), .Z(n31258) );
  XOR U44236 ( .A(n34366), .B(n31258), .Z(n34385) );
  IV U44237 ( .A(n34385), .Z(n34372) );
  IV U44238 ( .A(n31259), .Z(n31261) );
  NOR U44239 ( .A(n31261), .B(n31260), .Z(n34369) );
  NOR U44240 ( .A(n31262), .B(n34369), .Z(n31263) );
  XOR U44241 ( .A(n31264), .B(n31263), .Z(n34380) );
  NOR U44242 ( .A(n34372), .B(n34380), .Z(n31265) );
  IV U44243 ( .A(n31265), .Z(n34377) );
  IV U44244 ( .A(n31266), .Z(n31268) );
  NOR U44245 ( .A(n31268), .B(n31267), .Z(n34379) );
  IV U44246 ( .A(n34379), .Z(n31269) );
  NOR U44247 ( .A(n34377), .B(n31269), .Z(n34438) );
  IV U44248 ( .A(n31270), .Z(n31271) );
  NOR U44249 ( .A(n31272), .B(n31271), .Z(n31273) );
  NOR U44250 ( .A(n34450), .B(n31273), .Z(n34362) );
  IV U44251 ( .A(n31274), .Z(n31275) );
  NOR U44252 ( .A(n34360), .B(n31275), .Z(n34447) );
  IV U44253 ( .A(n31276), .Z(n34352) );
  IV U44254 ( .A(n31277), .Z(n37873) );
  NOR U44255 ( .A(n34352), .B(n37873), .Z(n31278) );
  IV U44256 ( .A(n31278), .Z(n34350) );
  IV U44257 ( .A(n31279), .Z(n31280) );
  NOR U44258 ( .A(n37870), .B(n31280), .Z(n37854) );
  IV U44259 ( .A(n31281), .Z(n31282) );
  NOR U44260 ( .A(n31283), .B(n31282), .Z(n37865) );
  NOR U44261 ( .A(n37854), .B(n37865), .Z(n31284) );
  IV U44262 ( .A(n31284), .Z(n34346) );
  IV U44263 ( .A(n31285), .Z(n31287) );
  NOR U44264 ( .A(n31287), .B(n31286), .Z(n37859) );
  IV U44265 ( .A(n31288), .Z(n31291) );
  NOR U44266 ( .A(n31289), .B(n34341), .Z(n31290) );
  IV U44267 ( .A(n31290), .Z(n34344) );
  NOR U44268 ( .A(n31291), .B(n34344), .Z(n37856) );
  IV U44269 ( .A(n31292), .Z(n31294) );
  NOR U44270 ( .A(n31294), .B(n31293), .Z(n31295) );
  IV U44271 ( .A(n31295), .Z(n34464) );
  IV U44272 ( .A(n31296), .Z(n31302) );
  NOR U44273 ( .A(n34328), .B(n34325), .Z(n31297) );
  XOR U44274 ( .A(n31307), .B(n31297), .Z(n31300) );
  IV U44275 ( .A(n31298), .Z(n31299) );
  NOR U44276 ( .A(n31300), .B(n31299), .Z(n31301) );
  IV U44277 ( .A(n31301), .Z(n31304) );
  NOR U44278 ( .A(n31302), .B(n31304), .Z(n37840) );
  IV U44279 ( .A(n31303), .Z(n31305) );
  NOR U44280 ( .A(n31305), .B(n31304), .Z(n37837) );
  IV U44281 ( .A(n31306), .Z(n31308) );
  IV U44282 ( .A(n31307), .Z(n34329) );
  NOR U44283 ( .A(n31308), .B(n34329), .Z(n37833) );
  IV U44284 ( .A(n31309), .Z(n31310) );
  NOR U44285 ( .A(n31310), .B(n37825), .Z(n34468) );
  IV U44286 ( .A(n31311), .Z(n31313) );
  NOR U44287 ( .A(n31313), .B(n31312), .Z(n34472) );
  IV U44288 ( .A(n31314), .Z(n31320) );
  IV U44289 ( .A(n31315), .Z(n34313) );
  XOR U44290 ( .A(n31316), .B(n34313), .Z(n31317) );
  NOR U44291 ( .A(n31318), .B(n31317), .Z(n31319) );
  IV U44292 ( .A(n31319), .Z(n31322) );
  NOR U44293 ( .A(n31320), .B(n31322), .Z(n34478) );
  IV U44294 ( .A(n31321), .Z(n31323) );
  NOR U44295 ( .A(n31323), .B(n31322), .Z(n34475) );
  NOR U44296 ( .A(n34489), .B(n34487), .Z(n31324) );
  IV U44297 ( .A(n31324), .Z(n34298) );
  IV U44298 ( .A(n31325), .Z(n31326) );
  NOR U44299 ( .A(n31327), .B(n31326), .Z(n37802) );
  IV U44300 ( .A(n31328), .Z(n31331) );
  IV U44301 ( .A(n31329), .Z(n31330) );
  NOR U44302 ( .A(n31331), .B(n31330), .Z(n31332) );
  IV U44303 ( .A(n31332), .Z(n37797) );
  IV U44304 ( .A(n31333), .Z(n31338) );
  IV U44305 ( .A(n31334), .Z(n31335) );
  NOR U44306 ( .A(n31336), .B(n31335), .Z(n31337) );
  IV U44307 ( .A(n31337), .Z(n31341) );
  NOR U44308 ( .A(n31338), .B(n31341), .Z(n31339) );
  IV U44309 ( .A(n31339), .Z(n34494) );
  IV U44310 ( .A(n31340), .Z(n31342) );
  NOR U44311 ( .A(n31342), .B(n31341), .Z(n34290) );
  IV U44312 ( .A(n31343), .Z(n31345) );
  NOR U44313 ( .A(n31345), .B(n31344), .Z(n34497) );
  IV U44314 ( .A(n31346), .Z(n31349) );
  NOR U44315 ( .A(n31347), .B(n34254), .Z(n31348) );
  IV U44316 ( .A(n31348), .Z(n34257) );
  NOR U44317 ( .A(n31349), .B(n34257), .Z(n34503) );
  NOR U44318 ( .A(n34513), .B(n31350), .Z(n34252) );
  IV U44319 ( .A(n31351), .Z(n31355) );
  IV U44320 ( .A(n31352), .Z(n31358) );
  NOR U44321 ( .A(n31353), .B(n31358), .Z(n31354) );
  IV U44322 ( .A(n31354), .Z(n34250) );
  NOR U44323 ( .A(n31355), .B(n34250), .Z(n37775) );
  NOR U44324 ( .A(n31356), .B(n38000), .Z(n37755) );
  IV U44325 ( .A(n31357), .Z(n31359) );
  NOR U44326 ( .A(n31359), .B(n31358), .Z(n34516) );
  NOR U44327 ( .A(n37755), .B(n34516), .Z(n31360) );
  IV U44328 ( .A(n31360), .Z(n34248) );
  IV U44329 ( .A(n31361), .Z(n34247) );
  IV U44330 ( .A(n31362), .Z(n31363) );
  NOR U44331 ( .A(n34247), .B(n31363), .Z(n37762) );
  IV U44332 ( .A(n31364), .Z(n31365) );
  NOR U44333 ( .A(n31370), .B(n31365), .Z(n37765) );
  NOR U44334 ( .A(n37762), .B(n37765), .Z(n34241) );
  IV U44335 ( .A(n31366), .Z(n31367) );
  NOR U44336 ( .A(n31370), .B(n31367), .Z(n34523) );
  IV U44337 ( .A(n31368), .Z(n31369) );
  NOR U44338 ( .A(n31370), .B(n31369), .Z(n34520) );
  IV U44339 ( .A(n31371), .Z(n31376) );
  IV U44340 ( .A(n31372), .Z(n31373) );
  NOR U44341 ( .A(n31374), .B(n31373), .Z(n31375) );
  IV U44342 ( .A(n31375), .Z(n31378) );
  NOR U44343 ( .A(n31376), .B(n31378), .Z(n37745) );
  IV U44344 ( .A(n31377), .Z(n31379) );
  NOR U44345 ( .A(n31379), .B(n31378), .Z(n37742) );
  IV U44346 ( .A(n31380), .Z(n31381) );
  NOR U44347 ( .A(n31381), .B(n34231), .Z(n31382) );
  IV U44348 ( .A(n31382), .Z(n34224) );
  IV U44349 ( .A(n31383), .Z(n31385) );
  IV U44350 ( .A(n31384), .Z(n34219) );
  NOR U44351 ( .A(n31385), .B(n34219), .Z(n37713) );
  NOR U44352 ( .A(n31386), .B(n40870), .Z(n31387) );
  NOR U44353 ( .A(n31387), .B(n40873), .Z(n37695) );
  IV U44354 ( .A(n31388), .Z(n31391) );
  NOR U44355 ( .A(n40873), .B(n31389), .Z(n31390) );
  IV U44356 ( .A(n31390), .Z(n31393) );
  NOR U44357 ( .A(n31391), .B(n31393), .Z(n37691) );
  IV U44358 ( .A(n31392), .Z(n31394) );
  NOR U44359 ( .A(n31394), .B(n31393), .Z(n37688) );
  IV U44360 ( .A(n31395), .Z(n31398) );
  IV U44361 ( .A(n31396), .Z(n31397) );
  NOR U44362 ( .A(n31398), .B(n31397), .Z(n37684) );
  IV U44363 ( .A(n31399), .Z(n34205) );
  IV U44364 ( .A(n31400), .Z(n31404) );
  IV U44365 ( .A(n31401), .Z(n31402) );
  NOR U44366 ( .A(n31404), .B(n31402), .Z(n34549) );
  IV U44367 ( .A(n31403), .Z(n37678) );
  NOR U44368 ( .A(n31404), .B(n37678), .Z(n34194) );
  IV U44369 ( .A(n31405), .Z(n31406) );
  NOR U44370 ( .A(n37681), .B(n31406), .Z(n37674) );
  IV U44371 ( .A(n31407), .Z(n31408) );
  NOR U44372 ( .A(n37681), .B(n31408), .Z(n34554) );
  IV U44373 ( .A(n31409), .Z(n31410) );
  NOR U44374 ( .A(n31411), .B(n31410), .Z(n34557) );
  NOR U44375 ( .A(n34563), .B(n34557), .Z(n31412) );
  IV U44376 ( .A(n31412), .Z(n34193) );
  NOR U44377 ( .A(n34559), .B(n34569), .Z(n31413) );
  NOR U44378 ( .A(n31413), .B(n34571), .Z(n34192) );
  IV U44379 ( .A(n31414), .Z(n31418) );
  NOR U44380 ( .A(n31416), .B(n31415), .Z(n31417) );
  IV U44381 ( .A(n31417), .Z(n31420) );
  NOR U44382 ( .A(n31418), .B(n31420), .Z(n34566) );
  IV U44383 ( .A(n31419), .Z(n31421) );
  NOR U44384 ( .A(n31421), .B(n31420), .Z(n34575) );
  IV U44385 ( .A(n31422), .Z(n31424) );
  IV U44386 ( .A(n31423), .Z(n31426) );
  NOR U44387 ( .A(n31424), .B(n31426), .Z(n34581) );
  IV U44388 ( .A(n31425), .Z(n31427) );
  NOR U44389 ( .A(n31427), .B(n31426), .Z(n34578) );
  IV U44390 ( .A(n31428), .Z(n31429) );
  NOR U44391 ( .A(n31430), .B(n31429), .Z(n31431) );
  IV U44392 ( .A(n31431), .Z(n37670) );
  XOR U44393 ( .A(n34584), .B(n37662), .Z(n31432) );
  NOR U44394 ( .A(n37665), .B(n31432), .Z(n34191) );
  IV U44395 ( .A(n31433), .Z(n37654) );
  IV U44396 ( .A(n31434), .Z(n31439) );
  XOR U44397 ( .A(n31435), .B(n31447), .Z(n31437) );
  NOR U44398 ( .A(n31437), .B(n31436), .Z(n31438) );
  IV U44399 ( .A(n31438), .Z(n34183) );
  NOR U44400 ( .A(n31439), .B(n34183), .Z(n37639) );
  IV U44401 ( .A(n31440), .Z(n31441) );
  NOR U44402 ( .A(n31442), .B(n31441), .Z(n37642) );
  IV U44403 ( .A(n31443), .Z(n31444) );
  NOR U44404 ( .A(n31447), .B(n31444), .Z(n34594) );
  IV U44405 ( .A(n31445), .Z(n31449) );
  NOR U44406 ( .A(n31447), .B(n31446), .Z(n31448) );
  IV U44407 ( .A(n31448), .Z(n31452) );
  NOR U44408 ( .A(n31449), .B(n31452), .Z(n34597) );
  NOR U44409 ( .A(n34594), .B(n34597), .Z(n31450) );
  IV U44410 ( .A(n31450), .Z(n34181) );
  IV U44411 ( .A(n31451), .Z(n31453) );
  NOR U44412 ( .A(n31453), .B(n31452), .Z(n34599) );
  IV U44413 ( .A(n31454), .Z(n31455) );
  NOR U44414 ( .A(n31455), .B(n31458), .Z(n31456) );
  IV U44415 ( .A(n31456), .Z(n37636) );
  IV U44416 ( .A(n31457), .Z(n31459) );
  NOR U44417 ( .A(n31459), .B(n31458), .Z(n38044) );
  NOR U44418 ( .A(n38049), .B(n38044), .Z(n37634) );
  IV U44419 ( .A(n37634), .Z(n34164) );
  IV U44420 ( .A(n31460), .Z(n31461) );
  NOR U44421 ( .A(n31464), .B(n31461), .Z(n34619) );
  IV U44422 ( .A(n31462), .Z(n31463) );
  NOR U44423 ( .A(n31464), .B(n31463), .Z(n34625) );
  IV U44424 ( .A(n31465), .Z(n31467) );
  NOR U44425 ( .A(n31467), .B(n31466), .Z(n37623) );
  IV U44426 ( .A(n31468), .Z(n31471) );
  NOR U44427 ( .A(n31469), .B(n31477), .Z(n31470) );
  IV U44428 ( .A(n31470), .Z(n31473) );
  NOR U44429 ( .A(n31471), .B(n31473), .Z(n37620) );
  IV U44430 ( .A(n31472), .Z(n31474) );
  NOR U44431 ( .A(n31474), .B(n31473), .Z(n37616) );
  IV U44432 ( .A(n31475), .Z(n31476) );
  NOR U44433 ( .A(n31477), .B(n31476), .Z(n37613) );
  IV U44434 ( .A(n31478), .Z(n31482) );
  IV U44435 ( .A(n31479), .Z(n31480) );
  NOR U44436 ( .A(n31482), .B(n31480), .Z(n34631) );
  IV U44437 ( .A(n31481), .Z(n31483) );
  NOR U44438 ( .A(n31483), .B(n31482), .Z(n34628) );
  NOR U44439 ( .A(n31485), .B(n31484), .Z(n34645) );
  IV U44440 ( .A(n31486), .Z(n31489) );
  IV U44441 ( .A(n31487), .Z(n31488) );
  NOR U44442 ( .A(n31489), .B(n31488), .Z(n34642) );
  IV U44443 ( .A(n31490), .Z(n31492) );
  NOR U44444 ( .A(n31492), .B(n31491), .Z(n34651) );
  IV U44445 ( .A(n31493), .Z(n31494) );
  NOR U44446 ( .A(n31494), .B(n34678), .Z(n34160) );
  IV U44447 ( .A(n31495), .Z(n34155) );
  IV U44448 ( .A(n31496), .Z(n31497) );
  NOR U44449 ( .A(n34155), .B(n31497), .Z(n37603) );
  NOR U44450 ( .A(n31499), .B(n31498), .Z(n37600) );
  IV U44451 ( .A(n31500), .Z(n31501) );
  NOR U44452 ( .A(n31507), .B(n31501), .Z(n37584) );
  NOR U44453 ( .A(n37600), .B(n37584), .Z(n31502) );
  IV U44454 ( .A(n31502), .Z(n34153) );
  IV U44455 ( .A(n31503), .Z(n31504) );
  NOR U44456 ( .A(n31507), .B(n31504), .Z(n34685) );
  IV U44457 ( .A(n31505), .Z(n31506) );
  NOR U44458 ( .A(n31507), .B(n31506), .Z(n37586) );
  NOR U44459 ( .A(n31513), .B(n31508), .Z(n37580) );
  IV U44460 ( .A(n31509), .Z(n31510) );
  NOR U44461 ( .A(n31513), .B(n31510), .Z(n37577) );
  IV U44462 ( .A(n31511), .Z(n31512) );
  NOR U44463 ( .A(n31513), .B(n31512), .Z(n37566) );
  IV U44464 ( .A(n31514), .Z(n31515) );
  NOR U44465 ( .A(n31516), .B(n31515), .Z(n34689) );
  IV U44466 ( .A(n31517), .Z(n31520) );
  NOR U44467 ( .A(n31518), .B(n34148), .Z(n31519) );
  IV U44468 ( .A(n31519), .Z(n31522) );
  NOR U44469 ( .A(n31520), .B(n31522), .Z(n37569) );
  IV U44470 ( .A(n31521), .Z(n31523) );
  NOR U44471 ( .A(n31523), .B(n31522), .Z(n37562) );
  IV U44472 ( .A(n31524), .Z(n34151) );
  IV U44473 ( .A(n31525), .Z(n31526) );
  NOR U44474 ( .A(n34151), .B(n31526), .Z(n34697) );
  NOR U44475 ( .A(n34699), .B(n34697), .Z(n31527) );
  IV U44476 ( .A(n31527), .Z(n34140) );
  IV U44477 ( .A(n31528), .Z(n31529) );
  NOR U44478 ( .A(n31533), .B(n31529), .Z(n37557) );
  IV U44479 ( .A(n31530), .Z(n31531) );
  NOR U44480 ( .A(n31531), .B(n31533), .Z(n37554) );
  IV U44481 ( .A(n31532), .Z(n31534) );
  NOR U44482 ( .A(n31534), .B(n31533), .Z(n37547) );
  IV U44483 ( .A(n31535), .Z(n31536) );
  NOR U44484 ( .A(n31536), .B(n50781), .Z(n44016) );
  IV U44485 ( .A(n31537), .Z(n44023) );
  IV U44486 ( .A(n31538), .Z(n44018) );
  NOR U44487 ( .A(n44023), .B(n44018), .Z(n34712) );
  NOR U44488 ( .A(n44016), .B(n34712), .Z(n31539) );
  IV U44489 ( .A(n31539), .Z(n34113) );
  IV U44490 ( .A(n31540), .Z(n31545) );
  IV U44491 ( .A(n31541), .Z(n31542) );
  NOR U44492 ( .A(n31543), .B(n31542), .Z(n31544) );
  IV U44493 ( .A(n31544), .Z(n31547) );
  NOR U44494 ( .A(n31545), .B(n31547), .Z(n34717) );
  IV U44495 ( .A(n31546), .Z(n31548) );
  NOR U44496 ( .A(n31548), .B(n31547), .Z(n34722) );
  XOR U44497 ( .A(n34721), .B(n34722), .Z(n31549) );
  NOR U44498 ( .A(n34717), .B(n31549), .Z(n34112) );
  IV U44499 ( .A(n31550), .Z(n31551) );
  NOR U44500 ( .A(n31551), .B(n34109), .Z(n37531) );
  IV U44501 ( .A(n31552), .Z(n31554) );
  NOR U44502 ( .A(n31554), .B(n31553), .Z(n37524) );
  IV U44503 ( .A(n31555), .Z(n31556) );
  NOR U44504 ( .A(n31557), .B(n31556), .Z(n37527) );
  NOR U44505 ( .A(n37524), .B(n37527), .Z(n34105) );
  NOR U44506 ( .A(n31559), .B(n31558), .Z(n34729) );
  IV U44507 ( .A(n31560), .Z(n31562) );
  NOR U44508 ( .A(n31562), .B(n31561), .Z(n34727) );
  NOR U44509 ( .A(n34729), .B(n34727), .Z(n34104) );
  NOR U44510 ( .A(n31563), .B(n34748), .Z(n31565) );
  NOR U44511 ( .A(n31565), .B(n31564), .Z(n34100) );
  IV U44512 ( .A(n31566), .Z(n31567) );
  NOR U44513 ( .A(n31568), .B(n31567), .Z(n34751) );
  NOR U44514 ( .A(n37519), .B(n34751), .Z(n31569) );
  IV U44515 ( .A(n31569), .Z(n34099) );
  IV U44516 ( .A(n31570), .Z(n31573) );
  IV U44517 ( .A(n31571), .Z(n31572) );
  NOR U44518 ( .A(n31573), .B(n31572), .Z(n37516) );
  NOR U44519 ( .A(n34754), .B(n37516), .Z(n34098) );
  IV U44520 ( .A(n31574), .Z(n31576) );
  NOR U44521 ( .A(n31576), .B(n31575), .Z(n34757) );
  IV U44522 ( .A(n31577), .Z(n31580) );
  NOR U44523 ( .A(n31578), .B(n34091), .Z(n31579) );
  IV U44524 ( .A(n31579), .Z(n34095) );
  NOR U44525 ( .A(n31580), .B(n34095), .Z(n37512) );
  NOR U44526 ( .A(n34757), .B(n37512), .Z(n34097) );
  NOR U44527 ( .A(n31582), .B(n31581), .Z(n31583) );
  IV U44528 ( .A(n31583), .Z(n34771) );
  IV U44529 ( .A(n31584), .Z(n31585) );
  NOR U44530 ( .A(n34071), .B(n31585), .Z(n37488) );
  IV U44531 ( .A(n31586), .Z(n31587) );
  NOR U44532 ( .A(n34071), .B(n31587), .Z(n37485) );
  IV U44533 ( .A(n31588), .Z(n31592) );
  IV U44534 ( .A(n31589), .Z(n34786) );
  NOR U44535 ( .A(n31590), .B(n34786), .Z(n31591) );
  IV U44536 ( .A(n31591), .Z(n31594) );
  NOR U44537 ( .A(n31592), .B(n31594), .Z(n34795) );
  IV U44538 ( .A(n31593), .Z(n31595) );
  NOR U44539 ( .A(n31595), .B(n31594), .Z(n34792) );
  IV U44540 ( .A(n31596), .Z(n31599) );
  IV U44541 ( .A(n31597), .Z(n31598) );
  NOR U44542 ( .A(n31599), .B(n31598), .Z(n34802) );
  NOR U44543 ( .A(n37475), .B(n34802), .Z(n31600) );
  IV U44544 ( .A(n31600), .Z(n34065) );
  IV U44545 ( .A(n31601), .Z(n31603) );
  NOR U44546 ( .A(n31603), .B(n31602), .Z(n34805) );
  NOR U44547 ( .A(n31605), .B(n31604), .Z(n37478) );
  NOR U44548 ( .A(n34805), .B(n37478), .Z(n34064) );
  IV U44549 ( .A(n31606), .Z(n31607) );
  NOR U44550 ( .A(n31608), .B(n31607), .Z(n37472) );
  IV U44551 ( .A(n31609), .Z(n31611) );
  NOR U44552 ( .A(n31611), .B(n31610), .Z(n34808) );
  NOR U44553 ( .A(n37472), .B(n34808), .Z(n34063) );
  IV U44554 ( .A(n34042), .Z(n34036) );
  IV U44555 ( .A(n31612), .Z(n31613) );
  NOR U44556 ( .A(n34039), .B(n31613), .Z(n34830) );
  IV U44557 ( .A(n31614), .Z(n31617) );
  NOR U44558 ( .A(n31615), .B(n47236), .Z(n31616) );
  IV U44559 ( .A(n31616), .Z(n31624) );
  NOR U44560 ( .A(n31617), .B(n31624), .Z(n31618) );
  IV U44561 ( .A(n31618), .Z(n37455) );
  IV U44562 ( .A(n31619), .Z(n31620) );
  NOR U44563 ( .A(n31620), .B(n47236), .Z(n31621) );
  IV U44564 ( .A(n31621), .Z(n31622) );
  NOR U44565 ( .A(n31627), .B(n31622), .Z(n37437) );
  IV U44566 ( .A(n31623), .Z(n31625) );
  NOR U44567 ( .A(n31625), .B(n31624), .Z(n37451) );
  NOR U44568 ( .A(n37437), .B(n37451), .Z(n31626) );
  IV U44569 ( .A(n31626), .Z(n34029) );
  IV U44570 ( .A(n31627), .Z(n31628) );
  NOR U44571 ( .A(n31629), .B(n31628), .Z(n31630) );
  NOR U44572 ( .A(n47244), .B(n31630), .Z(n31631) );
  NOR U44573 ( .A(n47246), .B(n31631), .Z(n37440) );
  IV U44574 ( .A(n31632), .Z(n34027) );
  IV U44575 ( .A(n31633), .Z(n31634) );
  NOR U44576 ( .A(n34027), .B(n31634), .Z(n34834) );
  NOR U44577 ( .A(n31636), .B(n31635), .Z(n31637) );
  IV U44578 ( .A(n31637), .Z(n37432) );
  NOR U44579 ( .A(n31638), .B(n41470), .Z(n40508) );
  NOR U44580 ( .A(n40508), .B(n40506), .Z(n34021) );
  IV U44581 ( .A(n31639), .Z(n31642) );
  NOR U44582 ( .A(n31640), .B(n31651), .Z(n31641) );
  IV U44583 ( .A(n31641), .Z(n31647) );
  NOR U44584 ( .A(n31642), .B(n31647), .Z(n37421) );
  IV U44585 ( .A(n31643), .Z(n31644) );
  NOR U44586 ( .A(n31645), .B(n31644), .Z(n37415) );
  IV U44587 ( .A(n31646), .Z(n31648) );
  NOR U44588 ( .A(n31648), .B(n31647), .Z(n37424) );
  NOR U44589 ( .A(n37415), .B(n37424), .Z(n31649) );
  IV U44590 ( .A(n31649), .Z(n34020) );
  IV U44591 ( .A(n31650), .Z(n31652) );
  NOR U44592 ( .A(n31652), .B(n31651), .Z(n37417) );
  NOR U44593 ( .A(n37408), .B(n37417), .Z(n34019) );
  IV U44594 ( .A(n31653), .Z(n31656) );
  IV U44595 ( .A(n31654), .Z(n31655) );
  NOR U44596 ( .A(n31656), .B(n31655), .Z(n37396) );
  NOR U44597 ( .A(n37402), .B(n37396), .Z(n34018) );
  IV U44598 ( .A(n31657), .Z(n31658) );
  NOR U44599 ( .A(n31659), .B(n31658), .Z(n34840) );
  IV U44600 ( .A(n31660), .Z(n31665) );
  IV U44601 ( .A(n31661), .Z(n31675) );
  XOR U44602 ( .A(n31674), .B(n31675), .Z(n31662) );
  NOR U44603 ( .A(n31663), .B(n31662), .Z(n31664) );
  IV U44604 ( .A(n31664), .Z(n31670) );
  NOR U44605 ( .A(n31665), .B(n31670), .Z(n34837) );
  IV U44606 ( .A(n31666), .Z(n31668) );
  NOR U44607 ( .A(n31668), .B(n31667), .Z(n34846) );
  IV U44608 ( .A(n31669), .Z(n31671) );
  NOR U44609 ( .A(n31671), .B(n31670), .Z(n34844) );
  NOR U44610 ( .A(n34846), .B(n34844), .Z(n34017) );
  IV U44611 ( .A(n31672), .Z(n31673) );
  NOR U44612 ( .A(n31675), .B(n31673), .Z(n34849) );
  IV U44613 ( .A(n31674), .Z(n31676) );
  NOR U44614 ( .A(n31676), .B(n31675), .Z(n37392) );
  NOR U44615 ( .A(n34849), .B(n37392), .Z(n34016) );
  NOR U44616 ( .A(n31678), .B(n31677), .Z(n37389) );
  IV U44617 ( .A(n31679), .Z(n31683) );
  IV U44618 ( .A(n31680), .Z(n31681) );
  NOR U44619 ( .A(n31683), .B(n31681), .Z(n37386) );
  IV U44620 ( .A(n31682), .Z(n31684) );
  NOR U44621 ( .A(n31684), .B(n31683), .Z(n34852) );
  NOR U44622 ( .A(n34870), .B(n34865), .Z(n33996) );
  NOR U44623 ( .A(n34874), .B(n34867), .Z(n33995) );
  IV U44624 ( .A(n31685), .Z(n31686) );
  NOR U44625 ( .A(n31691), .B(n31686), .Z(n37358) );
  IV U44626 ( .A(n31687), .Z(n31688) );
  NOR U44627 ( .A(n31688), .B(n31694), .Z(n34877) );
  IV U44628 ( .A(n31689), .Z(n31690) );
  NOR U44629 ( .A(n31691), .B(n31690), .Z(n37361) );
  NOR U44630 ( .A(n34877), .B(n37361), .Z(n33994) );
  IV U44631 ( .A(n31695), .Z(n31692) );
  NOR U44632 ( .A(n31692), .B(n31694), .Z(n34879) );
  IV U44633 ( .A(n31693), .Z(n31697) );
  XOR U44634 ( .A(n31695), .B(n31694), .Z(n31696) );
  NOR U44635 ( .A(n31697), .B(n31696), .Z(n34881) );
  NOR U44636 ( .A(n34879), .B(n34881), .Z(n33993) );
  IV U44637 ( .A(n31698), .Z(n31700) );
  NOR U44638 ( .A(n31700), .B(n31699), .Z(n34885) );
  IV U44639 ( .A(n31701), .Z(n33988) );
  IV U44640 ( .A(n31704), .Z(n31702) );
  NOR U44641 ( .A(n33988), .B(n31702), .Z(n34899) );
  IV U44642 ( .A(n31703), .Z(n31706) );
  XOR U44643 ( .A(n31704), .B(n33988), .Z(n31705) );
  NOR U44644 ( .A(n31706), .B(n31705), .Z(n34891) );
  NOR U44645 ( .A(n34899), .B(n34891), .Z(n33985) );
  IV U44646 ( .A(n31707), .Z(n31709) );
  NOR U44647 ( .A(n31709), .B(n31708), .Z(n34896) );
  IV U44648 ( .A(n31710), .Z(n31711) );
  NOR U44649 ( .A(n31714), .B(n31711), .Z(n34902) );
  IV U44650 ( .A(n31712), .Z(n31713) );
  NOR U44651 ( .A(n31714), .B(n31713), .Z(n34905) );
  IV U44652 ( .A(n31715), .Z(n31718) );
  NOR U44653 ( .A(n31716), .B(n33979), .Z(n31717) );
  IV U44654 ( .A(n31717), .Z(n31720) );
  NOR U44655 ( .A(n31718), .B(n31720), .Z(n37351) );
  IV U44656 ( .A(n31719), .Z(n31721) );
  NOR U44657 ( .A(n31721), .B(n31720), .Z(n37348) );
  IV U44658 ( .A(n31722), .Z(n31723) );
  NOR U44659 ( .A(n33976), .B(n31723), .Z(n38255) );
  IV U44660 ( .A(n31724), .Z(n33983) );
  IV U44661 ( .A(n31725), .Z(n31726) );
  NOR U44662 ( .A(n33983), .B(n31726), .Z(n38251) );
  NOR U44663 ( .A(n38255), .B(n38251), .Z(n34918) );
  IV U44664 ( .A(n31727), .Z(n31729) );
  NOR U44665 ( .A(n31729), .B(n31728), .Z(n37342) );
  IV U44666 ( .A(n31730), .Z(n31732) );
  NOR U44667 ( .A(n31732), .B(n31731), .Z(n37344) );
  NOR U44668 ( .A(n37342), .B(n37344), .Z(n33966) );
  IV U44669 ( .A(n31733), .Z(n31734) );
  NOR U44670 ( .A(n31735), .B(n31734), .Z(n34931) );
  IV U44671 ( .A(n31736), .Z(n31739) );
  NOR U44672 ( .A(n33950), .B(n31737), .Z(n31738) );
  IV U44673 ( .A(n31738), .Z(n33956) );
  NOR U44674 ( .A(n31739), .B(n33956), .Z(n34938) );
  IV U44675 ( .A(n31740), .Z(n31741) );
  NOR U44676 ( .A(n33938), .B(n31741), .Z(n34956) );
  IV U44677 ( .A(n31742), .Z(n31743) );
  NOR U44678 ( .A(n31743), .B(n34968), .Z(n33930) );
  IV U44679 ( .A(n31744), .Z(n31745) );
  NOR U44680 ( .A(n34968), .B(n31745), .Z(n37320) );
  IV U44681 ( .A(n31746), .Z(n37313) );
  NOR U44682 ( .A(n31747), .B(n37313), .Z(n33929) );
  IV U44683 ( .A(n31748), .Z(n31751) );
  IV U44684 ( .A(n31749), .Z(n31750) );
  NOR U44685 ( .A(n31751), .B(n31750), .Z(n31752) );
  IV U44686 ( .A(n31752), .Z(n33920) );
  IV U44687 ( .A(n31753), .Z(n31754) );
  NOR U44688 ( .A(n31754), .B(n34990), .Z(n33918) );
  IV U44689 ( .A(n31755), .Z(n31757) );
  NOR U44690 ( .A(n31757), .B(n31756), .Z(n35002) );
  IV U44691 ( .A(n31758), .Z(n31759) );
  NOR U44692 ( .A(n31759), .B(n34990), .Z(n35000) );
  NOR U44693 ( .A(n35002), .B(n35000), .Z(n33917) );
  IV U44694 ( .A(n31760), .Z(n31762) );
  NOR U44695 ( .A(n31762), .B(n31761), .Z(n35005) );
  IV U44696 ( .A(n31763), .Z(n31767) );
  IV U44697 ( .A(n31764), .Z(n31773) );
  NOR U44698 ( .A(n31765), .B(n31773), .Z(n31766) );
  IV U44699 ( .A(n31766), .Z(n31769) );
  NOR U44700 ( .A(n31767), .B(n31769), .Z(n37304) );
  NOR U44701 ( .A(n35005), .B(n37304), .Z(n33916) );
  IV U44702 ( .A(n31768), .Z(n31770) );
  NOR U44703 ( .A(n31770), .B(n31769), .Z(n37301) );
  IV U44704 ( .A(n31771), .Z(n31772) );
  NOR U44705 ( .A(n31773), .B(n31772), .Z(n35007) );
  NOR U44706 ( .A(n35016), .B(n31774), .Z(n33915) );
  IV U44707 ( .A(n31775), .Z(n31778) );
  NOR U44708 ( .A(n31776), .B(n33910), .Z(n31777) );
  IV U44709 ( .A(n31777), .Z(n33912) );
  NOR U44710 ( .A(n31778), .B(n33912), .Z(n35011) );
  IV U44711 ( .A(n31779), .Z(n31782) );
  IV U44712 ( .A(n31780), .Z(n31781) );
  NOR U44713 ( .A(n31782), .B(n31781), .Z(n31783) );
  IV U44714 ( .A(n31783), .Z(n35026) );
  NOR U44715 ( .A(n37282), .B(n31784), .Z(n38350) );
  IV U44716 ( .A(n31785), .Z(n31788) );
  IV U44717 ( .A(n31786), .Z(n31787) );
  NOR U44718 ( .A(n31788), .B(n31787), .Z(n38355) );
  NOR U44719 ( .A(n38350), .B(n38355), .Z(n37277) );
  IV U44720 ( .A(n37277), .Z(n33898) );
  IV U44721 ( .A(n31789), .Z(n31792) );
  IV U44722 ( .A(n31790), .Z(n31791) );
  NOR U44723 ( .A(n31792), .B(n31791), .Z(n43768) );
  NOR U44724 ( .A(n41627), .B(n43768), .Z(n40353) );
  IV U44725 ( .A(n31793), .Z(n37268) );
  NOR U44726 ( .A(n37268), .B(n35027), .Z(n31796) );
  IV U44727 ( .A(n31794), .Z(n35029) );
  NOR U44728 ( .A(n35029), .B(n33896), .Z(n31795) );
  NOR U44729 ( .A(n31796), .B(n31795), .Z(n33890) );
  IV U44730 ( .A(n31797), .Z(n31798) );
  NOR U44731 ( .A(n31808), .B(n31798), .Z(n31799) );
  IV U44732 ( .A(n31799), .Z(n35031) );
  IV U44733 ( .A(n31800), .Z(n31802) );
  XOR U44734 ( .A(n31806), .B(n31808), .Z(n31801) );
  NOR U44735 ( .A(n31802), .B(n31801), .Z(n37254) );
  IV U44736 ( .A(n31803), .Z(n31805) );
  NOR U44737 ( .A(n31805), .B(n31804), .Z(n35032) );
  IV U44738 ( .A(n31806), .Z(n31807) );
  NOR U44739 ( .A(n31808), .B(n31807), .Z(n37257) );
  NOR U44740 ( .A(n35032), .B(n37257), .Z(n31809) );
  IV U44741 ( .A(n31809), .Z(n33888) );
  IV U44742 ( .A(n31810), .Z(n31812) );
  IV U44743 ( .A(n31811), .Z(n33885) );
  NOR U44744 ( .A(n31812), .B(n33885), .Z(n35034) );
  IV U44745 ( .A(n31813), .Z(n35047) );
  NOR U44746 ( .A(n31815), .B(n31814), .Z(n35043) );
  IV U44747 ( .A(n31816), .Z(n31817) );
  NOR U44748 ( .A(n31819), .B(n31817), .Z(n37249) );
  IV U44749 ( .A(n31818), .Z(n31820) );
  NOR U44750 ( .A(n31820), .B(n31819), .Z(n37247) );
  NOR U44751 ( .A(n37249), .B(n37247), .Z(n31821) );
  IV U44752 ( .A(n31821), .Z(n33883) );
  IV U44753 ( .A(n31822), .Z(n33878) );
  IV U44754 ( .A(n31823), .Z(n31824) );
  NOR U44755 ( .A(n33878), .B(n31824), .Z(n35051) );
  IV U44756 ( .A(n31825), .Z(n31826) );
  NOR U44757 ( .A(n31828), .B(n31826), .Z(n35061) );
  IV U44758 ( .A(n31827), .Z(n31831) );
  NOR U44759 ( .A(n31829), .B(n31828), .Z(n31830) );
  IV U44760 ( .A(n31830), .Z(n33873) );
  NOR U44761 ( .A(n31831), .B(n33873), .Z(n35059) );
  NOR U44762 ( .A(n35061), .B(n35059), .Z(n31832) );
  IV U44763 ( .A(n31832), .Z(n33871) );
  IV U44764 ( .A(n31833), .Z(n31842) );
  IV U44765 ( .A(n31834), .Z(n31835) );
  NOR U44766 ( .A(n31842), .B(n31835), .Z(n31836) );
  IV U44767 ( .A(n31836), .Z(n35066) );
  NOR U44768 ( .A(n35066), .B(n31837), .Z(n33870) );
  IV U44769 ( .A(n31838), .Z(n31839) );
  NOR U44770 ( .A(n31839), .B(n35075), .Z(n35070) );
  IV U44771 ( .A(n31840), .Z(n31841) );
  NOR U44772 ( .A(n31842), .B(n31841), .Z(n37240) );
  NOR U44773 ( .A(n35070), .B(n37240), .Z(n33869) );
  NOR U44774 ( .A(n31843), .B(n35075), .Z(n31849) );
  IV U44775 ( .A(n31844), .Z(n31845) );
  NOR U44776 ( .A(n31846), .B(n31845), .Z(n31847) );
  IV U44777 ( .A(n31847), .Z(n31848) );
  NOR U44778 ( .A(n31850), .B(n31848), .Z(n35078) );
  NOR U44779 ( .A(n31849), .B(n35078), .Z(n33868) );
  IV U44780 ( .A(n31850), .Z(n31852) );
  IV U44781 ( .A(n31851), .Z(n35082) );
  NOR U44782 ( .A(n31852), .B(n35082), .Z(n33867) );
  NOR U44783 ( .A(n31854), .B(n31853), .Z(n35095) );
  IV U44784 ( .A(n31855), .Z(n31857) );
  NOR U44785 ( .A(n31857), .B(n31856), .Z(n40265) );
  IV U44786 ( .A(n31858), .Z(n31859) );
  NOR U44787 ( .A(n31859), .B(n33860), .Z(n38402) );
  NOR U44788 ( .A(n40265), .B(n38402), .Z(n35101) );
  IV U44789 ( .A(n31860), .Z(n31861) );
  NOR U44790 ( .A(n31862), .B(n31861), .Z(n37227) );
  IV U44791 ( .A(n31863), .Z(n31866) );
  IV U44792 ( .A(n31864), .Z(n31865) );
  NOR U44793 ( .A(n31866), .B(n31865), .Z(n37224) );
  IV U44794 ( .A(n31867), .Z(n31870) );
  IV U44795 ( .A(n31868), .Z(n31869) );
  NOR U44796 ( .A(n31870), .B(n31869), .Z(n35106) );
  IV U44797 ( .A(n31871), .Z(n31873) );
  NOR U44798 ( .A(n31873), .B(n31872), .Z(n35112) );
  IV U44799 ( .A(n31874), .Z(n31875) );
  NOR U44800 ( .A(n35117), .B(n31875), .Z(n33858) );
  IV U44801 ( .A(n31876), .Z(n31877) );
  NOR U44802 ( .A(n35117), .B(n31877), .Z(n37216) );
  IV U44803 ( .A(n31878), .Z(n31880) );
  IV U44804 ( .A(n31879), .Z(n31882) );
  NOR U44805 ( .A(n31880), .B(n31882), .Z(n37213) );
  IV U44806 ( .A(n31881), .Z(n31883) );
  NOR U44807 ( .A(n31883), .B(n31882), .Z(n37202) );
  IV U44808 ( .A(n31884), .Z(n31888) );
  NOR U44809 ( .A(n31886), .B(n31885), .Z(n31887) );
  IV U44810 ( .A(n31887), .Z(n31890) );
  NOR U44811 ( .A(n31888), .B(n31890), .Z(n35123) );
  IV U44812 ( .A(n31889), .Z(n31891) );
  NOR U44813 ( .A(n31891), .B(n31890), .Z(n37205) );
  IV U44814 ( .A(n31892), .Z(n31894) );
  IV U44815 ( .A(n31893), .Z(n31898) );
  NOR U44816 ( .A(n31894), .B(n31898), .Z(n37198) );
  IV U44817 ( .A(n31895), .Z(n31896) );
  NOR U44818 ( .A(n31896), .B(n31898), .Z(n37195) );
  IV U44819 ( .A(n31897), .Z(n31899) );
  NOR U44820 ( .A(n31899), .B(n31898), .Z(n35127) );
  NOR U44821 ( .A(n31901), .B(n31900), .Z(n31902) );
  IV U44822 ( .A(n31902), .Z(n35132) );
  NOR U44823 ( .A(n35132), .B(n31903), .Z(n33856) );
  NOR U44824 ( .A(n31905), .B(n31904), .Z(n31906) );
  IV U44825 ( .A(n31906), .Z(n31908) );
  IV U44826 ( .A(n31907), .Z(n35140) );
  NOR U44827 ( .A(n31908), .B(n35140), .Z(n33855) );
  IV U44828 ( .A(n31909), .Z(n31915) );
  IV U44829 ( .A(n31910), .Z(n33848) );
  XOR U44830 ( .A(n31911), .B(n33848), .Z(n31912) );
  NOR U44831 ( .A(n31913), .B(n31912), .Z(n31914) );
  IV U44832 ( .A(n31914), .Z(n31917) );
  NOR U44833 ( .A(n31915), .B(n31917), .Z(n37187) );
  IV U44834 ( .A(n31916), .Z(n31918) );
  NOR U44835 ( .A(n31918), .B(n31917), .Z(n37184) );
  NOR U44836 ( .A(n31920), .B(n31919), .Z(n35143) );
  IV U44837 ( .A(n31921), .Z(n31924) );
  NOR U44838 ( .A(n31922), .B(n33848), .Z(n31923) );
  IV U44839 ( .A(n31923), .Z(n33851) );
  NOR U44840 ( .A(n31924), .B(n33851), .Z(n40213) );
  NOR U44841 ( .A(n38437), .B(n40213), .Z(n37179) );
  IV U44842 ( .A(n31925), .Z(n35157) );
  IV U44843 ( .A(n31926), .Z(n31927) );
  NOR U44844 ( .A(n31929), .B(n31927), .Z(n35159) );
  IV U44845 ( .A(n31928), .Z(n31930) );
  NOR U44846 ( .A(n31930), .B(n31929), .Z(n37174) );
  NOR U44847 ( .A(n35159), .B(n37174), .Z(n33836) );
  IV U44848 ( .A(n31931), .Z(n31938) );
  IV U44849 ( .A(n31932), .Z(n31933) );
  NOR U44850 ( .A(n31938), .B(n31933), .Z(n37171) );
  IV U44851 ( .A(n31934), .Z(n31935) );
  NOR U44852 ( .A(n31935), .B(n31938), .Z(n35167) );
  IV U44853 ( .A(n31936), .Z(n31937) );
  NOR U44854 ( .A(n31938), .B(n31937), .Z(n35164) );
  IV U44855 ( .A(n31939), .Z(n31940) );
  NOR U44856 ( .A(n31940), .B(n33812), .Z(n35175) );
  IV U44857 ( .A(n31941), .Z(n31942) );
  NOR U44858 ( .A(n31943), .B(n31942), .Z(n35188) );
  IV U44859 ( .A(n31944), .Z(n31947) );
  IV U44860 ( .A(n31945), .Z(n31946) );
  NOR U44861 ( .A(n31947), .B(n31946), .Z(n37122) );
  IV U44862 ( .A(n31948), .Z(n31952) );
  NOR U44863 ( .A(n31950), .B(n31949), .Z(n31951) );
  IV U44864 ( .A(n31951), .Z(n33800) );
  NOR U44865 ( .A(n31952), .B(n33800), .Z(n35197) );
  IV U44866 ( .A(n31953), .Z(n31954) );
  NOR U44867 ( .A(n31957), .B(n31954), .Z(n37114) );
  IV U44868 ( .A(n31955), .Z(n31956) );
  NOR U44869 ( .A(n31957), .B(n31956), .Z(n35200) );
  NOR U44870 ( .A(n37114), .B(n35200), .Z(n31958) );
  IV U44871 ( .A(n31958), .Z(n33798) );
  IV U44872 ( .A(n31959), .Z(n31963) );
  IV U44873 ( .A(n31960), .Z(n31961) );
  NOR U44874 ( .A(n31963), .B(n31961), .Z(n37099) );
  IV U44875 ( .A(n31962), .Z(n31964) );
  NOR U44876 ( .A(n31964), .B(n31963), .Z(n37096) );
  IV U44877 ( .A(n31965), .Z(n31968) );
  NOR U44878 ( .A(n31966), .B(n33795), .Z(n31967) );
  IV U44879 ( .A(n31967), .Z(n31970) );
  NOR U44880 ( .A(n31968), .B(n31970), .Z(n35202) );
  IV U44881 ( .A(n31969), .Z(n31971) );
  NOR U44882 ( .A(n31971), .B(n31970), .Z(n37090) );
  IV U44883 ( .A(n31972), .Z(n31973) );
  NOR U44884 ( .A(n31974), .B(n31973), .Z(n37080) );
  IV U44885 ( .A(n31975), .Z(n31977) );
  NOR U44886 ( .A(n31977), .B(n31976), .Z(n35208) );
  NOR U44887 ( .A(n37080), .B(n35208), .Z(n33791) );
  IV U44888 ( .A(n31978), .Z(n31979) );
  NOR U44889 ( .A(n31985), .B(n31979), .Z(n35214) );
  NOR U44890 ( .A(n37083), .B(n35214), .Z(n33790) );
  IV U44891 ( .A(n31980), .Z(n31982) );
  NOR U44892 ( .A(n31982), .B(n31981), .Z(n35219) );
  IV U44893 ( .A(n31983), .Z(n31984) );
  NOR U44894 ( .A(n31985), .B(n31984), .Z(n35216) );
  NOR U44895 ( .A(n35219), .B(n35216), .Z(n33789) );
  NOR U44896 ( .A(n31986), .B(n31989), .Z(n31987) );
  IV U44897 ( .A(n31987), .Z(n35225) );
  NOR U44898 ( .A(n35225), .B(n35227), .Z(n33788) );
  IV U44899 ( .A(n31988), .Z(n31990) );
  NOR U44900 ( .A(n31990), .B(n31989), .Z(n31991) );
  IV U44901 ( .A(n31991), .Z(n31992) );
  NOR U44902 ( .A(n31993), .B(n31992), .Z(n35233) );
  IV U44903 ( .A(n31993), .Z(n31998) );
  NOR U44904 ( .A(n31995), .B(n31994), .Z(n31996) );
  IV U44905 ( .A(n31996), .Z(n31997) );
  NOR U44906 ( .A(n31998), .B(n31997), .Z(n35230) );
  IV U44907 ( .A(n31999), .Z(n32002) );
  NOR U44908 ( .A(n32000), .B(n33782), .Z(n32001) );
  IV U44909 ( .A(n32001), .Z(n33785) );
  NOR U44910 ( .A(n32002), .B(n33785), .Z(n35236) );
  IV U44911 ( .A(n32003), .Z(n32005) );
  IV U44912 ( .A(n32004), .Z(n32010) );
  NOR U44913 ( .A(n32005), .B(n32010), .Z(n32006) );
  IV U44914 ( .A(n32006), .Z(n35239) );
  NOR U44915 ( .A(n32007), .B(n35255), .Z(n32011) );
  IV U44916 ( .A(n32008), .Z(n32009) );
  NOR U44917 ( .A(n32010), .B(n32009), .Z(n35241) );
  NOR U44918 ( .A(n32011), .B(n35241), .Z(n32012) );
  IV U44919 ( .A(n32012), .Z(n33780) );
  IV U44920 ( .A(n32013), .Z(n32014) );
  NOR U44921 ( .A(n32014), .B(n35245), .Z(n35251) );
  NOR U44922 ( .A(n32018), .B(n32015), .Z(n32016) );
  IV U44923 ( .A(n32016), .Z(n37064) );
  IV U44924 ( .A(n32017), .Z(n32019) );
  NOR U44925 ( .A(n32019), .B(n32018), .Z(n37059) );
  IV U44926 ( .A(n32020), .Z(n32023) );
  NOR U44927 ( .A(n32021), .B(n32025), .Z(n32022) );
  IV U44928 ( .A(n32022), .Z(n33772) );
  NOR U44929 ( .A(n32023), .B(n33772), .Z(n35259) );
  IV U44930 ( .A(n32024), .Z(n32026) );
  NOR U44931 ( .A(n32026), .B(n32025), .Z(n35267) );
  IV U44932 ( .A(n32027), .Z(n32029) );
  NOR U44933 ( .A(n32029), .B(n32028), .Z(n35262) );
  NOR U44934 ( .A(n35267), .B(n35262), .Z(n33770) );
  IV U44935 ( .A(n32030), .Z(n32032) );
  NOR U44936 ( .A(n32032), .B(n32031), .Z(n32033) );
  IV U44937 ( .A(n32033), .Z(n33754) );
  NOR U44938 ( .A(n32034), .B(n35280), .Z(n33747) );
  IV U44939 ( .A(n32035), .Z(n32036) );
  NOR U44940 ( .A(n32037), .B(n32036), .Z(n40132) );
  IV U44941 ( .A(n32038), .Z(n32039) );
  NOR U44942 ( .A(n32040), .B(n32039), .Z(n40138) );
  NOR U44943 ( .A(n40132), .B(n40138), .Z(n37034) );
  IV U44944 ( .A(n32041), .Z(n32042) );
  NOR U44945 ( .A(n32044), .B(n32042), .Z(n37031) );
  IV U44946 ( .A(n32043), .Z(n32045) );
  NOR U44947 ( .A(n32045), .B(n32044), .Z(n37027) );
  IV U44948 ( .A(n32046), .Z(n32047) );
  NOR U44949 ( .A(n32048), .B(n32047), .Z(n37024) );
  IV U44950 ( .A(n32049), .Z(n38592) );
  IV U44951 ( .A(n32050), .Z(n32051) );
  NOR U44952 ( .A(n38592), .B(n32051), .Z(n37020) );
  NOR U44953 ( .A(n37024), .B(n37020), .Z(n32052) );
  IV U44954 ( .A(n32052), .Z(n33742) );
  IV U44955 ( .A(n32053), .Z(n32055) );
  NOR U44956 ( .A(n32055), .B(n32054), .Z(n32056) );
  IV U44957 ( .A(n32056), .Z(n33729) );
  IV U44958 ( .A(n32057), .Z(n32059) );
  IV U44959 ( .A(n32058), .Z(n33715) );
  NOR U44960 ( .A(n32059), .B(n33715), .Z(n35292) );
  IV U44961 ( .A(n32060), .Z(n32061) );
  NOR U44962 ( .A(n32061), .B(n33715), .Z(n32062) );
  IV U44963 ( .A(n32062), .Z(n32063) );
  NOR U44964 ( .A(n33714), .B(n32063), .Z(n35294) );
  NOR U44965 ( .A(n35292), .B(n35294), .Z(n33721) );
  IV U44966 ( .A(n32064), .Z(n32066) );
  IV U44967 ( .A(n32065), .Z(n33701) );
  NOR U44968 ( .A(n32066), .B(n33701), .Z(n37003) );
  IV U44969 ( .A(n32067), .Z(n32069) );
  IV U44970 ( .A(n32068), .Z(n33704) );
  NOR U44971 ( .A(n32069), .B(n33704), .Z(n40094) );
  IV U44972 ( .A(n33708), .Z(n32073) );
  NOR U44973 ( .A(n32070), .B(n33704), .Z(n32071) );
  IV U44974 ( .A(n32071), .Z(n32072) );
  NOR U44975 ( .A(n32073), .B(n32072), .Z(n40107) );
  NOR U44976 ( .A(n40094), .B(n40107), .Z(n35307) );
  IV U44977 ( .A(n32074), .Z(n32076) );
  IV U44978 ( .A(n32075), .Z(n35315) );
  NOR U44979 ( .A(n32076), .B(n35315), .Z(n33694) );
  IV U44980 ( .A(n32077), .Z(n32078) );
  NOR U44981 ( .A(n32078), .B(n32083), .Z(n35322) );
  NOR U44982 ( .A(n32079), .B(n35315), .Z(n36991) );
  NOR U44983 ( .A(n35322), .B(n36991), .Z(n33693) );
  IV U44984 ( .A(n32080), .Z(n35329) );
  XOR U44985 ( .A(n32082), .B(n32083), .Z(n32081) );
  NOR U44986 ( .A(n35329), .B(n32081), .Z(n33692) );
  IV U44987 ( .A(n32082), .Z(n32084) );
  NOR U44988 ( .A(n32084), .B(n32083), .Z(n33689) );
  IV U44989 ( .A(n33689), .Z(n33678) );
  IV U44990 ( .A(n32085), .Z(n32086) );
  NOR U44991 ( .A(n32086), .B(n35336), .Z(n33677) );
  IV U44992 ( .A(n32087), .Z(n32090) );
  NOR U44993 ( .A(n32088), .B(n32093), .Z(n32089) );
  IV U44994 ( .A(n32089), .Z(n33633) );
  NOR U44995 ( .A(n32090), .B(n33633), .Z(n35371) );
  IV U44996 ( .A(n32091), .Z(n32092) );
  NOR U44997 ( .A(n32093), .B(n32092), .Z(n36967) );
  IV U44998 ( .A(n32094), .Z(n32096) );
  NOR U44999 ( .A(n32096), .B(n32095), .Z(n35376) );
  IV U45000 ( .A(n32097), .Z(n32098) );
  NOR U45001 ( .A(n32099), .B(n32098), .Z(n35374) );
  NOR U45002 ( .A(n35376), .B(n35374), .Z(n32100) );
  IV U45003 ( .A(n32100), .Z(n33631) );
  IV U45004 ( .A(n32101), .Z(n32102) );
  NOR U45005 ( .A(n32105), .B(n32102), .Z(n35382) );
  IV U45006 ( .A(n32103), .Z(n32104) );
  NOR U45007 ( .A(n32105), .B(n32104), .Z(n35379) );
  IV U45008 ( .A(n32106), .Z(n32114) );
  XOR U45009 ( .A(n32108), .B(n32107), .Z(n32111) );
  IV U45010 ( .A(n32109), .Z(n33625) );
  XOR U45011 ( .A(n33616), .B(n33625), .Z(n32110) );
  NOR U45012 ( .A(n32111), .B(n32110), .Z(n32112) );
  IV U45013 ( .A(n32112), .Z(n32113) );
  NOR U45014 ( .A(n32114), .B(n32113), .Z(n33620) );
  IV U45015 ( .A(n32115), .Z(n32116) );
  NOR U45016 ( .A(n32116), .B(n35394), .Z(n33615) );
  IV U45017 ( .A(n32117), .Z(n32119) );
  NOR U45018 ( .A(n32119), .B(n32118), .Z(n35412) );
  IV U45019 ( .A(n32120), .Z(n32122) );
  NOR U45020 ( .A(n32122), .B(n32121), .Z(n36959) );
  NOR U45021 ( .A(n35412), .B(n36959), .Z(n33608) );
  NOR U45022 ( .A(n32124), .B(n32123), .Z(n35414) );
  IV U45023 ( .A(n32125), .Z(n35421) );
  IV U45024 ( .A(n32126), .Z(n32128) );
  NOR U45025 ( .A(n32128), .B(n32127), .Z(n35428) );
  IV U45026 ( .A(n32129), .Z(n32130) );
  NOR U45027 ( .A(n32130), .B(n32135), .Z(n32131) );
  IV U45028 ( .A(n32131), .Z(n35426) );
  IV U45029 ( .A(n32132), .Z(n32133) );
  NOR U45030 ( .A(n32133), .B(n33597), .Z(n35431) );
  IV U45031 ( .A(n32134), .Z(n32136) );
  NOR U45032 ( .A(n32136), .B(n32135), .Z(n36936) );
  NOR U45033 ( .A(n35431), .B(n36936), .Z(n33595) );
  IV U45034 ( .A(n32137), .Z(n32138) );
  NOR U45035 ( .A(n32138), .B(n33590), .Z(n35438) );
  IV U45036 ( .A(n32139), .Z(n32142) );
  IV U45037 ( .A(n32140), .Z(n32141) );
  NOR U45038 ( .A(n32142), .B(n32141), .Z(n35436) );
  NOR U45039 ( .A(n35438), .B(n35436), .Z(n33585) );
  IV U45040 ( .A(n32143), .Z(n32147) );
  IV U45041 ( .A(n32144), .Z(n33583) );
  NOR U45042 ( .A(n32145), .B(n33583), .Z(n32146) );
  IV U45043 ( .A(n32146), .Z(n32149) );
  NOR U45044 ( .A(n32147), .B(n32149), .Z(n35444) );
  IV U45045 ( .A(n32148), .Z(n32150) );
  NOR U45046 ( .A(n32150), .B(n32149), .Z(n35441) );
  IV U45047 ( .A(n33567), .Z(n32151) );
  NOR U45048 ( .A(n33580), .B(n32151), .Z(n32152) );
  IV U45049 ( .A(n32152), .Z(n33575) );
  IV U45050 ( .A(n32153), .Z(n32154) );
  NOR U45051 ( .A(n32159), .B(n32154), .Z(n35463) );
  IV U45052 ( .A(n32155), .Z(n32156) );
  NOR U45053 ( .A(n32159), .B(n32156), .Z(n35460) );
  IV U45054 ( .A(n32157), .Z(n32158) );
  NOR U45055 ( .A(n32159), .B(n32158), .Z(n35466) );
  IV U45056 ( .A(n32160), .Z(n32161) );
  NOR U45057 ( .A(n32161), .B(n32163), .Z(n35472) );
  IV U45058 ( .A(n32162), .Z(n32164) );
  NOR U45059 ( .A(n32164), .B(n32163), .Z(n35469) );
  IV U45060 ( .A(n32165), .Z(n32170) );
  IV U45061 ( .A(n32166), .Z(n32167) );
  NOR U45062 ( .A(n32168), .B(n32167), .Z(n32169) );
  IV U45063 ( .A(n32169), .Z(n33564) );
  NOR U45064 ( .A(n32170), .B(n33564), .Z(n33559) );
  IV U45065 ( .A(n32171), .Z(n32172) );
  NOR U45066 ( .A(n32172), .B(n32177), .Z(n35489) );
  NOR U45067 ( .A(n32174), .B(n32173), .Z(n35487) );
  NOR U45068 ( .A(n35489), .B(n35487), .Z(n33553) );
  NOR U45069 ( .A(n32175), .B(n35496), .Z(n32179) );
  IV U45070 ( .A(n32176), .Z(n32178) );
  NOR U45071 ( .A(n32178), .B(n32177), .Z(n35492) );
  NOR U45072 ( .A(n32179), .B(n35492), .Z(n33552) );
  IV U45073 ( .A(n32180), .Z(n32181) );
  NOR U45074 ( .A(n32182), .B(n32181), .Z(n36907) );
  IV U45075 ( .A(n32183), .Z(n32185) );
  NOR U45076 ( .A(n32185), .B(n32184), .Z(n32186) );
  IV U45077 ( .A(n32186), .Z(n35506) );
  IV U45078 ( .A(n32187), .Z(n32188) );
  NOR U45079 ( .A(n32188), .B(n32193), .Z(n35507) );
  IV U45080 ( .A(n32189), .Z(n32191) );
  NOR U45081 ( .A(n32191), .B(n32190), .Z(n35513) );
  IV U45082 ( .A(n32192), .Z(n32194) );
  NOR U45083 ( .A(n32194), .B(n32193), .Z(n35510) );
  NOR U45084 ( .A(n35513), .B(n35510), .Z(n32195) );
  IV U45085 ( .A(n32195), .Z(n33544) );
  IV U45086 ( .A(n32196), .Z(n33541) );
  IV U45087 ( .A(n32197), .Z(n32198) );
  NOR U45088 ( .A(n33541), .B(n32198), .Z(n35516) );
  NOR U45089 ( .A(n36893), .B(n35522), .Z(n33535) );
  IV U45090 ( .A(n32199), .Z(n32201) );
  NOR U45091 ( .A(n32201), .B(n32200), .Z(n36889) );
  IV U45092 ( .A(n32202), .Z(n32205) );
  NOR U45093 ( .A(n32203), .B(n33526), .Z(n32204) );
  IV U45094 ( .A(n32204), .Z(n33533) );
  NOR U45095 ( .A(n32205), .B(n33533), .Z(n36896) );
  IV U45096 ( .A(n32206), .Z(n32209) );
  NOR U45097 ( .A(n32207), .B(n32211), .Z(n32208) );
  IV U45098 ( .A(n32208), .Z(n32214) );
  NOR U45099 ( .A(n32209), .B(n32214), .Z(n36868) );
  IV U45100 ( .A(n32210), .Z(n32212) );
  NOR U45101 ( .A(n32212), .B(n32211), .Z(n36865) );
  IV U45102 ( .A(n32213), .Z(n32215) );
  NOR U45103 ( .A(n32215), .B(n32214), .Z(n36871) );
  NOR U45104 ( .A(n36865), .B(n36871), .Z(n32216) );
  IV U45105 ( .A(n32216), .Z(n33503) );
  IV U45106 ( .A(n32217), .Z(n32219) );
  NOR U45107 ( .A(n32219), .B(n32218), .Z(n35538) );
  IV U45108 ( .A(n32220), .Z(n32225) );
  IV U45109 ( .A(n32221), .Z(n32222) );
  NOR U45110 ( .A(n32225), .B(n32222), .Z(n35543) );
  IV U45111 ( .A(n32223), .Z(n32224) );
  NOR U45112 ( .A(n32225), .B(n32224), .Z(n35540) );
  IV U45113 ( .A(n32226), .Z(n32230) );
  NOR U45114 ( .A(n32228), .B(n32227), .Z(n32229) );
  IV U45115 ( .A(n32229), .Z(n32232) );
  NOR U45116 ( .A(n32230), .B(n32232), .Z(n35546) );
  IV U45117 ( .A(n32231), .Z(n32233) );
  NOR U45118 ( .A(n32233), .B(n32232), .Z(n36856) );
  XOR U45119 ( .A(n33491), .B(n33492), .Z(n32236) );
  IV U45120 ( .A(n32234), .Z(n32235) );
  NOR U45121 ( .A(n32236), .B(n32235), .Z(n33500) );
  IV U45122 ( .A(n33500), .Z(n42091) );
  IV U45123 ( .A(n32237), .Z(n32238) );
  NOR U45124 ( .A(n32238), .B(n33492), .Z(n36850) );
  IV U45125 ( .A(n32239), .Z(n32240) );
  NOR U45126 ( .A(n42096), .B(n32240), .Z(n32241) );
  IV U45127 ( .A(n32241), .Z(n33487) );
  IV U45128 ( .A(n32242), .Z(n32244) );
  IV U45129 ( .A(n32243), .Z(n33485) );
  NOR U45130 ( .A(n32244), .B(n33485), .Z(n39839) );
  NOR U45131 ( .A(n39834), .B(n39839), .Z(n36838) );
  IV U45132 ( .A(n32245), .Z(n32248) );
  NOR U45133 ( .A(n32253), .B(n32246), .Z(n32247) );
  IV U45134 ( .A(n32247), .Z(n32250) );
  NOR U45135 ( .A(n32248), .B(n32250), .Z(n35556) );
  NOR U45136 ( .A(n35553), .B(n35556), .Z(n33479) );
  IV U45137 ( .A(n32249), .Z(n32251) );
  NOR U45138 ( .A(n32251), .B(n32250), .Z(n35558) );
  IV U45139 ( .A(n32252), .Z(n32256) );
  NOR U45140 ( .A(n32254), .B(n32253), .Z(n32255) );
  IV U45141 ( .A(n32255), .Z(n32261) );
  NOR U45142 ( .A(n32256), .B(n32261), .Z(n35560) );
  NOR U45143 ( .A(n35558), .B(n35560), .Z(n33478) );
  IV U45144 ( .A(n32257), .Z(n32258) );
  NOR U45145 ( .A(n32259), .B(n32258), .Z(n36831) );
  IV U45146 ( .A(n32260), .Z(n32262) );
  NOR U45147 ( .A(n32262), .B(n32261), .Z(n36834) );
  NOR U45148 ( .A(n36831), .B(n36834), .Z(n33477) );
  IV U45149 ( .A(n32263), .Z(n32266) );
  IV U45150 ( .A(n32264), .Z(n32265) );
  NOR U45151 ( .A(n32266), .B(n32265), .Z(n36828) );
  NOR U45152 ( .A(n32267), .B(n32271), .Z(n32268) );
  IV U45153 ( .A(n32268), .Z(n36815) );
  NOR U45154 ( .A(n32269), .B(n36815), .Z(n33476) );
  NOR U45155 ( .A(n32271), .B(n32270), .Z(n36811) );
  IV U45156 ( .A(n32272), .Z(n32273) );
  NOR U45157 ( .A(n32275), .B(n32273), .Z(n36807) );
  IV U45158 ( .A(n32274), .Z(n32276) );
  NOR U45159 ( .A(n32276), .B(n32275), .Z(n36804) );
  IV U45160 ( .A(n32277), .Z(n32280) );
  NOR U45161 ( .A(n32278), .B(n33463), .Z(n32279) );
  IV U45162 ( .A(n32279), .Z(n33474) );
  NOR U45163 ( .A(n32280), .B(n33474), .Z(n35566) );
  IV U45164 ( .A(n32281), .Z(n32283) );
  XOR U45165 ( .A(n32284), .B(n33466), .Z(n32282) );
  NOR U45166 ( .A(n32283), .B(n32282), .Z(n35573) );
  IV U45167 ( .A(n32284), .Z(n32285) );
  NOR U45168 ( .A(n32285), .B(n33466), .Z(n33459) );
  IV U45169 ( .A(n33459), .Z(n33453) );
  IV U45170 ( .A(n32286), .Z(n32289) );
  IV U45171 ( .A(n32287), .Z(n33455) );
  XOR U45172 ( .A(n33450), .B(n33455), .Z(n32288) );
  NOR U45173 ( .A(n32289), .B(n32288), .Z(n35576) );
  IV U45174 ( .A(n32290), .Z(n32291) );
  NOR U45175 ( .A(n33438), .B(n32291), .Z(n32292) );
  IV U45176 ( .A(n32292), .Z(n35580) );
  IV U45177 ( .A(n32293), .Z(n32294) );
  NOR U45178 ( .A(n33432), .B(n32294), .Z(n35585) );
  IV U45179 ( .A(n32295), .Z(n32298) );
  NOR U45180 ( .A(n32296), .B(n32301), .Z(n32297) );
  IV U45181 ( .A(n32297), .Z(n33428) );
  NOR U45182 ( .A(n32298), .B(n33428), .Z(n32299) );
  IV U45183 ( .A(n32299), .Z(n36759) );
  NOR U45184 ( .A(n32301), .B(n32300), .Z(n35588) );
  IV U45185 ( .A(n32302), .Z(n36744) );
  IV U45186 ( .A(n32303), .Z(n32304) );
  NOR U45187 ( .A(n36744), .B(n32304), .Z(n35593) );
  NOR U45188 ( .A(n35588), .B(n35593), .Z(n33425) );
  IV U45189 ( .A(n32305), .Z(n32306) );
  NOR U45190 ( .A(n32306), .B(n36744), .Z(n36751) );
  IV U45191 ( .A(n32307), .Z(n32308) );
  NOR U45192 ( .A(n32308), .B(n33419), .Z(n35596) );
  IV U45193 ( .A(n32309), .Z(n32313) );
  IV U45194 ( .A(n32310), .Z(n32315) );
  NOR U45195 ( .A(n32311), .B(n32315), .Z(n32312) );
  IV U45196 ( .A(n32312), .Z(n33411) );
  NOR U45197 ( .A(n32313), .B(n33411), .Z(n36725) );
  IV U45198 ( .A(n32314), .Z(n32316) );
  NOR U45199 ( .A(n32316), .B(n32315), .Z(n32317) );
  IV U45200 ( .A(n32317), .Z(n32318) );
  NOR U45201 ( .A(n32319), .B(n32318), .Z(n36721) );
  IV U45202 ( .A(n32319), .Z(n32324) );
  IV U45203 ( .A(n32320), .Z(n32327) );
  NOR U45204 ( .A(n32321), .B(n32327), .Z(n32322) );
  IV U45205 ( .A(n32322), .Z(n32323) );
  NOR U45206 ( .A(n32324), .B(n32323), .Z(n36718) );
  IV U45207 ( .A(n32325), .Z(n32326) );
  NOR U45208 ( .A(n32327), .B(n32326), .Z(n36713) );
  NOR U45209 ( .A(n35601), .B(n36713), .Z(n33406) );
  NOR U45210 ( .A(n32328), .B(n33377), .Z(n43226) );
  IV U45211 ( .A(n32329), .Z(n32332) );
  IV U45212 ( .A(n32330), .Z(n32331) );
  NOR U45213 ( .A(n32332), .B(n32331), .Z(n42199) );
  NOR U45214 ( .A(n43226), .B(n42199), .Z(n35625) );
  IV U45215 ( .A(n32333), .Z(n32336) );
  NOR U45216 ( .A(n32334), .B(n32337), .Z(n32335) );
  IV U45217 ( .A(n32335), .Z(n32340) );
  NOR U45218 ( .A(n32336), .B(n32340), .Z(n35638) );
  NOR U45219 ( .A(n32338), .B(n32337), .Z(n35649) );
  IV U45220 ( .A(n32339), .Z(n32341) );
  NOR U45221 ( .A(n32341), .B(n32340), .Z(n35644) );
  NOR U45222 ( .A(n35649), .B(n35644), .Z(n32342) );
  IV U45223 ( .A(n32342), .Z(n33352) );
  IV U45224 ( .A(n32343), .Z(n32345) );
  XOR U45225 ( .A(n33337), .B(n33346), .Z(n32344) );
  NOR U45226 ( .A(n32345), .B(n32344), .Z(n33341) );
  IV U45227 ( .A(n32346), .Z(n32350) );
  NOR U45228 ( .A(n32348), .B(n32347), .Z(n32349) );
  IV U45229 ( .A(n32349), .Z(n33325) );
  NOR U45230 ( .A(n32350), .B(n33325), .Z(n32351) );
  IV U45231 ( .A(n32351), .Z(n35659) );
  IV U45232 ( .A(n32352), .Z(n32353) );
  NOR U45233 ( .A(n32354), .B(n32353), .Z(n32355) );
  IV U45234 ( .A(n32355), .Z(n32356) );
  NOR U45235 ( .A(n32356), .B(n32363), .Z(n35669) );
  IV U45236 ( .A(n32357), .Z(n32358) );
  NOR U45237 ( .A(n32358), .B(n32363), .Z(n35666) );
  IV U45238 ( .A(n32359), .Z(n43196) );
  NOR U45239 ( .A(n32360), .B(n43196), .Z(n38870) );
  IV U45240 ( .A(n32361), .Z(n32362) );
  NOR U45241 ( .A(n32363), .B(n32362), .Z(n38866) );
  NOR U45242 ( .A(n38870), .B(n38866), .Z(n35672) );
  IV U45243 ( .A(n35672), .Z(n33323) );
  IV U45244 ( .A(n32364), .Z(n32367) );
  NOR U45245 ( .A(n32365), .B(n32373), .Z(n32366) );
  IV U45246 ( .A(n32366), .Z(n32369) );
  NOR U45247 ( .A(n32367), .B(n32369), .Z(n35684) );
  IV U45248 ( .A(n32368), .Z(n32370) );
  NOR U45249 ( .A(n32370), .B(n32369), .Z(n36663) );
  IV U45250 ( .A(n32371), .Z(n32372) );
  NOR U45251 ( .A(n32373), .B(n32372), .Z(n36660) );
  IV U45252 ( .A(n32374), .Z(n32375) );
  NOR U45253 ( .A(n32376), .B(n32375), .Z(n35687) );
  IV U45254 ( .A(n32377), .Z(n32388) );
  IV U45255 ( .A(n32378), .Z(n32379) );
  NOR U45256 ( .A(n32380), .B(n32379), .Z(n32386) );
  IV U45257 ( .A(n32381), .Z(n35700) );
  XOR U45258 ( .A(n35700), .B(n32393), .Z(n32382) );
  NOR U45259 ( .A(n32383), .B(n32382), .Z(n32384) );
  IV U45260 ( .A(n32384), .Z(n32385) );
  NOR U45261 ( .A(n32386), .B(n32385), .Z(n32387) );
  IV U45262 ( .A(n32387), .Z(n32390) );
  NOR U45263 ( .A(n32388), .B(n32390), .Z(n36651) );
  IV U45264 ( .A(n32389), .Z(n32391) );
  NOR U45265 ( .A(n32391), .B(n32390), .Z(n36648) );
  IV U45266 ( .A(n32392), .Z(n32396) );
  IV U45267 ( .A(n32393), .Z(n33316) );
  NOR U45268 ( .A(n32394), .B(n33316), .Z(n32395) );
  IV U45269 ( .A(n32395), .Z(n33320) );
  NOR U45270 ( .A(n32396), .B(n33320), .Z(n35690) );
  IV U45271 ( .A(n33311), .Z(n48954) );
  IV U45272 ( .A(n32397), .Z(n32398) );
  NOR U45273 ( .A(n32398), .B(n33299), .Z(n35707) );
  IV U45274 ( .A(n32399), .Z(n32402) );
  IV U45275 ( .A(n32400), .Z(n32401) );
  NOR U45276 ( .A(n32402), .B(n32401), .Z(n38898) );
  NOR U45277 ( .A(n38902), .B(n38898), .Z(n36635) );
  IV U45278 ( .A(n32403), .Z(n32405) );
  NOR U45279 ( .A(n32405), .B(n32404), .Z(n35711) );
  IV U45280 ( .A(n32406), .Z(n32407) );
  NOR U45281 ( .A(n32414), .B(n32407), .Z(n32408) );
  IV U45282 ( .A(n32408), .Z(n35716) );
  IV U45283 ( .A(n32409), .Z(n32410) );
  NOR U45284 ( .A(n32411), .B(n32410), .Z(n35725) );
  IV U45285 ( .A(n32412), .Z(n32413) );
  NOR U45286 ( .A(n32414), .B(n32413), .Z(n35720) );
  NOR U45287 ( .A(n35725), .B(n35720), .Z(n32415) );
  IV U45288 ( .A(n32415), .Z(n33291) );
  IV U45289 ( .A(n32416), .Z(n32418) );
  IV U45290 ( .A(n32417), .Z(n33289) );
  NOR U45291 ( .A(n32418), .B(n33289), .Z(n35722) );
  NOR U45292 ( .A(n33281), .B(n39657), .Z(n32419) );
  NOR U45293 ( .A(n32419), .B(n38922), .Z(n32420) );
  IV U45294 ( .A(n32420), .Z(n36625) );
  IV U45295 ( .A(n32421), .Z(n32422) );
  NOR U45296 ( .A(n32423), .B(n32422), .Z(n32424) );
  IV U45297 ( .A(n32424), .Z(n33277) );
  NOR U45298 ( .A(n32425), .B(n42328), .Z(n35738) );
  NOR U45299 ( .A(n35736), .B(n35738), .Z(n33274) );
  IV U45300 ( .A(n32426), .Z(n32430) );
  NOR U45301 ( .A(n32428), .B(n32427), .Z(n32429) );
  IV U45302 ( .A(n32429), .Z(n33263) );
  NOR U45303 ( .A(n32430), .B(n33263), .Z(n35745) );
  IV U45304 ( .A(n32431), .Z(n32435) );
  NOR U45305 ( .A(n32433), .B(n32432), .Z(n32434) );
  IV U45306 ( .A(n32434), .Z(n33245) );
  NOR U45307 ( .A(n32435), .B(n33245), .Z(n36602) );
  IV U45308 ( .A(n32436), .Z(n32440) );
  IV U45309 ( .A(n32437), .Z(n33225) );
  NOR U45310 ( .A(n32438), .B(n33225), .Z(n32439) );
  IV U45311 ( .A(n32439), .Z(n32442) );
  NOR U45312 ( .A(n32440), .B(n32442), .Z(n35766) );
  IV U45313 ( .A(n32441), .Z(n32443) );
  NOR U45314 ( .A(n32443), .B(n32442), .Z(n35772) );
  NOR U45315 ( .A(n35766), .B(n35772), .Z(n33232) );
  IV U45316 ( .A(n32444), .Z(n32445) );
  NOR U45317 ( .A(n33222), .B(n32445), .Z(n36578) );
  IV U45318 ( .A(n32446), .Z(n32447) );
  NOR U45319 ( .A(n32447), .B(n36561), .Z(n33221) );
  IV U45320 ( .A(n32448), .Z(n32449) );
  NOR U45321 ( .A(n32449), .B(n36561), .Z(n35776) );
  IV U45322 ( .A(n32450), .Z(n32453) );
  NOR U45323 ( .A(n32451), .B(n33207), .Z(n32452) );
  IV U45324 ( .A(n32452), .Z(n32455) );
  NOR U45325 ( .A(n32453), .B(n32455), .Z(n35783) );
  IV U45326 ( .A(n32454), .Z(n32456) );
  NOR U45327 ( .A(n32456), .B(n32455), .Z(n32457) );
  IV U45328 ( .A(n32457), .Z(n35790) );
  IV U45329 ( .A(n33187), .Z(n32458) );
  NOR U45330 ( .A(n32458), .B(n33197), .Z(n32459) );
  IV U45331 ( .A(n32459), .Z(n33192) );
  IV U45332 ( .A(n32460), .Z(n42379) );
  IV U45333 ( .A(n32463), .Z(n32461) );
  NOR U45334 ( .A(n42379), .B(n32461), .Z(n38989) );
  IV U45335 ( .A(n32462), .Z(n32465) );
  XOR U45336 ( .A(n42379), .B(n32463), .Z(n32464) );
  NOR U45337 ( .A(n32465), .B(n32464), .Z(n38984) );
  NOR U45338 ( .A(n38989), .B(n38984), .Z(n36539) );
  IV U45339 ( .A(n36539), .Z(n33185) );
  IV U45340 ( .A(n32466), .Z(n32467) );
  NOR U45341 ( .A(n32467), .B(n33183), .Z(n35804) );
  IV U45342 ( .A(n32468), .Z(n32470) );
  NOR U45343 ( .A(n32470), .B(n32469), .Z(n39002) );
  IV U45344 ( .A(n32471), .Z(n32472) );
  NOR U45345 ( .A(n32472), .B(n33183), .Z(n38993) );
  NOR U45346 ( .A(n39002), .B(n38993), .Z(n35808) );
  IV U45347 ( .A(n32473), .Z(n35810) );
  NOR U45348 ( .A(n32474), .B(n35810), .Z(n33180) );
  IV U45349 ( .A(n32475), .Z(n32478) );
  NOR U45350 ( .A(n32476), .B(n32484), .Z(n32477) );
  IV U45351 ( .A(n32477), .Z(n32480) );
  NOR U45352 ( .A(n32478), .B(n32480), .Z(n35819) );
  IV U45353 ( .A(n32479), .Z(n32481) );
  NOR U45354 ( .A(n32481), .B(n32480), .Z(n35816) );
  IV U45355 ( .A(n32482), .Z(n32483) );
  NOR U45356 ( .A(n32484), .B(n32483), .Z(n36522) );
  XOR U45357 ( .A(n32492), .B(n35831), .Z(n32487) );
  IV U45358 ( .A(n32485), .Z(n32486) );
  NOR U45359 ( .A(n32487), .B(n32486), .Z(n36519) );
  IV U45360 ( .A(n32488), .Z(n32489) );
  NOR U45361 ( .A(n35831), .B(n32489), .Z(n35822) );
  IV U45362 ( .A(n32490), .Z(n32491) );
  NOR U45363 ( .A(n35831), .B(n32491), .Z(n35826) );
  IV U45364 ( .A(n32492), .Z(n32493) );
  NOR U45365 ( .A(n35831), .B(n32493), .Z(n33179) );
  IV U45366 ( .A(n32494), .Z(n32498) );
  IV U45367 ( .A(n32495), .Z(n33173) );
  NOR U45368 ( .A(n32496), .B(n33173), .Z(n32497) );
  IV U45369 ( .A(n32497), .Z(n32500) );
  NOR U45370 ( .A(n32498), .B(n32500), .Z(n35844) );
  IV U45371 ( .A(n32499), .Z(n32501) );
  NOR U45372 ( .A(n32501), .B(n32500), .Z(n35841) );
  IV U45373 ( .A(n32502), .Z(n32505) );
  NOR U45374 ( .A(n33177), .B(n32503), .Z(n32504) );
  IV U45375 ( .A(n32504), .Z(n33170) );
  NOR U45376 ( .A(n32505), .B(n33170), .Z(n33165) );
  IV U45377 ( .A(n32506), .Z(n33157) );
  IV U45378 ( .A(n32507), .Z(n32508) );
  NOR U45379 ( .A(n33157), .B(n32508), .Z(n35857) );
  NOR U45380 ( .A(n32510), .B(n32509), .Z(n33147) );
  NOR U45381 ( .A(n32512), .B(n32511), .Z(n32513) );
  IV U45382 ( .A(n32513), .Z(n33137) );
  IV U45383 ( .A(n32514), .Z(n33130) );
  NOR U45384 ( .A(n33130), .B(n35870), .Z(n33128) );
  IV U45385 ( .A(n32515), .Z(n32520) );
  IV U45386 ( .A(n32516), .Z(n32517) );
  NOR U45387 ( .A(n32518), .B(n32517), .Z(n32519) );
  IV U45388 ( .A(n32519), .Z(n33120) );
  NOR U45389 ( .A(n32520), .B(n33120), .Z(n35882) );
  IV U45390 ( .A(n32521), .Z(n32522) );
  NOR U45391 ( .A(n35892), .B(n32522), .Z(n32523) );
  NOR U45392 ( .A(n36504), .B(n32523), .Z(n32524) );
  IV U45393 ( .A(n32524), .Z(n33118) );
  IV U45394 ( .A(n32525), .Z(n32528) );
  NOR U45395 ( .A(n32526), .B(n32537), .Z(n32527) );
  IV U45396 ( .A(n32527), .Z(n32530) );
  NOR U45397 ( .A(n32528), .B(n32530), .Z(n36494) );
  IV U45398 ( .A(n32529), .Z(n32531) );
  NOR U45399 ( .A(n32531), .B(n32530), .Z(n35893) );
  IV U45400 ( .A(n32532), .Z(n32533) );
  NOR U45401 ( .A(n32533), .B(n32537), .Z(n32534) );
  IV U45402 ( .A(n32534), .Z(n32535) );
  NOR U45403 ( .A(n32536), .B(n32535), .Z(n36490) );
  IV U45404 ( .A(n32536), .Z(n32541) );
  NOR U45405 ( .A(n32538), .B(n32537), .Z(n32539) );
  IV U45406 ( .A(n32539), .Z(n32540) );
  NOR U45407 ( .A(n32541), .B(n32540), .Z(n36487) );
  IV U45408 ( .A(n32542), .Z(n35900) );
  IV U45409 ( .A(n32543), .Z(n32544) );
  NOR U45410 ( .A(n32546), .B(n32544), .Z(n35896) );
  IV U45411 ( .A(n32545), .Z(n32547) );
  NOR U45412 ( .A(n32547), .B(n32546), .Z(n36479) );
  NOR U45413 ( .A(n32548), .B(n35901), .Z(n32549) );
  NOR U45414 ( .A(n32549), .B(n36473), .Z(n32550) );
  IV U45415 ( .A(n32550), .Z(n33092) );
  IV U45416 ( .A(n32551), .Z(n32552) );
  NOR U45417 ( .A(n32552), .B(n32557), .Z(n32553) );
  IV U45418 ( .A(n32553), .Z(n35919) );
  IV U45419 ( .A(n32554), .Z(n32555) );
  NOR U45420 ( .A(n32555), .B(n32557), .Z(n35915) );
  IV U45421 ( .A(n32556), .Z(n32558) );
  NOR U45422 ( .A(n32558), .B(n32557), .Z(n36462) );
  IV U45423 ( .A(n32559), .Z(n32564) );
  NOR U45424 ( .A(n32561), .B(n32560), .Z(n32562) );
  IV U45425 ( .A(n32562), .Z(n32563) );
  NOR U45426 ( .A(n32564), .B(n32563), .Z(n35920) );
  NOR U45427 ( .A(n36462), .B(n35920), .Z(n32565) );
  IV U45428 ( .A(n32565), .Z(n33083) );
  IV U45429 ( .A(n32566), .Z(n32570) );
  IV U45430 ( .A(n32567), .Z(n32571) );
  NOR U45431 ( .A(n32571), .B(n33080), .Z(n32568) );
  IV U45432 ( .A(n32568), .Z(n32569) );
  NOR U45433 ( .A(n32570), .B(n32569), .Z(n35922) );
  NOR U45434 ( .A(n32572), .B(n32571), .Z(n32573) );
  IV U45435 ( .A(n32573), .Z(n32574) );
  NOR U45436 ( .A(n32574), .B(n33080), .Z(n36458) );
  IV U45437 ( .A(n32575), .Z(n32576) );
  NOR U45438 ( .A(n32576), .B(n32581), .Z(n36451) );
  IV U45439 ( .A(n32577), .Z(n32578) );
  NOR U45440 ( .A(n32579), .B(n32578), .Z(n35926) );
  IV U45441 ( .A(n32580), .Z(n32582) );
  NOR U45442 ( .A(n32582), .B(n32581), .Z(n36450) );
  NOR U45443 ( .A(n35926), .B(n36450), .Z(n32583) );
  IV U45444 ( .A(n32583), .Z(n32584) );
  NOR U45445 ( .A(n36451), .B(n32584), .Z(n33078) );
  IV U45446 ( .A(n32585), .Z(n32589) );
  IV U45447 ( .A(n32586), .Z(n32595) );
  NOR U45448 ( .A(n32595), .B(n32587), .Z(n32588) );
  IV U45449 ( .A(n32588), .Z(n32591) );
  NOR U45450 ( .A(n32589), .B(n32591), .Z(n35927) );
  IV U45451 ( .A(n32590), .Z(n32592) );
  NOR U45452 ( .A(n32592), .B(n32591), .Z(n35930) );
  IV U45453 ( .A(n32593), .Z(n32597) );
  NOR U45454 ( .A(n32595), .B(n32594), .Z(n32596) );
  IV U45455 ( .A(n32596), .Z(n32599) );
  NOR U45456 ( .A(n32597), .B(n32599), .Z(n35933) );
  IV U45457 ( .A(n32598), .Z(n32600) );
  NOR U45458 ( .A(n32600), .B(n32599), .Z(n36441) );
  IV U45459 ( .A(n32601), .Z(n32604) );
  NOR U45460 ( .A(n32602), .B(n32606), .Z(n32603) );
  IV U45461 ( .A(n32603), .Z(n33075) );
  NOR U45462 ( .A(n32604), .B(n33075), .Z(n36438) );
  IV U45463 ( .A(n32605), .Z(n32607) );
  NOR U45464 ( .A(n32607), .B(n32606), .Z(n33070) );
  NOR U45465 ( .A(n32608), .B(n33058), .Z(n32609) );
  IV U45466 ( .A(n32609), .Z(n35944) );
  NOR U45467 ( .A(n32610), .B(n35944), .Z(n33061) );
  IV U45468 ( .A(n32611), .Z(n32612) );
  NOR U45469 ( .A(n32613), .B(n32612), .Z(n33038) );
  IV U45470 ( .A(n33038), .Z(n33033) );
  IV U45471 ( .A(n32614), .Z(n32615) );
  NOR U45472 ( .A(n32623), .B(n32615), .Z(n35962) );
  IV U45473 ( .A(n32616), .Z(n32618) );
  IV U45474 ( .A(n32617), .Z(n35953) );
  NOR U45475 ( .A(n32618), .B(n35953), .Z(n36409) );
  NOR U45476 ( .A(n35962), .B(n36409), .Z(n33032) );
  IV U45477 ( .A(n32619), .Z(n32620) );
  NOR U45478 ( .A(n32621), .B(n32620), .Z(n35967) );
  IV U45479 ( .A(n32622), .Z(n32624) );
  NOR U45480 ( .A(n32624), .B(n32623), .Z(n35964) );
  NOR U45481 ( .A(n35967), .B(n35964), .Z(n33031) );
  NOR U45482 ( .A(n32626), .B(n32625), .Z(n35972) );
  IV U45483 ( .A(n32627), .Z(n32628) );
  NOR U45484 ( .A(n33025), .B(n32628), .Z(n36397) );
  IV U45485 ( .A(n32629), .Z(n32631) );
  NOR U45486 ( .A(n32631), .B(n32630), .Z(n35975) );
  IV U45487 ( .A(n32632), .Z(n32633) );
  NOR U45488 ( .A(n32634), .B(n32633), .Z(n36384) );
  IV U45489 ( .A(n32635), .Z(n32637) );
  NOR U45490 ( .A(n32637), .B(n32636), .Z(n36388) );
  NOR U45491 ( .A(n36384), .B(n36388), .Z(n36380) );
  NOR U45492 ( .A(n32641), .B(n32638), .Z(n35982) );
  IV U45493 ( .A(n32639), .Z(n32640) );
  NOR U45494 ( .A(n32641), .B(n32640), .Z(n36372) );
  IV U45495 ( .A(n32642), .Z(n32645) );
  NOR U45496 ( .A(n32643), .B(n33020), .Z(n32644) );
  IV U45497 ( .A(n32644), .Z(n33013) );
  NOR U45498 ( .A(n32645), .B(n33013), .Z(n35988) );
  IV U45499 ( .A(n32646), .Z(n32650) );
  IV U45500 ( .A(n32647), .Z(n32648) );
  NOR U45501 ( .A(n32648), .B(n32655), .Z(n32649) );
  IV U45502 ( .A(n32649), .Z(n33004) );
  NOR U45503 ( .A(n32650), .B(n33004), .Z(n35996) );
  IV U45504 ( .A(n32651), .Z(n32652) );
  NOR U45505 ( .A(n32653), .B(n32652), .Z(n36360) );
  IV U45506 ( .A(n32654), .Z(n32656) );
  NOR U45507 ( .A(n32656), .B(n32655), .Z(n36002) );
  NOR U45508 ( .A(n36360), .B(n36002), .Z(n32657) );
  IV U45509 ( .A(n32657), .Z(n33002) );
  IV U45510 ( .A(n32658), .Z(n32659) );
  NOR U45511 ( .A(n32660), .B(n32659), .Z(n36353) );
  IV U45512 ( .A(n32661), .Z(n32662) );
  NOR U45513 ( .A(n32662), .B(n36010), .Z(n33001) );
  IV U45514 ( .A(n32663), .Z(n32666) );
  NOR U45515 ( .A(n32664), .B(n32998), .Z(n32665) );
  IV U45516 ( .A(n32665), .Z(n32668) );
  NOR U45517 ( .A(n32666), .B(n32668), .Z(n36348) );
  IV U45518 ( .A(n32667), .Z(n32669) );
  NOR U45519 ( .A(n32669), .B(n32668), .Z(n36345) );
  IV U45520 ( .A(n32670), .Z(n32671) );
  NOR U45521 ( .A(n32672), .B(n32671), .Z(n32673) );
  IV U45522 ( .A(n32673), .Z(n36023) );
  NOR U45523 ( .A(n36031), .B(n36029), .Z(n32674) );
  IV U45524 ( .A(n32674), .Z(n32993) );
  IV U45525 ( .A(n32675), .Z(n32676) );
  NOR U45526 ( .A(n32676), .B(n36035), .Z(n36335) );
  IV U45527 ( .A(n32677), .Z(n32680) );
  IV U45528 ( .A(n32678), .Z(n32679) );
  NOR U45529 ( .A(n32680), .B(n32679), .Z(n36341) );
  NOR U45530 ( .A(n36335), .B(n36341), .Z(n32992) );
  NOR U45531 ( .A(n32681), .B(n36035), .Z(n32682) );
  NOR U45532 ( .A(n36044), .B(n32682), .Z(n32991) );
  IV U45533 ( .A(n32683), .Z(n32686) );
  IV U45534 ( .A(n32684), .Z(n32685) );
  NOR U45535 ( .A(n32686), .B(n32685), .Z(n36041) );
  IV U45536 ( .A(n32687), .Z(n32691) );
  IV U45537 ( .A(n32688), .Z(n32695) );
  NOR U45538 ( .A(n32695), .B(n32689), .Z(n32690) );
  IV U45539 ( .A(n32690), .Z(n32987) );
  NOR U45540 ( .A(n32691), .B(n32987), .Z(n32692) );
  IV U45541 ( .A(n32692), .Z(n36051) );
  IV U45542 ( .A(n32693), .Z(n32697) );
  NOR U45543 ( .A(n32695), .B(n32694), .Z(n32696) );
  IV U45544 ( .A(n32696), .Z(n32979) );
  NOR U45545 ( .A(n32697), .B(n32979), .Z(n36055) );
  IV U45546 ( .A(n32698), .Z(n32699) );
  NOR U45547 ( .A(n32977), .B(n32699), .Z(n36316) );
  IV U45548 ( .A(n32700), .Z(n32701) );
  NOR U45549 ( .A(n32977), .B(n32701), .Z(n36313) );
  IV U45550 ( .A(n32702), .Z(n32706) );
  IV U45551 ( .A(n32703), .Z(n32704) );
  NOR U45552 ( .A(n32706), .B(n32704), .Z(n36059) );
  IV U45553 ( .A(n32705), .Z(n32707) );
  NOR U45554 ( .A(n32707), .B(n32706), .Z(n42603) );
  NOR U45555 ( .A(n36059), .B(n42603), .Z(n32974) );
  IV U45556 ( .A(n32708), .Z(n32709) );
  NOR U45557 ( .A(n32712), .B(n32709), .Z(n36069) );
  IV U45558 ( .A(n32710), .Z(n32711) );
  NOR U45559 ( .A(n32712), .B(n32711), .Z(n36298) );
  IV U45560 ( .A(n32713), .Z(n32717) );
  IV U45561 ( .A(n32714), .Z(n36077) );
  NOR U45562 ( .A(n32715), .B(n36077), .Z(n32716) );
  IV U45563 ( .A(n32716), .Z(n32719) );
  NOR U45564 ( .A(n32717), .B(n32719), .Z(n36292) );
  IV U45565 ( .A(n32718), .Z(n32720) );
  NOR U45566 ( .A(n32720), .B(n32719), .Z(n36289) );
  IV U45567 ( .A(n32721), .Z(n32722) );
  NOR U45568 ( .A(n32722), .B(n32725), .Z(n32723) );
  IV U45569 ( .A(n32723), .Z(n36087) );
  IV U45570 ( .A(n32726), .Z(n32724) );
  NOR U45571 ( .A(n32725), .B(n32724), .Z(n39198) );
  XOR U45572 ( .A(n32726), .B(n32725), .Z(n32729) );
  IV U45573 ( .A(n32727), .Z(n32728) );
  NOR U45574 ( .A(n32729), .B(n32728), .Z(n39191) );
  NOR U45575 ( .A(n39198), .B(n39191), .Z(n36261) );
  IV U45576 ( .A(n36261), .Z(n32959) );
  NOR U45577 ( .A(n32731), .B(n32730), .Z(n36095) );
  NOR U45578 ( .A(n36253), .B(n36095), .Z(n32951) );
  IV U45579 ( .A(n32732), .Z(n32736) );
  NOR U45580 ( .A(n32734), .B(n32733), .Z(n32735) );
  IV U45581 ( .A(n32735), .Z(n32738) );
  NOR U45582 ( .A(n32736), .B(n32738), .Z(n36092) );
  IV U45583 ( .A(n32737), .Z(n32739) );
  NOR U45584 ( .A(n32739), .B(n32738), .Z(n36097) );
  IV U45585 ( .A(n32740), .Z(n32743) );
  NOR U45586 ( .A(n32741), .B(n32749), .Z(n32742) );
  IV U45587 ( .A(n32742), .Z(n32745) );
  NOR U45588 ( .A(n32743), .B(n32745), .Z(n36241) );
  IV U45589 ( .A(n32744), .Z(n32746) );
  NOR U45590 ( .A(n32746), .B(n32745), .Z(n36100) );
  IV U45591 ( .A(n32747), .Z(n32748) );
  NOR U45592 ( .A(n32749), .B(n32748), .Z(n36103) );
  IV U45593 ( .A(n32750), .Z(n32751) );
  NOR U45594 ( .A(n32754), .B(n32751), .Z(n36231) );
  IV U45595 ( .A(n32752), .Z(n32756) );
  NOR U45596 ( .A(n32754), .B(n32753), .Z(n32755) );
  IV U45597 ( .A(n32755), .Z(n32758) );
  NOR U45598 ( .A(n32756), .B(n32758), .Z(n36228) );
  IV U45599 ( .A(n32757), .Z(n32759) );
  NOR U45600 ( .A(n32759), .B(n32758), .Z(n36106) );
  IV U45601 ( .A(n32760), .Z(n32765) );
  IV U45602 ( .A(n32761), .Z(n32762) );
  NOR U45603 ( .A(n32763), .B(n32762), .Z(n32764) );
  IV U45604 ( .A(n32764), .Z(n32949) );
  NOR U45605 ( .A(n32765), .B(n32949), .Z(n36220) );
  IV U45606 ( .A(n32766), .Z(n32769) );
  NOR U45607 ( .A(n32921), .B(n32767), .Z(n32768) );
  IV U45608 ( .A(n32768), .Z(n32937) );
  NOR U45609 ( .A(n32769), .B(n32937), .Z(n36116) );
  IV U45610 ( .A(n32770), .Z(n32772) );
  NOR U45611 ( .A(n32772), .B(n32771), .Z(n32918) );
  IV U45612 ( .A(n32918), .Z(n32913) );
  IV U45613 ( .A(n32773), .Z(n32775) );
  NOR U45614 ( .A(n32775), .B(n32774), .Z(n36129) );
  IV U45615 ( .A(n32776), .Z(n32778) );
  NOR U45616 ( .A(n32778), .B(n32777), .Z(n32779) );
  IV U45617 ( .A(n32779), .Z(n32900) );
  IV U45618 ( .A(n32780), .Z(n32784) );
  IV U45619 ( .A(n32781), .Z(n32890) );
  NOR U45620 ( .A(n32782), .B(n32890), .Z(n32783) );
  IV U45621 ( .A(n32783), .Z(n32786) );
  NOR U45622 ( .A(n32784), .B(n32786), .Z(n36190) );
  IV U45623 ( .A(n32785), .Z(n32787) );
  NOR U45624 ( .A(n32787), .B(n32786), .Z(n36187) );
  IV U45625 ( .A(n32788), .Z(n32789) );
  NOR U45626 ( .A(n32789), .B(n32867), .Z(n36145) );
  IV U45627 ( .A(n32790), .Z(n32792) );
  XOR U45628 ( .A(n32866), .B(n32867), .Z(n32791) );
  NOR U45629 ( .A(n32792), .B(n32791), .Z(n36142) );
  IV U45630 ( .A(n32793), .Z(n32794) );
  NOR U45631 ( .A(n32795), .B(n32794), .Z(n36165) );
  IV U45632 ( .A(n32796), .Z(n32797) );
  NOR U45633 ( .A(n32798), .B(n32797), .Z(n36171) );
  NOR U45634 ( .A(n36165), .B(n36171), .Z(n32837) );
  IV U45635 ( .A(n32799), .Z(n32802) );
  IV U45636 ( .A(n32800), .Z(n32801) );
  NOR U45637 ( .A(n32802), .B(n32801), .Z(n32826) );
  IV U45638 ( .A(n32803), .Z(n32804) );
  NOR U45639 ( .A(n32804), .B(n32808), .Z(n32805) );
  IV U45640 ( .A(n32805), .Z(n36162) );
  IV U45641 ( .A(n32806), .Z(n32807) );
  NOR U45642 ( .A(n32808), .B(n32807), .Z(n32809) );
  NOR U45643 ( .A(n32810), .B(n32809), .Z(n36160) );
  NOR U45644 ( .A(n32812), .B(n32811), .Z(n32818) );
  IV U45645 ( .A(n32818), .Z(n36159) );
  XOR U45646 ( .A(n36160), .B(n36159), .Z(n32820) );
  IV U45647 ( .A(n32813), .Z(n32815) );
  NOR U45648 ( .A(n32815), .B(n32814), .Z(n32816) );
  IV U45649 ( .A(n32816), .Z(n32817) );
  NOR U45650 ( .A(n32818), .B(n32817), .Z(n32819) );
  NOR U45651 ( .A(n32820), .B(n32819), .Z(n36161) );
  XOR U45652 ( .A(n36162), .B(n36161), .Z(n32827) );
  NOR U45653 ( .A(n32826), .B(n32827), .Z(n32821) );
  IV U45654 ( .A(n32821), .Z(n32825) );
  IV U45655 ( .A(n32822), .Z(n32823) );
  NOR U45656 ( .A(n32824), .B(n32823), .Z(n32830) );
  NOR U45657 ( .A(n32825), .B(n32830), .Z(n32836) );
  IV U45658 ( .A(n32826), .Z(n32831) );
  XOR U45659 ( .A(n32830), .B(n32831), .Z(n32829) );
  IV U45660 ( .A(n32827), .Z(n32828) );
  NOR U45661 ( .A(n32829), .B(n32828), .Z(n32834) );
  IV U45662 ( .A(n32830), .Z(n32832) );
  NOR U45663 ( .A(n32832), .B(n32831), .Z(n32833) );
  NOR U45664 ( .A(n32834), .B(n32833), .Z(n39247) );
  IV U45665 ( .A(n39247), .Z(n32835) );
  NOR U45666 ( .A(n32836), .B(n32835), .Z(n36166) );
  XOR U45667 ( .A(n32837), .B(n36166), .Z(n36175) );
  IV U45668 ( .A(n36175), .Z(n32845) );
  IV U45669 ( .A(n32838), .Z(n32839) );
  NOR U45670 ( .A(n32840), .B(n32839), .Z(n36174) );
  IV U45671 ( .A(n32841), .Z(n32843) );
  NOR U45672 ( .A(n32843), .B(n32842), .Z(n36155) );
  NOR U45673 ( .A(n36174), .B(n36155), .Z(n32844) );
  XOR U45674 ( .A(n32845), .B(n32844), .Z(n36153) );
  IV U45675 ( .A(n32851), .Z(n32846) );
  NOR U45676 ( .A(n32846), .B(n32849), .Z(n32854) );
  IV U45677 ( .A(n32860), .Z(n32847) );
  NOR U45678 ( .A(n32848), .B(n32847), .Z(n32852) );
  IV U45679 ( .A(n32849), .Z(n32850) );
  NOR U45680 ( .A(n32851), .B(n32850), .Z(n36152) );
  NOR U45681 ( .A(n32852), .B(n36152), .Z(n32853) );
  NOR U45682 ( .A(n32854), .B(n32853), .Z(n32855) );
  XOR U45683 ( .A(n36153), .B(n32855), .Z(n32862) );
  IV U45684 ( .A(n32856), .Z(n32858) );
  NOR U45685 ( .A(n32858), .B(n32857), .Z(n32859) );
  IV U45686 ( .A(n32859), .Z(n36151) );
  NOR U45687 ( .A(n32860), .B(n36151), .Z(n32861) );
  XOR U45688 ( .A(n32862), .B(n32861), .Z(n36150) );
  IV U45689 ( .A(n36150), .Z(n32871) );
  IV U45690 ( .A(n32863), .Z(n32865) );
  NOR U45691 ( .A(n32865), .B(n32864), .Z(n32870) );
  IV U45692 ( .A(n32866), .Z(n32868) );
  NOR U45693 ( .A(n32868), .B(n32867), .Z(n32869) );
  NOR U45694 ( .A(n32870), .B(n32869), .Z(n36149) );
  XOR U45695 ( .A(n32871), .B(n36149), .Z(n36143) );
  XOR U45696 ( .A(n36142), .B(n36143), .Z(n36146) );
  XOR U45697 ( .A(n36145), .B(n36146), .Z(n36182) );
  IV U45698 ( .A(n32872), .Z(n32874) );
  NOR U45699 ( .A(n32874), .B(n32873), .Z(n36140) );
  IV U45700 ( .A(n32875), .Z(n32877) );
  NOR U45701 ( .A(n32877), .B(n32876), .Z(n36181) );
  NOR U45702 ( .A(n36140), .B(n36181), .Z(n32878) );
  XOR U45703 ( .A(n36182), .B(n32878), .Z(n36137) );
  IV U45704 ( .A(n32879), .Z(n32880) );
  NOR U45705 ( .A(n32881), .B(n32880), .Z(n36138) );
  IV U45706 ( .A(n32882), .Z(n32884) );
  NOR U45707 ( .A(n32884), .B(n32883), .Z(n36184) );
  NOR U45708 ( .A(n36138), .B(n36184), .Z(n32885) );
  XOR U45709 ( .A(n36137), .B(n32885), .Z(n36135) );
  NOR U45710 ( .A(n32887), .B(n32886), .Z(n36134) );
  IV U45711 ( .A(n32888), .Z(n32889) );
  NOR U45712 ( .A(n32890), .B(n32889), .Z(n36132) );
  NOR U45713 ( .A(n36134), .B(n36132), .Z(n32891) );
  XOR U45714 ( .A(n36135), .B(n32891), .Z(n32892) );
  IV U45715 ( .A(n32892), .Z(n36188) );
  XOR U45716 ( .A(n36187), .B(n36188), .Z(n36191) );
  XOR U45717 ( .A(n36190), .B(n36191), .Z(n36194) );
  NOR U45718 ( .A(n32900), .B(n36194), .Z(n42724) );
  IV U45719 ( .A(n32893), .Z(n32894) );
  NOR U45720 ( .A(n32895), .B(n32894), .Z(n36196) );
  IV U45721 ( .A(n32896), .Z(n32897) );
  NOR U45722 ( .A(n32898), .B(n32897), .Z(n32899) );
  IV U45723 ( .A(n32899), .Z(n36195) );
  XOR U45724 ( .A(n36195), .B(n36194), .Z(n36197) );
  XOR U45725 ( .A(n36196), .B(n36197), .Z(n32902) );
  NOR U45726 ( .A(n36197), .B(n32900), .Z(n32901) );
  NOR U45727 ( .A(n32902), .B(n32901), .Z(n32903) );
  NOR U45728 ( .A(n42724), .B(n32903), .Z(n36201) );
  IV U45729 ( .A(n32904), .Z(n32905) );
  NOR U45730 ( .A(n32910), .B(n32905), .Z(n36200) );
  IV U45731 ( .A(n32906), .Z(n32907) );
  NOR U45732 ( .A(n32907), .B(n32910), .Z(n36208) );
  NOR U45733 ( .A(n36200), .B(n36208), .Z(n32908) );
  XOR U45734 ( .A(n36201), .B(n32908), .Z(n36207) );
  IV U45735 ( .A(n32909), .Z(n32911) );
  NOR U45736 ( .A(n32911), .B(n32910), .Z(n36205) );
  XOR U45737 ( .A(n36207), .B(n36205), .Z(n36130) );
  XOR U45738 ( .A(n36129), .B(n36130), .Z(n32912) );
  NOR U45739 ( .A(n32913), .B(n32912), .Z(n39224) );
  IV U45740 ( .A(n32914), .Z(n32915) );
  NOR U45741 ( .A(n32916), .B(n32915), .Z(n36126) );
  NOR U45742 ( .A(n36126), .B(n36129), .Z(n32917) );
  XOR U45743 ( .A(n32917), .B(n36130), .Z(n32927) );
  NOR U45744 ( .A(n32918), .B(n32927), .Z(n32919) );
  NOR U45745 ( .A(n39224), .B(n32919), .Z(n32934) );
  IV U45746 ( .A(n32934), .Z(n32926) );
  IV U45747 ( .A(n32920), .Z(n32924) );
  NOR U45748 ( .A(n32922), .B(n32921), .Z(n32923) );
  IV U45749 ( .A(n32923), .Z(n32929) );
  NOR U45750 ( .A(n32924), .B(n32929), .Z(n32925) );
  IV U45751 ( .A(n32925), .Z(n42672) );
  NOR U45752 ( .A(n32926), .B(n42672), .Z(n39216) );
  IV U45753 ( .A(n32927), .Z(n32932) );
  IV U45754 ( .A(n32928), .Z(n32930) );
  NOR U45755 ( .A(n32930), .B(n32929), .Z(n32933) );
  IV U45756 ( .A(n32933), .Z(n32931) );
  NOR U45757 ( .A(n32932), .B(n32931), .Z(n39227) );
  NOR U45758 ( .A(n32934), .B(n32933), .Z(n32935) );
  NOR U45759 ( .A(n39227), .B(n32935), .Z(n36123) );
  IV U45760 ( .A(n32936), .Z(n32938) );
  NOR U45761 ( .A(n32938), .B(n32937), .Z(n36124) );
  XOR U45762 ( .A(n36123), .B(n36124), .Z(n32940) );
  NOR U45763 ( .A(n36124), .B(n42672), .Z(n32939) );
  NOR U45764 ( .A(n32940), .B(n32939), .Z(n32941) );
  NOR U45765 ( .A(n39216), .B(n32941), .Z(n36117) );
  XOR U45766 ( .A(n36116), .B(n36117), .Z(n36112) );
  IV U45767 ( .A(n32942), .Z(n32943) );
  NOR U45768 ( .A(n32946), .B(n32943), .Z(n36120) );
  IV U45769 ( .A(n32944), .Z(n32945) );
  NOR U45770 ( .A(n32946), .B(n32945), .Z(n36113) );
  NOR U45771 ( .A(n36120), .B(n36113), .Z(n32947) );
  XOR U45772 ( .A(n36112), .B(n32947), .Z(n36111) );
  IV U45773 ( .A(n32948), .Z(n32950) );
  NOR U45774 ( .A(n32950), .B(n32949), .Z(n36109) );
  XOR U45775 ( .A(n36111), .B(n36109), .Z(n36222) );
  XOR U45776 ( .A(n36220), .B(n36222), .Z(n36108) );
  XOR U45777 ( .A(n36106), .B(n36108), .Z(n36229) );
  XOR U45778 ( .A(n36228), .B(n36229), .Z(n36233) );
  XOR U45779 ( .A(n36231), .B(n36233), .Z(n36104) );
  XOR U45780 ( .A(n36103), .B(n36104), .Z(n36101) );
  XOR U45781 ( .A(n36100), .B(n36101), .Z(n36242) );
  XOR U45782 ( .A(n36241), .B(n36242), .Z(n36098) );
  XOR U45783 ( .A(n36097), .B(n36098), .Z(n36094) );
  XOR U45784 ( .A(n36092), .B(n36094), .Z(n36254) );
  XOR U45785 ( .A(n32951), .B(n36254), .Z(n36090) );
  IV U45786 ( .A(n32952), .Z(n32954) );
  NOR U45787 ( .A(n32954), .B(n32953), .Z(n36256) );
  IV U45788 ( .A(n32955), .Z(n32956) );
  NOR U45789 ( .A(n32957), .B(n32956), .Z(n36089) );
  NOR U45790 ( .A(n36256), .B(n36089), .Z(n32958) );
  XOR U45791 ( .A(n36090), .B(n32958), .Z(n39192) );
  XOR U45792 ( .A(n32959), .B(n39192), .Z(n36086) );
  XOR U45793 ( .A(n36087), .B(n36086), .Z(n36265) );
  IV U45794 ( .A(n32960), .Z(n32963) );
  IV U45795 ( .A(n32961), .Z(n32962) );
  NOR U45796 ( .A(n32963), .B(n32962), .Z(n36275) );
  NOR U45797 ( .A(n36264), .B(n36275), .Z(n32964) );
  XOR U45798 ( .A(n36265), .B(n32964), .Z(n36084) );
  XOR U45799 ( .A(n36082), .B(n36084), .Z(n36273) );
  XOR U45800 ( .A(n36272), .B(n36273), .Z(n36284) );
  XOR U45801 ( .A(n36283), .B(n36284), .Z(n36290) );
  XOR U45802 ( .A(n36289), .B(n36290), .Z(n36293) );
  XOR U45803 ( .A(n36292), .B(n36293), .Z(n36299) );
  XOR U45804 ( .A(n36298), .B(n36299), .Z(n36071) );
  XOR U45805 ( .A(n36069), .B(n36071), .Z(n36063) );
  IV U45806 ( .A(n32965), .Z(n32966) );
  NOR U45807 ( .A(n32967), .B(n32966), .Z(n32968) );
  IV U45808 ( .A(n32968), .Z(n32970) );
  NOR U45809 ( .A(n36063), .B(n32970), .Z(n42608) );
  IV U45810 ( .A(n32969), .Z(n36064) );
  XOR U45811 ( .A(n36064), .B(n36063), .Z(n36066) );
  XOR U45812 ( .A(n36065), .B(n36066), .Z(n32972) );
  NOR U45813 ( .A(n36066), .B(n32970), .Z(n32971) );
  NOR U45814 ( .A(n32972), .B(n32971), .Z(n32973) );
  NOR U45815 ( .A(n42608), .B(n32973), .Z(n36058) );
  XOR U45816 ( .A(n32974), .B(n36058), .Z(n36062) );
  IV U45817 ( .A(n32975), .Z(n32976) );
  NOR U45818 ( .A(n32977), .B(n32976), .Z(n36060) );
  XOR U45819 ( .A(n36062), .B(n36060), .Z(n36314) );
  XOR U45820 ( .A(n36313), .B(n36314), .Z(n36317) );
  XOR U45821 ( .A(n36316), .B(n36317), .Z(n36054) );
  IV U45822 ( .A(n32978), .Z(n32980) );
  NOR U45823 ( .A(n32980), .B(n32979), .Z(n36052) );
  XOR U45824 ( .A(n36054), .B(n36052), .Z(n36056) );
  XOR U45825 ( .A(n36055), .B(n36056), .Z(n36050) );
  XOR U45826 ( .A(n36051), .B(n36050), .Z(n36048) );
  IV U45827 ( .A(n32981), .Z(n32982) );
  NOR U45828 ( .A(n32982), .B(n32984), .Z(n36047) );
  IV U45829 ( .A(n32983), .Z(n32985) );
  NOR U45830 ( .A(n32985), .B(n32984), .Z(n39164) );
  IV U45831 ( .A(n32986), .Z(n32988) );
  NOR U45832 ( .A(n32988), .B(n32987), .Z(n39170) );
  NOR U45833 ( .A(n39164), .B(n39170), .Z(n36325) );
  IV U45834 ( .A(n36325), .Z(n32989) );
  NOR U45835 ( .A(n36047), .B(n32989), .Z(n32990) );
  XOR U45836 ( .A(n36048), .B(n32990), .Z(n36042) );
  XOR U45837 ( .A(n36041), .B(n36042), .Z(n36045) );
  XOR U45838 ( .A(n32991), .B(n36045), .Z(n36334) );
  XOR U45839 ( .A(n32992), .B(n36334), .Z(n36032) );
  XOR U45840 ( .A(n32993), .B(n36032), .Z(n36024) );
  XOR U45841 ( .A(n36023), .B(n36024), .Z(n36020) );
  IV U45842 ( .A(n32994), .Z(n32996) );
  NOR U45843 ( .A(n32996), .B(n32995), .Z(n36025) );
  IV U45844 ( .A(n32997), .Z(n32999) );
  NOR U45845 ( .A(n32999), .B(n32998), .Z(n36019) );
  NOR U45846 ( .A(n36025), .B(n36019), .Z(n33000) );
  XOR U45847 ( .A(n36020), .B(n33000), .Z(n36346) );
  XOR U45848 ( .A(n36345), .B(n36346), .Z(n36349) );
  XOR U45849 ( .A(n36348), .B(n36349), .Z(n36009) );
  XOR U45850 ( .A(n33001), .B(n36009), .Z(n36361) );
  XOR U45851 ( .A(n36353), .B(n36361), .Z(n36003) );
  XOR U45852 ( .A(n33002), .B(n36003), .Z(n35998) );
  XOR U45853 ( .A(n35996), .B(n35998), .Z(n36001) );
  IV U45854 ( .A(n33003), .Z(n33005) );
  NOR U45855 ( .A(n33005), .B(n33004), .Z(n35999) );
  XOR U45856 ( .A(n36001), .B(n35999), .Z(n35992) );
  IV U45857 ( .A(n33006), .Z(n33010) );
  NOR U45858 ( .A(n33008), .B(n33007), .Z(n33009) );
  IV U45859 ( .A(n33009), .Z(n33016) );
  NOR U45860 ( .A(n33010), .B(n33016), .Z(n33011) );
  IV U45861 ( .A(n33011), .Z(n35991) );
  XOR U45862 ( .A(n35992), .B(n35991), .Z(n35986) );
  IV U45863 ( .A(n33012), .Z(n33014) );
  NOR U45864 ( .A(n33014), .B(n33013), .Z(n35985) );
  IV U45865 ( .A(n33015), .Z(n33017) );
  NOR U45866 ( .A(n33017), .B(n33016), .Z(n35993) );
  NOR U45867 ( .A(n35985), .B(n35993), .Z(n33018) );
  XOR U45868 ( .A(n35986), .B(n33018), .Z(n35989) );
  XOR U45869 ( .A(n35988), .B(n35989), .Z(n36368) );
  NOR U45870 ( .A(n33020), .B(n33019), .Z(n33021) );
  IV U45871 ( .A(n33021), .Z(n36367) );
  NOR U45872 ( .A(n33022), .B(n36367), .Z(n33023) );
  XOR U45873 ( .A(n36368), .B(n33023), .Z(n36374) );
  XOR U45874 ( .A(n36372), .B(n36374), .Z(n35983) );
  XOR U45875 ( .A(n35982), .B(n35983), .Z(n36385) );
  XOR U45876 ( .A(n36380), .B(n36385), .Z(n35980) );
  IV U45877 ( .A(n33024), .Z(n33026) );
  NOR U45878 ( .A(n33026), .B(n33025), .Z(n35979) );
  IV U45879 ( .A(n33027), .Z(n33029) );
  NOR U45880 ( .A(n33029), .B(n33028), .Z(n36400) );
  NOR U45881 ( .A(n35979), .B(n36400), .Z(n33030) );
  XOR U45882 ( .A(n35980), .B(n33030), .Z(n35977) );
  XOR U45883 ( .A(n35975), .B(n35977), .Z(n36399) );
  XOR U45884 ( .A(n36397), .B(n36399), .Z(n35970) );
  XOR U45885 ( .A(n35969), .B(n35970), .Z(n35973) );
  XOR U45886 ( .A(n35972), .B(n35973), .Z(n35965) );
  XOR U45887 ( .A(n33031), .B(n35965), .Z(n35961) );
  XOR U45888 ( .A(n33032), .B(n35961), .Z(n35952) );
  NOR U45889 ( .A(n33033), .B(n35952), .Z(n39095) );
  IV U45890 ( .A(n33034), .Z(n33035) );
  NOR U45891 ( .A(n35953), .B(n33035), .Z(n33036) );
  XOR U45892 ( .A(n35952), .B(n33036), .Z(n36417) );
  IV U45893 ( .A(n36417), .Z(n33037) );
  NOR U45894 ( .A(n33038), .B(n33037), .Z(n33039) );
  NOR U45895 ( .A(n39095), .B(n33039), .Z(n36420) );
  IV U45896 ( .A(n33040), .Z(n33042) );
  NOR U45897 ( .A(n33042), .B(n33041), .Z(n36416) );
  IV U45898 ( .A(n33043), .Z(n33045) );
  NOR U45899 ( .A(n33045), .B(n33044), .Z(n36419) );
  NOR U45900 ( .A(n36416), .B(n36419), .Z(n33046) );
  XOR U45901 ( .A(n36420), .B(n33046), .Z(n36427) );
  IV U45902 ( .A(n33047), .Z(n33049) );
  NOR U45903 ( .A(n33049), .B(n33048), .Z(n36423) );
  IV U45904 ( .A(n33050), .Z(n33052) );
  NOR U45905 ( .A(n33052), .B(n33051), .Z(n36425) );
  NOR U45906 ( .A(n36423), .B(n36425), .Z(n33053) );
  XOR U45907 ( .A(n36427), .B(n33053), .Z(n35950) );
  IV U45908 ( .A(n33054), .Z(n33056) );
  NOR U45909 ( .A(n33056), .B(n33055), .Z(n35949) );
  IV U45910 ( .A(n33057), .Z(n33059) );
  NOR U45911 ( .A(n33059), .B(n33058), .Z(n36428) );
  NOR U45912 ( .A(n35949), .B(n36428), .Z(n33060) );
  XOR U45913 ( .A(n35950), .B(n33060), .Z(n35945) );
  XOR U45914 ( .A(n33061), .B(n35945), .Z(n36433) );
  IV U45915 ( .A(n33062), .Z(n33063) );
  NOR U45916 ( .A(n33064), .B(n33063), .Z(n36431) );
  IV U45917 ( .A(n33065), .Z(n33067) );
  NOR U45918 ( .A(n33067), .B(n33066), .Z(n35942) );
  NOR U45919 ( .A(n36431), .B(n35942), .Z(n33068) );
  XOR U45920 ( .A(n36433), .B(n33068), .Z(n33069) );
  NOR U45921 ( .A(n33070), .B(n33069), .Z(n33073) );
  IV U45922 ( .A(n33070), .Z(n33072) );
  XOR U45923 ( .A(n36431), .B(n36433), .Z(n33071) );
  NOR U45924 ( .A(n33072), .B(n33071), .Z(n39067) );
  NOR U45925 ( .A(n33073), .B(n39067), .Z(n35939) );
  IV U45926 ( .A(n33074), .Z(n33076) );
  NOR U45927 ( .A(n33076), .B(n33075), .Z(n33077) );
  IV U45928 ( .A(n33077), .Z(n35940) );
  XOR U45929 ( .A(n35939), .B(n35940), .Z(n36439) );
  XOR U45930 ( .A(n36438), .B(n36439), .Z(n36443) );
  XOR U45931 ( .A(n36441), .B(n36443), .Z(n35934) );
  XOR U45932 ( .A(n35933), .B(n35934), .Z(n35931) );
  XOR U45933 ( .A(n35930), .B(n35931), .Z(n35929) );
  XOR U45934 ( .A(n35927), .B(n35929), .Z(n36447) );
  XOR U45935 ( .A(n33078), .B(n36447), .Z(n36455) );
  IV U45936 ( .A(n33079), .Z(n33081) );
  NOR U45937 ( .A(n33081), .B(n33080), .Z(n33082) );
  IV U45938 ( .A(n33082), .Z(n36457) );
  XOR U45939 ( .A(n36455), .B(n36457), .Z(n36459) );
  XOR U45940 ( .A(n36458), .B(n36459), .Z(n35923) );
  XOR U45941 ( .A(n35922), .B(n35923), .Z(n36464) );
  XOR U45942 ( .A(n33083), .B(n36464), .Z(n35917) );
  XOR U45943 ( .A(n35915), .B(n35917), .Z(n35918) );
  XOR U45944 ( .A(n35919), .B(n35918), .Z(n35908) );
  IV U45945 ( .A(n33084), .Z(n33085) );
  NOR U45946 ( .A(n33086), .B(n33085), .Z(n35913) );
  IV U45947 ( .A(n33087), .Z(n33088) );
  NOR U45948 ( .A(n35904), .B(n33088), .Z(n35909) );
  NOR U45949 ( .A(n35913), .B(n35909), .Z(n33089) );
  XOR U45950 ( .A(n35908), .B(n33089), .Z(n35907) );
  IV U45951 ( .A(n33090), .Z(n33091) );
  NOR U45952 ( .A(n35904), .B(n33091), .Z(n35905) );
  XOR U45953 ( .A(n35907), .B(n35905), .Z(n36474) );
  XOR U45954 ( .A(n33092), .B(n36474), .Z(n36478) );
  XOR U45955 ( .A(n36476), .B(n36478), .Z(n36480) );
  XOR U45956 ( .A(n36479), .B(n36480), .Z(n35897) );
  XOR U45957 ( .A(n35896), .B(n35897), .Z(n35899) );
  XOR U45958 ( .A(n35900), .B(n35899), .Z(n33104) );
  IV U45959 ( .A(n33095), .Z(n33094) );
  IV U45960 ( .A(n33093), .Z(n33112) );
  NOR U45961 ( .A(n33094), .B(n33112), .Z(n33107) );
  IV U45962 ( .A(n33116), .Z(n33100) );
  XOR U45963 ( .A(n33095), .B(n33112), .Z(n33096) );
  NOR U45964 ( .A(n33097), .B(n33096), .Z(n33098) );
  IV U45965 ( .A(n33098), .Z(n33099) );
  NOR U45966 ( .A(n33100), .B(n33099), .Z(n33103) );
  NOR U45967 ( .A(n33107), .B(n33103), .Z(n33101) );
  IV U45968 ( .A(n33101), .Z(n33102) );
  NOR U45969 ( .A(n33104), .B(n33102), .Z(n33110) );
  IV U45970 ( .A(n33103), .Z(n33106) );
  IV U45971 ( .A(n33104), .Z(n33105) );
  NOR U45972 ( .A(n33106), .B(n33105), .Z(n42945) );
  IV U45973 ( .A(n33107), .Z(n33108) );
  NOR U45974 ( .A(n33108), .B(n35899), .Z(n42457) );
  NOR U45975 ( .A(n42945), .B(n42457), .Z(n39043) );
  IV U45976 ( .A(n39043), .Z(n33109) );
  NOR U45977 ( .A(n33110), .B(n33109), .Z(n36483) );
  IV U45978 ( .A(n33111), .Z(n33113) );
  NOR U45979 ( .A(n33113), .B(n33112), .Z(n33114) );
  IV U45980 ( .A(n33114), .Z(n33115) );
  NOR U45981 ( .A(n33116), .B(n33115), .Z(n33117) );
  IV U45982 ( .A(n33117), .Z(n36484) );
  XOR U45983 ( .A(n36483), .B(n36484), .Z(n36489) );
  XOR U45984 ( .A(n36487), .B(n36489), .Z(n36491) );
  XOR U45985 ( .A(n36490), .B(n36491), .Z(n35895) );
  XOR U45986 ( .A(n35893), .B(n35895), .Z(n36496) );
  XOR U45987 ( .A(n36494), .B(n36496), .Z(n36498) );
  XOR U45988 ( .A(n36497), .B(n36498), .Z(n36502) );
  XOR U45989 ( .A(n36501), .B(n36502), .Z(n36505) );
  XOR U45990 ( .A(n33118), .B(n36505), .Z(n35884) );
  XOR U45991 ( .A(n35882), .B(n35884), .Z(n35887) );
  IV U45992 ( .A(n33119), .Z(n33121) );
  NOR U45993 ( .A(n33121), .B(n33120), .Z(n35885) );
  NOR U45994 ( .A(n35880), .B(n35885), .Z(n33122) );
  XOR U45995 ( .A(n35887), .B(n33122), .Z(n35874) );
  IV U45996 ( .A(n33123), .Z(n33126) );
  IV U45997 ( .A(n33124), .Z(n33125) );
  NOR U45998 ( .A(n33126), .B(n33125), .Z(n35877) );
  NOR U45999 ( .A(n35875), .B(n35877), .Z(n33127) );
  XOR U46000 ( .A(n35874), .B(n33127), .Z(n35869) );
  XOR U46001 ( .A(n33128), .B(n35869), .Z(n33134) );
  NOR U46002 ( .A(n33137), .B(n33134), .Z(n39554) );
  IV U46003 ( .A(n33129), .Z(n33131) );
  NOR U46004 ( .A(n33131), .B(n33130), .Z(n33135) );
  IV U46005 ( .A(n33135), .Z(n33132) );
  NOR U46006 ( .A(n33132), .B(n35869), .Z(n39547) );
  NOR U46007 ( .A(n39554), .B(n39547), .Z(n33133) );
  IV U46008 ( .A(n33133), .Z(n36508) );
  IV U46009 ( .A(n33134), .Z(n33138) );
  NOR U46010 ( .A(n33135), .B(n33138), .Z(n33136) );
  NOR U46011 ( .A(n36508), .B(n33136), .Z(n33140) );
  NOR U46012 ( .A(n33138), .B(n33137), .Z(n33139) );
  NOR U46013 ( .A(n33140), .B(n33139), .Z(n39551) );
  IV U46014 ( .A(n33141), .Z(n33142) );
  NOR U46015 ( .A(n33142), .B(n33144), .Z(n35866) );
  IV U46016 ( .A(n33143), .Z(n33145) );
  NOR U46017 ( .A(n33145), .B(n33144), .Z(n39562) );
  NOR U46018 ( .A(n39549), .B(n39562), .Z(n35868) );
  IV U46019 ( .A(n35868), .Z(n33148) );
  NOR U46020 ( .A(n35866), .B(n33148), .Z(n33146) );
  XOR U46021 ( .A(n39551), .B(n33146), .Z(n33151) );
  NOR U46022 ( .A(n33147), .B(n33151), .Z(n35865) );
  IV U46023 ( .A(n33147), .Z(n33150) );
  XOR U46024 ( .A(n33148), .B(n39551), .Z(n33149) );
  NOR U46025 ( .A(n33150), .B(n33149), .Z(n42424) );
  NOR U46026 ( .A(n35865), .B(n42424), .Z(n42987) );
  NOR U46027 ( .A(n42987), .B(n35863), .Z(n33155) );
  IV U46028 ( .A(n35863), .Z(n33153) );
  IV U46029 ( .A(n33151), .Z(n33152) );
  NOR U46030 ( .A(n33153), .B(n33152), .Z(n33154) );
  NOR U46031 ( .A(n33155), .B(n33154), .Z(n35856) );
  XOR U46032 ( .A(n35857), .B(n35856), .Z(n35860) );
  IV U46033 ( .A(n33156), .Z(n33160) );
  NOR U46034 ( .A(n33158), .B(n33157), .Z(n33159) );
  IV U46035 ( .A(n33159), .Z(n33162) );
  NOR U46036 ( .A(n33160), .B(n33162), .Z(n35861) );
  IV U46037 ( .A(n33161), .Z(n33163) );
  NOR U46038 ( .A(n33163), .B(n33162), .Z(n36511) );
  NOR U46039 ( .A(n35861), .B(n36511), .Z(n33164) );
  XOR U46040 ( .A(n35860), .B(n33164), .Z(n36515) );
  NOR U46041 ( .A(n33165), .B(n36515), .Z(n33168) );
  XOR U46042 ( .A(n35860), .B(n35861), .Z(n33166) );
  IV U46043 ( .A(n33165), .Z(n36514) );
  NOR U46044 ( .A(n33166), .B(n36514), .Z(n33167) );
  NOR U46045 ( .A(n33168), .B(n33167), .Z(n35851) );
  IV U46046 ( .A(n33169), .Z(n33171) );
  NOR U46047 ( .A(n33171), .B(n33170), .Z(n35849) );
  XOR U46048 ( .A(n35851), .B(n35849), .Z(n35854) );
  IV U46049 ( .A(n33172), .Z(n33174) );
  NOR U46050 ( .A(n33174), .B(n33173), .Z(n35847) );
  IV U46051 ( .A(n33175), .Z(n33176) );
  NOR U46052 ( .A(n33177), .B(n33176), .Z(n35852) );
  XOR U46053 ( .A(n35847), .B(n35852), .Z(n33178) );
  XOR U46054 ( .A(n35854), .B(n33178), .Z(n35843) );
  XOR U46055 ( .A(n35841), .B(n35843), .Z(n35846) );
  XOR U46056 ( .A(n35844), .B(n35846), .Z(n35830) );
  XOR U46057 ( .A(n33179), .B(n35830), .Z(n35827) );
  XOR U46058 ( .A(n35826), .B(n35827), .Z(n35824) );
  XOR U46059 ( .A(n35822), .B(n35824), .Z(n36521) );
  XOR U46060 ( .A(n36519), .B(n36521), .Z(n36524) );
  XOR U46061 ( .A(n36522), .B(n36524), .Z(n35818) );
  XOR U46062 ( .A(n35816), .B(n35818), .Z(n35821) );
  XOR U46063 ( .A(n35819), .B(n35821), .Z(n39004) );
  XOR U46064 ( .A(n33180), .B(n39004), .Z(n35807) );
  XOR U46065 ( .A(n35808), .B(n35807), .Z(n33181) );
  IV U46066 ( .A(n33181), .Z(n35803) );
  IV U46067 ( .A(n33182), .Z(n33184) );
  NOR U46068 ( .A(n33184), .B(n33183), .Z(n35801) );
  XOR U46069 ( .A(n35803), .B(n35801), .Z(n35805) );
  XOR U46070 ( .A(n35804), .B(n35805), .Z(n38986) );
  XOR U46071 ( .A(n33185), .B(n38986), .Z(n36537) );
  NOR U46072 ( .A(n33192), .B(n36537), .Z(n36545) );
  IV U46073 ( .A(n33186), .Z(n33189) );
  XOR U46074 ( .A(n33187), .B(n33197), .Z(n33188) );
  NOR U46075 ( .A(n33189), .B(n33188), .Z(n35797) );
  NOR U46076 ( .A(n42379), .B(n33190), .Z(n33191) );
  IV U46077 ( .A(n33191), .Z(n36538) );
  XOR U46078 ( .A(n36538), .B(n36537), .Z(n35798) );
  XOR U46079 ( .A(n35797), .B(n35798), .Z(n33194) );
  NOR U46080 ( .A(n35798), .B(n33192), .Z(n33193) );
  NOR U46081 ( .A(n33194), .B(n33193), .Z(n33195) );
  NOR U46082 ( .A(n36545), .B(n33195), .Z(n35792) );
  IV U46083 ( .A(n33196), .Z(n33198) );
  NOR U46084 ( .A(n33198), .B(n33197), .Z(n35794) );
  IV U46085 ( .A(n33199), .Z(n33201) );
  NOR U46086 ( .A(n33201), .B(n33200), .Z(n35791) );
  NOR U46087 ( .A(n35794), .B(n35791), .Z(n33202) );
  XOR U46088 ( .A(n35792), .B(n33202), .Z(n43068) );
  IV U46089 ( .A(n33203), .Z(n33204) );
  NOR U46090 ( .A(n33205), .B(n33204), .Z(n43064) );
  IV U46091 ( .A(n33206), .Z(n33208) );
  NOR U46092 ( .A(n33208), .B(n33207), .Z(n43075) );
  NOR U46093 ( .A(n43064), .B(n43075), .Z(n36547) );
  XOR U46094 ( .A(n43068), .B(n36547), .Z(n35781) );
  XOR U46095 ( .A(n35790), .B(n35781), .Z(n35784) );
  XOR U46096 ( .A(n35783), .B(n35784), .Z(n35788) );
  IV U46097 ( .A(n33209), .Z(n33218) );
  IV U46098 ( .A(n33210), .Z(n33211) );
  NOR U46099 ( .A(n33218), .B(n33211), .Z(n35780) );
  IV U46100 ( .A(n33212), .Z(n33213) );
  NOR U46101 ( .A(n33214), .B(n33213), .Z(n35786) );
  NOR U46102 ( .A(n35780), .B(n35786), .Z(n33215) );
  XOR U46103 ( .A(n35788), .B(n33215), .Z(n36556) );
  IV U46104 ( .A(n33216), .Z(n33217) );
  NOR U46105 ( .A(n33218), .B(n33217), .Z(n39611) );
  NOR U46106 ( .A(n33220), .B(n33219), .Z(n38968) );
  NOR U46107 ( .A(n39611), .B(n38968), .Z(n36557) );
  XOR U46108 ( .A(n36556), .B(n36557), .Z(n35777) );
  XOR U46109 ( .A(n35776), .B(n35777), .Z(n36560) );
  XOR U46110 ( .A(n33221), .B(n36560), .Z(n36582) );
  IV U46111 ( .A(n33222), .Z(n33229) );
  NOR U46112 ( .A(n33224), .B(n33223), .Z(n33226) );
  NOR U46113 ( .A(n33226), .B(n33225), .Z(n33227) );
  IV U46114 ( .A(n33227), .Z(n33228) );
  NOR U46115 ( .A(n33229), .B(n33228), .Z(n36581) );
  NOR U46116 ( .A(n36572), .B(n36581), .Z(n33230) );
  XOR U46117 ( .A(n36582), .B(n33230), .Z(n33231) );
  IV U46118 ( .A(n33231), .Z(n36580) );
  XOR U46119 ( .A(n36578), .B(n36580), .Z(n35774) );
  XOR U46120 ( .A(n33232), .B(n35774), .Z(n35769) );
  IV U46121 ( .A(n33233), .Z(n33234) );
  NOR U46122 ( .A(n33239), .B(n33234), .Z(n35768) );
  IV U46123 ( .A(n33235), .Z(n33237) );
  NOR U46124 ( .A(n33237), .B(n33236), .Z(n35762) );
  NOR U46125 ( .A(n35768), .B(n35762), .Z(n33238) );
  XOR U46126 ( .A(n35769), .B(n33238), .Z(n36587) );
  NOR U46127 ( .A(n33240), .B(n33239), .Z(n33241) );
  IV U46128 ( .A(n33241), .Z(n36586) );
  NOR U46129 ( .A(n33242), .B(n36586), .Z(n33243) );
  XOR U46130 ( .A(n36587), .B(n33243), .Z(n36593) );
  IV U46131 ( .A(n33244), .Z(n33246) );
  NOR U46132 ( .A(n33246), .B(n33245), .Z(n36591) );
  XOR U46133 ( .A(n36593), .B(n36591), .Z(n36603) );
  XOR U46134 ( .A(n36602), .B(n36603), .Z(n36606) );
  IV U46135 ( .A(n33247), .Z(n33248) );
  NOR U46136 ( .A(n35756), .B(n33248), .Z(n36605) );
  IV U46137 ( .A(n33249), .Z(n33250) );
  NOR U46138 ( .A(n35756), .B(n33250), .Z(n33251) );
  XOR U46139 ( .A(n36605), .B(n33251), .Z(n33252) );
  XOR U46140 ( .A(n36606), .B(n33252), .Z(n35748) );
  XOR U46141 ( .A(n33253), .B(n35748), .Z(n35743) );
  XOR U46142 ( .A(n35742), .B(n35743), .Z(n36616) );
  XOR U46143 ( .A(n35745), .B(n36616), .Z(n33260) );
  IV U46144 ( .A(n33254), .Z(n33258) );
  NOR U46145 ( .A(n33256), .B(n33255), .Z(n33257) );
  IV U46146 ( .A(n33257), .Z(n33271) );
  NOR U46147 ( .A(n33258), .B(n33271), .Z(n33268) );
  IV U46148 ( .A(n33268), .Z(n33259) );
  NOR U46149 ( .A(n33260), .B(n33259), .Z(n38931) );
  IV U46150 ( .A(n33261), .Z(n35740) );
  IV U46151 ( .A(n33262), .Z(n33264) );
  NOR U46152 ( .A(n33264), .B(n33263), .Z(n36614) );
  NOR U46153 ( .A(n35745), .B(n36614), .Z(n33265) );
  IV U46154 ( .A(n33265), .Z(n33266) );
  XOR U46155 ( .A(n33266), .B(n36616), .Z(n35739) );
  XOR U46156 ( .A(n35740), .B(n35739), .Z(n33267) );
  NOR U46157 ( .A(n33268), .B(n33267), .Z(n33269) );
  NOR U46158 ( .A(n38931), .B(n33269), .Z(n35733) );
  IV U46159 ( .A(n33270), .Z(n33272) );
  NOR U46160 ( .A(n33272), .B(n33271), .Z(n33273) );
  IV U46161 ( .A(n33273), .Z(n35734) );
  XOR U46162 ( .A(n35733), .B(n35734), .Z(n42316) );
  XOR U46163 ( .A(n33274), .B(n42316), .Z(n33276) );
  NOR U46164 ( .A(n33277), .B(n33276), .Z(n33275) );
  IV U46165 ( .A(n33275), .Z(n38914) );
  NOR U46166 ( .A(n33278), .B(n38914), .Z(n39667) );
  IV U46167 ( .A(n33276), .Z(n33280) );
  NOR U46168 ( .A(n33278), .B(n33277), .Z(n33279) );
  NOR U46169 ( .A(n33280), .B(n33279), .Z(n38919) );
  NOR U46170 ( .A(n39667), .B(n38919), .Z(n36623) );
  XOR U46171 ( .A(n36625), .B(n36623), .Z(n35729) );
  XOR U46172 ( .A(n33281), .B(n38922), .Z(n33284) );
  IV U46173 ( .A(n33282), .Z(n33283) );
  NOR U46174 ( .A(n33284), .B(n33283), .Z(n33285) );
  IV U46175 ( .A(n33285), .Z(n35728) );
  XOR U46176 ( .A(n35729), .B(n35728), .Z(n35730) );
  IV U46177 ( .A(n33286), .Z(n33287) );
  NOR U46178 ( .A(n38922), .B(n33287), .Z(n39660) );
  IV U46179 ( .A(n33288), .Z(n33290) );
  NOR U46180 ( .A(n33290), .B(n33289), .Z(n39675) );
  NOR U46181 ( .A(n39660), .B(n39675), .Z(n35731) );
  XOR U46182 ( .A(n35730), .B(n35731), .Z(n35724) );
  XOR U46183 ( .A(n35722), .B(n35724), .Z(n35726) );
  XOR U46184 ( .A(n33291), .B(n35726), .Z(n35715) );
  XOR U46185 ( .A(n35716), .B(n35715), .Z(n35718) );
  IV U46186 ( .A(n33292), .Z(n33293) );
  NOR U46187 ( .A(n33296), .B(n33293), .Z(n35717) );
  IV U46188 ( .A(n33294), .Z(n33295) );
  NOR U46189 ( .A(n33296), .B(n33295), .Z(n36632) );
  NOR U46190 ( .A(n35717), .B(n36632), .Z(n33297) );
  XOR U46191 ( .A(n35718), .B(n33297), .Z(n35713) );
  XOR U46192 ( .A(n35711), .B(n35713), .Z(n38899) );
  XOR U46193 ( .A(n36635), .B(n38899), .Z(n36637) );
  IV U46194 ( .A(n33298), .Z(n33302) );
  NOR U46195 ( .A(n33300), .B(n33299), .Z(n33301) );
  IV U46196 ( .A(n33301), .Z(n33305) );
  NOR U46197 ( .A(n33302), .B(n33305), .Z(n36641) );
  NOR U46198 ( .A(n36636), .B(n36641), .Z(n33303) );
  XOR U46199 ( .A(n36637), .B(n33303), .Z(n35706) );
  IV U46200 ( .A(n33304), .Z(n33306) );
  NOR U46201 ( .A(n33306), .B(n33305), .Z(n35704) );
  XOR U46202 ( .A(n35706), .B(n35704), .Z(n35708) );
  XOR U46203 ( .A(n35707), .B(n35708), .Z(n33307) );
  NOR U46204 ( .A(n48954), .B(n33307), .Z(n45431) );
  NOR U46205 ( .A(n33309), .B(n33308), .Z(n35701) );
  NOR U46206 ( .A(n35707), .B(n35701), .Z(n33310) );
  XOR U46207 ( .A(n33310), .B(n35708), .Z(n48956) );
  NOR U46208 ( .A(n33311), .B(n48956), .Z(n33312) );
  NOR U46209 ( .A(n45431), .B(n33312), .Z(n35696) );
  IV U46210 ( .A(n33313), .Z(n33315) );
  IV U46211 ( .A(n33314), .Z(n35697) );
  NOR U46212 ( .A(n33315), .B(n35697), .Z(n36645) );
  NOR U46213 ( .A(n35700), .B(n33316), .Z(n33317) );
  NOR U46214 ( .A(n36645), .B(n33317), .Z(n33318) );
  XOR U46215 ( .A(n35696), .B(n33318), .Z(n35695) );
  IV U46216 ( .A(n33319), .Z(n33321) );
  NOR U46217 ( .A(n33321), .B(n33320), .Z(n35693) );
  XOR U46218 ( .A(n35695), .B(n35693), .Z(n35692) );
  XOR U46219 ( .A(n35690), .B(n35692), .Z(n36649) );
  XOR U46220 ( .A(n36648), .B(n36649), .Z(n36652) );
  XOR U46221 ( .A(n36651), .B(n36652), .Z(n35688) );
  XOR U46222 ( .A(n35687), .B(n35688), .Z(n36661) );
  XOR U46223 ( .A(n36660), .B(n36661), .Z(n36664) );
  XOR U46224 ( .A(n36663), .B(n36664), .Z(n35685) );
  XOR U46225 ( .A(n35684), .B(n35685), .Z(n35676) );
  XOR U46226 ( .A(n33322), .B(n35676), .Z(n43189) );
  XOR U46227 ( .A(n35673), .B(n43189), .Z(n38867) );
  XOR U46228 ( .A(n33323), .B(n38867), .Z(n35667) );
  XOR U46229 ( .A(n35666), .B(n35667), .Z(n35670) );
  XOR U46230 ( .A(n35669), .B(n35670), .Z(n35665) );
  IV U46231 ( .A(n33324), .Z(n33326) );
  NOR U46232 ( .A(n33326), .B(n33325), .Z(n35663) );
  XOR U46233 ( .A(n35665), .B(n35663), .Z(n35658) );
  XOR U46234 ( .A(n35659), .B(n35658), .Z(n35661) );
  IV U46235 ( .A(n33327), .Z(n33328) );
  NOR U46236 ( .A(n33329), .B(n33328), .Z(n35660) );
  IV U46237 ( .A(n33330), .Z(n33332) );
  NOR U46238 ( .A(n33332), .B(n33331), .Z(n36673) );
  NOR U46239 ( .A(n35660), .B(n36673), .Z(n33333) );
  XOR U46240 ( .A(n35661), .B(n33333), .Z(n35657) );
  IV U46241 ( .A(n33334), .Z(n33336) );
  NOR U46242 ( .A(n33336), .B(n33335), .Z(n35655) );
  IV U46243 ( .A(n33337), .Z(n33338) );
  NOR U46244 ( .A(n33338), .B(n33346), .Z(n35653) );
  NOR U46245 ( .A(n35655), .B(n35653), .Z(n33339) );
  XOR U46246 ( .A(n35657), .B(n33339), .Z(n33340) );
  NOR U46247 ( .A(n33341), .B(n33340), .Z(n33344) );
  IV U46248 ( .A(n33341), .Z(n33343) );
  XOR U46249 ( .A(n35655), .B(n35657), .Z(n33342) );
  NOR U46250 ( .A(n33343), .B(n33342), .Z(n42231) );
  NOR U46251 ( .A(n33344), .B(n42231), .Z(n35647) );
  IV U46252 ( .A(n33345), .Z(n33347) );
  NOR U46253 ( .A(n33347), .B(n33346), .Z(n36676) );
  IV U46254 ( .A(n33348), .Z(n33349) );
  NOR U46255 ( .A(n33350), .B(n33349), .Z(n35646) );
  NOR U46256 ( .A(n36676), .B(n35646), .Z(n33351) );
  XOR U46257 ( .A(n35647), .B(n33351), .Z(n35650) );
  XOR U46258 ( .A(n33352), .B(n35650), .Z(n35640) );
  XOR U46259 ( .A(n35638), .B(n35640), .Z(n35637) );
  IV U46260 ( .A(n33353), .Z(n33356) );
  IV U46261 ( .A(n33354), .Z(n33355) );
  NOR U46262 ( .A(n33356), .B(n33355), .Z(n35635) );
  XOR U46263 ( .A(n35637), .B(n35635), .Z(n35631) );
  IV U46264 ( .A(n33357), .Z(n33358) );
  NOR U46265 ( .A(n33359), .B(n33358), .Z(n35633) );
  IV U46266 ( .A(n33360), .Z(n33361) );
  NOR U46267 ( .A(n33365), .B(n33361), .Z(n35630) );
  NOR U46268 ( .A(n35633), .B(n35630), .Z(n33362) );
  XOR U46269 ( .A(n35631), .B(n33362), .Z(n36681) );
  IV U46270 ( .A(n33363), .Z(n33364) );
  NOR U46271 ( .A(n33365), .B(n33364), .Z(n36684) );
  NOR U46272 ( .A(n33367), .B(n33366), .Z(n36682) );
  NOR U46273 ( .A(n36684), .B(n36682), .Z(n33368) );
  XOR U46274 ( .A(n36681), .B(n33368), .Z(n43227) );
  IV U46275 ( .A(n33369), .Z(n33370) );
  NOR U46276 ( .A(n33371), .B(n33370), .Z(n35627) );
  NOR U46277 ( .A(n43228), .B(n35627), .Z(n33372) );
  XOR U46278 ( .A(n43227), .B(n33372), .Z(n35623) );
  XOR U46279 ( .A(n35625), .B(n35623), .Z(n35622) );
  IV U46280 ( .A(n33373), .Z(n33374) );
  NOR U46281 ( .A(n33375), .B(n33374), .Z(n35618) );
  IV U46282 ( .A(n33376), .Z(n33378) );
  NOR U46283 ( .A(n33378), .B(n33377), .Z(n35620) );
  NOR U46284 ( .A(n35618), .B(n35620), .Z(n33379) );
  XOR U46285 ( .A(n35622), .B(n33379), .Z(n36696) );
  IV U46286 ( .A(n33380), .Z(n33381) );
  NOR U46287 ( .A(n33388), .B(n33381), .Z(n36699) );
  IV U46288 ( .A(n33382), .Z(n33383) );
  NOR U46289 ( .A(n33384), .B(n33383), .Z(n36697) );
  NOR U46290 ( .A(n36699), .B(n36697), .Z(n33385) );
  XOR U46291 ( .A(n36696), .B(n33385), .Z(n35616) );
  IV U46292 ( .A(n33386), .Z(n33391) );
  IV U46293 ( .A(n33387), .Z(n33389) );
  NOR U46294 ( .A(n33389), .B(n33388), .Z(n33390) );
  IV U46295 ( .A(n33390), .Z(n33393) );
  NOR U46296 ( .A(n33391), .B(n33393), .Z(n35614) );
  XOR U46297 ( .A(n35616), .B(n35614), .Z(n36709) );
  IV U46298 ( .A(n33392), .Z(n33394) );
  NOR U46299 ( .A(n33394), .B(n33393), .Z(n36707) );
  XOR U46300 ( .A(n36709), .B(n36707), .Z(n35608) );
  NOR U46301 ( .A(n33396), .B(n33395), .Z(n33397) );
  IV U46302 ( .A(n33397), .Z(n35607) );
  NOR U46303 ( .A(n33398), .B(n35607), .Z(n33399) );
  XOR U46304 ( .A(n35608), .B(n33399), .Z(n36714) );
  IV U46305 ( .A(n33400), .Z(n33401) );
  NOR U46306 ( .A(n33402), .B(n33401), .Z(n36715) );
  NOR U46307 ( .A(n33404), .B(n33403), .Z(n35599) );
  NOR U46308 ( .A(n36715), .B(n35599), .Z(n33405) );
  XOR U46309 ( .A(n36714), .B(n33405), .Z(n35602) );
  XOR U46310 ( .A(n33406), .B(n35602), .Z(n36720) );
  XOR U46311 ( .A(n36718), .B(n36720), .Z(n36722) );
  XOR U46312 ( .A(n36721), .B(n36722), .Z(n36726) );
  XOR U46313 ( .A(n36725), .B(n36726), .Z(n36732) );
  IV U46314 ( .A(n33407), .Z(n33408) );
  NOR U46315 ( .A(n33409), .B(n33408), .Z(n36731) );
  IV U46316 ( .A(n33410), .Z(n33412) );
  NOR U46317 ( .A(n33412), .B(n33411), .Z(n36728) );
  NOR U46318 ( .A(n36731), .B(n36728), .Z(n33413) );
  XOR U46319 ( .A(n36732), .B(n33413), .Z(n36734) );
  IV U46320 ( .A(n33414), .Z(n33416) );
  NOR U46321 ( .A(n33416), .B(n33415), .Z(n36735) );
  IV U46322 ( .A(n33417), .Z(n33418) );
  NOR U46323 ( .A(n33419), .B(n33418), .Z(n36737) );
  NOR U46324 ( .A(n36735), .B(n36737), .Z(n33420) );
  XOR U46325 ( .A(n36734), .B(n33420), .Z(n35597) );
  XOR U46326 ( .A(n35596), .B(n35597), .Z(n36743) );
  NOR U46327 ( .A(n33421), .B(n36740), .Z(n33422) );
  NOR U46328 ( .A(n33423), .B(n33422), .Z(n33424) );
  XOR U46329 ( .A(n36743), .B(n33424), .Z(n36752) );
  XOR U46330 ( .A(n36751), .B(n36752), .Z(n35595) );
  XOR U46331 ( .A(n33425), .B(n35595), .Z(n33426) );
  IV U46332 ( .A(n33426), .Z(n35592) );
  IV U46333 ( .A(n33427), .Z(n33429) );
  NOR U46334 ( .A(n33429), .B(n33428), .Z(n35590) );
  XOR U46335 ( .A(n35592), .B(n35590), .Z(n36758) );
  XOR U46336 ( .A(n36759), .B(n36758), .Z(n36760) );
  IV U46337 ( .A(n33430), .Z(n33431) );
  NOR U46338 ( .A(n33432), .B(n33431), .Z(n36766) );
  IV U46339 ( .A(n33433), .Z(n33436) );
  IV U46340 ( .A(n33434), .Z(n33435) );
  NOR U46341 ( .A(n33436), .B(n33435), .Z(n36761) );
  NOR U46342 ( .A(n36766), .B(n36761), .Z(n33437) );
  XOR U46343 ( .A(n36760), .B(n33437), .Z(n35586) );
  XOR U46344 ( .A(n35585), .B(n35586), .Z(n36781) );
  IV U46345 ( .A(n33438), .Z(n33443) );
  NOR U46346 ( .A(n33440), .B(n33439), .Z(n33441) );
  IV U46347 ( .A(n33441), .Z(n33442) );
  NOR U46348 ( .A(n33443), .B(n33442), .Z(n36779) );
  NOR U46349 ( .A(n35583), .B(n36779), .Z(n33444) );
  XOR U46350 ( .A(n36781), .B(n33444), .Z(n35579) );
  XOR U46351 ( .A(n35580), .B(n35579), .Z(n36785) );
  XOR U46352 ( .A(n33445), .B(n36785), .Z(n38781) );
  IV U46353 ( .A(n33446), .Z(n33449) );
  IV U46354 ( .A(n33447), .Z(n33448) );
  NOR U46355 ( .A(n33449), .B(n33448), .Z(n39798) );
  IV U46356 ( .A(n33450), .Z(n33451) );
  NOR U46357 ( .A(n33451), .B(n33455), .Z(n38779) );
  NOR U46358 ( .A(n39798), .B(n38779), .Z(n36797) );
  XOR U46359 ( .A(n38781), .B(n36797), .Z(n33452) );
  IV U46360 ( .A(n33452), .Z(n35577) );
  XOR U46361 ( .A(n35576), .B(n35577), .Z(n39808) );
  NOR U46362 ( .A(n33453), .B(n39808), .Z(n38773) );
  IV U46363 ( .A(n33454), .Z(n33456) );
  NOR U46364 ( .A(n33456), .B(n33455), .Z(n35575) );
  NOR U46365 ( .A(n35576), .B(n35575), .Z(n33457) );
  XOR U46366 ( .A(n35577), .B(n33457), .Z(n33458) );
  NOR U46367 ( .A(n33459), .B(n33458), .Z(n33460) );
  NOR U46368 ( .A(n38773), .B(n33460), .Z(n33461) );
  XOR U46369 ( .A(n35573), .B(n33461), .Z(n35570) );
  IV U46370 ( .A(n33462), .Z(n33464) );
  NOR U46371 ( .A(n33464), .B(n33463), .Z(n35569) );
  IV U46372 ( .A(n33465), .Z(n33467) );
  NOR U46373 ( .A(n33467), .B(n33466), .Z(n43297) );
  IV U46374 ( .A(n33468), .Z(n33469) );
  NOR U46375 ( .A(n33470), .B(n33469), .Z(n42127) );
  NOR U46376 ( .A(n43297), .B(n42127), .Z(n35572) );
  IV U46377 ( .A(n35572), .Z(n33471) );
  NOR U46378 ( .A(n35569), .B(n33471), .Z(n33472) );
  XOR U46379 ( .A(n35570), .B(n33472), .Z(n35565) );
  IV U46380 ( .A(n33473), .Z(n33475) );
  NOR U46381 ( .A(n33475), .B(n33474), .Z(n35563) );
  XOR U46382 ( .A(n35565), .B(n35563), .Z(n35568) );
  XOR U46383 ( .A(n35566), .B(n35568), .Z(n36806) );
  XOR U46384 ( .A(n36804), .B(n36806), .Z(n36808) );
  XOR U46385 ( .A(n36807), .B(n36808), .Z(n36812) );
  XOR U46386 ( .A(n36811), .B(n36812), .Z(n36816) );
  XOR U46387 ( .A(n33476), .B(n36816), .Z(n36830) );
  XOR U46388 ( .A(n36828), .B(n36830), .Z(n36836) );
  XOR U46389 ( .A(n33477), .B(n36836), .Z(n35555) );
  XOR U46390 ( .A(n33478), .B(n35555), .Z(n42104) );
  XOR U46391 ( .A(n33479), .B(n42104), .Z(n36837) );
  XOR U46392 ( .A(n36838), .B(n36837), .Z(n36839) );
  NOR U46393 ( .A(n33487), .B(n36839), .Z(n36841) );
  IV U46394 ( .A(n33480), .Z(n33482) );
  NOR U46395 ( .A(n33482), .B(n33481), .Z(n35549) );
  IV U46396 ( .A(n33483), .Z(n33484) );
  NOR U46397 ( .A(n33485), .B(n33484), .Z(n33486) );
  IV U46398 ( .A(n33486), .Z(n36840) );
  XOR U46399 ( .A(n36840), .B(n36839), .Z(n35550) );
  XOR U46400 ( .A(n35549), .B(n35550), .Z(n33489) );
  NOR U46401 ( .A(n35550), .B(n33487), .Z(n33488) );
  NOR U46402 ( .A(n33489), .B(n33488), .Z(n33490) );
  NOR U46403 ( .A(n36841), .B(n33490), .Z(n36847) );
  IV U46404 ( .A(n33491), .Z(n33493) );
  NOR U46405 ( .A(n33493), .B(n33492), .Z(n33494) );
  IV U46406 ( .A(n33494), .Z(n36849) );
  XOR U46407 ( .A(n36847), .B(n36849), .Z(n36851) );
  XOR U46408 ( .A(n36850), .B(n36851), .Z(n33495) );
  NOR U46409 ( .A(n42091), .B(n33495), .Z(n38724) );
  IV U46410 ( .A(n33496), .Z(n33497) );
  NOR U46411 ( .A(n33498), .B(n33497), .Z(n36845) );
  NOR U46412 ( .A(n36850), .B(n36845), .Z(n33499) );
  XOR U46413 ( .A(n33499), .B(n36851), .Z(n42085) );
  NOR U46414 ( .A(n33500), .B(n42085), .Z(n33501) );
  NOR U46415 ( .A(n38724), .B(n33501), .Z(n33502) );
  IV U46416 ( .A(n33502), .Z(n36857) );
  XOR U46417 ( .A(n36856), .B(n36857), .Z(n35548) );
  XOR U46418 ( .A(n35546), .B(n35548), .Z(n35541) );
  XOR U46419 ( .A(n35540), .B(n35541), .Z(n35544) );
  XOR U46420 ( .A(n35543), .B(n35544), .Z(n36866) );
  XOR U46421 ( .A(n35538), .B(n36866), .Z(n36873) );
  XOR U46422 ( .A(n33503), .B(n36873), .Z(n36870) );
  XOR U46423 ( .A(n36868), .B(n36870), .Z(n36877) );
  IV U46424 ( .A(n33504), .Z(n33508) );
  NOR U46425 ( .A(n33506), .B(n33505), .Z(n33507) );
  IV U46426 ( .A(n33507), .Z(n33515) );
  NOR U46427 ( .A(n33508), .B(n33515), .Z(n36875) );
  XOR U46428 ( .A(n36877), .B(n36875), .Z(n36880) );
  IV U46429 ( .A(n33509), .Z(n33513) );
  IV U46430 ( .A(n33510), .Z(n33529) );
  NOR U46431 ( .A(n33529), .B(n33511), .Z(n33512) );
  IV U46432 ( .A(n33512), .Z(n33521) );
  NOR U46433 ( .A(n33513), .B(n33521), .Z(n35536) );
  IV U46434 ( .A(n33514), .Z(n33516) );
  NOR U46435 ( .A(n33516), .B(n33515), .Z(n36878) );
  NOR U46436 ( .A(n35536), .B(n36878), .Z(n33517) );
  XOR U46437 ( .A(n36880), .B(n33517), .Z(n35529) );
  IV U46438 ( .A(n33518), .Z(n33519) );
  NOR U46439 ( .A(n33529), .B(n33519), .Z(n35530) );
  IV U46440 ( .A(n33520), .Z(n33522) );
  NOR U46441 ( .A(n33522), .B(n33521), .Z(n35533) );
  NOR U46442 ( .A(n35530), .B(n35533), .Z(n33523) );
  XOR U46443 ( .A(n35529), .B(n33523), .Z(n36886) );
  IV U46444 ( .A(n33524), .Z(n33525) );
  NOR U46445 ( .A(n33526), .B(n33525), .Z(n36885) );
  IV U46446 ( .A(n33527), .Z(n33528) );
  NOR U46447 ( .A(n33529), .B(n33528), .Z(n35527) );
  NOR U46448 ( .A(n36885), .B(n35527), .Z(n33530) );
  XOR U46449 ( .A(n36886), .B(n33530), .Z(n33531) );
  IV U46450 ( .A(n33531), .Z(n36884) );
  IV U46451 ( .A(n33532), .Z(n33534) );
  NOR U46452 ( .A(n33534), .B(n33533), .Z(n36882) );
  XOR U46453 ( .A(n36884), .B(n36882), .Z(n36898) );
  XOR U46454 ( .A(n36896), .B(n36898), .Z(n36890) );
  XOR U46455 ( .A(n36889), .B(n36890), .Z(n36894) );
  XOR U46456 ( .A(n33535), .B(n36894), .Z(n35520) );
  IV U46457 ( .A(n33536), .Z(n33539) );
  IV U46458 ( .A(n33537), .Z(n33538) );
  NOR U46459 ( .A(n33539), .B(n33538), .Z(n35524) );
  IV U46460 ( .A(n33540), .Z(n33542) );
  NOR U46461 ( .A(n33542), .B(n33541), .Z(n35519) );
  NOR U46462 ( .A(n35524), .B(n35519), .Z(n33543) );
  XOR U46463 ( .A(n35520), .B(n33543), .Z(n35518) );
  XOR U46464 ( .A(n35516), .B(n35518), .Z(n35514) );
  XOR U46465 ( .A(n33544), .B(n35514), .Z(n35509) );
  XOR U46466 ( .A(n35507), .B(n35509), .Z(n35505) );
  XOR U46467 ( .A(n35506), .B(n35505), .Z(n36911) );
  IV U46468 ( .A(n33545), .Z(n33547) );
  NOR U46469 ( .A(n33547), .B(n33546), .Z(n35502) );
  IV U46470 ( .A(n33548), .Z(n33549) );
  NOR U46471 ( .A(n33550), .B(n33549), .Z(n36910) );
  NOR U46472 ( .A(n35502), .B(n36910), .Z(n33551) );
  XOR U46473 ( .A(n36911), .B(n33551), .Z(n36909) );
  XOR U46474 ( .A(n36907), .B(n36909), .Z(n35493) );
  XOR U46475 ( .A(n33552), .B(n35493), .Z(n35486) );
  XOR U46476 ( .A(n33553), .B(n35486), .Z(n35484) );
  IV U46477 ( .A(n33554), .Z(n33556) );
  NOR U46478 ( .A(n33556), .B(n33555), .Z(n35483) );
  NOR U46479 ( .A(n35481), .B(n35483), .Z(n33557) );
  XOR U46480 ( .A(n35484), .B(n33557), .Z(n33558) );
  NOR U46481 ( .A(n33559), .B(n33558), .Z(n33562) );
  IV U46482 ( .A(n33559), .Z(n33561) );
  XOR U46483 ( .A(n35481), .B(n35484), .Z(n33560) );
  NOR U46484 ( .A(n33561), .B(n33560), .Z(n42023) );
  NOR U46485 ( .A(n33562), .B(n42023), .Z(n36916) );
  IV U46486 ( .A(n33563), .Z(n33565) );
  NOR U46487 ( .A(n33565), .B(n33564), .Z(n33566) );
  IV U46488 ( .A(n33566), .Z(n36917) );
  XOR U46489 ( .A(n36916), .B(n36917), .Z(n35476) );
  XOR U46490 ( .A(n35475), .B(n35476), .Z(n35479) );
  XOR U46491 ( .A(n35478), .B(n35479), .Z(n35470) );
  XOR U46492 ( .A(n35469), .B(n35470), .Z(n35473) );
  XOR U46493 ( .A(n35472), .B(n35473), .Z(n35468) );
  XOR U46494 ( .A(n35466), .B(n35468), .Z(n35461) );
  XOR U46495 ( .A(n35460), .B(n35461), .Z(n35465) );
  XOR U46496 ( .A(n35463), .B(n35465), .Z(n35458) );
  NOR U46497 ( .A(n33575), .B(n35458), .Z(n39961) );
  XOR U46498 ( .A(n33567), .B(n33580), .Z(n33570) );
  IV U46499 ( .A(n33568), .Z(n33569) );
  NOR U46500 ( .A(n33570), .B(n33569), .Z(n35450) );
  IV U46501 ( .A(n33571), .Z(n33572) );
  NOR U46502 ( .A(n33573), .B(n33572), .Z(n33574) );
  IV U46503 ( .A(n33574), .Z(n35459) );
  XOR U46504 ( .A(n35459), .B(n35458), .Z(n35451) );
  XOR U46505 ( .A(n35450), .B(n35451), .Z(n33577) );
  NOR U46506 ( .A(n35451), .B(n33575), .Z(n33576) );
  NOR U46507 ( .A(n33577), .B(n33576), .Z(n33578) );
  NOR U46508 ( .A(n39961), .B(n33578), .Z(n35448) );
  IV U46509 ( .A(n33579), .Z(n33581) );
  NOR U46510 ( .A(n33581), .B(n33580), .Z(n35454) );
  NOR U46511 ( .A(n33583), .B(n33582), .Z(n35447) );
  NOR U46512 ( .A(n35454), .B(n35447), .Z(n33584) );
  XOR U46513 ( .A(n35448), .B(n33584), .Z(n35443) );
  XOR U46514 ( .A(n35441), .B(n35443), .Z(n35446) );
  XOR U46515 ( .A(n35444), .B(n35446), .Z(n35439) );
  XOR U46516 ( .A(n33585), .B(n35439), .Z(n35435) );
  IV U46517 ( .A(n33586), .Z(n33587) );
  NOR U46518 ( .A(n33588), .B(n33587), .Z(n35434) );
  IV U46519 ( .A(n33589), .Z(n33593) );
  XOR U46520 ( .A(n33591), .B(n33590), .Z(n33592) );
  NOR U46521 ( .A(n33593), .B(n33592), .Z(n36929) );
  NOR U46522 ( .A(n35434), .B(n36929), .Z(n33594) );
  XOR U46523 ( .A(n35435), .B(n33594), .Z(n36937) );
  XOR U46524 ( .A(n33595), .B(n36937), .Z(n36939) );
  IV U46525 ( .A(n33596), .Z(n33598) );
  NOR U46526 ( .A(n33598), .B(n33597), .Z(n33599) );
  NOR U46527 ( .A(n36939), .B(n33599), .Z(n33602) );
  IV U46528 ( .A(n33599), .Z(n36940) );
  XOR U46529 ( .A(n35431), .B(n36937), .Z(n33600) );
  NOR U46530 ( .A(n36940), .B(n33600), .Z(n33601) );
  NOR U46531 ( .A(n33602), .B(n33601), .Z(n35425) );
  XOR U46532 ( .A(n35426), .B(n35425), .Z(n35429) );
  XOR U46533 ( .A(n35428), .B(n35429), .Z(n35420) );
  XOR U46534 ( .A(n35421), .B(n35420), .Z(n35418) );
  IV U46535 ( .A(n33603), .Z(n33606) );
  IV U46536 ( .A(n33604), .Z(n33605) );
  NOR U46537 ( .A(n33606), .B(n33605), .Z(n35417) );
  NOR U46538 ( .A(n35422), .B(n35417), .Z(n33607) );
  XOR U46539 ( .A(n35418), .B(n33607), .Z(n36949) );
  XOR U46540 ( .A(n36947), .B(n36949), .Z(n35416) );
  XOR U46541 ( .A(n35414), .B(n35416), .Z(n36960) );
  XOR U46542 ( .A(n33608), .B(n36960), .Z(n35402) );
  IV U46543 ( .A(n33609), .Z(n33610) );
  NOR U46544 ( .A(n33611), .B(n33610), .Z(n35409) );
  IV U46545 ( .A(n33612), .Z(n33613) );
  NOR U46546 ( .A(n35394), .B(n33613), .Z(n35401) );
  NOR U46547 ( .A(n35409), .B(n35401), .Z(n33614) );
  XOR U46548 ( .A(n35402), .B(n33614), .Z(n35395) );
  XOR U46549 ( .A(n33615), .B(n35395), .Z(n35392) );
  IV U46550 ( .A(n33616), .Z(n33617) );
  NOR U46551 ( .A(n33617), .B(n33625), .Z(n35390) );
  NOR U46552 ( .A(n35388), .B(n35390), .Z(n33618) );
  XOR U46553 ( .A(n35392), .B(n33618), .Z(n33619) );
  NOR U46554 ( .A(n33620), .B(n33619), .Z(n33623) );
  XOR U46555 ( .A(n35388), .B(n35392), .Z(n33622) );
  IV U46556 ( .A(n33620), .Z(n33621) );
  NOR U46557 ( .A(n33622), .B(n33621), .Z(n41955) );
  NOR U46558 ( .A(n33623), .B(n41955), .Z(n35385) );
  IV U46559 ( .A(n33624), .Z(n33629) );
  NOR U46560 ( .A(n33626), .B(n33625), .Z(n33627) );
  IV U46561 ( .A(n33627), .Z(n33628) );
  NOR U46562 ( .A(n33629), .B(n33628), .Z(n33630) );
  IV U46563 ( .A(n33630), .Z(n35386) );
  XOR U46564 ( .A(n35385), .B(n35386), .Z(n35380) );
  XOR U46565 ( .A(n35379), .B(n35380), .Z(n35383) );
  XOR U46566 ( .A(n35382), .B(n35383), .Z(n35377) );
  XOR U46567 ( .A(n33631), .B(n35377), .Z(n36968) );
  XOR U46568 ( .A(n36967), .B(n36968), .Z(n35372) );
  XOR U46569 ( .A(n35371), .B(n35372), .Z(n36976) );
  IV U46570 ( .A(n33632), .Z(n33634) );
  NOR U46571 ( .A(n33634), .B(n33633), .Z(n33635) );
  IV U46572 ( .A(n33635), .Z(n36975) );
  XOR U46573 ( .A(n36976), .B(n36975), .Z(n35368) );
  NOR U46574 ( .A(n33646), .B(n33636), .Z(n36977) );
  IV U46575 ( .A(n33637), .Z(n33638) );
  NOR U46576 ( .A(n33646), .B(n33638), .Z(n35369) );
  NOR U46577 ( .A(n36977), .B(n35369), .Z(n33639) );
  XOR U46578 ( .A(n35368), .B(n33639), .Z(n35367) );
  IV U46579 ( .A(n33640), .Z(n33643) );
  IV U46580 ( .A(n33641), .Z(n33642) );
  NOR U46581 ( .A(n33643), .B(n33642), .Z(n35363) );
  IV U46582 ( .A(n33644), .Z(n33645) );
  NOR U46583 ( .A(n33646), .B(n33645), .Z(n35365) );
  NOR U46584 ( .A(n35363), .B(n35365), .Z(n33647) );
  XOR U46585 ( .A(n35367), .B(n33647), .Z(n35357) );
  IV U46586 ( .A(n33648), .Z(n33649) );
  NOR U46587 ( .A(n33650), .B(n33649), .Z(n35360) );
  IV U46588 ( .A(n33651), .Z(n33652) );
  NOR U46589 ( .A(n33653), .B(n33652), .Z(n35356) );
  NOR U46590 ( .A(n35360), .B(n35356), .Z(n33654) );
  XOR U46591 ( .A(n35357), .B(n33654), .Z(n35355) );
  IV U46592 ( .A(n33655), .Z(n33656) );
  NOR U46593 ( .A(n33657), .B(n33656), .Z(n35353) );
  IV U46594 ( .A(n33658), .Z(n33660) );
  NOR U46595 ( .A(n33660), .B(n33659), .Z(n35351) );
  NOR U46596 ( .A(n35353), .B(n35351), .Z(n33661) );
  XOR U46597 ( .A(n35355), .B(n33661), .Z(n35349) );
  IV U46598 ( .A(n33662), .Z(n33663) );
  NOR U46599 ( .A(n33664), .B(n33663), .Z(n35348) );
  NOR U46600 ( .A(n33666), .B(n33665), .Z(n36980) );
  NOR U46601 ( .A(n35348), .B(n36980), .Z(n33667) );
  XOR U46602 ( .A(n35349), .B(n33667), .Z(n36983) );
  IV U46603 ( .A(n33668), .Z(n33669) );
  NOR U46604 ( .A(n33669), .B(n35336), .Z(n33674) );
  IV U46605 ( .A(n33674), .Z(n33670) );
  NOR U46606 ( .A(n36983), .B(n33670), .Z(n38626) );
  IV U46607 ( .A(n33671), .Z(n33672) );
  NOR U46608 ( .A(n33672), .B(n35336), .Z(n35346) );
  NOR U46609 ( .A(n36982), .B(n35346), .Z(n33673) );
  XOR U46610 ( .A(n33673), .B(n36983), .Z(n35335) );
  NOR U46611 ( .A(n33674), .B(n35335), .Z(n33675) );
  NOR U46612 ( .A(n38626), .B(n33675), .Z(n33676) );
  IV U46613 ( .A(n33676), .Z(n33685) );
  XOR U46614 ( .A(n33677), .B(n33685), .Z(n35332) );
  XOR U46615 ( .A(n35331), .B(n35332), .Z(n33682) );
  NOR U46616 ( .A(n33678), .B(n33682), .Z(n38617) );
  IV U46617 ( .A(n33679), .Z(n33680) );
  NOR U46618 ( .A(n33681), .B(n33680), .Z(n33684) );
  IV U46619 ( .A(n33682), .Z(n33683) );
  NOR U46620 ( .A(n33684), .B(n33683), .Z(n33687) );
  IV U46621 ( .A(n33684), .Z(n33686) );
  NOR U46622 ( .A(n33686), .B(n33685), .Z(n40062) );
  NOR U46623 ( .A(n33687), .B(n40062), .Z(n33688) );
  NOR U46624 ( .A(n33689), .B(n33688), .Z(n33690) );
  NOR U46625 ( .A(n38617), .B(n33690), .Z(n33691) );
  IV U46626 ( .A(n33691), .Z(n35325) );
  XOR U46627 ( .A(n33692), .B(n35325), .Z(n36992) );
  XOR U46628 ( .A(n33693), .B(n36992), .Z(n35320) );
  XOR U46629 ( .A(n33694), .B(n35320), .Z(n36999) );
  IV U46630 ( .A(n33695), .Z(n33698) );
  IV U46631 ( .A(n33696), .Z(n33697) );
  NOR U46632 ( .A(n33698), .B(n33697), .Z(n35310) );
  NOR U46633 ( .A(n35313), .B(n35310), .Z(n33699) );
  XOR U46634 ( .A(n36999), .B(n33699), .Z(n35306) );
  XOR U46635 ( .A(n35304), .B(n35306), .Z(n40096) );
  XOR U46636 ( .A(n35307), .B(n40096), .Z(n35298) );
  IV U46637 ( .A(n33700), .Z(n33702) );
  NOR U46638 ( .A(n33702), .B(n33701), .Z(n35297) );
  IV U46639 ( .A(n33703), .Z(n33705) );
  NOR U46640 ( .A(n33705), .B(n33704), .Z(n33706) );
  IV U46641 ( .A(n33706), .Z(n33707) );
  NOR U46642 ( .A(n33708), .B(n33707), .Z(n35301) );
  NOR U46643 ( .A(n35297), .B(n35301), .Z(n33709) );
  XOR U46644 ( .A(n35298), .B(n33709), .Z(n37005) );
  XOR U46645 ( .A(n37003), .B(n37005), .Z(n37007) );
  XOR U46646 ( .A(n37006), .B(n37007), .Z(n37013) );
  IV U46647 ( .A(n33710), .Z(n33713) );
  IV U46648 ( .A(n33711), .Z(n33712) );
  NOR U46649 ( .A(n33713), .B(n33712), .Z(n37001) );
  IV U46650 ( .A(n33714), .Z(n33719) );
  NOR U46651 ( .A(n33716), .B(n33715), .Z(n33717) );
  IV U46652 ( .A(n33717), .Z(n33718) );
  NOR U46653 ( .A(n33719), .B(n33718), .Z(n37011) );
  NOR U46654 ( .A(n37001), .B(n37011), .Z(n33720) );
  XOR U46655 ( .A(n37013), .B(n33720), .Z(n35291) );
  XOR U46656 ( .A(n33721), .B(n35291), .Z(n35289) );
  NOR U46657 ( .A(n33729), .B(n35289), .Z(n41876) );
  IV U46658 ( .A(n33722), .Z(n33723) );
  NOR U46659 ( .A(n33726), .B(n33723), .Z(n35288) );
  XOR U46660 ( .A(n35288), .B(n35289), .Z(n35287) );
  IV U46661 ( .A(n33724), .Z(n33728) );
  NOR U46662 ( .A(n33726), .B(n33725), .Z(n33727) );
  IV U46663 ( .A(n33727), .Z(n33738) );
  NOR U46664 ( .A(n33728), .B(n33738), .Z(n33730) );
  IV U46665 ( .A(n33730), .Z(n35286) );
  XOR U46666 ( .A(n35287), .B(n35286), .Z(n33732) );
  NOR U46667 ( .A(n33730), .B(n33729), .Z(n33731) );
  NOR U46668 ( .A(n33732), .B(n33731), .Z(n33733) );
  NOR U46669 ( .A(n41876), .B(n33733), .Z(n35284) );
  IV U46670 ( .A(n33734), .Z(n33735) );
  NOR U46671 ( .A(n33736), .B(n33735), .Z(n37015) );
  IV U46672 ( .A(n33737), .Z(n33739) );
  NOR U46673 ( .A(n33739), .B(n33738), .Z(n35283) );
  NOR U46674 ( .A(n37015), .B(n35283), .Z(n33740) );
  XOR U46675 ( .A(n35284), .B(n33740), .Z(n38589) );
  NOR U46676 ( .A(n33741), .B(n38592), .Z(n37018) );
  XOR U46677 ( .A(n38589), .B(n37018), .Z(n37025) );
  XOR U46678 ( .A(n33742), .B(n37025), .Z(n37028) );
  XOR U46679 ( .A(n37027), .B(n37028), .Z(n37032) );
  XOR U46680 ( .A(n37031), .B(n37032), .Z(n40134) );
  XOR U46681 ( .A(n37034), .B(n40134), .Z(n33748) );
  IV U46682 ( .A(n33748), .Z(n37045) );
  XOR U46683 ( .A(n33747), .B(n37045), .Z(n33743) );
  NOR U46684 ( .A(n33754), .B(n33743), .Z(n38570) );
  IV U46685 ( .A(n33744), .Z(n33746) );
  NOR U46686 ( .A(n33746), .B(n33745), .Z(n37044) );
  NOR U46687 ( .A(n33747), .B(n37044), .Z(n33749) );
  XOR U46688 ( .A(n33749), .B(n33748), .Z(n35277) );
  IV U46689 ( .A(n33765), .Z(n33753) );
  NOR U46690 ( .A(n33750), .B(n33761), .Z(n33751) );
  IV U46691 ( .A(n33751), .Z(n33752) );
  NOR U46692 ( .A(n33753), .B(n33752), .Z(n33755) );
  IV U46693 ( .A(n33755), .Z(n35276) );
  XOR U46694 ( .A(n35277), .B(n35276), .Z(n33757) );
  NOR U46695 ( .A(n33755), .B(n33754), .Z(n33756) );
  NOR U46696 ( .A(n33757), .B(n33756), .Z(n33758) );
  NOR U46697 ( .A(n38570), .B(n33758), .Z(n33759) );
  IV U46698 ( .A(n33759), .Z(n37043) );
  IV U46699 ( .A(n33760), .Z(n33762) );
  NOR U46700 ( .A(n33762), .B(n33761), .Z(n33763) );
  IV U46701 ( .A(n33763), .Z(n33764) );
  NOR U46702 ( .A(n33765), .B(n33764), .Z(n37041) );
  XOR U46703 ( .A(n37043), .B(n37041), .Z(n37053) );
  XOR U46704 ( .A(n37052), .B(n37053), .Z(n35271) );
  XOR U46705 ( .A(n35270), .B(n35271), .Z(n35274) );
  IV U46706 ( .A(n33766), .Z(n33767) );
  NOR U46707 ( .A(n33768), .B(n33767), .Z(n35265) );
  NOR U46708 ( .A(n35273), .B(n35265), .Z(n33769) );
  XOR U46709 ( .A(n35274), .B(n33769), .Z(n35263) );
  XOR U46710 ( .A(n33770), .B(n35263), .Z(n35261) );
  XOR U46711 ( .A(n35259), .B(n35261), .Z(n37058) );
  IV U46712 ( .A(n33771), .Z(n33773) );
  NOR U46713 ( .A(n33773), .B(n33772), .Z(n37056) );
  XOR U46714 ( .A(n37058), .B(n37056), .Z(n37060) );
  XOR U46715 ( .A(n37059), .B(n37060), .Z(n37063) );
  XOR U46716 ( .A(n37064), .B(n37063), .Z(n37065) );
  IV U46717 ( .A(n33774), .Z(n33775) );
  NOR U46718 ( .A(n33776), .B(n33775), .Z(n38544) );
  IV U46719 ( .A(n33777), .Z(n33779) );
  NOR U46720 ( .A(n33779), .B(n33778), .Z(n38540) );
  NOR U46721 ( .A(n38544), .B(n38540), .Z(n37066) );
  XOR U46722 ( .A(n37065), .B(n37066), .Z(n35254) );
  XOR U46723 ( .A(n35251), .B(n35254), .Z(n35244) );
  XOR U46724 ( .A(n33780), .B(n35244), .Z(n35240) );
  XOR U46725 ( .A(n35239), .B(n35240), .Z(n37070) );
  IV U46726 ( .A(n33781), .Z(n33783) );
  NOR U46727 ( .A(n33783), .B(n33782), .Z(n37073) );
  IV U46728 ( .A(n33784), .Z(n33786) );
  NOR U46729 ( .A(n33786), .B(n33785), .Z(n37074) );
  NOR U46730 ( .A(n37073), .B(n37074), .Z(n33787) );
  XOR U46731 ( .A(n37070), .B(n33787), .Z(n35238) );
  XOR U46732 ( .A(n35236), .B(n35238), .Z(n35231) );
  XOR U46733 ( .A(n35230), .B(n35231), .Z(n35234) );
  XOR U46734 ( .A(n35233), .B(n35234), .Z(n35224) );
  XOR U46735 ( .A(n33788), .B(n35224), .Z(n35222) );
  XOR U46736 ( .A(n35221), .B(n35222), .Z(n35217) );
  XOR U46737 ( .A(n33789), .B(n35217), .Z(n35213) );
  XOR U46738 ( .A(n33790), .B(n35213), .Z(n37081) );
  XOR U46739 ( .A(n33791), .B(n37081), .Z(n35206) );
  IV U46740 ( .A(n33792), .Z(n33793) );
  NOR U46741 ( .A(n33794), .B(n33793), .Z(n35210) );
  NOR U46742 ( .A(n33796), .B(n33795), .Z(n35205) );
  NOR U46743 ( .A(n35210), .B(n35205), .Z(n33797) );
  XOR U46744 ( .A(n35206), .B(n33797), .Z(n37091) );
  XOR U46745 ( .A(n37090), .B(n37091), .Z(n35203) );
  XOR U46746 ( .A(n35202), .B(n35203), .Z(n37098) );
  XOR U46747 ( .A(n37096), .B(n37098), .Z(n37101) );
  XOR U46748 ( .A(n37099), .B(n37101), .Z(n37115) );
  XOR U46749 ( .A(n33798), .B(n37115), .Z(n35195) );
  XOR U46750 ( .A(n35194), .B(n35195), .Z(n35198) );
  XOR U46751 ( .A(n35197), .B(n35198), .Z(n37121) );
  IV U46752 ( .A(n33799), .Z(n33801) );
  NOR U46753 ( .A(n33801), .B(n33800), .Z(n37119) );
  XOR U46754 ( .A(n37121), .B(n37119), .Z(n37123) );
  XOR U46755 ( .A(n37122), .B(n37123), .Z(n35189) );
  XOR U46756 ( .A(n35188), .B(n35189), .Z(n35182) );
  NOR U46757 ( .A(n33802), .B(n35185), .Z(n33806) );
  IV U46758 ( .A(n33803), .Z(n33805) );
  IV U46759 ( .A(n33804), .Z(n33809) );
  NOR U46760 ( .A(n33805), .B(n33809), .Z(n35181) );
  NOR U46761 ( .A(n33806), .B(n35181), .Z(n33807) );
  XOR U46762 ( .A(n35182), .B(n33807), .Z(n35178) );
  IV U46763 ( .A(n33808), .Z(n33810) );
  NOR U46764 ( .A(n33810), .B(n33809), .Z(n35179) );
  IV U46765 ( .A(n33811), .Z(n33813) );
  NOR U46766 ( .A(n33813), .B(n33812), .Z(n37128) );
  NOR U46767 ( .A(n35179), .B(n37128), .Z(n33814) );
  XOR U46768 ( .A(n35178), .B(n33814), .Z(n37132) );
  XOR U46769 ( .A(n35175), .B(n37132), .Z(n35172) );
  IV U46770 ( .A(n33815), .Z(n33816) );
  NOR U46771 ( .A(n33817), .B(n33816), .Z(n35171) );
  NOR U46772 ( .A(n37131), .B(n35171), .Z(n33818) );
  XOR U46773 ( .A(n35172), .B(n33818), .Z(n37139) );
  IV U46774 ( .A(n33819), .Z(n33821) );
  NOR U46775 ( .A(n33821), .B(n33820), .Z(n37140) );
  IV U46776 ( .A(n33822), .Z(n33823) );
  NOR U46777 ( .A(n33823), .B(n33825), .Z(n37147) );
  NOR U46778 ( .A(n37140), .B(n37147), .Z(n33824) );
  XOR U46779 ( .A(n37139), .B(n33824), .Z(n37143) );
  NOR U46780 ( .A(n33826), .B(n33825), .Z(n33827) );
  IV U46781 ( .A(n33827), .Z(n37144) );
  NOR U46782 ( .A(n33828), .B(n37144), .Z(n33829) );
  XOR U46783 ( .A(n37143), .B(n33829), .Z(n37162) );
  NOR U46784 ( .A(n33831), .B(n33830), .Z(n35170) );
  IV U46785 ( .A(n33832), .Z(n33834) );
  NOR U46786 ( .A(n33834), .B(n33833), .Z(n37158) );
  NOR U46787 ( .A(n35170), .B(n37158), .Z(n37163) );
  XOR U46788 ( .A(n37162), .B(n37163), .Z(n33835) );
  IV U46789 ( .A(n33835), .Z(n35165) );
  XOR U46790 ( .A(n35164), .B(n35165), .Z(n35168) );
  XOR U46791 ( .A(n35167), .B(n35168), .Z(n37173) );
  XOR U46792 ( .A(n37171), .B(n37173), .Z(n37175) );
  XOR U46793 ( .A(n33836), .B(n37175), .Z(n35161) );
  NOR U46794 ( .A(n35161), .B(n33837), .Z(n33840) );
  IV U46795 ( .A(n33837), .Z(n35163) );
  XOR U46796 ( .A(n37174), .B(n37175), .Z(n33838) );
  NOR U46797 ( .A(n35163), .B(n33838), .Z(n33839) );
  NOR U46798 ( .A(n33840), .B(n33839), .Z(n35156) );
  XOR U46799 ( .A(n35157), .B(n35156), .Z(n37181) );
  IV U46800 ( .A(n33841), .Z(n33844) );
  IV U46801 ( .A(n33842), .Z(n33843) );
  NOR U46802 ( .A(n33844), .B(n33843), .Z(n37180) );
  NOR U46803 ( .A(n33845), .B(n37180), .Z(n33846) );
  XOR U46804 ( .A(n37181), .B(n33846), .Z(n37178) );
  XOR U46805 ( .A(n37179), .B(n37178), .Z(n35150) );
  IV U46806 ( .A(n33847), .Z(n33849) );
  NOR U46807 ( .A(n33849), .B(n33848), .Z(n35146) );
  IV U46808 ( .A(n33850), .Z(n33852) );
  NOR U46809 ( .A(n33852), .B(n33851), .Z(n35148) );
  NOR U46810 ( .A(n35146), .B(n35148), .Z(n33853) );
  XOR U46811 ( .A(n35150), .B(n33853), .Z(n33854) );
  IV U46812 ( .A(n33854), .Z(n35145) );
  XOR U46813 ( .A(n35143), .B(n35145), .Z(n37186) );
  XOR U46814 ( .A(n37184), .B(n37186), .Z(n37188) );
  XOR U46815 ( .A(n37187), .B(n37188), .Z(n35139) );
  XOR U46816 ( .A(n33855), .B(n35139), .Z(n35131) );
  XOR U46817 ( .A(n33856), .B(n35131), .Z(n35129) );
  XOR U46818 ( .A(n35127), .B(n35129), .Z(n37197) );
  XOR U46819 ( .A(n37195), .B(n37197), .Z(n37199) );
  XOR U46820 ( .A(n37198), .B(n37199), .Z(n37206) );
  XOR U46821 ( .A(n37205), .B(n37206), .Z(n35124) );
  XOR U46822 ( .A(n35123), .B(n35124), .Z(n37204) );
  XOR U46823 ( .A(n37202), .B(n37204), .Z(n37214) );
  XOR U46824 ( .A(n37213), .B(n37214), .Z(n37217) );
  XOR U46825 ( .A(n37216), .B(n37217), .Z(n33857) );
  XOR U46826 ( .A(n33858), .B(n33857), .Z(n35110) );
  XOR U46827 ( .A(n35109), .B(n35110), .Z(n35114) );
  XOR U46828 ( .A(n35112), .B(n35114), .Z(n35107) );
  XOR U46829 ( .A(n35106), .B(n35107), .Z(n37226) );
  XOR U46830 ( .A(n37224), .B(n37226), .Z(n37229) );
  XOR U46831 ( .A(n37227), .B(n37229), .Z(n38404) );
  XOR U46832 ( .A(n35101), .B(n38404), .Z(n35099) );
  IV U46833 ( .A(n33859), .Z(n33861) );
  NOR U46834 ( .A(n33861), .B(n33860), .Z(n35102) );
  IV U46835 ( .A(n33862), .Z(n33864) );
  NOR U46836 ( .A(n33864), .B(n33863), .Z(n35098) );
  NOR U46837 ( .A(n35102), .B(n35098), .Z(n33865) );
  XOR U46838 ( .A(n35099), .B(n33865), .Z(n35097) );
  XOR U46839 ( .A(n35095), .B(n35097), .Z(n35091) );
  XOR U46840 ( .A(n33866), .B(n35091), .Z(n35079) );
  XOR U46841 ( .A(n33867), .B(n35079), .Z(n35074) );
  XOR U46842 ( .A(n33868), .B(n35074), .Z(n35069) );
  XOR U46843 ( .A(n33869), .B(n35069), .Z(n35065) );
  XOR U46844 ( .A(n33870), .B(n35065), .Z(n35062) );
  XOR U46845 ( .A(n33871), .B(n35062), .Z(n35055) );
  IV U46846 ( .A(n33872), .Z(n33874) );
  NOR U46847 ( .A(n33874), .B(n33873), .Z(n33875) );
  IV U46848 ( .A(n33875), .Z(n35054) );
  XOR U46849 ( .A(n35055), .B(n35054), .Z(n35049) );
  IV U46850 ( .A(n33876), .Z(n33877) );
  NOR U46851 ( .A(n33878), .B(n33877), .Z(n35048) );
  IV U46852 ( .A(n33879), .Z(n33881) );
  NOR U46853 ( .A(n33881), .B(n33880), .Z(n35056) );
  NOR U46854 ( .A(n35048), .B(n35056), .Z(n33882) );
  XOR U46855 ( .A(n35049), .B(n33882), .Z(n35052) );
  XOR U46856 ( .A(n35051), .B(n35052), .Z(n37248) );
  XOR U46857 ( .A(n33883), .B(n37248), .Z(n35044) );
  XOR U46858 ( .A(n35043), .B(n35044), .Z(n35046) );
  XOR U46859 ( .A(n35047), .B(n35046), .Z(n35038) );
  IV U46860 ( .A(n33884), .Z(n33886) );
  NOR U46861 ( .A(n33886), .B(n33885), .Z(n35037) );
  NOR U46862 ( .A(n35040), .B(n35037), .Z(n33887) );
  XOR U46863 ( .A(n35038), .B(n33887), .Z(n35036) );
  XOR U46864 ( .A(n35034), .B(n35036), .Z(n37258) );
  XOR U46865 ( .A(n33888), .B(n37258), .Z(n37256) );
  XOR U46866 ( .A(n37254), .B(n37256), .Z(n35030) );
  XOR U46867 ( .A(n35031), .B(n35030), .Z(n33889) );
  XOR U46868 ( .A(n33890), .B(n33889), .Z(n37271) );
  IV U46869 ( .A(n33891), .Z(n33892) );
  NOR U46870 ( .A(n33893), .B(n33892), .Z(n37272) );
  IV U46871 ( .A(n33894), .Z(n33895) );
  NOR U46872 ( .A(n33896), .B(n33895), .Z(n37270) );
  NOR U46873 ( .A(n37272), .B(n37270), .Z(n33897) );
  XOR U46874 ( .A(n37271), .B(n33897), .Z(n37276) );
  XOR U46875 ( .A(n40353), .B(n37276), .Z(n38352) );
  XOR U46876 ( .A(n33898), .B(n38352), .Z(n37281) );
  XOR U46877 ( .A(n33899), .B(n37281), .Z(n37291) );
  IV U46878 ( .A(n33900), .Z(n33904) );
  NOR U46879 ( .A(n33902), .B(n33901), .Z(n33903) );
  IV U46880 ( .A(n33903), .Z(n33906) );
  NOR U46881 ( .A(n33904), .B(n33906), .Z(n37289) );
  XOR U46882 ( .A(n37291), .B(n37289), .Z(n37294) );
  IV U46883 ( .A(n33905), .Z(n33907) );
  NOR U46884 ( .A(n33907), .B(n33906), .Z(n37292) );
  XOR U46885 ( .A(n37294), .B(n37292), .Z(n35025) );
  XOR U46886 ( .A(n35026), .B(n35025), .Z(n35019) );
  IV U46887 ( .A(n33908), .Z(n33909) );
  NOR U46888 ( .A(n33910), .B(n33909), .Z(n35022) );
  IV U46889 ( .A(n33911), .Z(n33913) );
  NOR U46890 ( .A(n33913), .B(n33912), .Z(n35020) );
  NOR U46891 ( .A(n35022), .B(n35020), .Z(n33914) );
  XOR U46892 ( .A(n35019), .B(n33914), .Z(n35013) );
  XOR U46893 ( .A(n35011), .B(n35013), .Z(n35015) );
  XOR U46894 ( .A(n33915), .B(n35015), .Z(n35008) );
  XOR U46895 ( .A(n35007), .B(n35008), .Z(n37302) );
  XOR U46896 ( .A(n37301), .B(n37302), .Z(n37306) );
  XOR U46897 ( .A(n33916), .B(n37306), .Z(n34999) );
  XOR U46898 ( .A(n33917), .B(n34999), .Z(n34989) );
  XOR U46899 ( .A(n33918), .B(n34989), .Z(n34986) );
  NOR U46900 ( .A(n33920), .B(n34986), .Z(n41588) );
  IV U46901 ( .A(n33919), .Z(n34987) );
  XOR U46902 ( .A(n34987), .B(n34986), .Z(n34983) );
  XOR U46903 ( .A(n34982), .B(n34983), .Z(n33922) );
  NOR U46904 ( .A(n34983), .B(n33920), .Z(n33921) );
  NOR U46905 ( .A(n33922), .B(n33921), .Z(n33923) );
  NOR U46906 ( .A(n41588), .B(n33923), .Z(n33924) );
  IV U46907 ( .A(n33924), .Z(n34975) );
  IV U46908 ( .A(n33925), .Z(n34976) );
  IV U46909 ( .A(n33926), .Z(n33927) );
  NOR U46910 ( .A(n34976), .B(n33927), .Z(n33928) );
  XOR U46911 ( .A(n34975), .B(n33928), .Z(n37312) );
  XOR U46912 ( .A(n33929), .B(n37312), .Z(n37321) );
  XOR U46913 ( .A(n37320), .B(n37321), .Z(n34967) );
  XOR U46914 ( .A(n33930), .B(n34967), .Z(n34964) );
  NOR U46915 ( .A(n33932), .B(n33931), .Z(n33933) );
  XOR U46916 ( .A(n34964), .B(n33933), .Z(n34955) );
  IV U46917 ( .A(n33934), .Z(n33935) );
  NOR U46918 ( .A(n33938), .B(n33935), .Z(n34953) );
  XOR U46919 ( .A(n34955), .B(n34953), .Z(n34957) );
  XOR U46920 ( .A(n34956), .B(n34957), .Z(n37328) );
  IV U46921 ( .A(n33936), .Z(n33940) );
  NOR U46922 ( .A(n33938), .B(n33937), .Z(n33939) );
  IV U46923 ( .A(n33939), .Z(n33945) );
  NOR U46924 ( .A(n33940), .B(n33945), .Z(n37326) );
  XOR U46925 ( .A(n37328), .B(n37326), .Z(n37334) );
  IV U46926 ( .A(n33941), .Z(n33943) );
  IV U46927 ( .A(n33942), .Z(n33952) );
  NOR U46928 ( .A(n33943), .B(n33952), .Z(n37332) );
  IV U46929 ( .A(n33944), .Z(n33946) );
  NOR U46930 ( .A(n33946), .B(n33945), .Z(n37329) );
  NOR U46931 ( .A(n37332), .B(n37329), .Z(n33947) );
  XOR U46932 ( .A(n37334), .B(n33947), .Z(n34947) );
  IV U46933 ( .A(n33948), .Z(n33949) );
  NOR U46934 ( .A(n33950), .B(n33949), .Z(n34948) );
  IV U46935 ( .A(n33951), .Z(n33953) );
  NOR U46936 ( .A(n33953), .B(n33952), .Z(n34950) );
  NOR U46937 ( .A(n34948), .B(n34950), .Z(n33954) );
  XOR U46938 ( .A(n34947), .B(n33954), .Z(n34946) );
  IV U46939 ( .A(n33955), .Z(n33957) );
  NOR U46940 ( .A(n33957), .B(n33956), .Z(n34944) );
  XOR U46941 ( .A(n34946), .B(n34944), .Z(n34939) );
  XOR U46942 ( .A(n34938), .B(n34939), .Z(n34942) );
  XOR U46943 ( .A(n34941), .B(n34942), .Z(n37336) );
  XOR U46944 ( .A(n37335), .B(n37336), .Z(n37339) );
  XOR U46945 ( .A(n37338), .B(n37339), .Z(n34932) );
  XOR U46946 ( .A(n34931), .B(n34932), .Z(n34936) );
  IV U46947 ( .A(n33958), .Z(n33959) );
  NOR U46948 ( .A(n33960), .B(n33959), .Z(n34928) );
  IV U46949 ( .A(n33961), .Z(n33964) );
  IV U46950 ( .A(n33962), .Z(n33963) );
  NOR U46951 ( .A(n33964), .B(n33963), .Z(n34934) );
  NOR U46952 ( .A(n34928), .B(n34934), .Z(n33965) );
  XOR U46953 ( .A(n34936), .B(n33965), .Z(n34925) );
  XOR U46954 ( .A(n33966), .B(n34925), .Z(n34922) );
  IV U46955 ( .A(n33967), .Z(n33968) );
  NOR U46956 ( .A(n33969), .B(n33968), .Z(n34924) );
  IV U46957 ( .A(n33970), .Z(n33972) );
  NOR U46958 ( .A(n33972), .B(n33971), .Z(n34921) );
  NOR U46959 ( .A(n34924), .B(n34921), .Z(n33973) );
  XOR U46960 ( .A(n34922), .B(n33973), .Z(n33974) );
  IV U46961 ( .A(n33974), .Z(n34917) );
  IV U46962 ( .A(n33975), .Z(n33977) );
  NOR U46963 ( .A(n33977), .B(n33976), .Z(n34915) );
  XOR U46964 ( .A(n34917), .B(n34915), .Z(n38252) );
  XOR U46965 ( .A(n34918), .B(n38252), .Z(n34908) );
  IV U46966 ( .A(n33978), .Z(n33980) );
  NOR U46967 ( .A(n33980), .B(n33979), .Z(n34909) );
  IV U46968 ( .A(n33981), .Z(n33982) );
  NOR U46969 ( .A(n33983), .B(n33982), .Z(n34912) );
  NOR U46970 ( .A(n34909), .B(n34912), .Z(n33984) );
  XOR U46971 ( .A(n34908), .B(n33984), .Z(n37350) );
  XOR U46972 ( .A(n37348), .B(n37350), .Z(n37352) );
  XOR U46973 ( .A(n37351), .B(n37352), .Z(n34906) );
  XOR U46974 ( .A(n34905), .B(n34906), .Z(n34904) );
  XOR U46975 ( .A(n34902), .B(n34904), .Z(n34897) );
  XOR U46976 ( .A(n34896), .B(n34897), .Z(n34900) );
  XOR U46977 ( .A(n33985), .B(n34900), .Z(n34889) );
  IV U46978 ( .A(n33986), .Z(n33987) );
  NOR U46979 ( .A(n33988), .B(n33987), .Z(n34893) );
  IV U46980 ( .A(n33989), .Z(n33991) );
  NOR U46981 ( .A(n33991), .B(n33990), .Z(n34888) );
  NOR U46982 ( .A(n34893), .B(n34888), .Z(n33992) );
  XOR U46983 ( .A(n34889), .B(n33992), .Z(n34886) );
  XOR U46984 ( .A(n34885), .B(n34886), .Z(n34882) );
  XOR U46985 ( .A(n33993), .B(n34882), .Z(n34876) );
  XOR U46986 ( .A(n33994), .B(n34876), .Z(n37360) );
  XOR U46987 ( .A(n37358), .B(n37360), .Z(n34868) );
  XOR U46988 ( .A(n33995), .B(n34868), .Z(n34864) );
  XOR U46989 ( .A(n33996), .B(n34864), .Z(n37366) );
  XOR U46990 ( .A(n37365), .B(n37366), .Z(n37374) );
  XOR U46991 ( .A(n37368), .B(n33997), .Z(n33998) );
  XOR U46992 ( .A(n37374), .B(n33998), .Z(n34002) );
  IV U46993 ( .A(n34002), .Z(n33999) );
  NOR U46994 ( .A(n34000), .B(n33999), .Z(n34014) );
  IV U46995 ( .A(n34001), .Z(n34008) );
  NOR U46996 ( .A(n34003), .B(n34002), .Z(n34004) );
  IV U46997 ( .A(n34004), .Z(n34005) );
  NOR U46998 ( .A(n34006), .B(n34005), .Z(n34007) );
  IV U46999 ( .A(n34007), .Z(n34010) );
  NOR U47000 ( .A(n34008), .B(n34010), .Z(n38223) );
  IV U47001 ( .A(n34009), .Z(n34011) );
  NOR U47002 ( .A(n34011), .B(n34010), .Z(n38220) );
  NOR U47003 ( .A(n38223), .B(n38220), .Z(n34012) );
  IV U47004 ( .A(n34012), .Z(n34013) );
  NOR U47005 ( .A(n34014), .B(n34013), .Z(n34015) );
  IV U47006 ( .A(n34015), .Z(n34853) );
  XOR U47007 ( .A(n34852), .B(n34853), .Z(n37387) );
  XOR U47008 ( .A(n37386), .B(n37387), .Z(n37393) );
  XOR U47009 ( .A(n37389), .B(n37393), .Z(n34850) );
  XOR U47010 ( .A(n34016), .B(n34850), .Z(n34843) );
  XOR U47011 ( .A(n34017), .B(n34843), .Z(n34838) );
  XOR U47012 ( .A(n34837), .B(n34838), .Z(n34841) );
  XOR U47013 ( .A(n34840), .B(n34841), .Z(n37400) );
  XOR U47014 ( .A(n37399), .B(n37400), .Z(n37403) );
  XOR U47015 ( .A(n34018), .B(n37403), .Z(n37407) );
  XOR U47016 ( .A(n34019), .B(n37407), .Z(n37425) );
  XOR U47017 ( .A(n34020), .B(n37425), .Z(n37423) );
  XOR U47018 ( .A(n37421), .B(n37423), .Z(n40503) );
  XOR U47019 ( .A(n34021), .B(n40503), .Z(n37431) );
  XOR U47020 ( .A(n37432), .B(n37431), .Z(n37433) );
  IV U47021 ( .A(n34022), .Z(n34025) );
  IV U47022 ( .A(n34023), .Z(n34024) );
  NOR U47023 ( .A(n34025), .B(n34024), .Z(n40514) );
  IV U47024 ( .A(n34026), .Z(n34028) );
  NOR U47025 ( .A(n34028), .B(n34027), .Z(n40523) );
  NOR U47026 ( .A(n40514), .B(n40523), .Z(n37434) );
  XOR U47027 ( .A(n37433), .B(n37434), .Z(n34836) );
  XOR U47028 ( .A(n34834), .B(n34836), .Z(n37442) );
  XOR U47029 ( .A(n37440), .B(n37442), .Z(n37453) );
  XOR U47030 ( .A(n34029), .B(n37453), .Z(n37456) );
  XOR U47031 ( .A(n37455), .B(n37456), .Z(n37457) );
  IV U47032 ( .A(n34030), .Z(n34031) );
  NOR U47033 ( .A(n34039), .B(n34031), .Z(n40532) );
  IV U47034 ( .A(n34032), .Z(n34034) );
  NOR U47035 ( .A(n34034), .B(n34033), .Z(n38187) );
  NOR U47036 ( .A(n40532), .B(n38187), .Z(n37458) );
  XOR U47037 ( .A(n37457), .B(n37458), .Z(n34832) );
  XOR U47038 ( .A(n34830), .B(n34832), .Z(n34035) );
  NOR U47039 ( .A(n34036), .B(n34035), .Z(n47271) );
  IV U47040 ( .A(n34037), .Z(n34038) );
  NOR U47041 ( .A(n34039), .B(n34038), .Z(n34827) );
  NOR U47042 ( .A(n34827), .B(n34830), .Z(n34040) );
  XOR U47043 ( .A(n34832), .B(n34040), .Z(n34041) );
  NOR U47044 ( .A(n34042), .B(n34041), .Z(n34043) );
  NOR U47045 ( .A(n47271), .B(n34043), .Z(n34818) );
  NOR U47046 ( .A(n34045), .B(n34044), .Z(n34822) );
  IV U47047 ( .A(n34046), .Z(n34051) );
  IV U47048 ( .A(n34047), .Z(n34058) );
  NOR U47049 ( .A(n34048), .B(n34058), .Z(n34049) );
  IV U47050 ( .A(n34049), .Z(n34050) );
  NOR U47051 ( .A(n34051), .B(n34050), .Z(n34819) );
  NOR U47052 ( .A(n34822), .B(n34819), .Z(n34052) );
  XOR U47053 ( .A(n34818), .B(n34052), .Z(n34817) );
  IV U47054 ( .A(n34053), .Z(n34057) );
  NOR U47055 ( .A(n34054), .B(n34058), .Z(n34055) );
  IV U47056 ( .A(n34055), .Z(n34056) );
  NOR U47057 ( .A(n34057), .B(n34056), .Z(n34815) );
  XOR U47058 ( .A(n34817), .B(n34815), .Z(n34812) );
  NOR U47059 ( .A(n34059), .B(n34058), .Z(n34060) );
  IV U47060 ( .A(n34060), .Z(n34811) );
  NOR U47061 ( .A(n34061), .B(n34811), .Z(n34062) );
  XOR U47062 ( .A(n34812), .B(n34062), .Z(n37473) );
  XOR U47063 ( .A(n34063), .B(n37473), .Z(n34804) );
  XOR U47064 ( .A(n34064), .B(n34804), .Z(n37476) );
  XOR U47065 ( .A(n34065), .B(n37476), .Z(n34801) );
  XOR U47066 ( .A(n34799), .B(n34801), .Z(n34793) );
  XOR U47067 ( .A(n34792), .B(n34793), .Z(n34796) );
  XOR U47068 ( .A(n34795), .B(n34796), .Z(n34785) );
  IV U47069 ( .A(n34066), .Z(n34067) );
  NOR U47070 ( .A(n34786), .B(n34067), .Z(n34068) );
  XOR U47071 ( .A(n34785), .B(n34068), .Z(n37486) );
  XOR U47072 ( .A(n37485), .B(n37486), .Z(n37489) );
  XOR U47073 ( .A(n37488), .B(n37489), .Z(n34780) );
  IV U47074 ( .A(n34069), .Z(n34070) );
  NOR U47075 ( .A(n34071), .B(n34070), .Z(n34778) );
  XOR U47076 ( .A(n34780), .B(n34778), .Z(n34782) );
  IV U47077 ( .A(n34072), .Z(n34073) );
  NOR U47078 ( .A(n34074), .B(n34073), .Z(n34781) );
  IV U47079 ( .A(n34075), .Z(n34076) );
  NOR U47080 ( .A(n34076), .B(n34080), .Z(n34775) );
  NOR U47081 ( .A(n34781), .B(n34775), .Z(n34077) );
  XOR U47082 ( .A(n34782), .B(n34077), .Z(n37492) );
  IV U47083 ( .A(n34081), .Z(n34078) );
  NOR U47084 ( .A(n34078), .B(n34080), .Z(n40577) );
  IV U47085 ( .A(n34079), .Z(n34083) );
  XOR U47086 ( .A(n34081), .B(n34080), .Z(n34082) );
  NOR U47087 ( .A(n34083), .B(n34082), .Z(n40589) );
  NOR U47088 ( .A(n40577), .B(n40589), .Z(n37493) );
  XOR U47089 ( .A(n37492), .B(n37493), .Z(n37499) );
  IV U47090 ( .A(n34084), .Z(n34086) );
  IV U47091 ( .A(n34085), .Z(n37500) );
  NOR U47092 ( .A(n34086), .B(n37500), .Z(n37494) );
  XOR U47093 ( .A(n37499), .B(n37494), .Z(n34770) );
  XOR U47094 ( .A(n34771), .B(n34770), .Z(n37506) );
  IV U47095 ( .A(n34087), .Z(n34764) );
  NOR U47096 ( .A(n34088), .B(n34764), .Z(n34092) );
  IV U47097 ( .A(n34089), .Z(n34090) );
  NOR U47098 ( .A(n34091), .B(n34090), .Z(n37505) );
  NOR U47099 ( .A(n34092), .B(n37505), .Z(n34093) );
  XOR U47100 ( .A(n37506), .B(n34093), .Z(n37514) );
  IV U47101 ( .A(n34094), .Z(n34096) );
  NOR U47102 ( .A(n34096), .B(n34095), .Z(n34761) );
  XOR U47103 ( .A(n37514), .B(n34761), .Z(n34759) );
  XOR U47104 ( .A(n34097), .B(n34759), .Z(n34753) );
  XOR U47105 ( .A(n34098), .B(n34753), .Z(n37520) );
  XOR U47106 ( .A(n34099), .B(n37520), .Z(n34750) );
  XOR U47107 ( .A(n34100), .B(n34750), .Z(n34734) );
  NOR U47108 ( .A(n34101), .B(n34735), .Z(n34102) );
  NOR U47109 ( .A(n34102), .B(n34736), .Z(n34103) );
  XOR U47110 ( .A(n34734), .B(n34103), .Z(n34731) );
  XOR U47111 ( .A(n34104), .B(n34731), .Z(n37525) );
  XOR U47112 ( .A(n34105), .B(n37525), .Z(n37533) );
  XOR U47113 ( .A(n37531), .B(n37533), .Z(n37536) );
  IV U47114 ( .A(n34106), .Z(n34107) );
  NOR U47115 ( .A(n34109), .B(n34107), .Z(n34725) );
  IV U47116 ( .A(n34108), .Z(n34110) );
  NOR U47117 ( .A(n34110), .B(n34109), .Z(n37534) );
  NOR U47118 ( .A(n34725), .B(n37534), .Z(n34111) );
  XOR U47119 ( .A(n37536), .B(n34111), .Z(n34716) );
  XOR U47120 ( .A(n34112), .B(n34716), .Z(n44015) );
  XOR U47121 ( .A(n34113), .B(n44015), .Z(n34709) );
  IV U47122 ( .A(n34114), .Z(n34117) );
  NOR U47123 ( .A(n34115), .B(n44023), .Z(n34116) );
  IV U47124 ( .A(n34116), .Z(n34122) );
  NOR U47125 ( .A(n34117), .B(n34122), .Z(n34707) );
  XOR U47126 ( .A(n34709), .B(n34707), .Z(n37544) );
  IV U47127 ( .A(n34118), .Z(n34119) );
  NOR U47128 ( .A(n34120), .B(n34119), .Z(n37543) );
  IV U47129 ( .A(n34121), .Z(n34123) );
  NOR U47130 ( .A(n34123), .B(n34122), .Z(n34710) );
  NOR U47131 ( .A(n37543), .B(n34710), .Z(n34124) );
  XOR U47132 ( .A(n37544), .B(n34124), .Z(n34702) );
  IV U47133 ( .A(n34125), .Z(n34127) );
  NOR U47134 ( .A(n34127), .B(n34126), .Z(n37540) );
  IV U47135 ( .A(n34128), .Z(n34130) );
  NOR U47136 ( .A(n34130), .B(n34129), .Z(n34703) );
  NOR U47137 ( .A(n37540), .B(n34703), .Z(n34131) );
  XOR U47138 ( .A(n34702), .B(n34131), .Z(n37551) );
  IV U47139 ( .A(n34132), .Z(n34134) );
  NOR U47140 ( .A(n34134), .B(n34133), .Z(n34705) );
  IV U47141 ( .A(n34135), .Z(n34136) );
  NOR U47142 ( .A(n34137), .B(n34136), .Z(n37550) );
  NOR U47143 ( .A(n34705), .B(n37550), .Z(n34138) );
  XOR U47144 ( .A(n37551), .B(n34138), .Z(n34139) );
  IV U47145 ( .A(n34139), .Z(n37549) );
  XOR U47146 ( .A(n37547), .B(n37549), .Z(n37555) );
  XOR U47147 ( .A(n37554), .B(n37555), .Z(n37558) );
  XOR U47148 ( .A(n37557), .B(n37558), .Z(n34700) );
  XOR U47149 ( .A(n34140), .B(n34700), .Z(n34696) );
  IV U47150 ( .A(n34141), .Z(n34144) );
  IV U47151 ( .A(n34142), .Z(n34143) );
  NOR U47152 ( .A(n34144), .B(n34143), .Z(n34145) );
  IV U47153 ( .A(n34145), .Z(n34695) );
  XOR U47154 ( .A(n34696), .B(n34695), .Z(n34693) );
  IV U47155 ( .A(n34146), .Z(n34147) );
  NOR U47156 ( .A(n34148), .B(n34147), .Z(n37561) );
  IV U47157 ( .A(n34149), .Z(n34150) );
  NOR U47158 ( .A(n34151), .B(n34150), .Z(n51653) );
  NOR U47159 ( .A(n37561), .B(n51653), .Z(n34152) );
  XOR U47160 ( .A(n34693), .B(n34152), .Z(n37564) );
  XOR U47161 ( .A(n37562), .B(n37564), .Z(n37571) );
  XOR U47162 ( .A(n37569), .B(n37571), .Z(n34690) );
  XOR U47163 ( .A(n34689), .B(n34690), .Z(n37568) );
  XOR U47164 ( .A(n37566), .B(n37568), .Z(n37579) );
  XOR U47165 ( .A(n37577), .B(n37579), .Z(n37581) );
  XOR U47166 ( .A(n37580), .B(n37581), .Z(n37587) );
  XOR U47167 ( .A(n37586), .B(n37587), .Z(n34686) );
  XOR U47168 ( .A(n34685), .B(n34686), .Z(n37601) );
  XOR U47169 ( .A(n34153), .B(n37601), .Z(n37604) );
  XOR U47170 ( .A(n37603), .B(n37604), .Z(n38091) );
  IV U47171 ( .A(n38091), .Z(n34159) );
  IV U47172 ( .A(n34154), .Z(n34156) );
  NOR U47173 ( .A(n34156), .B(n34155), .Z(n38090) );
  IV U47174 ( .A(n34157), .Z(n34158) );
  NOR U47175 ( .A(n34158), .B(n34678), .Z(n40706) );
  NOR U47176 ( .A(n38090), .B(n40706), .Z(n34684) );
  XOR U47177 ( .A(n34159), .B(n34684), .Z(n34677) );
  XOR U47178 ( .A(n34160), .B(n34677), .Z(n34666) );
  XOR U47179 ( .A(n34161), .B(n34666), .Z(n34655) );
  XOR U47180 ( .A(n34162), .B(n34655), .Z(n34649) );
  XOR U47181 ( .A(n34648), .B(n34649), .Z(n34653) );
  XOR U47182 ( .A(n34651), .B(n34653), .Z(n34644) );
  XOR U47183 ( .A(n34642), .B(n34644), .Z(n34646) );
  XOR U47184 ( .A(n34645), .B(n34646), .Z(n34635) );
  XOR U47185 ( .A(n34163), .B(n34635), .Z(n34629) );
  XOR U47186 ( .A(n34628), .B(n34629), .Z(n34632) );
  XOR U47187 ( .A(n34631), .B(n34632), .Z(n37614) );
  XOR U47188 ( .A(n37613), .B(n37614), .Z(n37618) );
  XOR U47189 ( .A(n37616), .B(n37618), .Z(n37621) );
  XOR U47190 ( .A(n37620), .B(n37621), .Z(n37625) );
  XOR U47191 ( .A(n37623), .B(n37625), .Z(n34626) );
  XOR U47192 ( .A(n34625), .B(n34626), .Z(n34620) );
  XOR U47193 ( .A(n34619), .B(n34620), .Z(n34623) );
  XOR U47194 ( .A(n34622), .B(n34623), .Z(n38046) );
  XOR U47195 ( .A(n34164), .B(n38046), .Z(n37635) );
  XOR U47196 ( .A(n37636), .B(n37635), .Z(n34613) );
  IV U47197 ( .A(n34165), .Z(n34170) );
  IV U47198 ( .A(n34166), .Z(n34168) );
  NOR U47199 ( .A(n34168), .B(n34167), .Z(n34169) );
  IV U47200 ( .A(n34169), .Z(n34173) );
  NOR U47201 ( .A(n34170), .B(n34173), .Z(n34614) );
  NOR U47202 ( .A(n34617), .B(n34614), .Z(n34171) );
  XOR U47203 ( .A(n34613), .B(n34171), .Z(n34612) );
  IV U47204 ( .A(n34172), .Z(n34174) );
  NOR U47205 ( .A(n34174), .B(n34173), .Z(n34610) );
  XOR U47206 ( .A(n34612), .B(n34610), .Z(n34604) );
  IV U47207 ( .A(n34175), .Z(n34176) );
  NOR U47208 ( .A(n34177), .B(n34176), .Z(n34178) );
  IV U47209 ( .A(n34178), .Z(n34603) );
  NOR U47210 ( .A(n34179), .B(n34603), .Z(n34180) );
  XOR U47211 ( .A(n34604), .B(n34180), .Z(n34601) );
  XOR U47212 ( .A(n34599), .B(n34601), .Z(n34595) );
  XOR U47213 ( .A(n34181), .B(n34595), .Z(n37644) );
  XOR U47214 ( .A(n37642), .B(n37644), .Z(n34592) );
  IV U47215 ( .A(n34182), .Z(n34184) );
  NOR U47216 ( .A(n34184), .B(n34183), .Z(n34590) );
  XOR U47217 ( .A(n34592), .B(n34590), .Z(n37640) );
  XOR U47218 ( .A(n37639), .B(n37640), .Z(n37653) );
  XOR U47219 ( .A(n37654), .B(n37653), .Z(n34587) );
  IV U47220 ( .A(n34185), .Z(n34186) );
  NOR U47221 ( .A(n34187), .B(n34186), .Z(n37650) );
  IV U47222 ( .A(n34187), .Z(n34189) );
  NOR U47223 ( .A(n34189), .B(n34188), .Z(n34588) );
  NOR U47224 ( .A(n37650), .B(n34588), .Z(n34190) );
  XOR U47225 ( .A(n34587), .B(n34190), .Z(n37660) );
  XOR U47226 ( .A(n37659), .B(n37660), .Z(n37666) );
  XOR U47227 ( .A(n34191), .B(n37666), .Z(n37668) );
  XOR U47228 ( .A(n37670), .B(n37668), .Z(n34580) );
  XOR U47229 ( .A(n34578), .B(n34580), .Z(n34583) );
  XOR U47230 ( .A(n34581), .B(n34583), .Z(n34577) );
  XOR U47231 ( .A(n34575), .B(n34577), .Z(n34568) );
  XOR U47232 ( .A(n34566), .B(n34568), .Z(n34570) );
  XOR U47233 ( .A(n34192), .B(n34570), .Z(n34564) );
  XOR U47234 ( .A(n34193), .B(n34564), .Z(n34556) );
  XOR U47235 ( .A(n34554), .B(n34556), .Z(n37675) );
  XOR U47236 ( .A(n37674), .B(n37675), .Z(n37677) );
  XOR U47237 ( .A(n34194), .B(n37677), .Z(n34550) );
  XOR U47238 ( .A(n34549), .B(n34550), .Z(n34547) );
  IV U47239 ( .A(n34195), .Z(n34196) );
  NOR U47240 ( .A(n34197), .B(n34196), .Z(n34552) );
  NOR U47241 ( .A(n34211), .B(n34198), .Z(n34546) );
  NOR U47242 ( .A(n34552), .B(n34546), .Z(n34199) );
  XOR U47243 ( .A(n34547), .B(n34199), .Z(n34213) );
  IV U47244 ( .A(n34213), .Z(n34200) );
  NOR U47245 ( .A(n34200), .B(n34211), .Z(n34201) );
  IV U47246 ( .A(n34201), .Z(n34202) );
  NOR U47247 ( .A(n34203), .B(n34202), .Z(n34204) );
  IV U47248 ( .A(n34204), .Z(n34207) );
  NOR U47249 ( .A(n34205), .B(n34207), .Z(n40860) );
  IV U47250 ( .A(n34206), .Z(n34208) );
  NOR U47251 ( .A(n34208), .B(n34207), .Z(n40857) );
  NOR U47252 ( .A(n40860), .B(n40857), .Z(n34209) );
  IV U47253 ( .A(n34209), .Z(n34216) );
  IV U47254 ( .A(n34210), .Z(n34212) );
  NOR U47255 ( .A(n34212), .B(n34211), .Z(n34214) );
  NOR U47256 ( .A(n34214), .B(n34213), .Z(n34215) );
  NOR U47257 ( .A(n34216), .B(n34215), .Z(n34217) );
  IV U47258 ( .A(n34217), .Z(n37685) );
  XOR U47259 ( .A(n37684), .B(n37685), .Z(n37690) );
  XOR U47260 ( .A(n37688), .B(n37690), .Z(n37692) );
  XOR U47261 ( .A(n37691), .B(n37692), .Z(n40871) );
  XOR U47262 ( .A(n37695), .B(n40871), .Z(n37708) );
  XOR U47263 ( .A(n37707), .B(n37708), .Z(n37714) );
  XOR U47264 ( .A(n37713), .B(n37714), .Z(n37717) );
  NOR U47265 ( .A(n34224), .B(n37717), .Z(n34545) );
  IV U47266 ( .A(n34218), .Z(n34220) );
  NOR U47267 ( .A(n34220), .B(n34219), .Z(n37716) );
  XOR U47268 ( .A(n37716), .B(n37717), .Z(n34544) );
  IV U47269 ( .A(n34221), .Z(n34223) );
  NOR U47270 ( .A(n34223), .B(n34222), .Z(n34225) );
  IV U47271 ( .A(n34225), .Z(n34543) );
  XOR U47272 ( .A(n34544), .B(n34543), .Z(n34227) );
  NOR U47273 ( .A(n34225), .B(n34224), .Z(n34226) );
  NOR U47274 ( .A(n34227), .B(n34226), .Z(n34228) );
  NOR U47275 ( .A(n34545), .B(n34228), .Z(n34229) );
  IV U47276 ( .A(n34229), .Z(n34542) );
  IV U47277 ( .A(n34230), .Z(n34232) );
  NOR U47278 ( .A(n34232), .B(n34231), .Z(n34540) );
  XOR U47279 ( .A(n34542), .B(n34540), .Z(n37721) );
  IV U47280 ( .A(n37721), .Z(n34236) );
  NOR U47281 ( .A(n34234), .B(n34233), .Z(n34235) );
  XOR U47282 ( .A(n34236), .B(n34235), .Z(n34529) );
  IV U47283 ( .A(n34237), .Z(n34528) );
  IV U47284 ( .A(n34238), .Z(n34239) );
  NOR U47285 ( .A(n34528), .B(n34239), .Z(n34240) );
  XOR U47286 ( .A(n34529), .B(n34240), .Z(n37744) );
  XOR U47287 ( .A(n37742), .B(n37744), .Z(n37746) );
  XOR U47288 ( .A(n37745), .B(n37746), .Z(n34521) );
  XOR U47289 ( .A(n34520), .B(n34521), .Z(n34524) );
  XOR U47290 ( .A(n34523), .B(n34524), .Z(n37767) );
  XOR U47291 ( .A(n34241), .B(n37767), .Z(n37749) );
  IV U47292 ( .A(n34242), .Z(n34243) );
  NOR U47293 ( .A(n34244), .B(n34243), .Z(n34519) );
  IV U47294 ( .A(n34245), .Z(n34246) );
  NOR U47295 ( .A(n34247), .B(n34246), .Z(n37752) );
  NOR U47296 ( .A(n34519), .B(n37752), .Z(n37761) );
  XOR U47297 ( .A(n37749), .B(n37761), .Z(n37997) );
  XOR U47298 ( .A(n34248), .B(n37997), .Z(n37777) );
  XOR U47299 ( .A(n37775), .B(n37777), .Z(n37780) );
  IV U47300 ( .A(n34249), .Z(n34251) );
  NOR U47301 ( .A(n34251), .B(n34250), .Z(n37778) );
  XOR U47302 ( .A(n37780), .B(n37778), .Z(n34512) );
  XOR U47303 ( .A(n34252), .B(n34512), .Z(n34507) );
  IV U47304 ( .A(n34253), .Z(n34255) );
  NOR U47305 ( .A(n34255), .B(n34254), .Z(n34509) );
  IV U47306 ( .A(n34256), .Z(n34258) );
  NOR U47307 ( .A(n34258), .B(n34257), .Z(n34506) );
  NOR U47308 ( .A(n34509), .B(n34506), .Z(n34259) );
  XOR U47309 ( .A(n34507), .B(n34259), .Z(n34260) );
  IV U47310 ( .A(n34260), .Z(n34505) );
  XOR U47311 ( .A(n34503), .B(n34505), .Z(n34498) );
  XOR U47312 ( .A(n34497), .B(n34498), .Z(n37788) );
  IV U47313 ( .A(n34261), .Z(n34262) );
  NOR U47314 ( .A(n34262), .B(n34273), .Z(n34495) );
  IV U47315 ( .A(n34277), .Z(n34266) );
  NOR U47316 ( .A(n34263), .B(n34273), .Z(n34264) );
  IV U47317 ( .A(n34264), .Z(n34265) );
  NOR U47318 ( .A(n34266), .B(n34265), .Z(n37786) );
  NOR U47319 ( .A(n34495), .B(n37786), .Z(n34267) );
  XOR U47320 ( .A(n34500), .B(n34267), .Z(n34268) );
  XOR U47321 ( .A(n37788), .B(n34268), .Z(n34279) );
  IV U47322 ( .A(n34279), .Z(n37791) );
  IV U47323 ( .A(n34269), .Z(n34270) );
  NOR U47324 ( .A(n34280), .B(n34270), .Z(n34287) );
  IV U47325 ( .A(n34287), .Z(n34271) );
  NOR U47326 ( .A(n37791), .B(n34271), .Z(n37974) );
  IV U47327 ( .A(n34272), .Z(n34274) );
  NOR U47328 ( .A(n34274), .B(n34273), .Z(n34275) );
  IV U47329 ( .A(n34275), .Z(n34276) );
  NOR U47330 ( .A(n34277), .B(n34276), .Z(n34278) );
  IV U47331 ( .A(n34278), .Z(n37790) );
  XOR U47332 ( .A(n37790), .B(n34279), .Z(n37793) );
  IV U47333 ( .A(n34280), .Z(n34285) );
  NOR U47334 ( .A(n34282), .B(n34281), .Z(n34283) );
  IV U47335 ( .A(n34283), .Z(n34284) );
  NOR U47336 ( .A(n34285), .B(n34284), .Z(n34286) );
  IV U47337 ( .A(n34286), .Z(n37792) );
  XOR U47338 ( .A(n37793), .B(n37792), .Z(n34291) );
  NOR U47339 ( .A(n34291), .B(n34287), .Z(n34288) );
  NOR U47340 ( .A(n37974), .B(n34288), .Z(n34289) );
  NOR U47341 ( .A(n34290), .B(n34289), .Z(n34294) );
  IV U47342 ( .A(n34290), .Z(n34293) );
  IV U47343 ( .A(n34291), .Z(n34292) );
  NOR U47344 ( .A(n34293), .B(n34292), .Z(n40960) );
  NOR U47345 ( .A(n34294), .B(n40960), .Z(n34492) );
  XOR U47346 ( .A(n34494), .B(n34492), .Z(n37796) );
  XOR U47347 ( .A(n37797), .B(n37796), .Z(n37798) );
  NOR U47348 ( .A(n34296), .B(n34295), .Z(n40970) );
  NOR U47349 ( .A(n37801), .B(n40970), .Z(n34297) );
  XOR U47350 ( .A(n37798), .B(n34297), .Z(n37803) );
  XOR U47351 ( .A(n37802), .B(n37803), .Z(n34490) );
  XOR U47352 ( .A(n34298), .B(n34490), .Z(n37814) );
  XOR U47353 ( .A(n37812), .B(n37814), .Z(n37816) );
  IV U47354 ( .A(n34299), .Z(n34302) );
  NOR U47355 ( .A(n34300), .B(n34313), .Z(n34301) );
  IV U47356 ( .A(n34301), .Z(n34309) );
  NOR U47357 ( .A(n34302), .B(n34309), .Z(n34303) );
  IV U47358 ( .A(n34303), .Z(n37815) );
  XOR U47359 ( .A(n37816), .B(n37815), .Z(n34484) );
  IV U47360 ( .A(n34317), .Z(n34307) );
  NOR U47361 ( .A(n34304), .B(n34313), .Z(n34305) );
  IV U47362 ( .A(n34305), .Z(n34306) );
  NOR U47363 ( .A(n34307), .B(n34306), .Z(n34485) );
  IV U47364 ( .A(n34308), .Z(n34310) );
  NOR U47365 ( .A(n34310), .B(n34309), .Z(n37818) );
  NOR U47366 ( .A(n34485), .B(n37818), .Z(n34311) );
  XOR U47367 ( .A(n34484), .B(n34311), .Z(n34483) );
  IV U47368 ( .A(n34312), .Z(n34314) );
  NOR U47369 ( .A(n34314), .B(n34313), .Z(n34315) );
  IV U47370 ( .A(n34315), .Z(n34316) );
  NOR U47371 ( .A(n34317), .B(n34316), .Z(n34481) );
  XOR U47372 ( .A(n34483), .B(n34481), .Z(n34477) );
  XOR U47373 ( .A(n34475), .B(n34477), .Z(n34480) );
  XOR U47374 ( .A(n34478), .B(n34480), .Z(n34473) );
  XOR U47375 ( .A(n34472), .B(n34473), .Z(n37823) );
  IV U47376 ( .A(n34318), .Z(n34319) );
  NOR U47377 ( .A(n34320), .B(n34319), .Z(n34470) );
  IV U47378 ( .A(n34321), .Z(n34322) );
  NOR U47379 ( .A(n37825), .B(n34322), .Z(n37822) );
  NOR U47380 ( .A(n34470), .B(n37822), .Z(n34323) );
  XOR U47381 ( .A(n37823), .B(n34323), .Z(n34324) );
  IV U47382 ( .A(n34324), .Z(n37826) );
  XOR U47383 ( .A(n34468), .B(n37826), .Z(n34327) );
  IV U47384 ( .A(n34325), .Z(n37829) );
  NOR U47385 ( .A(n34329), .B(n37829), .Z(n34326) );
  XOR U47386 ( .A(n34327), .B(n34326), .Z(n37832) );
  IV U47387 ( .A(n34328), .Z(n34330) );
  NOR U47388 ( .A(n34330), .B(n34329), .Z(n37830) );
  XOR U47389 ( .A(n37832), .B(n37830), .Z(n37834) );
  XOR U47390 ( .A(n37833), .B(n37834), .Z(n37838) );
  XOR U47391 ( .A(n37837), .B(n37838), .Z(n37841) );
  XOR U47392 ( .A(n37840), .B(n37841), .Z(n37846) );
  NOR U47393 ( .A(n34332), .B(n34331), .Z(n34333) );
  IV U47394 ( .A(n34333), .Z(n37845) );
  NOR U47395 ( .A(n34334), .B(n37845), .Z(n34335) );
  XOR U47396 ( .A(n37846), .B(n34335), .Z(n34466) );
  XOR U47397 ( .A(n34464), .B(n34466), .Z(n34461) );
  IV U47398 ( .A(n34336), .Z(n34337) );
  NOR U47399 ( .A(n34338), .B(n34337), .Z(n34465) );
  IV U47400 ( .A(n34339), .Z(n34340) );
  NOR U47401 ( .A(n34341), .B(n34340), .Z(n34460) );
  NOR U47402 ( .A(n34465), .B(n34460), .Z(n34342) );
  XOR U47403 ( .A(n34461), .B(n34342), .Z(n34459) );
  IV U47404 ( .A(n34343), .Z(n34345) );
  NOR U47405 ( .A(n34345), .B(n34344), .Z(n34457) );
  XOR U47406 ( .A(n34459), .B(n34457), .Z(n37857) );
  XOR U47407 ( .A(n37856), .B(n37857), .Z(n37861) );
  XOR U47408 ( .A(n37859), .B(n37861), .Z(n37866) );
  XOR U47409 ( .A(n34346), .B(n37866), .Z(n37869) );
  NOR U47410 ( .A(n37870), .B(n34347), .Z(n34348) );
  IV U47411 ( .A(n34348), .Z(n37864) );
  XOR U47412 ( .A(n37869), .B(n37864), .Z(n34349) );
  XOR U47413 ( .A(n34350), .B(n34349), .Z(n37876) );
  IV U47414 ( .A(n34351), .Z(n34353) );
  NOR U47415 ( .A(n34353), .B(n34352), .Z(n34354) );
  IV U47416 ( .A(n34354), .Z(n37875) );
  XOR U47417 ( .A(n37876), .B(n37875), .Z(n34455) );
  IV U47418 ( .A(n34355), .Z(n34356) );
  NOR U47419 ( .A(n34357), .B(n34356), .Z(n37877) );
  IV U47420 ( .A(n34358), .Z(n34359) );
  NOR U47421 ( .A(n34360), .B(n34359), .Z(n34454) );
  NOR U47422 ( .A(n37877), .B(n34454), .Z(n34361) );
  XOR U47423 ( .A(n34455), .B(n34361), .Z(n34449) );
  XOR U47424 ( .A(n34447), .B(n34449), .Z(n34451) );
  XOR U47425 ( .A(n34362), .B(n34451), .Z(n34363) );
  IV U47426 ( .A(n34363), .Z(n37886) );
  IV U47427 ( .A(n34364), .Z(n34365) );
  NOR U47428 ( .A(n34366), .B(n34365), .Z(n37884) );
  XOR U47429 ( .A(n37886), .B(n37884), .Z(n41073) );
  NOR U47430 ( .A(n34370), .B(n34366), .Z(n34367) );
  IV U47431 ( .A(n34367), .Z(n41066) );
  NOR U47432 ( .A(n34368), .B(n41066), .Z(n37887) );
  XOR U47433 ( .A(n41073), .B(n37887), .Z(n37893) );
  IV U47434 ( .A(n34369), .Z(n41064) );
  NOR U47435 ( .A(n34370), .B(n41064), .Z(n34383) );
  IV U47436 ( .A(n34383), .Z(n34371) );
  NOR U47437 ( .A(n34372), .B(n34371), .Z(n37891) );
  XOR U47438 ( .A(n37893), .B(n37891), .Z(n34439) );
  XOR U47439 ( .A(n34438), .B(n34439), .Z(n37904) );
  IV U47440 ( .A(n34373), .Z(n34375) );
  NOR U47441 ( .A(n34375), .B(n34374), .Z(n34378) );
  IV U47442 ( .A(n34378), .Z(n34376) );
  NOR U47443 ( .A(n34377), .B(n34376), .Z(n37902) );
  XOR U47444 ( .A(n37904), .B(n37902), .Z(n34437) );
  NOR U47445 ( .A(n34379), .B(n34378), .Z(n34381) );
  XOR U47446 ( .A(n34380), .B(n34381), .Z(n34398) );
  IV U47447 ( .A(n34398), .Z(n34409) );
  NOR U47448 ( .A(n34381), .B(n34380), .Z(n34382) );
  NOR U47449 ( .A(n34383), .B(n34382), .Z(n34384) );
  XOR U47450 ( .A(n34385), .B(n34384), .Z(n34414) );
  NOR U47451 ( .A(n34409), .B(n34414), .Z(n34386) );
  IV U47452 ( .A(n34386), .Z(n34395) );
  IV U47453 ( .A(n34387), .Z(n34389) );
  NOR U47454 ( .A(n34389), .B(n34388), .Z(n34397) );
  IV U47455 ( .A(n34397), .Z(n34390) );
  NOR U47456 ( .A(n34395), .B(n34390), .Z(n34435) );
  XOR U47457 ( .A(n34437), .B(n34435), .Z(n37916) );
  IV U47458 ( .A(n34391), .Z(n34393) );
  NOR U47459 ( .A(n34393), .B(n34392), .Z(n34396) );
  IV U47460 ( .A(n34396), .Z(n34394) );
  NOR U47461 ( .A(n34395), .B(n34394), .Z(n37914) );
  XOR U47462 ( .A(n37916), .B(n37914), .Z(n37919) );
  NOR U47463 ( .A(n34397), .B(n34396), .Z(n34410) );
  XOR U47464 ( .A(n34398), .B(n34410), .Z(n34415) );
  IV U47465 ( .A(n34399), .Z(n34401) );
  NOR U47466 ( .A(n34401), .B(n34400), .Z(n34417) );
  IV U47467 ( .A(n34417), .Z(n34402) );
  NOR U47468 ( .A(n34415), .B(n34402), .Z(n34411) );
  IV U47469 ( .A(n34411), .Z(n34403) );
  NOR U47470 ( .A(n34414), .B(n34403), .Z(n37917) );
  XOR U47471 ( .A(n37919), .B(n37917), .Z(n34433) );
  IV U47472 ( .A(n34404), .Z(n34406) );
  NOR U47473 ( .A(n34406), .B(n34405), .Z(n34416) );
  IV U47474 ( .A(n34416), .Z(n34407) );
  NOR U47475 ( .A(n34415), .B(n34407), .Z(n44354) );
  IV U47476 ( .A(n44354), .Z(n34408) );
  NOR U47477 ( .A(n34414), .B(n34408), .Z(n44356) );
  XOR U47478 ( .A(n34433), .B(n44356), .Z(n41054) );
  NOR U47479 ( .A(n34410), .B(n34409), .Z(n34412) );
  NOR U47480 ( .A(n34412), .B(n34411), .Z(n34413) );
  XOR U47481 ( .A(n34414), .B(n34413), .Z(n44353) );
  IV U47482 ( .A(n44353), .Z(n44386) );
  IV U47483 ( .A(n34415), .Z(n34419) );
  NOR U47484 ( .A(n34417), .B(n34416), .Z(n34418) );
  XOR U47485 ( .A(n34419), .B(n34418), .Z(n44348) );
  IV U47486 ( .A(n34420), .Z(n34422) );
  NOR U47487 ( .A(n34422), .B(n34421), .Z(n44347) );
  IV U47488 ( .A(n44347), .Z(n34423) );
  NOR U47489 ( .A(n44348), .B(n34423), .Z(n44383) );
  IV U47490 ( .A(n44383), .Z(n34424) );
  NOR U47491 ( .A(n44386), .B(n34424), .Z(n34425) );
  IV U47492 ( .A(n34425), .Z(n41053) );
  XOR U47493 ( .A(n41054), .B(n41053), .Z(n44377) );
  IV U47494 ( .A(n44377), .Z(n44346) );
  IV U47495 ( .A(n34426), .Z(n34428) );
  NOR U47496 ( .A(n34428), .B(n34427), .Z(n44379) );
  IV U47497 ( .A(n44379), .Z(n34429) );
  NOR U47498 ( .A(n44348), .B(n34429), .Z(n44382) );
  IV U47499 ( .A(n44382), .Z(n34430) );
  NOR U47500 ( .A(n44386), .B(n34430), .Z(n44375) );
  IV U47501 ( .A(n44375), .Z(n34431) );
  NOR U47502 ( .A(n44346), .B(n34431), .Z(n44340) );
  IV U47503 ( .A(n44340), .Z(n37922) );
  IV U47504 ( .A(n44356), .Z(n34432) );
  NOR U47505 ( .A(n34433), .B(n34432), .Z(n34434) );
  IV U47506 ( .A(n34434), .Z(n44336) );
  IV U47507 ( .A(n34435), .Z(n34436) );
  NOR U47508 ( .A(n34437), .B(n34436), .Z(n37912) );
  IV U47509 ( .A(n37912), .Z(n37901) );
  IV U47510 ( .A(n34438), .Z(n34440) );
  NOR U47511 ( .A(n34440), .B(n34439), .Z(n37898) );
  IV U47512 ( .A(n37898), .Z(n37890) );
  IV U47513 ( .A(n34441), .Z(n34446) );
  IV U47514 ( .A(n34442), .Z(n34444) );
  XOR U47515 ( .A(n34450), .B(n34451), .Z(n34443) );
  NOR U47516 ( .A(n34444), .B(n34443), .Z(n34445) );
  IV U47517 ( .A(n34445), .Z(n37882) );
  NOR U47518 ( .A(n34446), .B(n37882), .Z(n41030) );
  IV U47519 ( .A(n34447), .Z(n34448) );
  NOR U47520 ( .A(n34449), .B(n34448), .Z(n37927) );
  IV U47521 ( .A(n34450), .Z(n34452) );
  NOR U47522 ( .A(n34452), .B(n34451), .Z(n41033) );
  NOR U47523 ( .A(n37927), .B(n41033), .Z(n34453) );
  IV U47524 ( .A(n34453), .Z(n37880) );
  IV U47525 ( .A(n34454), .Z(n34456) );
  IV U47526 ( .A(n34455), .Z(n37878) );
  NOR U47527 ( .A(n34456), .B(n37878), .Z(n37930) );
  IV U47528 ( .A(n34457), .Z(n34458) );
  NOR U47529 ( .A(n34459), .B(n34458), .Z(n41016) );
  IV U47530 ( .A(n34460), .Z(n34463) );
  IV U47531 ( .A(n34461), .Z(n34462) );
  NOR U47532 ( .A(n34463), .B(n34462), .Z(n41012) );
  NOR U47533 ( .A(n34464), .B(n34466), .Z(n41008) );
  IV U47534 ( .A(n34465), .Z(n34467) );
  NOR U47535 ( .A(n34467), .B(n34466), .Z(n41019) );
  NOR U47536 ( .A(n41008), .B(n41019), .Z(n37853) );
  IV U47537 ( .A(n34468), .Z(n34469) );
  NOR U47538 ( .A(n37826), .B(n34469), .Z(n37952) );
  IV U47539 ( .A(n34470), .Z(n34471) );
  NOR U47540 ( .A(n34471), .B(n37823), .Z(n37958) );
  IV U47541 ( .A(n34472), .Z(n34474) );
  NOR U47542 ( .A(n34474), .B(n34473), .Z(n37965) );
  IV U47543 ( .A(n34475), .Z(n34476) );
  NOR U47544 ( .A(n34477), .B(n34476), .Z(n44279) );
  IV U47545 ( .A(n34478), .Z(n34479) );
  NOR U47546 ( .A(n34480), .B(n34479), .Z(n44286) );
  NOR U47547 ( .A(n44279), .B(n44286), .Z(n37964) );
  IV U47548 ( .A(n37964), .Z(n37821) );
  IV U47549 ( .A(n34481), .Z(n34482) );
  NOR U47550 ( .A(n34483), .B(n34482), .Z(n40994) );
  IV U47551 ( .A(n34484), .Z(n37820) );
  IV U47552 ( .A(n34485), .Z(n34486) );
  NOR U47553 ( .A(n37820), .B(n34486), .Z(n40991) );
  IV U47554 ( .A(n34487), .Z(n34488) );
  NOR U47555 ( .A(n34488), .B(n34490), .Z(n40976) );
  IV U47556 ( .A(n34489), .Z(n34491) );
  NOR U47557 ( .A(n34491), .B(n34490), .Z(n37807) );
  IV U47558 ( .A(n34492), .Z(n34493) );
  NOR U47559 ( .A(n34494), .B(n34493), .Z(n40963) );
  NOR U47560 ( .A(n40960), .B(n40963), .Z(n37795) );
  IV U47561 ( .A(n34495), .Z(n34496) );
  NOR U47562 ( .A(n34496), .B(n37788), .Z(n40938) );
  IV U47563 ( .A(n34497), .Z(n34499) );
  NOR U47564 ( .A(n34499), .B(n34498), .Z(n40935) );
  IV U47565 ( .A(n34500), .Z(n34501) );
  NOR U47566 ( .A(n34501), .B(n37788), .Z(n37976) );
  NOR U47567 ( .A(n40935), .B(n37976), .Z(n34502) );
  IV U47568 ( .A(n34502), .Z(n37785) );
  IV U47569 ( .A(n34503), .Z(n34504) );
  NOR U47570 ( .A(n34505), .B(n34504), .Z(n40932) );
  IV U47571 ( .A(n34506), .Z(n34508) );
  NOR U47572 ( .A(n34508), .B(n34507), .Z(n40929) );
  IV U47573 ( .A(n34509), .Z(n34510) );
  NOR U47574 ( .A(n34510), .B(n34512), .Z(n37979) );
  IV U47575 ( .A(n34511), .Z(n34515) );
  NOR U47576 ( .A(n34513), .B(n34512), .Z(n34514) );
  IV U47577 ( .A(n34514), .Z(n37783) );
  NOR U47578 ( .A(n34515), .B(n37783), .Z(n37986) );
  IV U47579 ( .A(n34516), .Z(n34517) );
  NOR U47580 ( .A(n37997), .B(n34517), .Z(n34518) );
  IV U47581 ( .A(n34518), .Z(n40920) );
  IV U47582 ( .A(n34519), .Z(n37751) );
  IV U47583 ( .A(n34520), .Z(n34522) );
  NOR U47584 ( .A(n34522), .B(n34521), .Z(n38006) );
  IV U47585 ( .A(n34523), .Z(n34525) );
  NOR U47586 ( .A(n34525), .B(n34524), .Z(n40915) );
  NOR U47587 ( .A(n38006), .B(n40915), .Z(n34526) );
  IV U47588 ( .A(n34526), .Z(n37748) );
  IV U47589 ( .A(n34527), .Z(n34534) );
  NOR U47590 ( .A(n34529), .B(n34528), .Z(n34530) );
  IV U47591 ( .A(n34530), .Z(n34531) );
  NOR U47592 ( .A(n34532), .B(n34531), .Z(n34533) );
  IV U47593 ( .A(n34533), .Z(n37737) );
  NOR U47594 ( .A(n34534), .B(n37737), .Z(n37740) );
  IV U47595 ( .A(n37740), .Z(n47611) );
  IV U47596 ( .A(n34535), .Z(n34538) );
  NOR U47597 ( .A(n34536), .B(n37721), .Z(n34537) );
  IV U47598 ( .A(n34537), .Z(n37729) );
  NOR U47599 ( .A(n34538), .B(n37729), .Z(n34539) );
  IV U47600 ( .A(n34539), .Z(n38021) );
  IV U47601 ( .A(n34540), .Z(n34541) );
  NOR U47602 ( .A(n34542), .B(n34541), .Z(n38017) );
  NOR U47603 ( .A(n34544), .B(n34543), .Z(n38022) );
  IV U47604 ( .A(n34545), .Z(n40898) );
  IV U47605 ( .A(n34546), .Z(n34548) );
  NOR U47606 ( .A(n34548), .B(n34547), .Z(n38029) );
  IV U47607 ( .A(n34549), .Z(n34551) );
  NOR U47608 ( .A(n34551), .B(n34550), .Z(n44169) );
  IV U47609 ( .A(n34552), .Z(n34553) );
  NOR U47610 ( .A(n34553), .B(n37677), .Z(n41226) );
  NOR U47611 ( .A(n44169), .B(n41226), .Z(n38028) );
  IV U47612 ( .A(n38028), .Z(n37683) );
  IV U47613 ( .A(n34554), .Z(n34555) );
  NOR U47614 ( .A(n34556), .B(n34555), .Z(n40831) );
  IV U47615 ( .A(n34557), .Z(n34558) );
  NOR U47616 ( .A(n34558), .B(n34564), .Z(n40842) );
  NOR U47617 ( .A(n40831), .B(n40842), .Z(n40828) );
  IV U47618 ( .A(n34559), .Z(n34560) );
  NOR U47619 ( .A(n34571), .B(n34560), .Z(n34561) );
  IV U47620 ( .A(n34561), .Z(n34562) );
  NOR U47621 ( .A(n34562), .B(n34570), .Z(n44151) );
  IV U47622 ( .A(n34563), .Z(n34565) );
  NOR U47623 ( .A(n34565), .B(n34564), .Z(n44164) );
  NOR U47624 ( .A(n44151), .B(n44164), .Z(n40832) );
  IV U47625 ( .A(n34566), .Z(n34567) );
  NOR U47626 ( .A(n34568), .B(n34567), .Z(n38035) );
  IV U47627 ( .A(n34569), .Z(n34574) );
  NOR U47628 ( .A(n34571), .B(n34570), .Z(n34572) );
  IV U47629 ( .A(n34572), .Z(n34573) );
  NOR U47630 ( .A(n34574), .B(n34573), .Z(n38032) );
  NOR U47631 ( .A(n38035), .B(n38032), .Z(n37673) );
  IV U47632 ( .A(n34575), .Z(n34576) );
  NOR U47633 ( .A(n34577), .B(n34576), .Z(n40815) );
  IV U47634 ( .A(n34578), .Z(n34579) );
  NOR U47635 ( .A(n34580), .B(n34579), .Z(n40809) );
  IV U47636 ( .A(n34581), .Z(n34582) );
  NOR U47637 ( .A(n34583), .B(n34582), .Z(n40818) );
  NOR U47638 ( .A(n40809), .B(n40818), .Z(n37672) );
  IV U47639 ( .A(n34584), .Z(n34586) );
  XOR U47640 ( .A(n37662), .B(n37666), .Z(n34585) );
  NOR U47641 ( .A(n34586), .B(n34585), .Z(n40802) );
  IV U47642 ( .A(n34587), .Z(n37651) );
  IV U47643 ( .A(n34588), .Z(n34589) );
  NOR U47644 ( .A(n37651), .B(n34589), .Z(n41242) );
  IV U47645 ( .A(n41242), .Z(n44600) );
  IV U47646 ( .A(n34590), .Z(n34591) );
  NOR U47647 ( .A(n34592), .B(n34591), .Z(n34593) );
  IV U47648 ( .A(n34593), .Z(n37646) );
  IV U47649 ( .A(n34594), .Z(n34596) );
  NOR U47650 ( .A(n34596), .B(n34595), .Z(n40781) );
  IV U47651 ( .A(n34597), .Z(n34598) );
  NOR U47652 ( .A(n34604), .B(n34598), .Z(n40777) );
  IV U47653 ( .A(n34599), .Z(n34600) );
  NOR U47654 ( .A(n34601), .B(n34600), .Z(n40774) );
  IV U47655 ( .A(n34602), .Z(n34606) );
  NOR U47656 ( .A(n34604), .B(n34603), .Z(n34605) );
  IV U47657 ( .A(n34605), .Z(n34608) );
  NOR U47658 ( .A(n34606), .B(n34608), .Z(n40770) );
  IV U47659 ( .A(n34607), .Z(n34609) );
  NOR U47660 ( .A(n34609), .B(n34608), .Z(n40767) );
  IV U47661 ( .A(n34610), .Z(n34611) );
  NOR U47662 ( .A(n34612), .B(n34611), .Z(n40763) );
  IV U47663 ( .A(n34613), .Z(n34616) );
  IV U47664 ( .A(n34614), .Z(n34615) );
  NOR U47665 ( .A(n34616), .B(n34615), .Z(n40760) );
  IV U47666 ( .A(n34617), .Z(n34618) );
  NOR U47667 ( .A(n34618), .B(n38046), .Z(n38041) );
  IV U47668 ( .A(n34619), .Z(n34621) );
  NOR U47669 ( .A(n34621), .B(n34620), .Z(n38054) );
  IV U47670 ( .A(n34622), .Z(n34624) );
  NOR U47671 ( .A(n34624), .B(n34623), .Z(n38052) );
  NOR U47672 ( .A(n38054), .B(n38052), .Z(n37633) );
  IV U47673 ( .A(n34625), .Z(n34627) );
  NOR U47674 ( .A(n34627), .B(n34626), .Z(n37628) );
  IV U47675 ( .A(n34628), .Z(n34630) );
  NOR U47676 ( .A(n34630), .B(n34629), .Z(n40743) );
  IV U47677 ( .A(n34631), .Z(n34633) );
  NOR U47678 ( .A(n34633), .B(n34632), .Z(n38062) );
  NOR U47679 ( .A(n40743), .B(n38062), .Z(n37612) );
  IV U47680 ( .A(n34634), .Z(n34638) );
  NOR U47681 ( .A(n34636), .B(n34635), .Z(n34637) );
  IV U47682 ( .A(n34637), .Z(n34640) );
  NOR U47683 ( .A(n34638), .B(n34640), .Z(n40725) );
  IV U47684 ( .A(n34639), .Z(n34641) );
  NOR U47685 ( .A(n34641), .B(n34640), .Z(n40728) );
  IV U47686 ( .A(n34642), .Z(n34643) );
  NOR U47687 ( .A(n34644), .B(n34643), .Z(n40719) );
  IV U47688 ( .A(n34645), .Z(n34647) );
  NOR U47689 ( .A(n34647), .B(n34646), .Z(n40715) );
  NOR U47690 ( .A(n40719), .B(n40715), .Z(n38069) );
  IV U47691 ( .A(n34648), .Z(n34650) );
  NOR U47692 ( .A(n34650), .B(n34649), .Z(n38075) );
  IV U47693 ( .A(n34651), .Z(n34652) );
  NOR U47694 ( .A(n34653), .B(n34652), .Z(n38070) );
  NOR U47695 ( .A(n38075), .B(n38070), .Z(n37611) );
  IV U47696 ( .A(n34654), .Z(n34661) );
  NOR U47697 ( .A(n34656), .B(n34655), .Z(n34657) );
  IV U47698 ( .A(n34657), .Z(n34658) );
  NOR U47699 ( .A(n34659), .B(n34658), .Z(n34660) );
  IV U47700 ( .A(n34660), .Z(n34663) );
  NOR U47701 ( .A(n34661), .B(n34663), .Z(n38072) );
  IV U47702 ( .A(n34662), .Z(n34664) );
  NOR U47703 ( .A(n34664), .B(n34663), .Z(n38081) );
  IV U47704 ( .A(n34665), .Z(n34672) );
  NOR U47705 ( .A(n34667), .B(n34666), .Z(n34668) );
  IV U47706 ( .A(n34668), .Z(n34669) );
  NOR U47707 ( .A(n34670), .B(n34669), .Z(n34671) );
  IV U47708 ( .A(n34671), .Z(n34674) );
  NOR U47709 ( .A(n34672), .B(n34674), .Z(n38078) );
  IV U47710 ( .A(n34673), .Z(n34675) );
  NOR U47711 ( .A(n34675), .B(n34674), .Z(n38087) );
  IV U47712 ( .A(n34676), .Z(n34683) );
  NOR U47713 ( .A(n34678), .B(n34677), .Z(n34679) );
  IV U47714 ( .A(n34679), .Z(n34680) );
  NOR U47715 ( .A(n34681), .B(n34680), .Z(n34682) );
  IV U47716 ( .A(n34682), .Z(n37609) );
  NOR U47717 ( .A(n34683), .B(n37609), .Z(n38084) );
  NOR U47718 ( .A(n34684), .B(n38091), .Z(n37607) );
  IV U47719 ( .A(n34685), .Z(n34687) );
  NOR U47720 ( .A(n34687), .B(n34686), .Z(n34688) );
  IV U47721 ( .A(n34688), .Z(n37596) );
  IV U47722 ( .A(n34689), .Z(n34691) );
  NOR U47723 ( .A(n34691), .B(n34690), .Z(n34692) );
  IV U47724 ( .A(n34692), .Z(n37573) );
  IV U47725 ( .A(n34693), .Z(n51652) );
  IV U47726 ( .A(n51653), .Z(n34694) );
  NOR U47727 ( .A(n51652), .B(n34694), .Z(n40658) );
  NOR U47728 ( .A(n34696), .B(n34695), .Z(n40643) );
  IV U47729 ( .A(n34697), .Z(n34698) );
  NOR U47730 ( .A(n34698), .B(n34700), .Z(n40640) );
  IV U47731 ( .A(n34699), .Z(n34701) );
  NOR U47732 ( .A(n34701), .B(n34700), .Z(n38097) );
  IV U47733 ( .A(n34702), .Z(n37542) );
  IV U47734 ( .A(n34703), .Z(n34704) );
  NOR U47735 ( .A(n37542), .B(n34704), .Z(n41326) );
  IV U47736 ( .A(n34705), .Z(n34706) );
  NOR U47737 ( .A(n34706), .B(n37551), .Z(n41320) );
  NOR U47738 ( .A(n41326), .B(n41320), .Z(n38105) );
  IV U47739 ( .A(n34707), .Z(n34708) );
  NOR U47740 ( .A(n34709), .B(n34708), .Z(n38116) );
  IV U47741 ( .A(n34710), .Z(n34711) );
  NOR U47742 ( .A(n37544), .B(n34711), .Z(n38113) );
  NOR U47743 ( .A(n38116), .B(n38113), .Z(n37539) );
  IV U47744 ( .A(n34712), .Z(n34713) );
  NOR U47745 ( .A(n44015), .B(n34713), .Z(n34715) );
  IV U47746 ( .A(n44016), .Z(n34714) );
  NOR U47747 ( .A(n34714), .B(n44015), .Z(n44007) );
  NOR U47748 ( .A(n34715), .B(n44007), .Z(n38121) );
  IV U47749 ( .A(n34716), .Z(n34720) );
  IV U47750 ( .A(n34717), .Z(n34718) );
  NOR U47751 ( .A(n34720), .B(n34718), .Z(n38119) );
  IV U47752 ( .A(n34721), .Z(n34719) );
  NOR U47753 ( .A(n34719), .B(n34720), .Z(n43999) );
  XOR U47754 ( .A(n34721), .B(n34720), .Z(n34724) );
  IV U47755 ( .A(n34722), .Z(n34723) );
  NOR U47756 ( .A(n34724), .B(n34723), .Z(n44004) );
  NOR U47757 ( .A(n43999), .B(n44004), .Z(n38126) );
  IV U47758 ( .A(n38126), .Z(n37538) );
  IV U47759 ( .A(n34725), .Z(n34726) );
  NOR U47760 ( .A(n37536), .B(n34726), .Z(n38123) );
  IV U47761 ( .A(n34727), .Z(n34728) );
  NOR U47762 ( .A(n34731), .B(n34728), .Z(n40617) );
  IV U47763 ( .A(n34729), .Z(n34730) );
  NOR U47764 ( .A(n34731), .B(n34730), .Z(n40612) );
  IV U47765 ( .A(n34732), .Z(n34733) );
  NOR U47766 ( .A(n34734), .B(n34733), .Z(n40611) );
  IV U47767 ( .A(n34735), .Z(n34738) );
  NOR U47768 ( .A(n34750), .B(n34736), .Z(n34737) );
  IV U47769 ( .A(n34737), .Z(n34741) );
  NOR U47770 ( .A(n34738), .B(n34741), .Z(n41355) );
  NOR U47771 ( .A(n40611), .B(n41355), .Z(n34739) );
  IV U47772 ( .A(n34739), .Z(n37523) );
  IV U47773 ( .A(n34740), .Z(n34744) );
  NOR U47774 ( .A(n34742), .B(n34741), .Z(n34743) );
  IV U47775 ( .A(n34743), .Z(n34746) );
  NOR U47776 ( .A(n34744), .B(n34746), .Z(n38135) );
  IV U47777 ( .A(n34745), .Z(n34747) );
  NOR U47778 ( .A(n34747), .B(n34746), .Z(n38132) );
  IV U47779 ( .A(n34748), .Z(n34749) );
  NOR U47780 ( .A(n34750), .B(n34749), .Z(n40606) );
  IV U47781 ( .A(n34751), .Z(n34752) );
  NOR U47782 ( .A(n34752), .B(n37520), .Z(n40603) );
  IV U47783 ( .A(n34753), .Z(n37518) );
  IV U47784 ( .A(n34754), .Z(n34755) );
  NOR U47785 ( .A(n37518), .B(n34755), .Z(n34756) );
  IV U47786 ( .A(n34756), .Z(n38148) );
  IV U47787 ( .A(n34757), .Z(n34758) );
  NOR U47788 ( .A(n34759), .B(n34758), .Z(n34760) );
  IV U47789 ( .A(n34760), .Z(n38146) );
  IV U47790 ( .A(n34761), .Z(n34762) );
  NOR U47791 ( .A(n37514), .B(n34762), .Z(n37511) );
  IV U47792 ( .A(n37511), .Z(n37504) );
  IV U47793 ( .A(n34763), .Z(n34766) );
  NOR U47794 ( .A(n34764), .B(n34770), .Z(n34765) );
  IV U47795 ( .A(n34765), .Z(n34768) );
  NOR U47796 ( .A(n34766), .B(n34768), .Z(n38153) );
  IV U47797 ( .A(n34767), .Z(n34769) );
  NOR U47798 ( .A(n34769), .B(n34768), .Z(n38158) );
  NOR U47799 ( .A(n34771), .B(n34770), .Z(n34772) );
  IV U47800 ( .A(n34772), .Z(n34773) );
  NOR U47801 ( .A(n34774), .B(n34773), .Z(n40596) );
  IV U47802 ( .A(n34775), .Z(n34776) );
  NOR U47803 ( .A(n34776), .B(n34782), .Z(n34777) );
  IV U47804 ( .A(n34777), .Z(n40576) );
  IV U47805 ( .A(n34778), .Z(n34779) );
  NOR U47806 ( .A(n34780), .B(n34779), .Z(n40579) );
  IV U47807 ( .A(n34781), .Z(n34783) );
  NOR U47808 ( .A(n34783), .B(n34782), .Z(n40571) );
  NOR U47809 ( .A(n40579), .B(n40571), .Z(n37491) );
  IV U47810 ( .A(n34784), .Z(n34791) );
  NOR U47811 ( .A(n34786), .B(n34785), .Z(n34787) );
  IV U47812 ( .A(n34787), .Z(n34788) );
  NOR U47813 ( .A(n34789), .B(n34788), .Z(n34790) );
  IV U47814 ( .A(n34790), .Z(n37483) );
  NOR U47815 ( .A(n34791), .B(n37483), .Z(n38161) );
  IV U47816 ( .A(n34792), .Z(n34794) );
  NOR U47817 ( .A(n34794), .B(n34793), .Z(n38170) );
  IV U47818 ( .A(n34795), .Z(n34797) );
  NOR U47819 ( .A(n34797), .B(n34796), .Z(n38165) );
  NOR U47820 ( .A(n38170), .B(n38165), .Z(n34798) );
  IV U47821 ( .A(n34798), .Z(n37481) );
  IV U47822 ( .A(n34799), .Z(n34800) );
  NOR U47823 ( .A(n34801), .B(n34800), .Z(n38168) );
  IV U47824 ( .A(n34802), .Z(n34803) );
  NOR U47825 ( .A(n34803), .B(n37476), .Z(n38176) );
  IV U47826 ( .A(n34804), .Z(n37480) );
  IV U47827 ( .A(n34805), .Z(n34806) );
  NOR U47828 ( .A(n37480), .B(n34806), .Z(n34807) );
  IV U47829 ( .A(n34807), .Z(n38183) );
  IV U47830 ( .A(n34808), .Z(n34809) );
  NOR U47831 ( .A(n34809), .B(n37473), .Z(n38179) );
  IV U47832 ( .A(n34810), .Z(n34814) );
  NOR U47833 ( .A(n34812), .B(n34811), .Z(n34813) );
  IV U47834 ( .A(n34813), .Z(n37470) );
  NOR U47835 ( .A(n34814), .B(n37470), .Z(n40554) );
  IV U47836 ( .A(n34815), .Z(n34816) );
  NOR U47837 ( .A(n34817), .B(n34816), .Z(n40550) );
  IV U47838 ( .A(n34818), .Z(n37463) );
  IV U47839 ( .A(n34819), .Z(n34820) );
  NOR U47840 ( .A(n37463), .B(n34820), .Z(n40540) );
  NOR U47841 ( .A(n40550), .B(n40540), .Z(n34821) );
  IV U47842 ( .A(n34821), .Z(n37468) );
  IV U47843 ( .A(n34822), .Z(n34823) );
  NOR U47844 ( .A(n34823), .B(n37463), .Z(n34824) );
  IV U47845 ( .A(n34824), .Z(n34825) );
  NOR U47846 ( .A(n34826), .B(n34825), .Z(n40544) );
  IV U47847 ( .A(n34827), .Z(n34828) );
  NOR U47848 ( .A(n34828), .B(n34832), .Z(n34829) );
  IV U47849 ( .A(n34829), .Z(n41442) );
  IV U47850 ( .A(n34830), .Z(n34831) );
  NOR U47851 ( .A(n34832), .B(n34831), .Z(n34833) );
  IV U47852 ( .A(n34833), .Z(n40536) );
  IV U47853 ( .A(n34834), .Z(n34835) );
  NOR U47854 ( .A(n34836), .B(n34835), .Z(n40520) );
  IV U47855 ( .A(n34837), .Z(n34839) );
  NOR U47856 ( .A(n34839), .B(n34838), .Z(n41487) );
  IV U47857 ( .A(n34840), .Z(n34842) );
  NOR U47858 ( .A(n34842), .B(n34841), .Z(n43909) );
  NOR U47859 ( .A(n41487), .B(n43909), .Z(n40487) );
  IV U47860 ( .A(n34843), .Z(n34848) );
  IV U47861 ( .A(n34844), .Z(n34845) );
  NOR U47862 ( .A(n34848), .B(n34845), .Z(n40479) );
  IV U47863 ( .A(n34846), .Z(n34847) );
  NOR U47864 ( .A(n34848), .B(n34847), .Z(n41495) );
  IV U47865 ( .A(n34849), .Z(n34851) );
  NOR U47866 ( .A(n34851), .B(n34850), .Z(n41503) );
  NOR U47867 ( .A(n41495), .B(n41503), .Z(n40478) );
  IV U47868 ( .A(n40478), .Z(n37395) );
  IV U47869 ( .A(n34852), .Z(n34854) );
  NOR U47870 ( .A(n34854), .B(n34853), .Z(n34855) );
  IV U47871 ( .A(n34855), .Z(n38216) );
  IV U47872 ( .A(n34856), .Z(n34862) );
  NOR U47873 ( .A(n34857), .B(n37374), .Z(n34858) );
  IV U47874 ( .A(n34858), .Z(n34859) );
  NOR U47875 ( .A(n34860), .B(n34859), .Z(n34861) );
  IV U47876 ( .A(n34861), .Z(n37381) );
  NOR U47877 ( .A(n34862), .B(n37381), .Z(n38226) );
  NOR U47878 ( .A(n38220), .B(n38226), .Z(n37385) );
  IV U47879 ( .A(n34863), .Z(n37380) );
  IV U47880 ( .A(n34864), .Z(n34872) );
  IV U47881 ( .A(n34865), .Z(n34866) );
  NOR U47882 ( .A(n34872), .B(n34866), .Z(n38230) );
  IV U47883 ( .A(n34867), .Z(n34869) );
  NOR U47884 ( .A(n34869), .B(n34868), .Z(n40469) );
  IV U47885 ( .A(n34870), .Z(n34871) );
  NOR U47886 ( .A(n34872), .B(n34871), .Z(n38233) );
  NOR U47887 ( .A(n40469), .B(n38233), .Z(n34873) );
  IV U47888 ( .A(n34873), .Z(n37364) );
  IV U47889 ( .A(n34874), .Z(n34875) );
  NOR U47890 ( .A(n34875), .B(n37360), .Z(n40464) );
  IV U47891 ( .A(n34876), .Z(n37363) );
  IV U47892 ( .A(n34877), .Z(n34878) );
  NOR U47893 ( .A(n37363), .B(n34878), .Z(n38236) );
  IV U47894 ( .A(n34879), .Z(n34880) );
  NOR U47895 ( .A(n34880), .B(n34886), .Z(n40457) );
  IV U47896 ( .A(n34881), .Z(n34883) );
  NOR U47897 ( .A(n34883), .B(n34882), .Z(n40458) );
  XOR U47898 ( .A(n40457), .B(n40458), .Z(n34884) );
  NOR U47899 ( .A(n38236), .B(n34884), .Z(n37357) );
  IV U47900 ( .A(n34885), .Z(n34887) );
  NOR U47901 ( .A(n34887), .B(n34886), .Z(n40451) );
  IV U47902 ( .A(n34888), .Z(n34890) );
  IV U47903 ( .A(n34889), .Z(n34894) );
  NOR U47904 ( .A(n34890), .B(n34894), .Z(n40448) );
  IV U47905 ( .A(n34891), .Z(n34892) );
  NOR U47906 ( .A(n34892), .B(n34900), .Z(n40443) );
  IV U47907 ( .A(n34893), .Z(n34895) );
  NOR U47908 ( .A(n34895), .B(n34894), .Z(n40445) );
  NOR U47909 ( .A(n40443), .B(n40445), .Z(n37356) );
  IV U47910 ( .A(n34896), .Z(n34898) );
  NOR U47911 ( .A(n34898), .B(n34897), .Z(n38239) );
  IV U47912 ( .A(n34899), .Z(n34901) );
  NOR U47913 ( .A(n34901), .B(n34900), .Z(n40439) );
  NOR U47914 ( .A(n38239), .B(n40439), .Z(n37355) );
  IV U47915 ( .A(n34902), .Z(n34903) );
  NOR U47916 ( .A(n34904), .B(n34903), .Z(n38244) );
  IV U47917 ( .A(n34905), .Z(n34907) );
  NOR U47918 ( .A(n34907), .B(n34906), .Z(n38241) );
  IV U47919 ( .A(n34908), .Z(n34914) );
  IV U47920 ( .A(n34909), .Z(n34910) );
  NOR U47921 ( .A(n34914), .B(n34910), .Z(n34911) );
  IV U47922 ( .A(n34911), .Z(n40429) );
  IV U47923 ( .A(n34912), .Z(n34913) );
  NOR U47924 ( .A(n34914), .B(n34913), .Z(n38248) );
  IV U47925 ( .A(n34915), .Z(n34916) );
  NOR U47926 ( .A(n34917), .B(n34916), .Z(n38262) );
  NOR U47927 ( .A(n34918), .B(n38252), .Z(n34919) );
  NOR U47928 ( .A(n38262), .B(n34919), .Z(n34920) );
  IV U47929 ( .A(n34920), .Z(n37347) );
  IV U47930 ( .A(n34921), .Z(n34923) );
  NOR U47931 ( .A(n34923), .B(n34922), .Z(n38259) );
  IV U47932 ( .A(n34924), .Z(n34927) );
  IV U47933 ( .A(n34925), .Z(n37345) );
  XOR U47934 ( .A(n37342), .B(n37345), .Z(n34926) );
  NOR U47935 ( .A(n34927), .B(n34926), .Z(n38267) );
  IV U47936 ( .A(n34928), .Z(n34929) );
  NOR U47937 ( .A(n34929), .B(n34936), .Z(n34930) );
  IV U47938 ( .A(n34930), .Z(n38272) );
  IV U47939 ( .A(n34931), .Z(n34933) );
  NOR U47940 ( .A(n34933), .B(n34932), .Z(n38275) );
  IV U47941 ( .A(n34934), .Z(n34935) );
  NOR U47942 ( .A(n34936), .B(n34935), .Z(n40416) );
  NOR U47943 ( .A(n38275), .B(n40416), .Z(n34937) );
  IV U47944 ( .A(n34937), .Z(n37341) );
  IV U47945 ( .A(n34938), .Z(n34940) );
  NOR U47946 ( .A(n34940), .B(n34939), .Z(n41560) );
  IV U47947 ( .A(n34941), .Z(n34943) );
  NOR U47948 ( .A(n34943), .B(n34942), .Z(n41556) );
  NOR U47949 ( .A(n41560), .B(n41556), .Z(n38281) );
  IV U47950 ( .A(n34944), .Z(n34945) );
  NOR U47951 ( .A(n34946), .B(n34945), .Z(n38278) );
  IV U47952 ( .A(n34947), .Z(n34952) );
  IV U47953 ( .A(n34948), .Z(n34949) );
  NOR U47954 ( .A(n34952), .B(n34949), .Z(n38287) );
  IV U47955 ( .A(n34950), .Z(n34951) );
  NOR U47956 ( .A(n34952), .B(n34951), .Z(n38284) );
  IV U47957 ( .A(n34953), .Z(n34954) );
  NOR U47958 ( .A(n34955), .B(n34954), .Z(n43801) );
  IV U47959 ( .A(n34956), .Z(n34958) );
  NOR U47960 ( .A(n34958), .B(n34957), .Z(n43810) );
  NOR U47961 ( .A(n43801), .B(n43810), .Z(n40404) );
  NOR U47962 ( .A(n34959), .B(n34964), .Z(n34960) );
  IV U47963 ( .A(n34960), .Z(n34961) );
  NOR U47964 ( .A(n34962), .B(n34961), .Z(n40401) );
  IV U47965 ( .A(n34963), .Z(n34965) );
  NOR U47966 ( .A(n34965), .B(n34964), .Z(n38299) );
  IV U47967 ( .A(n34966), .Z(n34973) );
  NOR U47968 ( .A(n34968), .B(n34967), .Z(n34969) );
  IV U47969 ( .A(n34969), .Z(n34970) );
  NOR U47970 ( .A(n34971), .B(n34970), .Z(n34972) );
  IV U47971 ( .A(n34972), .Z(n37324) );
  NOR U47972 ( .A(n34973), .B(n37324), .Z(n38296) );
  IV U47973 ( .A(n34974), .Z(n34981) );
  NOR U47974 ( .A(n34976), .B(n34975), .Z(n34977) );
  IV U47975 ( .A(n34977), .Z(n34978) );
  NOR U47976 ( .A(n34979), .B(n34978), .Z(n34980) );
  IV U47977 ( .A(n34980), .Z(n37309) );
  NOR U47978 ( .A(n34981), .B(n37309), .Z(n38307) );
  IV U47979 ( .A(n34982), .Z(n34985) );
  IV U47980 ( .A(n34983), .Z(n34984) );
  NOR U47981 ( .A(n34985), .B(n34984), .Z(n40392) );
  NOR U47982 ( .A(n34987), .B(n34986), .Z(n41592) );
  NOR U47983 ( .A(n41592), .B(n41588), .Z(n38316) );
  IV U47984 ( .A(n38316), .Z(n37307) );
  IV U47985 ( .A(n34988), .Z(n34995) );
  NOR U47986 ( .A(n34990), .B(n34989), .Z(n34991) );
  IV U47987 ( .A(n34991), .Z(n34992) );
  NOR U47988 ( .A(n34993), .B(n34992), .Z(n34994) );
  IV U47989 ( .A(n34994), .Z(n34997) );
  NOR U47990 ( .A(n34995), .B(n34997), .Z(n38313) );
  IV U47991 ( .A(n34996), .Z(n34998) );
  NOR U47992 ( .A(n34998), .B(n34997), .Z(n38321) );
  IV U47993 ( .A(n34999), .Z(n35004) );
  IV U47994 ( .A(n35000), .Z(n35001) );
  NOR U47995 ( .A(n35004), .B(n35001), .Z(n38318) );
  IV U47996 ( .A(n35002), .Z(n35003) );
  NOR U47997 ( .A(n35004), .B(n35003), .Z(n38327) );
  IV U47998 ( .A(n35005), .Z(n35006) );
  NOR U47999 ( .A(n35006), .B(n37306), .Z(n38324) );
  IV U48000 ( .A(n35007), .Z(n35009) );
  NOR U48001 ( .A(n35009), .B(n35008), .Z(n35010) );
  IV U48002 ( .A(n35010), .Z(n38331) );
  IV U48003 ( .A(n35011), .Z(n35012) );
  NOR U48004 ( .A(n35013), .B(n35012), .Z(n38335) );
  IV U48005 ( .A(n35014), .Z(n35018) );
  NOR U48006 ( .A(n35016), .B(n35015), .Z(n35017) );
  IV U48007 ( .A(n35017), .Z(n37299) );
  NOR U48008 ( .A(n35018), .B(n37299), .Z(n40381) );
  NOR U48009 ( .A(n38335), .B(n40381), .Z(n37296) );
  IV U48010 ( .A(n35019), .Z(n35023) );
  IV U48011 ( .A(n35020), .Z(n35021) );
  NOR U48012 ( .A(n35023), .B(n35021), .Z(n38338) );
  IV U48013 ( .A(n35022), .Z(n35024) );
  NOR U48014 ( .A(n35024), .B(n35023), .Z(n40370) );
  NOR U48015 ( .A(n35026), .B(n35025), .Z(n40364) );
  NOR U48016 ( .A(n35027), .B(n35030), .Z(n35028) );
  IV U48017 ( .A(n35028), .Z(n37267) );
  NOR U48018 ( .A(n35029), .B(n37267), .Z(n40339) );
  NOR U48019 ( .A(n35031), .B(n35030), .Z(n37262) );
  IV U48020 ( .A(n35032), .Z(n35033) );
  NOR U48021 ( .A(n35036), .B(n35033), .Z(n38360) );
  IV U48022 ( .A(n35034), .Z(n35035) );
  NOR U48023 ( .A(n35036), .B(n35035), .Z(n38371) );
  IV U48024 ( .A(n35037), .Z(n35039) );
  IV U48025 ( .A(n35038), .Z(n35041) );
  NOR U48026 ( .A(n35039), .B(n35041), .Z(n38368) );
  IV U48027 ( .A(n35040), .Z(n35042) );
  NOR U48028 ( .A(n35042), .B(n35041), .Z(n40318) );
  IV U48029 ( .A(n35043), .Z(n35045) );
  NOR U48030 ( .A(n35045), .B(n35044), .Z(n40321) );
  NOR U48031 ( .A(n35047), .B(n35046), .Z(n38374) );
  NOR U48032 ( .A(n40321), .B(n38374), .Z(n37253) );
  IV U48033 ( .A(n35048), .Z(n35050) );
  IV U48034 ( .A(n35049), .Z(n35058) );
  NOR U48035 ( .A(n35050), .B(n35058), .Z(n40310) );
  IV U48036 ( .A(n35051), .Z(n35053) );
  NOR U48037 ( .A(n35053), .B(n35052), .Z(n40306) );
  NOR U48038 ( .A(n40310), .B(n40306), .Z(n37245) );
  NOR U48039 ( .A(n35055), .B(n35054), .Z(n40297) );
  IV U48040 ( .A(n35056), .Z(n35057) );
  NOR U48041 ( .A(n35058), .B(n35057), .Z(n40302) );
  NOR U48042 ( .A(n40297), .B(n40302), .Z(n37244) );
  IV U48043 ( .A(n35059), .Z(n35060) );
  NOR U48044 ( .A(n35062), .B(n35060), .Z(n40294) );
  IV U48045 ( .A(n35061), .Z(n35063) );
  NOR U48046 ( .A(n35063), .B(n35062), .Z(n38379) );
  IV U48047 ( .A(n35064), .Z(n35068) );
  NOR U48048 ( .A(n35066), .B(n35065), .Z(n35067) );
  IV U48049 ( .A(n35067), .Z(n37238) );
  NOR U48050 ( .A(n35068), .B(n37238), .Z(n38376) );
  IV U48051 ( .A(n35069), .Z(n37242) );
  IV U48052 ( .A(n35070), .Z(n35071) );
  NOR U48053 ( .A(n37242), .B(n35071), .Z(n35072) );
  IV U48054 ( .A(n35072), .Z(n40288) );
  IV U48055 ( .A(n35073), .Z(n35077) );
  NOR U48056 ( .A(n35075), .B(n35074), .Z(n35076) );
  IV U48057 ( .A(n35076), .Z(n37236) );
  NOR U48058 ( .A(n35077), .B(n37236), .Z(n38389) );
  IV U48059 ( .A(n35078), .Z(n35080) );
  NOR U48060 ( .A(n35080), .B(n35079), .Z(n38394) );
  NOR U48061 ( .A(n38389), .B(n38394), .Z(n37233) );
  IV U48062 ( .A(n35081), .Z(n35087) );
  NOR U48063 ( .A(n35097), .B(n35082), .Z(n35083) );
  IV U48064 ( .A(n35083), .Z(n35084) );
  NOR U48065 ( .A(n35085), .B(n35084), .Z(n35086) );
  IV U48066 ( .A(n35086), .Z(n35089) );
  NOR U48067 ( .A(n35087), .B(n35089), .Z(n38391) );
  IV U48068 ( .A(n35088), .Z(n35090) );
  NOR U48069 ( .A(n35090), .B(n35089), .Z(n40277) );
  NOR U48070 ( .A(n35092), .B(n35091), .Z(n35093) );
  IV U48071 ( .A(n35093), .Z(n40269) );
  NOR U48072 ( .A(n35094), .B(n40269), .Z(n40280) );
  IV U48073 ( .A(n35095), .Z(n35096) );
  NOR U48074 ( .A(n35097), .B(n35096), .Z(n40273) );
  IV U48075 ( .A(n35098), .Z(n35100) );
  IV U48076 ( .A(n35099), .Z(n35103) );
  NOR U48077 ( .A(n35100), .B(n35103), .Z(n38397) );
  NOR U48078 ( .A(n40273), .B(n38397), .Z(n37231) );
  NOR U48079 ( .A(n35101), .B(n38404), .Z(n35105) );
  IV U48080 ( .A(n35102), .Z(n35104) );
  NOR U48081 ( .A(n35104), .B(n35103), .Z(n38400) );
  NOR U48082 ( .A(n35105), .B(n38400), .Z(n37230) );
  IV U48083 ( .A(n35106), .Z(n35108) );
  NOR U48084 ( .A(n35108), .B(n35107), .Z(n40257) );
  IV U48085 ( .A(n35109), .Z(n35111) );
  NOR U48086 ( .A(n35111), .B(n35110), .Z(n40254) );
  IV U48087 ( .A(n35112), .Z(n35113) );
  NOR U48088 ( .A(n35114), .B(n35113), .Z(n40260) );
  NOR U48089 ( .A(n40254), .B(n40260), .Z(n35115) );
  IV U48090 ( .A(n35115), .Z(n37223) );
  IV U48091 ( .A(n35116), .Z(n35122) );
  NOR U48092 ( .A(n35117), .B(n37217), .Z(n35118) );
  IV U48093 ( .A(n35118), .Z(n35119) );
  NOR U48094 ( .A(n35120), .B(n35119), .Z(n35121) );
  IV U48095 ( .A(n35121), .Z(n37221) );
  NOR U48096 ( .A(n35122), .B(n37221), .Z(n40251) );
  IV U48097 ( .A(n35123), .Z(n35125) );
  NOR U48098 ( .A(n35125), .B(n35124), .Z(n35126) );
  IV U48099 ( .A(n35126), .Z(n37209) );
  IV U48100 ( .A(n35127), .Z(n35128) );
  NOR U48101 ( .A(n35129), .B(n35128), .Z(n38420) );
  IV U48102 ( .A(n35130), .Z(n35134) );
  NOR U48103 ( .A(n35132), .B(n35131), .Z(n35133) );
  IV U48104 ( .A(n35133), .Z(n35136) );
  NOR U48105 ( .A(n35134), .B(n35136), .Z(n38428) );
  NOR U48106 ( .A(n38420), .B(n38428), .Z(n37194) );
  IV U48107 ( .A(n35135), .Z(n35137) );
  NOR U48108 ( .A(n35137), .B(n35136), .Z(n38425) );
  IV U48109 ( .A(n35138), .Z(n35142) );
  NOR U48110 ( .A(n35140), .B(n35139), .Z(n35141) );
  IV U48111 ( .A(n35141), .Z(n37192) );
  NOR U48112 ( .A(n35142), .B(n37192), .Z(n40230) );
  IV U48113 ( .A(n35143), .Z(n35144) );
  NOR U48114 ( .A(n35145), .B(n35144), .Z(n43684) );
  IV U48115 ( .A(n35146), .Z(n35147) );
  NOR U48116 ( .A(n35147), .B(n35150), .Z(n43675) );
  NOR U48117 ( .A(n43684), .B(n43675), .Z(n40223) );
  IV U48118 ( .A(n35148), .Z(n35149) );
  NOR U48119 ( .A(n35150), .B(n35149), .Z(n40220) );
  NOR U48120 ( .A(n35151), .B(n37181), .Z(n35152) );
  IV U48121 ( .A(n35152), .Z(n35153) );
  NOR U48122 ( .A(n35154), .B(n35153), .Z(n35155) );
  IV U48123 ( .A(n35155), .Z(n40205) );
  IV U48124 ( .A(n35156), .Z(n35158) );
  NOR U48125 ( .A(n35158), .B(n35157), .Z(n38444) );
  IV U48126 ( .A(n35159), .Z(n35160) );
  NOR U48127 ( .A(n35160), .B(n37175), .Z(n43652) );
  IV U48128 ( .A(n35161), .Z(n35162) );
  NOR U48129 ( .A(n35163), .B(n35162), .Z(n43658) );
  NOR U48130 ( .A(n43652), .B(n43658), .Z(n40207) );
  IV U48131 ( .A(n35164), .Z(n35166) );
  NOR U48132 ( .A(n35166), .B(n35165), .Z(n40200) );
  IV U48133 ( .A(n35167), .Z(n35169) );
  NOR U48134 ( .A(n35169), .B(n35168), .Z(n38453) );
  NOR U48135 ( .A(n40200), .B(n38453), .Z(n37170) );
  IV U48136 ( .A(n35170), .Z(n37157) );
  IV U48137 ( .A(n35171), .Z(n35173) );
  NOR U48138 ( .A(n35173), .B(n35172), .Z(n35174) );
  IV U48139 ( .A(n35174), .Z(n38462) );
  IV U48140 ( .A(n35175), .Z(n35176) );
  NOR U48141 ( .A(n35176), .B(n37132), .Z(n35177) );
  IV U48142 ( .A(n35177), .Z(n37134) );
  IV U48143 ( .A(n35178), .Z(n37130) );
  IV U48144 ( .A(n35179), .Z(n35180) );
  NOR U48145 ( .A(n37130), .B(n35180), .Z(n38474) );
  IV U48146 ( .A(n35181), .Z(n35183) );
  NOR U48147 ( .A(n35183), .B(n35182), .Z(n38472) );
  IV U48148 ( .A(n35184), .Z(n35187) );
  NOR U48149 ( .A(n35185), .B(n35189), .Z(n35186) );
  IV U48150 ( .A(n35186), .Z(n35192) );
  NOR U48151 ( .A(n35187), .B(n35192), .Z(n40184) );
  NOR U48152 ( .A(n38472), .B(n40184), .Z(n37127) );
  IV U48153 ( .A(n35188), .Z(n35190) );
  NOR U48154 ( .A(n35190), .B(n35189), .Z(n38480) );
  IV U48155 ( .A(n35191), .Z(n35193) );
  NOR U48156 ( .A(n35193), .B(n35192), .Z(n40187) );
  NOR U48157 ( .A(n38480), .B(n40187), .Z(n37126) );
  IV U48158 ( .A(n35194), .Z(n35196) );
  NOR U48159 ( .A(n35196), .B(n35195), .Z(n38490) );
  IV U48160 ( .A(n35197), .Z(n35199) );
  NOR U48161 ( .A(n35199), .B(n35198), .Z(n38482) );
  NOR U48162 ( .A(n38490), .B(n38482), .Z(n37118) );
  IV U48163 ( .A(n35200), .Z(n35201) );
  NOR U48164 ( .A(n35201), .B(n37115), .Z(n38487) );
  IV U48165 ( .A(n35202), .Z(n35204) );
  NOR U48166 ( .A(n35204), .B(n35203), .Z(n37094) );
  IV U48167 ( .A(n37094), .Z(n37089) );
  IV U48168 ( .A(n35205), .Z(n35207) );
  IV U48169 ( .A(n35206), .Z(n35211) );
  NOR U48170 ( .A(n35207), .B(n35211), .Z(n40176) );
  IV U48171 ( .A(n35208), .Z(n35209) );
  NOR U48172 ( .A(n35209), .B(n37081), .Z(n38500) );
  IV U48173 ( .A(n35210), .Z(n35212) );
  NOR U48174 ( .A(n35212), .B(n35211), .Z(n40173) );
  NOR U48175 ( .A(n38500), .B(n40173), .Z(n37087) );
  IV U48176 ( .A(n35213), .Z(n37085) );
  IV U48177 ( .A(n35214), .Z(n35215) );
  NOR U48178 ( .A(n37085), .B(n35215), .Z(n38507) );
  IV U48179 ( .A(n35216), .Z(n35218) );
  NOR U48180 ( .A(n35218), .B(n35217), .Z(n38504) );
  IV U48181 ( .A(n35219), .Z(n35220) );
  NOR U48182 ( .A(n35220), .B(n35222), .Z(n38512) );
  IV U48183 ( .A(n35221), .Z(n35223) );
  NOR U48184 ( .A(n35223), .B(n35222), .Z(n38514) );
  NOR U48185 ( .A(n35225), .B(n35224), .Z(n35226) );
  IV U48186 ( .A(n35226), .Z(n38521) );
  NOR U48187 ( .A(n35227), .B(n38521), .Z(n38516) );
  NOR U48188 ( .A(n38514), .B(n38516), .Z(n35228) );
  IV U48189 ( .A(n35228), .Z(n35229) );
  NOR U48190 ( .A(n38512), .B(n35229), .Z(n37079) );
  IV U48191 ( .A(n35230), .Z(n35232) );
  NOR U48192 ( .A(n35232), .B(n35231), .Z(n38529) );
  IV U48193 ( .A(n35233), .Z(n35235) );
  NOR U48194 ( .A(n35235), .B(n35234), .Z(n38526) );
  NOR U48195 ( .A(n38529), .B(n38526), .Z(n37078) );
  IV U48196 ( .A(n35236), .Z(n35237) );
  NOR U48197 ( .A(n35238), .B(n35237), .Z(n40162) );
  NOR U48198 ( .A(n35240), .B(n35239), .Z(n38531) );
  IV U48199 ( .A(n35241), .Z(n35242) );
  NOR U48200 ( .A(n35242), .B(n35244), .Z(n40157) );
  NOR U48201 ( .A(n38531), .B(n40157), .Z(n37069) );
  IV U48202 ( .A(n35243), .Z(n35247) );
  NOR U48203 ( .A(n35245), .B(n35244), .Z(n35246) );
  IV U48204 ( .A(n35246), .Z(n35249) );
  NOR U48205 ( .A(n35247), .B(n35249), .Z(n40147) );
  IV U48206 ( .A(n35248), .Z(n35250) );
  NOR U48207 ( .A(n35250), .B(n35249), .Z(n38536) );
  IV U48208 ( .A(n35251), .Z(n35252) );
  NOR U48209 ( .A(n35252), .B(n35254), .Z(n41835) );
  IV U48210 ( .A(n35253), .Z(n35258) );
  NOR U48211 ( .A(n35255), .B(n35254), .Z(n35256) );
  IV U48212 ( .A(n35256), .Z(n35257) );
  NOR U48213 ( .A(n35258), .B(n35257), .Z(n41827) );
  NOR U48214 ( .A(n41835), .B(n41827), .Z(n40151) );
  IV U48215 ( .A(n35259), .Z(n35260) );
  NOR U48216 ( .A(n35261), .B(n35260), .Z(n43576) );
  IV U48217 ( .A(n35262), .Z(n35264) );
  IV U48218 ( .A(n35263), .Z(n35268) );
  NOR U48219 ( .A(n35264), .B(n35268), .Z(n43570) );
  NOR U48220 ( .A(n43576), .B(n43570), .Z(n38553) );
  IV U48221 ( .A(n35265), .Z(n35266) );
  NOR U48222 ( .A(n35266), .B(n35274), .Z(n43562) );
  IV U48223 ( .A(n35267), .Z(n35269) );
  NOR U48224 ( .A(n35269), .B(n35268), .Z(n43567) );
  NOR U48225 ( .A(n43562), .B(n43567), .Z(n38559) );
  IV U48226 ( .A(n35270), .Z(n35272) );
  NOR U48227 ( .A(n35272), .B(n35271), .Z(n43554) );
  IV U48228 ( .A(n35273), .Z(n35275) );
  NOR U48229 ( .A(n35275), .B(n35274), .Z(n43559) );
  NOR U48230 ( .A(n43554), .B(n43559), .Z(n38563) );
  NOR U48231 ( .A(n35277), .B(n35276), .Z(n35278) );
  IV U48232 ( .A(n35278), .Z(n37048) );
  IV U48233 ( .A(n35279), .Z(n35282) );
  NOR U48234 ( .A(n35280), .B(n37045), .Z(n35281) );
  IV U48235 ( .A(n35281), .Z(n37039) );
  NOR U48236 ( .A(n35282), .B(n37039), .Z(n38572) );
  IV U48237 ( .A(n35283), .Z(n35285) );
  IV U48238 ( .A(n35284), .Z(n37016) );
  NOR U48239 ( .A(n35285), .B(n37016), .Z(n38604) );
  NOR U48240 ( .A(n35287), .B(n35286), .Z(n38601) );
  IV U48241 ( .A(n35288), .Z(n35290) );
  NOR U48242 ( .A(n35290), .B(n35289), .Z(n43515) );
  NOR U48243 ( .A(n43515), .B(n41876), .Z(n38607) );
  IV U48244 ( .A(n38607), .Z(n37014) );
  IV U48245 ( .A(n35291), .Z(n35296) );
  IV U48246 ( .A(n35292), .Z(n35293) );
  NOR U48247 ( .A(n35296), .B(n35293), .Z(n38611) );
  IV U48248 ( .A(n35294), .Z(n35295) );
  NOR U48249 ( .A(n35296), .B(n35295), .Z(n38608) );
  IV U48250 ( .A(n35297), .Z(n35299) );
  IV U48251 ( .A(n35298), .Z(n35302) );
  NOR U48252 ( .A(n35299), .B(n35302), .Z(n35300) );
  IV U48253 ( .A(n35300), .Z(n40115) );
  IV U48254 ( .A(n35301), .Z(n35303) );
  NOR U48255 ( .A(n35303), .B(n35302), .Z(n40111) );
  IV U48256 ( .A(n35304), .Z(n35305) );
  NOR U48257 ( .A(n35306), .B(n35305), .Z(n40091) );
  NOR U48258 ( .A(n35307), .B(n40096), .Z(n35308) );
  NOR U48259 ( .A(n40091), .B(n35308), .Z(n35309) );
  IV U48260 ( .A(n35309), .Z(n37000) );
  IV U48261 ( .A(n35310), .Z(n35312) );
  IV U48262 ( .A(n36999), .Z(n35311) );
  NOR U48263 ( .A(n35312), .B(n35311), .Z(n40099) );
  IV U48264 ( .A(n35313), .Z(n35321) );
  IV U48265 ( .A(n35314), .Z(n35319) );
  NOR U48266 ( .A(n35316), .B(n35315), .Z(n35317) );
  IV U48267 ( .A(n35317), .Z(n35318) );
  NOR U48268 ( .A(n35319), .B(n35318), .Z(n36994) );
  IV U48269 ( .A(n35320), .Z(n36996) );
  XOR U48270 ( .A(n36994), .B(n36996), .Z(n36998) );
  NOR U48271 ( .A(n35321), .B(n36998), .Z(n40087) );
  IV U48272 ( .A(n35322), .Z(n35323) );
  NOR U48273 ( .A(n35323), .B(n36992), .Z(n40076) );
  IV U48274 ( .A(n40076), .Z(n41900) );
  IV U48275 ( .A(n35324), .Z(n35326) );
  NOR U48276 ( .A(n35326), .B(n35325), .Z(n35327) );
  IV U48277 ( .A(n35327), .Z(n35328) );
  NOR U48278 ( .A(n35329), .B(n35328), .Z(n40073) );
  NOR U48279 ( .A(n38617), .B(n40073), .Z(n35330) );
  IV U48280 ( .A(n35330), .Z(n36990) );
  IV U48281 ( .A(n35331), .Z(n35333) );
  NOR U48282 ( .A(n35333), .B(n35332), .Z(n40056) );
  IV U48283 ( .A(n35334), .Z(n35345) );
  IV U48284 ( .A(n35335), .Z(n35340) );
  NOR U48285 ( .A(n35337), .B(n35336), .Z(n35338) );
  IV U48286 ( .A(n35338), .Z(n35339) );
  NOR U48287 ( .A(n35340), .B(n35339), .Z(n35341) );
  IV U48288 ( .A(n35341), .Z(n35342) );
  NOR U48289 ( .A(n35343), .B(n35342), .Z(n35344) );
  IV U48290 ( .A(n35344), .Z(n36987) );
  NOR U48291 ( .A(n35345), .B(n36987), .Z(n40053) );
  IV U48292 ( .A(n35346), .Z(n35347) );
  NOR U48293 ( .A(n36983), .B(n35347), .Z(n38623) );
  IV U48294 ( .A(n35348), .Z(n35350) );
  IV U48295 ( .A(n35349), .Z(n36981) );
  NOR U48296 ( .A(n35350), .B(n36981), .Z(n40047) );
  IV U48297 ( .A(n35351), .Z(n35352) );
  NOR U48298 ( .A(n35355), .B(n35352), .Z(n38633) );
  IV U48299 ( .A(n35353), .Z(n35354) );
  NOR U48300 ( .A(n35355), .B(n35354), .Z(n38640) );
  IV U48301 ( .A(n35356), .Z(n35359) );
  IV U48302 ( .A(n35357), .Z(n35358) );
  NOR U48303 ( .A(n35359), .B(n35358), .Z(n38637) );
  IV U48304 ( .A(n35360), .Z(n35362) );
  XOR U48305 ( .A(n35367), .B(n35365), .Z(n35361) );
  NOR U48306 ( .A(n35362), .B(n35361), .Z(n38647) );
  IV U48307 ( .A(n35363), .Z(n35364) );
  NOR U48308 ( .A(n35367), .B(n35364), .Z(n38644) );
  IV U48309 ( .A(n35365), .Z(n35366) );
  NOR U48310 ( .A(n35367), .B(n35366), .Z(n38653) );
  IV U48311 ( .A(n35368), .Z(n36978) );
  IV U48312 ( .A(n35369), .Z(n35370) );
  NOR U48313 ( .A(n36978), .B(n35370), .Z(n38650) );
  IV U48314 ( .A(n35371), .Z(n35373) );
  NOR U48315 ( .A(n35373), .B(n35372), .Z(n36973) );
  IV U48316 ( .A(n36973), .Z(n36966) );
  IV U48317 ( .A(n35374), .Z(n35375) );
  NOR U48318 ( .A(n35375), .B(n35377), .Z(n40035) );
  IV U48319 ( .A(n35376), .Z(n35378) );
  NOR U48320 ( .A(n35378), .B(n35377), .Z(n40032) );
  IV U48321 ( .A(n35379), .Z(n35381) );
  NOR U48322 ( .A(n35381), .B(n35380), .Z(n41946) );
  IV U48323 ( .A(n35382), .Z(n35384) );
  NOR U48324 ( .A(n35384), .B(n35383), .Z(n41944) );
  NOR U48325 ( .A(n41946), .B(n41944), .Z(n40029) );
  IV U48326 ( .A(n35385), .Z(n35387) );
  NOR U48327 ( .A(n35387), .B(n35386), .Z(n41949) );
  NOR U48328 ( .A(n41955), .B(n41949), .Z(n38662) );
  IV U48329 ( .A(n35388), .Z(n35389) );
  NOR U48330 ( .A(n35392), .B(n35389), .Z(n43452) );
  IV U48331 ( .A(n35390), .Z(n35391) );
  NOR U48332 ( .A(n35392), .B(n35391), .Z(n41961) );
  NOR U48333 ( .A(n43452), .B(n41961), .Z(n38660) );
  IV U48334 ( .A(n35393), .Z(n35400) );
  NOR U48335 ( .A(n35395), .B(n35394), .Z(n35396) );
  IV U48336 ( .A(n35396), .Z(n35397) );
  NOR U48337 ( .A(n35398), .B(n35397), .Z(n35399) );
  IV U48338 ( .A(n35399), .Z(n35406) );
  NOR U48339 ( .A(n35400), .B(n35406), .Z(n38663) );
  IV U48340 ( .A(n35401), .Z(n35404) );
  IV U48341 ( .A(n35402), .Z(n35403) );
  NOR U48342 ( .A(n35404), .B(n35403), .Z(n40012) );
  IV U48343 ( .A(n35405), .Z(n35407) );
  NOR U48344 ( .A(n35407), .B(n35406), .Z(n40016) );
  NOR U48345 ( .A(n40012), .B(n40016), .Z(n35408) );
  IV U48346 ( .A(n35408), .Z(n36963) );
  IV U48347 ( .A(n35409), .Z(n35411) );
  XOR U48348 ( .A(n35412), .B(n36960), .Z(n35410) );
  NOR U48349 ( .A(n35411), .B(n35410), .Z(n38666) );
  IV U48350 ( .A(n35412), .Z(n35413) );
  NOR U48351 ( .A(n35413), .B(n36960), .Z(n36954) );
  IV U48352 ( .A(n35414), .Z(n35415) );
  NOR U48353 ( .A(n35416), .B(n35415), .Z(n36951) );
  IV U48354 ( .A(n36951), .Z(n36946) );
  IV U48355 ( .A(n35417), .Z(n35419) );
  IV U48356 ( .A(n35418), .Z(n35423) );
  NOR U48357 ( .A(n35419), .B(n35423), .Z(n39997) );
  NOR U48358 ( .A(n35421), .B(n35420), .Z(n39992) );
  IV U48359 ( .A(n35422), .Z(n35424) );
  NOR U48360 ( .A(n35424), .B(n35423), .Z(n39999) );
  NOR U48361 ( .A(n39992), .B(n39999), .Z(n36943) );
  IV U48362 ( .A(n35425), .Z(n35427) );
  NOR U48363 ( .A(n35427), .B(n35426), .Z(n39987) );
  IV U48364 ( .A(n35428), .Z(n35430) );
  NOR U48365 ( .A(n35430), .B(n35429), .Z(n39994) );
  NOR U48366 ( .A(n39987), .B(n39994), .Z(n36942) );
  IV U48367 ( .A(n35431), .Z(n35432) );
  NOR U48368 ( .A(n35432), .B(n36937), .Z(n35433) );
  IV U48369 ( .A(n35433), .Z(n39984) );
  IV U48370 ( .A(n35434), .Z(n36928) );
  IV U48371 ( .A(n35435), .Z(n36931) );
  XOR U48372 ( .A(n36929), .B(n36931), .Z(n36925) );
  IV U48373 ( .A(n35436), .Z(n35437) );
  NOR U48374 ( .A(n35437), .B(n35439), .Z(n39976) );
  IV U48375 ( .A(n35438), .Z(n35440) );
  NOR U48376 ( .A(n35440), .B(n35439), .Z(n39972) );
  IV U48377 ( .A(n35441), .Z(n35442) );
  NOR U48378 ( .A(n35443), .B(n35442), .Z(n42000) );
  IV U48379 ( .A(n35444), .Z(n35445) );
  NOR U48380 ( .A(n35446), .B(n35445), .Z(n41994) );
  NOR U48381 ( .A(n42000), .B(n41994), .Z(n39971) );
  IV U48382 ( .A(n35447), .Z(n35449) );
  IV U48383 ( .A(n35448), .Z(n35455) );
  NOR U48384 ( .A(n35449), .B(n35455), .Z(n39964) );
  IV U48385 ( .A(n35450), .Z(n35453) );
  IV U48386 ( .A(n35451), .Z(n35452) );
  NOR U48387 ( .A(n35453), .B(n35452), .Z(n38669) );
  IV U48388 ( .A(n35454), .Z(n35456) );
  NOR U48389 ( .A(n35456), .B(n35455), .Z(n39966) );
  NOR U48390 ( .A(n38669), .B(n39966), .Z(n35457) );
  IV U48391 ( .A(n35457), .Z(n36923) );
  NOR U48392 ( .A(n35459), .B(n35458), .Z(n39955) );
  NOR U48393 ( .A(n39955), .B(n39961), .Z(n36922) );
  IV U48394 ( .A(n35460), .Z(n35462) );
  NOR U48395 ( .A(n35462), .B(n35461), .Z(n39951) );
  IV U48396 ( .A(n35463), .Z(n35464) );
  NOR U48397 ( .A(n35465), .B(n35464), .Z(n39957) );
  NOR U48398 ( .A(n39951), .B(n39957), .Z(n36921) );
  IV U48399 ( .A(n35466), .Z(n35467) );
  NOR U48400 ( .A(n35468), .B(n35467), .Z(n39948) );
  IV U48401 ( .A(n35469), .Z(n35471) );
  NOR U48402 ( .A(n35471), .B(n35470), .Z(n39937) );
  IV U48403 ( .A(n35472), .Z(n35474) );
  NOR U48404 ( .A(n35474), .B(n35473), .Z(n39945) );
  NOR U48405 ( .A(n39937), .B(n39945), .Z(n36920) );
  IV U48406 ( .A(n35475), .Z(n35477) );
  NOR U48407 ( .A(n35477), .B(n35476), .Z(n39930) );
  IV U48408 ( .A(n35478), .Z(n35480) );
  NOR U48409 ( .A(n35480), .B(n35479), .Z(n39926) );
  NOR U48410 ( .A(n39930), .B(n39926), .Z(n36919) );
  IV U48411 ( .A(n35481), .Z(n35482) );
  NOR U48412 ( .A(n35482), .B(n35484), .Z(n38676) );
  IV U48413 ( .A(n35483), .Z(n35485) );
  NOR U48414 ( .A(n35485), .B(n35484), .Z(n38671) );
  NOR U48415 ( .A(n38676), .B(n38671), .Z(n36915) );
  IV U48416 ( .A(n35486), .Z(n35491) );
  IV U48417 ( .A(n35487), .Z(n35488) );
  NOR U48418 ( .A(n35491), .B(n35488), .Z(n38673) );
  IV U48419 ( .A(n35489), .Z(n35490) );
  NOR U48420 ( .A(n35491), .B(n35490), .Z(n38682) );
  IV U48421 ( .A(n35492), .Z(n35494) );
  NOR U48422 ( .A(n35494), .B(n35493), .Z(n38679) );
  IV U48423 ( .A(n35495), .Z(n35498) );
  NOR U48424 ( .A(n36909), .B(n35496), .Z(n35497) );
  IV U48425 ( .A(n35497), .Z(n35500) );
  NOR U48426 ( .A(n35498), .B(n35500), .Z(n39921) );
  IV U48427 ( .A(n35499), .Z(n35501) );
  NOR U48428 ( .A(n35501), .B(n35500), .Z(n39918) );
  IV U48429 ( .A(n35502), .Z(n35503) );
  NOR U48430 ( .A(n35503), .B(n35505), .Z(n35504) );
  IV U48431 ( .A(n35504), .Z(n38689) );
  NOR U48432 ( .A(n35506), .B(n35505), .Z(n38694) );
  IV U48433 ( .A(n35507), .Z(n35508) );
  NOR U48434 ( .A(n35509), .B(n35508), .Z(n39913) );
  IV U48435 ( .A(n35510), .Z(n35511) );
  NOR U48436 ( .A(n35511), .B(n35514), .Z(n39905) );
  NOR U48437 ( .A(n39913), .B(n39905), .Z(n35512) );
  IV U48438 ( .A(n35512), .Z(n36906) );
  IV U48439 ( .A(n35513), .Z(n35515) );
  NOR U48440 ( .A(n35515), .B(n35514), .Z(n38697) );
  IV U48441 ( .A(n35516), .Z(n35517) );
  NOR U48442 ( .A(n35518), .B(n35517), .Z(n46553) );
  IV U48443 ( .A(n35519), .Z(n35521) );
  IV U48444 ( .A(n35520), .Z(n35525) );
  NOR U48445 ( .A(n35521), .B(n35525), .Z(n46564) );
  NOR U48446 ( .A(n46553), .B(n46564), .Z(n39907) );
  IV U48447 ( .A(n35522), .Z(n35523) );
  NOR U48448 ( .A(n35523), .B(n36894), .Z(n39898) );
  IV U48449 ( .A(n35524), .Z(n35526) );
  NOR U48450 ( .A(n35526), .B(n35525), .Z(n39902) );
  NOR U48451 ( .A(n39898), .B(n39902), .Z(n36904) );
  IV U48452 ( .A(n35527), .Z(n35528) );
  NOR U48453 ( .A(n36886), .B(n35528), .Z(n39880) );
  IV U48454 ( .A(n39880), .Z(n39878) );
  IV U48455 ( .A(n35529), .Z(n35535) );
  IV U48456 ( .A(n35530), .Z(n35531) );
  NOR U48457 ( .A(n35535), .B(n35531), .Z(n35532) );
  IV U48458 ( .A(n35532), .Z(n38709) );
  IV U48459 ( .A(n35533), .Z(n35534) );
  NOR U48460 ( .A(n35535), .B(n35534), .Z(n38705) );
  IV U48461 ( .A(n35536), .Z(n35537) );
  NOR U48462 ( .A(n36880), .B(n35537), .Z(n38713) );
  IV U48463 ( .A(n35538), .Z(n35539) );
  NOR U48464 ( .A(n35539), .B(n36866), .Z(n39858) );
  IV U48465 ( .A(n35540), .Z(n35542) );
  NOR U48466 ( .A(n35542), .B(n35541), .Z(n42079) );
  IV U48467 ( .A(n35543), .Z(n35545) );
  NOR U48468 ( .A(n35545), .B(n35544), .Z(n42074) );
  NOR U48469 ( .A(n42079), .B(n42074), .Z(n38721) );
  IV U48470 ( .A(n35546), .Z(n35547) );
  NOR U48471 ( .A(n35548), .B(n35547), .Z(n36861) );
  IV U48472 ( .A(n35549), .Z(n35552) );
  IV U48473 ( .A(n35550), .Z(n35551) );
  NOR U48474 ( .A(n35552), .B(n35551), .Z(n38729) );
  IV U48475 ( .A(n35553), .Z(n35554) );
  NOR U48476 ( .A(n35554), .B(n42104), .Z(n39831) );
  IV U48477 ( .A(n35555), .Z(n35562) );
  IV U48478 ( .A(n35556), .Z(n35557) );
  NOR U48479 ( .A(n35562), .B(n35557), .Z(n38734) );
  IV U48480 ( .A(n35558), .Z(n35559) );
  NOR U48481 ( .A(n35562), .B(n35559), .Z(n38741) );
  IV U48482 ( .A(n35560), .Z(n35561) );
  NOR U48483 ( .A(n35562), .B(n35561), .Z(n38738) );
  IV U48484 ( .A(n35563), .Z(n35564) );
  NOR U48485 ( .A(n35565), .B(n35564), .Z(n38768) );
  IV U48486 ( .A(n35566), .Z(n35567) );
  NOR U48487 ( .A(n35568), .B(n35567), .Z(n38760) );
  NOR U48488 ( .A(n38768), .B(n38760), .Z(n36803) );
  IV U48489 ( .A(n35569), .Z(n35571) );
  IV U48490 ( .A(n35570), .Z(n43298) );
  NOR U48491 ( .A(n35571), .B(n43298), .Z(n38765) );
  NOR U48492 ( .A(n35572), .B(n43298), .Z(n38771) );
  IV U48493 ( .A(n35573), .Z(n35574) );
  NOR U48494 ( .A(n35574), .B(n39808), .Z(n38776) );
  IV U48495 ( .A(n35575), .Z(n39807) );
  NOR U48496 ( .A(n35577), .B(n39807), .Z(n39812) );
  IV U48497 ( .A(n35576), .Z(n35578) );
  NOR U48498 ( .A(n35578), .B(n35577), .Z(n39815) );
  IV U48499 ( .A(n35579), .Z(n35581) );
  NOR U48500 ( .A(n35581), .B(n35580), .Z(n35582) );
  IV U48501 ( .A(n35582), .Z(n36792) );
  IV U48502 ( .A(n35583), .Z(n35584) );
  NOR U48503 ( .A(n35584), .B(n36781), .Z(n36774) );
  IV U48504 ( .A(n35585), .Z(n35587) );
  NOR U48505 ( .A(n35587), .B(n35586), .Z(n36771) );
  IV U48506 ( .A(n36771), .Z(n36764) );
  IV U48507 ( .A(n35588), .Z(n35589) );
  NOR U48508 ( .A(n35589), .B(n35595), .Z(n42163) );
  IV U48509 ( .A(n35590), .Z(n35591) );
  NOR U48510 ( .A(n35592), .B(n35591), .Z(n42158) );
  NOR U48511 ( .A(n42163), .B(n42158), .Z(n38790) );
  IV U48512 ( .A(n35593), .Z(n35594) );
  NOR U48513 ( .A(n35595), .B(n35594), .Z(n39791) );
  IV U48514 ( .A(n35596), .Z(n35598) );
  NOR U48515 ( .A(n35598), .B(n35597), .Z(n39780) );
  IV U48516 ( .A(n35599), .Z(n35600) );
  NOR U48517 ( .A(n35600), .B(n36714), .Z(n38815) );
  IV U48518 ( .A(n35601), .Z(n35604) );
  IV U48519 ( .A(n35602), .Z(n35603) );
  NOR U48520 ( .A(n35604), .B(n35603), .Z(n38807) );
  NOR U48521 ( .A(n38815), .B(n38807), .Z(n36711) );
  IV U48522 ( .A(n36715), .Z(n35605) );
  NOR U48523 ( .A(n35605), .B(n36714), .Z(n38812) );
  IV U48524 ( .A(n35606), .Z(n35610) );
  NOR U48525 ( .A(n35608), .B(n35607), .Z(n35609) );
  IV U48526 ( .A(n35609), .Z(n35612) );
  NOR U48527 ( .A(n35610), .B(n35612), .Z(n39759) );
  IV U48528 ( .A(n35611), .Z(n35613) );
  NOR U48529 ( .A(n35613), .B(n35612), .Z(n39756) );
  IV U48530 ( .A(n35614), .Z(n35615) );
  NOR U48531 ( .A(n35616), .B(n35615), .Z(n35617) );
  IV U48532 ( .A(n35617), .Z(n36703) );
  IV U48533 ( .A(n35618), .Z(n35619) );
  NOR U48534 ( .A(n35619), .B(n35622), .Z(n36692) );
  IV U48535 ( .A(n35620), .Z(n35621) );
  NOR U48536 ( .A(n35622), .B(n35621), .Z(n36689) );
  IV U48537 ( .A(n35623), .Z(n35624) );
  NOR U48538 ( .A(n35625), .B(n35624), .Z(n35626) );
  IV U48539 ( .A(n35626), .Z(n38825) );
  IV U48540 ( .A(n35627), .Z(n35628) );
  NOR U48541 ( .A(n35628), .B(n43227), .Z(n39747) );
  IV U48542 ( .A(n43228), .Z(n35629) );
  NOR U48543 ( .A(n35629), .B(n43227), .Z(n38826) );
  NOR U48544 ( .A(n39747), .B(n38826), .Z(n36687) );
  IV U48545 ( .A(n35630), .Z(n35632) );
  NOR U48546 ( .A(n35632), .B(n35631), .Z(n38830) );
  IV U48547 ( .A(n35633), .Z(n35634) );
  NOR U48548 ( .A(n35634), .B(n35637), .Z(n38833) );
  IV U48549 ( .A(n35635), .Z(n35636) );
  NOR U48550 ( .A(n35637), .B(n35636), .Z(n38836) );
  IV U48551 ( .A(n35638), .Z(n35639) );
  NOR U48552 ( .A(n35640), .B(n35639), .Z(n39742) );
  NOR U48553 ( .A(n38836), .B(n39742), .Z(n35641) );
  IV U48554 ( .A(n35641), .Z(n35642) );
  NOR U48555 ( .A(n38833), .B(n35642), .Z(n35643) );
  IV U48556 ( .A(n35643), .Z(n36680) );
  IV U48557 ( .A(n35644), .Z(n35645) );
  NOR U48558 ( .A(n35645), .B(n35650), .Z(n39739) );
  IV U48559 ( .A(n35646), .Z(n35648) );
  IV U48560 ( .A(n35647), .Z(n36677) );
  NOR U48561 ( .A(n35648), .B(n36677), .Z(n38840) );
  IV U48562 ( .A(n35649), .Z(n35651) );
  NOR U48563 ( .A(n35651), .B(n35650), .Z(n38841) );
  XOR U48564 ( .A(n38840), .B(n38841), .Z(n35652) );
  NOR U48565 ( .A(n39739), .B(n35652), .Z(n36679) );
  IV U48566 ( .A(n35653), .Z(n35654) );
  NOR U48567 ( .A(n35657), .B(n35654), .Z(n38845) );
  IV U48568 ( .A(n35655), .Z(n35656) );
  NOR U48569 ( .A(n35657), .B(n35656), .Z(n39724) );
  NOR U48570 ( .A(n35659), .B(n35658), .Z(n38857) );
  IV U48571 ( .A(n35660), .Z(n35662) );
  IV U48572 ( .A(n35661), .Z(n36674) );
  NOR U48573 ( .A(n35662), .B(n36674), .Z(n38852) );
  NOR U48574 ( .A(n38857), .B(n38852), .Z(n36671) );
  IV U48575 ( .A(n35663), .Z(n35664) );
  NOR U48576 ( .A(n35665), .B(n35664), .Z(n38854) );
  IV U48577 ( .A(n35666), .Z(n35668) );
  NOR U48578 ( .A(n35668), .B(n35667), .Z(n38864) );
  IV U48579 ( .A(n35669), .Z(n35671) );
  NOR U48580 ( .A(n35671), .B(n35670), .Z(n38861) );
  NOR U48581 ( .A(n38864), .B(n38861), .Z(n36669) );
  NOR U48582 ( .A(n35672), .B(n38867), .Z(n36668) );
  IV U48583 ( .A(n35673), .Z(n35674) );
  NOR U48584 ( .A(n35674), .B(n43189), .Z(n39718) );
  IV U48585 ( .A(n35675), .Z(n35679) );
  NOR U48586 ( .A(n35677), .B(n35676), .Z(n35678) );
  IV U48587 ( .A(n35678), .Z(n35682) );
  NOR U48588 ( .A(n35679), .B(n35682), .Z(n39715) );
  NOR U48589 ( .A(n39718), .B(n39715), .Z(n35680) );
  IV U48590 ( .A(n35680), .Z(n36667) );
  IV U48591 ( .A(n35681), .Z(n35683) );
  NOR U48592 ( .A(n35683), .B(n35682), .Z(n39712) );
  IV U48593 ( .A(n35684), .Z(n35686) );
  NOR U48594 ( .A(n35686), .B(n35685), .Z(n38873) );
  IV U48595 ( .A(n35687), .Z(n35689) );
  NOR U48596 ( .A(n35689), .B(n35688), .Z(n36656) );
  IV U48597 ( .A(n35690), .Z(n35691) );
  NOR U48598 ( .A(n35692), .B(n35691), .Z(n39694) );
  IV U48599 ( .A(n35693), .Z(n35694) );
  NOR U48600 ( .A(n35695), .B(n35694), .Z(n39700) );
  IV U48601 ( .A(n35696), .Z(n36646) );
  NOR U48602 ( .A(n35697), .B(n36646), .Z(n35698) );
  IV U48603 ( .A(n35698), .Z(n35699) );
  NOR U48604 ( .A(n35700), .B(n35699), .Z(n39690) );
  IV U48605 ( .A(n35701), .Z(n35702) );
  NOR U48606 ( .A(n35702), .B(n35708), .Z(n35703) );
  IV U48607 ( .A(n35703), .Z(n38887) );
  IV U48608 ( .A(n35704), .Z(n35705) );
  NOR U48609 ( .A(n35706), .B(n35705), .Z(n38891) );
  IV U48610 ( .A(n35707), .Z(n35709) );
  NOR U48611 ( .A(n35709), .B(n35708), .Z(n38884) );
  NOR U48612 ( .A(n38891), .B(n38884), .Z(n35710) );
  IV U48613 ( .A(n35710), .Z(n36644) );
  IV U48614 ( .A(n35711), .Z(n35712) );
  NOR U48615 ( .A(n35713), .B(n35712), .Z(n35714) );
  IV U48616 ( .A(n35714), .Z(n38906) );
  NOR U48617 ( .A(n35716), .B(n35715), .Z(n43142) );
  IV U48618 ( .A(n35717), .Z(n35719) );
  IV U48619 ( .A(n35718), .Z(n36633) );
  NOR U48620 ( .A(n35719), .B(n36633), .Z(n43148) );
  NOR U48621 ( .A(n43142), .B(n43148), .Z(n39679) );
  IV U48622 ( .A(n35720), .Z(n35721) );
  NOR U48623 ( .A(n35721), .B(n35726), .Z(n38907) );
  IV U48624 ( .A(n35722), .Z(n35723) );
  NOR U48625 ( .A(n35724), .B(n35723), .Z(n39672) );
  IV U48626 ( .A(n35725), .Z(n35727) );
  NOR U48627 ( .A(n35727), .B(n35726), .Z(n38911) );
  NOR U48628 ( .A(n39672), .B(n38911), .Z(n36629) );
  NOR U48629 ( .A(n35729), .B(n35728), .Z(n39668) );
  IV U48630 ( .A(n35730), .Z(n39663) );
  NOR U48631 ( .A(n35731), .B(n39663), .Z(n35732) );
  NOR U48632 ( .A(n39668), .B(n35732), .Z(n36628) );
  IV U48633 ( .A(n35733), .Z(n35735) );
  NOR U48634 ( .A(n35735), .B(n35734), .Z(n42322) );
  NOR U48635 ( .A(n35736), .B(n42316), .Z(n35737) );
  IV U48636 ( .A(n35737), .Z(n42329) );
  NOR U48637 ( .A(n35738), .B(n42329), .Z(n38925) );
  NOR U48638 ( .A(n42322), .B(n38925), .Z(n36622) );
  NOR U48639 ( .A(n35740), .B(n35739), .Z(n35741) );
  IV U48640 ( .A(n35741), .Z(n36618) );
  IV U48641 ( .A(n35742), .Z(n35744) );
  NOR U48642 ( .A(n35744), .B(n35743), .Z(n45461) );
  IV U48643 ( .A(n35745), .Z(n35746) );
  NOR U48644 ( .A(n35746), .B(n36616), .Z(n45454) );
  NOR U48645 ( .A(n45461), .B(n45454), .Z(n39649) );
  IV U48646 ( .A(n39649), .Z(n36613) );
  IV U48647 ( .A(n35747), .Z(n35751) );
  NOR U48648 ( .A(n35749), .B(n35748), .Z(n35750) );
  IV U48649 ( .A(n35750), .Z(n35753) );
  NOR U48650 ( .A(n35751), .B(n35753), .Z(n39642) );
  IV U48651 ( .A(n35752), .Z(n35754) );
  NOR U48652 ( .A(n35754), .B(n35753), .Z(n39645) );
  IV U48653 ( .A(n35755), .Z(n35760) );
  NOR U48654 ( .A(n35756), .B(n36606), .Z(n35757) );
  IV U48655 ( .A(n35757), .Z(n38943) );
  NOR U48656 ( .A(n35758), .B(n38943), .Z(n35759) );
  IV U48657 ( .A(n35759), .Z(n36610) );
  NOR U48658 ( .A(n35760), .B(n36610), .Z(n38936) );
  NOR U48659 ( .A(n39645), .B(n38936), .Z(n35761) );
  IV U48660 ( .A(n35761), .Z(n36612) );
  IV U48661 ( .A(n35762), .Z(n35764) );
  XOR U48662 ( .A(n35772), .B(n35774), .Z(n35763) );
  NOR U48663 ( .A(n35764), .B(n35763), .Z(n35765) );
  IV U48664 ( .A(n35765), .Z(n38957) );
  IV U48665 ( .A(n35766), .Z(n35767) );
  NOR U48666 ( .A(n35774), .B(n35767), .Z(n43099) );
  IV U48667 ( .A(n35768), .Z(n35771) );
  IV U48668 ( .A(n35769), .Z(n35770) );
  NOR U48669 ( .A(n35771), .B(n35770), .Z(n43106) );
  NOR U48670 ( .A(n43099), .B(n43106), .Z(n38962) );
  IV U48671 ( .A(n35772), .Z(n35773) );
  NOR U48672 ( .A(n35774), .B(n35773), .Z(n35775) );
  IV U48673 ( .A(n35775), .Z(n39631) );
  IV U48674 ( .A(n35776), .Z(n35778) );
  NOR U48675 ( .A(n35778), .B(n35777), .Z(n35779) );
  IV U48676 ( .A(n35779), .Z(n36567) );
  IV U48677 ( .A(n35780), .Z(n35782) );
  IV U48678 ( .A(n35781), .Z(n35789) );
  NOR U48679 ( .A(n35782), .B(n35789), .Z(n39606) );
  IV U48680 ( .A(n35783), .Z(n35785) );
  NOR U48681 ( .A(n35785), .B(n35784), .Z(n43080) );
  IV U48682 ( .A(n35786), .Z(n35787) );
  NOR U48683 ( .A(n35788), .B(n35787), .Z(n42369) );
  NOR U48684 ( .A(n43080), .B(n42369), .Z(n39605) );
  NOR U48685 ( .A(n35790), .B(n35789), .Z(n36554) );
  IV U48686 ( .A(n36554), .Z(n36546) );
  IV U48687 ( .A(n35791), .Z(n35793) );
  IV U48688 ( .A(n35792), .Z(n35795) );
  NOR U48689 ( .A(n35793), .B(n35795), .Z(n38975) );
  IV U48690 ( .A(n35794), .Z(n35796) );
  NOR U48691 ( .A(n35796), .B(n35795), .Z(n38973) );
  IV U48692 ( .A(n35797), .Z(n35800) );
  IV U48693 ( .A(n35798), .Z(n35799) );
  NOR U48694 ( .A(n35800), .B(n35799), .Z(n38981) );
  IV U48695 ( .A(n35801), .Z(n35802) );
  NOR U48696 ( .A(n35803), .B(n35802), .Z(n43034) );
  IV U48697 ( .A(n35804), .Z(n35806) );
  NOR U48698 ( .A(n35806), .B(n35805), .Z(n43041) );
  NOR U48699 ( .A(n43034), .B(n43041), .Z(n38992) );
  NOR U48700 ( .A(n35808), .B(n35807), .Z(n38994) );
  IV U48701 ( .A(n35809), .Z(n35812) );
  NOR U48702 ( .A(n35810), .B(n35821), .Z(n35811) );
  IV U48703 ( .A(n35811), .Z(n35814) );
  NOR U48704 ( .A(n35812), .B(n35814), .Z(n38999) );
  IV U48705 ( .A(n35813), .Z(n35815) );
  NOR U48706 ( .A(n35815), .B(n35814), .Z(n39008) );
  IV U48707 ( .A(n35816), .Z(n35817) );
  NOR U48708 ( .A(n35818), .B(n35817), .Z(n39014) );
  IV U48709 ( .A(n35819), .Z(n35820) );
  NOR U48710 ( .A(n35821), .B(n35820), .Z(n39011) );
  NOR U48711 ( .A(n39014), .B(n39011), .Z(n36535) );
  IV U48712 ( .A(n35822), .Z(n35823) );
  NOR U48713 ( .A(n35824), .B(n35823), .Z(n35825) );
  IV U48714 ( .A(n35825), .Z(n39592) );
  IV U48715 ( .A(n35826), .Z(n35828) );
  NOR U48716 ( .A(n35828), .B(n35827), .Z(n39594) );
  IV U48717 ( .A(n35829), .Z(n35836) );
  NOR U48718 ( .A(n35831), .B(n35830), .Z(n35832) );
  IV U48719 ( .A(n35832), .Z(n35833) );
  NOR U48720 ( .A(n35834), .B(n35833), .Z(n35835) );
  IV U48721 ( .A(n35835), .Z(n35839) );
  NOR U48722 ( .A(n35836), .B(n35839), .Z(n39590) );
  NOR U48723 ( .A(n39594), .B(n39590), .Z(n35837) );
  IV U48724 ( .A(n35837), .Z(n36518) );
  IV U48725 ( .A(n35838), .Z(n35840) );
  NOR U48726 ( .A(n35840), .B(n35839), .Z(n39587) );
  IV U48727 ( .A(n35841), .Z(n35842) );
  NOR U48728 ( .A(n35843), .B(n35842), .Z(n42412) );
  IV U48729 ( .A(n35844), .Z(n35845) );
  NOR U48730 ( .A(n35846), .B(n35845), .Z(n42408) );
  NOR U48731 ( .A(n42412), .B(n42408), .Z(n39584) );
  IV U48732 ( .A(n35847), .Z(n35848) );
  NOR U48733 ( .A(n35851), .B(n35848), .Z(n39581) );
  IV U48734 ( .A(n35849), .Z(n35850) );
  NOR U48735 ( .A(n35851), .B(n35850), .Z(n39576) );
  IV U48736 ( .A(n35852), .Z(n35853) );
  NOR U48737 ( .A(n35854), .B(n35853), .Z(n39018) );
  NOR U48738 ( .A(n39576), .B(n39018), .Z(n35855) );
  IV U48739 ( .A(n35855), .Z(n36516) );
  IV U48740 ( .A(n35856), .Z(n35859) );
  IV U48741 ( .A(n35857), .Z(n35858) );
  NOR U48742 ( .A(n35859), .B(n35858), .Z(n39570) );
  IV U48743 ( .A(n35860), .Z(n36513) );
  IV U48744 ( .A(n35861), .Z(n35862) );
  NOR U48745 ( .A(n36513), .B(n35862), .Z(n39021) );
  NOR U48746 ( .A(n39570), .B(n39021), .Z(n36510) );
  NOR U48747 ( .A(n35863), .B(n42424), .Z(n35864) );
  NOR U48748 ( .A(n35865), .B(n35864), .Z(n39568) );
  IV U48749 ( .A(n35866), .Z(n35867) );
  NOR U48750 ( .A(n39551), .B(n35867), .Z(n39558) );
  NOR U48751 ( .A(n39551), .B(n35868), .Z(n36509) );
  NOR U48752 ( .A(n35870), .B(n35869), .Z(n35871) );
  IV U48753 ( .A(n35871), .Z(n35872) );
  NOR U48754 ( .A(n35873), .B(n35872), .Z(n39023) );
  IV U48755 ( .A(n35874), .Z(n35879) );
  IV U48756 ( .A(n35875), .Z(n35876) );
  NOR U48757 ( .A(n35879), .B(n35876), .Z(n39026) );
  IV U48758 ( .A(n35877), .Z(n35878) );
  NOR U48759 ( .A(n35879), .B(n35878), .Z(n39528) );
  IV U48760 ( .A(n35880), .Z(n35881) );
  NOR U48761 ( .A(n35881), .B(n35887), .Z(n39532) );
  NOR U48762 ( .A(n39528), .B(n39532), .Z(n39524) );
  IV U48763 ( .A(n35882), .Z(n35883) );
  NOR U48764 ( .A(n35884), .B(n35883), .Z(n42446) );
  IV U48765 ( .A(n35885), .Z(n35886) );
  NOR U48766 ( .A(n35887), .B(n35886), .Z(n42439) );
  NOR U48767 ( .A(n42446), .B(n42439), .Z(n39029) );
  XOR U48768 ( .A(n36504), .B(n36505), .Z(n35888) );
  NOR U48769 ( .A(n35889), .B(n35888), .Z(n35890) );
  IV U48770 ( .A(n35890), .Z(n35891) );
  NOR U48771 ( .A(n35892), .B(n35891), .Z(n39517) );
  IV U48772 ( .A(n35893), .Z(n35894) );
  NOR U48773 ( .A(n35895), .B(n35894), .Z(n39506) );
  IV U48774 ( .A(n35896), .Z(n35898) );
  NOR U48775 ( .A(n35898), .B(n35897), .Z(n39496) );
  NOR U48776 ( .A(n35900), .B(n35899), .Z(n39501) );
  NOR U48777 ( .A(n39496), .B(n39501), .Z(n36482) );
  NOR U48778 ( .A(n35901), .B(n36474), .Z(n35902) );
  IV U48779 ( .A(n35902), .Z(n35903) );
  NOR U48780 ( .A(n35904), .B(n35903), .Z(n39489) );
  IV U48781 ( .A(n35905), .Z(n35906) );
  NOR U48782 ( .A(n35907), .B(n35906), .Z(n39044) );
  IV U48783 ( .A(n35908), .Z(n35911) );
  IV U48784 ( .A(n35909), .Z(n35910) );
  NOR U48785 ( .A(n35911), .B(n35910), .Z(n39485) );
  NOR U48786 ( .A(n39044), .B(n39485), .Z(n35912) );
  IV U48787 ( .A(n35912), .Z(n36472) );
  IV U48788 ( .A(n35913), .Z(n35914) );
  NOR U48789 ( .A(n35914), .B(n35918), .Z(n39482) );
  IV U48790 ( .A(n35915), .Z(n35916) );
  NOR U48791 ( .A(n35917), .B(n35916), .Z(n42471) );
  NOR U48792 ( .A(n35919), .B(n35918), .Z(n42927) );
  NOR U48793 ( .A(n42471), .B(n42927), .Z(n39479) );
  IV U48794 ( .A(n35920), .Z(n35921) );
  NOR U48795 ( .A(n36464), .B(n35921), .Z(n36466) );
  IV U48796 ( .A(n35922), .Z(n35924) );
  NOR U48797 ( .A(n35924), .B(n35923), .Z(n35925) );
  IV U48798 ( .A(n35925), .Z(n39475) );
  IV U48799 ( .A(n35926), .Z(n36448) );
  NOR U48800 ( .A(n36448), .B(n36447), .Z(n39046) );
  IV U48801 ( .A(n35927), .Z(n35928) );
  NOR U48802 ( .A(n35929), .B(n35928), .Z(n39051) );
  IV U48803 ( .A(n35930), .Z(n35932) );
  NOR U48804 ( .A(n35932), .B(n35931), .Z(n39053) );
  IV U48805 ( .A(n35933), .Z(n35935) );
  NOR U48806 ( .A(n35935), .B(n35934), .Z(n39055) );
  NOR U48807 ( .A(n39053), .B(n39055), .Z(n35936) );
  IV U48808 ( .A(n35936), .Z(n35937) );
  NOR U48809 ( .A(n39051), .B(n35937), .Z(n35938) );
  IV U48810 ( .A(n35938), .Z(n36445) );
  IV U48811 ( .A(n35939), .Z(n35941) );
  NOR U48812 ( .A(n35941), .B(n35940), .Z(n39069) );
  NOR U48813 ( .A(n39067), .B(n39069), .Z(n36437) );
  IV U48814 ( .A(n35942), .Z(n35943) );
  NOR U48815 ( .A(n36433), .B(n35943), .Z(n39064) );
  NOR U48816 ( .A(n35945), .B(n35944), .Z(n35946) );
  IV U48817 ( .A(n35946), .Z(n36434) );
  NOR U48818 ( .A(n35947), .B(n36434), .Z(n35948) );
  IV U48819 ( .A(n35948), .Z(n39080) );
  IV U48820 ( .A(n35949), .Z(n35951) );
  IV U48821 ( .A(n35950), .Z(n36429) );
  NOR U48822 ( .A(n35951), .B(n36429), .Z(n39081) );
  NOR U48823 ( .A(n35953), .B(n35952), .Z(n35954) );
  IV U48824 ( .A(n35954), .Z(n35955) );
  NOR U48825 ( .A(n35956), .B(n35955), .Z(n35957) );
  IV U48826 ( .A(n35957), .Z(n36413) );
  NOR U48827 ( .A(n35958), .B(n36413), .Z(n35959) );
  IV U48828 ( .A(n35959), .Z(n35960) );
  NOR U48829 ( .A(n36412), .B(n35960), .Z(n39098) );
  NOR U48830 ( .A(n39095), .B(n39098), .Z(n36415) );
  IV U48831 ( .A(n35961), .Z(n36411) );
  IV U48832 ( .A(n35962), .Z(n35963) );
  NOR U48833 ( .A(n36411), .B(n35963), .Z(n39102) );
  IV U48834 ( .A(n35964), .Z(n35966) );
  NOR U48835 ( .A(n35966), .B(n35965), .Z(n39443) );
  IV U48836 ( .A(n35967), .Z(n35968) );
  NOR U48837 ( .A(n35968), .B(n35973), .Z(n39440) );
  IV U48838 ( .A(n35969), .Z(n35971) );
  NOR U48839 ( .A(n35971), .B(n35970), .Z(n39110) );
  IV U48840 ( .A(n35972), .Z(n35974) );
  NOR U48841 ( .A(n35974), .B(n35973), .Z(n39107) );
  NOR U48842 ( .A(n39110), .B(n39107), .Z(n36408) );
  IV U48843 ( .A(n35975), .Z(n35976) );
  NOR U48844 ( .A(n35977), .B(n35976), .Z(n35978) );
  IV U48845 ( .A(n35978), .Z(n36404) );
  IV U48846 ( .A(n35979), .Z(n35981) );
  IV U48847 ( .A(n35980), .Z(n36401) );
  NOR U48848 ( .A(n35981), .B(n36401), .Z(n36395) );
  IV U48849 ( .A(n36395), .Z(n36379) );
  IV U48850 ( .A(n35982), .Z(n35984) );
  NOR U48851 ( .A(n35984), .B(n35983), .Z(n39428) );
  IV U48852 ( .A(n35985), .Z(n35987) );
  IV U48853 ( .A(n35986), .Z(n35995) );
  NOR U48854 ( .A(n35987), .B(n35995), .Z(n42858) );
  IV U48855 ( .A(n35988), .Z(n35990) );
  NOR U48856 ( .A(n35990), .B(n35989), .Z(n42557) );
  NOR U48857 ( .A(n42858), .B(n42557), .Z(n39123) );
  IV U48858 ( .A(n39123), .Z(n36365) );
  NOR U48859 ( .A(n35992), .B(n35991), .Z(n39125) );
  IV U48860 ( .A(n35993), .Z(n35994) );
  NOR U48861 ( .A(n35995), .B(n35994), .Z(n39423) );
  NOR U48862 ( .A(n39125), .B(n39423), .Z(n36364) );
  IV U48863 ( .A(n35996), .Z(n35997) );
  NOR U48864 ( .A(n35998), .B(n35997), .Z(n39129) );
  IV U48865 ( .A(n35999), .Z(n36000) );
  NOR U48866 ( .A(n36001), .B(n36000), .Z(n39127) );
  NOR U48867 ( .A(n39129), .B(n39127), .Z(n36363) );
  IV U48868 ( .A(n36002), .Z(n36004) );
  NOR U48869 ( .A(n36004), .B(n36003), .Z(n39135) );
  IV U48870 ( .A(n36005), .Z(n36007) );
  NOR U48871 ( .A(n36007), .B(n36006), .Z(n36008) );
  IV U48872 ( .A(n36008), .Z(n36015) );
  NOR U48873 ( .A(n36010), .B(n36009), .Z(n36011) );
  IV U48874 ( .A(n36011), .Z(n36012) );
  NOR U48875 ( .A(n36013), .B(n36012), .Z(n36014) );
  IV U48876 ( .A(n36014), .Z(n36017) );
  NOR U48877 ( .A(n36015), .B(n36017), .Z(n39138) );
  IV U48878 ( .A(n36016), .Z(n36018) );
  NOR U48879 ( .A(n36018), .B(n36017), .Z(n39143) );
  NOR U48880 ( .A(n39138), .B(n39143), .Z(n36352) );
  IV U48881 ( .A(n36019), .Z(n36021) );
  IV U48882 ( .A(n36020), .Z(n36026) );
  NOR U48883 ( .A(n36021), .B(n36026), .Z(n36022) );
  IV U48884 ( .A(n36022), .Z(n39417) );
  NOR U48885 ( .A(n36024), .B(n36023), .Z(n39155) );
  IV U48886 ( .A(n36025), .Z(n36027) );
  NOR U48887 ( .A(n36027), .B(n36026), .Z(n39413) );
  NOR U48888 ( .A(n39155), .B(n39413), .Z(n36028) );
  IV U48889 ( .A(n36028), .Z(n36344) );
  IV U48890 ( .A(n36029), .Z(n36030) );
  NOR U48891 ( .A(n36030), .B(n36032), .Z(n39152) );
  IV U48892 ( .A(n36031), .Z(n36033) );
  NOR U48893 ( .A(n36033), .B(n36032), .Z(n39399) );
  IV U48894 ( .A(n36034), .Z(n36039) );
  NOR U48895 ( .A(n36035), .B(n36045), .Z(n36036) );
  IV U48896 ( .A(n36036), .Z(n36338) );
  NOR U48897 ( .A(n36037), .B(n36338), .Z(n36038) );
  IV U48898 ( .A(n36038), .Z(n36332) );
  NOR U48899 ( .A(n36039), .B(n36332), .Z(n36040) );
  IV U48900 ( .A(n36040), .Z(n39158) );
  IV U48901 ( .A(n36041), .Z(n36043) );
  NOR U48902 ( .A(n36043), .B(n36042), .Z(n39373) );
  IV U48903 ( .A(n36044), .Z(n36046) );
  NOR U48904 ( .A(n36046), .B(n36045), .Z(n39162) );
  NOR U48905 ( .A(n39373), .B(n39162), .Z(n36329) );
  IV U48906 ( .A(n36047), .Z(n36049) );
  IV U48907 ( .A(n36048), .Z(n39167) );
  NOR U48908 ( .A(n36049), .B(n39167), .Z(n39370) );
  NOR U48909 ( .A(n36051), .B(n36050), .Z(n36321) );
  IV U48910 ( .A(n36052), .Z(n36053) );
  NOR U48911 ( .A(n36054), .B(n36053), .Z(n39364) );
  IV U48912 ( .A(n36055), .Z(n36057) );
  NOR U48913 ( .A(n36057), .B(n36056), .Z(n39366) );
  NOR U48914 ( .A(n39364), .B(n39366), .Z(n36320) );
  IV U48915 ( .A(n36058), .Z(n42602) );
  IV U48916 ( .A(n36059), .Z(n42605) );
  NOR U48917 ( .A(n42602), .B(n42605), .Z(n39353) );
  IV U48918 ( .A(n36060), .Z(n36061) );
  NOR U48919 ( .A(n36062), .B(n36061), .Z(n39358) );
  NOR U48920 ( .A(n39353), .B(n39358), .Z(n36312) );
  NOR U48921 ( .A(n36064), .B(n36063), .Z(n42800) );
  IV U48922 ( .A(n36065), .Z(n36068) );
  IV U48923 ( .A(n36066), .Z(n36067) );
  NOR U48924 ( .A(n36068), .B(n36067), .Z(n39173) );
  NOR U48925 ( .A(n42800), .B(n39173), .Z(n36309) );
  IV U48926 ( .A(n36069), .Z(n36070) );
  NOR U48927 ( .A(n36071), .B(n36070), .Z(n36307) );
  IV U48928 ( .A(n36307), .Z(n36297) );
  IV U48929 ( .A(n36288), .Z(n36072) );
  NOR U48930 ( .A(n36284), .B(n36072), .Z(n36073) );
  IV U48931 ( .A(n36073), .Z(n36080) );
  XOR U48932 ( .A(n36075), .B(n36074), .Z(n36076) );
  NOR U48933 ( .A(n36077), .B(n36076), .Z(n36078) );
  IV U48934 ( .A(n36078), .Z(n36079) );
  NOR U48935 ( .A(n36080), .B(n36079), .Z(n36081) );
  IV U48936 ( .A(n36081), .Z(n39331) );
  IV U48937 ( .A(n36082), .Z(n36083) );
  NOR U48938 ( .A(n36084), .B(n36083), .Z(n36085) );
  IV U48939 ( .A(n36085), .Z(n36279) );
  NOR U48940 ( .A(n36087), .B(n36086), .Z(n36088) );
  IV U48941 ( .A(n36088), .Z(n36267) );
  IV U48942 ( .A(n36089), .Z(n36091) );
  IV U48943 ( .A(n36090), .Z(n36257) );
  NOR U48944 ( .A(n36091), .B(n36257), .Z(n39195) );
  IV U48945 ( .A(n36092), .Z(n36093) );
  NOR U48946 ( .A(n36094), .B(n36093), .Z(n42649) );
  IV U48947 ( .A(n36095), .Z(n36096) );
  NOR U48948 ( .A(n36096), .B(n36254), .Z(n42644) );
  NOR U48949 ( .A(n42649), .B(n42644), .Z(n39318) );
  IV U48950 ( .A(n36097), .Z(n36099) );
  NOR U48951 ( .A(n36099), .B(n36098), .Z(n36248) );
  IV U48952 ( .A(n36100), .Z(n36102) );
  NOR U48953 ( .A(n36102), .B(n36101), .Z(n39313) );
  IV U48954 ( .A(n36103), .Z(n36105) );
  NOR U48955 ( .A(n36105), .B(n36104), .Z(n36236) );
  IV U48956 ( .A(n36106), .Z(n36107) );
  NOR U48957 ( .A(n36108), .B(n36107), .Z(n36225) );
  IV U48958 ( .A(n36225), .Z(n36219) );
  IV U48959 ( .A(n36109), .Z(n36110) );
  NOR U48960 ( .A(n36111), .B(n36110), .Z(n39211) );
  IV U48961 ( .A(n36112), .Z(n36122) );
  IV U48962 ( .A(n36113), .Z(n36114) );
  NOR U48963 ( .A(n36122), .B(n36114), .Z(n36115) );
  IV U48964 ( .A(n36115), .Z(n39214) );
  IV U48965 ( .A(n36116), .Z(n36119) );
  IV U48966 ( .A(n36117), .Z(n36118) );
  NOR U48967 ( .A(n36119), .B(n36118), .Z(n42664) );
  IV U48968 ( .A(n36120), .Z(n36121) );
  NOR U48969 ( .A(n36122), .B(n36121), .Z(n42659) );
  NOR U48970 ( .A(n42664), .B(n42659), .Z(n39215) );
  IV U48971 ( .A(n36123), .Z(n42673) );
  IV U48972 ( .A(n36124), .Z(n36125) );
  NOR U48973 ( .A(n42673), .B(n36125), .Z(n39219) );
  IV U48974 ( .A(n36126), .Z(n36127) );
  NOR U48975 ( .A(n36127), .B(n36130), .Z(n36128) );
  IV U48976 ( .A(n36128), .Z(n39308) );
  IV U48977 ( .A(n36129), .Z(n36131) );
  NOR U48978 ( .A(n36131), .B(n36130), .Z(n36213) );
  IV U48979 ( .A(n36132), .Z(n36133) );
  NOR U48980 ( .A(n36135), .B(n36133), .Z(n39280) );
  IV U48981 ( .A(n36134), .Z(n36136) );
  NOR U48982 ( .A(n36136), .B(n36135), .Z(n39276) );
  IV U48983 ( .A(n36137), .Z(n36186) );
  IV U48984 ( .A(n36138), .Z(n36139) );
  NOR U48985 ( .A(n36186), .B(n36139), .Z(n39229) );
  IV U48986 ( .A(n36140), .Z(n36141) );
  NOR U48987 ( .A(n36141), .B(n36146), .Z(n39260) );
  IV U48988 ( .A(n36142), .Z(n36144) );
  NOR U48989 ( .A(n36144), .B(n36143), .Z(n39235) );
  IV U48990 ( .A(n36145), .Z(n36147) );
  NOR U48991 ( .A(n36147), .B(n36146), .Z(n39232) );
  NOR U48992 ( .A(n39235), .B(n39232), .Z(n36148) );
  IV U48993 ( .A(n36148), .Z(n36180) );
  NOR U48994 ( .A(n36150), .B(n36149), .Z(n39236) );
  NOR U48995 ( .A(n36153), .B(n36151), .Z(n39241) );
  IV U48996 ( .A(n36152), .Z(n36154) );
  NOR U48997 ( .A(n36154), .B(n36153), .Z(n36158) );
  IV U48998 ( .A(n36155), .Z(n36156) );
  NOR U48999 ( .A(n36156), .B(n36175), .Z(n36157) );
  NOR U49000 ( .A(n36158), .B(n36157), .Z(n39240) );
  NOR U49001 ( .A(n36160), .B(n36159), .Z(n36164) );
  NOR U49002 ( .A(n36162), .B(n36161), .Z(n36163) );
  NOR U49003 ( .A(n36164), .B(n36163), .Z(n39246) );
  IV U49004 ( .A(n36165), .Z(n36167) );
  IV U49005 ( .A(n36166), .Z(n36172) );
  NOR U49006 ( .A(n36167), .B(n36172), .Z(n36170) );
  IV U49007 ( .A(n36170), .Z(n36168) );
  NOR U49008 ( .A(n39246), .B(n36168), .Z(n39249) );
  XOR U49009 ( .A(n39247), .B(n39246), .Z(n36169) );
  NOR U49010 ( .A(n36170), .B(n36169), .Z(n39254) );
  NOR U49011 ( .A(n39249), .B(n39254), .Z(n36178) );
  IV U49012 ( .A(n36171), .Z(n36173) );
  NOR U49013 ( .A(n36173), .B(n36172), .Z(n39250) );
  IV U49014 ( .A(n36174), .Z(n36176) );
  NOR U49015 ( .A(n36176), .B(n36175), .Z(n36177) );
  NOR U49016 ( .A(n39250), .B(n36177), .Z(n39248) );
  XOR U49017 ( .A(n36178), .B(n39248), .Z(n39239) );
  XOR U49018 ( .A(n39240), .B(n39239), .Z(n36179) );
  IV U49019 ( .A(n36179), .Z(n39243) );
  XOR U49020 ( .A(n39241), .B(n39243), .Z(n39238) );
  XOR U49021 ( .A(n39236), .B(n39238), .Z(n39233) );
  XOR U49022 ( .A(n36180), .B(n39233), .Z(n39262) );
  XOR U49023 ( .A(n39260), .B(n39262), .Z(n39265) );
  IV U49024 ( .A(n36181), .Z(n36183) );
  NOR U49025 ( .A(n36183), .B(n36182), .Z(n39263) );
  XOR U49026 ( .A(n39265), .B(n39263), .Z(n39230) );
  XOR U49027 ( .A(n39229), .B(n39230), .Z(n39275) );
  IV U49028 ( .A(n36184), .Z(n36185) );
  NOR U49029 ( .A(n36186), .B(n36185), .Z(n39273) );
  XOR U49030 ( .A(n39275), .B(n39273), .Z(n39277) );
  XOR U49031 ( .A(n39276), .B(n39277), .Z(n39281) );
  XOR U49032 ( .A(n39280), .B(n39281), .Z(n39287) );
  IV U49033 ( .A(n36187), .Z(n36189) );
  NOR U49034 ( .A(n36189), .B(n36188), .Z(n39283) );
  IV U49035 ( .A(n36190), .Z(n36192) );
  NOR U49036 ( .A(n36192), .B(n36191), .Z(n39286) );
  NOR U49037 ( .A(n39283), .B(n39286), .Z(n36193) );
  XOR U49038 ( .A(n39287), .B(n36193), .Z(n39289) );
  NOR U49039 ( .A(n36195), .B(n36194), .Z(n42688) );
  NOR U49040 ( .A(n42688), .B(n42724), .Z(n39290) );
  XOR U49041 ( .A(n39289), .B(n39290), .Z(n39297) );
  IV U49042 ( .A(n36196), .Z(n36199) );
  IV U49043 ( .A(n36197), .Z(n36198) );
  NOR U49044 ( .A(n36199), .B(n36198), .Z(n39291) );
  IV U49045 ( .A(n36200), .Z(n36202) );
  IV U49046 ( .A(n36201), .Z(n36209) );
  NOR U49047 ( .A(n36202), .B(n36209), .Z(n39295) );
  NOR U49048 ( .A(n39291), .B(n39295), .Z(n36203) );
  XOR U49049 ( .A(n39297), .B(n36203), .Z(n36204) );
  IV U49050 ( .A(n36204), .Z(n39302) );
  IV U49051 ( .A(n36205), .Z(n36206) );
  NOR U49052 ( .A(n36207), .B(n36206), .Z(n39300) );
  IV U49053 ( .A(n36208), .Z(n36210) );
  NOR U49054 ( .A(n36210), .B(n36209), .Z(n39298) );
  NOR U49055 ( .A(n39300), .B(n39298), .Z(n36211) );
  XOR U49056 ( .A(n39302), .B(n36211), .Z(n36212) );
  NOR U49057 ( .A(n36213), .B(n36212), .Z(n36216) );
  IV U49058 ( .A(n36213), .Z(n36215) );
  XOR U49059 ( .A(n39302), .B(n39298), .Z(n36214) );
  NOR U49060 ( .A(n36215), .B(n36214), .Z(n45787) );
  NOR U49061 ( .A(n36216), .B(n45787), .Z(n39306) );
  XOR U49062 ( .A(n39308), .B(n39306), .Z(n39225) );
  XOR U49063 ( .A(n39224), .B(n39225), .Z(n42669) );
  XOR U49064 ( .A(n39227), .B(n42669), .Z(n39217) );
  XOR U49065 ( .A(n39216), .B(n39217), .Z(n39220) );
  XOR U49066 ( .A(n39219), .B(n39220), .Z(n42661) );
  XOR U49067 ( .A(n39215), .B(n42661), .Z(n36217) );
  XOR U49068 ( .A(n39214), .B(n36217), .Z(n39213) );
  XOR U49069 ( .A(n39211), .B(n39213), .Z(n36218) );
  NOR U49070 ( .A(n36219), .B(n36218), .Z(n42751) );
  IV U49071 ( .A(n36220), .Z(n36221) );
  NOR U49072 ( .A(n36222), .B(n36221), .Z(n39209) );
  NOR U49073 ( .A(n39211), .B(n39209), .Z(n36223) );
  XOR U49074 ( .A(n39213), .B(n36223), .Z(n36224) );
  NOR U49075 ( .A(n36225), .B(n36224), .Z(n36226) );
  NOR U49076 ( .A(n42751), .B(n36226), .Z(n36227) );
  IV U49077 ( .A(n36227), .Z(n39206) );
  IV U49078 ( .A(n36228), .Z(n36230) );
  NOR U49079 ( .A(n36230), .B(n36229), .Z(n39205) );
  IV U49080 ( .A(n36231), .Z(n36232) );
  NOR U49081 ( .A(n36233), .B(n36232), .Z(n39203) );
  NOR U49082 ( .A(n39205), .B(n39203), .Z(n36234) );
  XOR U49083 ( .A(n39206), .B(n36234), .Z(n36235) );
  NOR U49084 ( .A(n36236), .B(n36235), .Z(n36239) );
  IV U49085 ( .A(n36236), .Z(n36238) );
  XOR U49086 ( .A(n39205), .B(n39206), .Z(n36237) );
  NOR U49087 ( .A(n36238), .B(n36237), .Z(n42759) );
  NOR U49088 ( .A(n36239), .B(n42759), .Z(n36246) );
  XOR U49089 ( .A(n39313), .B(n36246), .Z(n36249) );
  NOR U49090 ( .A(n36248), .B(n36249), .Z(n36240) );
  IV U49091 ( .A(n36240), .Z(n36244) );
  IV U49092 ( .A(n36241), .Z(n36243) );
  NOR U49093 ( .A(n36243), .B(n36242), .Z(n36245) );
  NOR U49094 ( .A(n36244), .B(n36245), .Z(n36252) );
  IV U49095 ( .A(n36245), .Z(n36247) );
  IV U49096 ( .A(n36246), .Z(n39314) );
  NOR U49097 ( .A(n36247), .B(n39314), .Z(n45877) );
  IV U49098 ( .A(n36248), .Z(n36251) );
  IV U49099 ( .A(n36249), .Z(n36250) );
  NOR U49100 ( .A(n36251), .B(n36250), .Z(n45769) );
  NOR U49101 ( .A(n45877), .B(n45769), .Z(n42652) );
  IV U49102 ( .A(n42652), .Z(n39319) );
  NOR U49103 ( .A(n36252), .B(n39319), .Z(n39317) );
  XOR U49104 ( .A(n39318), .B(n39317), .Z(n39323) );
  IV U49105 ( .A(n39323), .Z(n36260) );
  IV U49106 ( .A(n36253), .Z(n36255) );
  NOR U49107 ( .A(n36255), .B(n36254), .Z(n39322) );
  IV U49108 ( .A(n36256), .Z(n36258) );
  NOR U49109 ( .A(n36258), .B(n36257), .Z(n39201) );
  NOR U49110 ( .A(n39322), .B(n39201), .Z(n36259) );
  XOR U49111 ( .A(n36260), .B(n36259), .Z(n39197) );
  XOR U49112 ( .A(n39195), .B(n39197), .Z(n36262) );
  NOR U49113 ( .A(n36267), .B(n36262), .Z(n42637) );
  NOR U49114 ( .A(n36261), .B(n39192), .Z(n36263) );
  XOR U49115 ( .A(n36263), .B(n36262), .Z(n39187) );
  IV U49116 ( .A(n36264), .Z(n36266) );
  IV U49117 ( .A(n36265), .Z(n36276) );
  NOR U49118 ( .A(n36266), .B(n36276), .Z(n36268) );
  IV U49119 ( .A(n36268), .Z(n39186) );
  XOR U49120 ( .A(n39187), .B(n39186), .Z(n36270) );
  NOR U49121 ( .A(n36268), .B(n36267), .Z(n36269) );
  NOR U49122 ( .A(n36270), .B(n36269), .Z(n36271) );
  NOR U49123 ( .A(n42637), .B(n36271), .Z(n36278) );
  IV U49124 ( .A(n36278), .Z(n39190) );
  NOR U49125 ( .A(n36279), .B(n39190), .Z(n42625) );
  IV U49126 ( .A(n36272), .Z(n36274) );
  NOR U49127 ( .A(n36274), .B(n36273), .Z(n39182) );
  IV U49128 ( .A(n36275), .Z(n36277) );
  NOR U49129 ( .A(n36277), .B(n36276), .Z(n39188) );
  XOR U49130 ( .A(n36278), .B(n39188), .Z(n39183) );
  XOR U49131 ( .A(n39182), .B(n39183), .Z(n36281) );
  NOR U49132 ( .A(n39183), .B(n36279), .Z(n36280) );
  NOR U49133 ( .A(n36281), .B(n36280), .Z(n36282) );
  NOR U49134 ( .A(n42625), .B(n36282), .Z(n39329) );
  XOR U49135 ( .A(n39331), .B(n39329), .Z(n39181) );
  IV U49136 ( .A(n36283), .Z(n36285) );
  NOR U49137 ( .A(n36285), .B(n36284), .Z(n36286) );
  IV U49138 ( .A(n36286), .Z(n36287) );
  NOR U49139 ( .A(n36288), .B(n36287), .Z(n39179) );
  XOR U49140 ( .A(n39181), .B(n39179), .Z(n39342) );
  IV U49141 ( .A(n36289), .Z(n36291) );
  NOR U49142 ( .A(n36291), .B(n36290), .Z(n39341) );
  IV U49143 ( .A(n36292), .Z(n36294) );
  NOR U49144 ( .A(n36294), .B(n36293), .Z(n39339) );
  NOR U49145 ( .A(n39341), .B(n39339), .Z(n36295) );
  XOR U49146 ( .A(n39342), .B(n36295), .Z(n36301) );
  IV U49147 ( .A(n36301), .Z(n36296) );
  NOR U49148 ( .A(n36297), .B(n36296), .Z(n42786) );
  IV U49149 ( .A(n36298), .Z(n36300) );
  NOR U49150 ( .A(n36300), .B(n36299), .Z(n36302) );
  NOR U49151 ( .A(n36302), .B(n36301), .Z(n36305) );
  IV U49152 ( .A(n36302), .Z(n36304) );
  XOR U49153 ( .A(n39341), .B(n39342), .Z(n36303) );
  NOR U49154 ( .A(n36304), .B(n36303), .Z(n42783) );
  NOR U49155 ( .A(n36305), .B(n42783), .Z(n36306) );
  NOR U49156 ( .A(n36307), .B(n36306), .Z(n36308) );
  NOR U49157 ( .A(n42786), .B(n36308), .Z(n39174) );
  XOR U49158 ( .A(n36309), .B(n39174), .Z(n42607) );
  IV U49159 ( .A(n42603), .Z(n36310) );
  NOR U49160 ( .A(n42602), .B(n36310), .Z(n39351) );
  NOR U49161 ( .A(n42608), .B(n39351), .Z(n36311) );
  XOR U49162 ( .A(n42607), .B(n36311), .Z(n39354) );
  XOR U49163 ( .A(n36312), .B(n39354), .Z(n42596) );
  IV U49164 ( .A(n36313), .Z(n36315) );
  NOR U49165 ( .A(n36315), .B(n36314), .Z(n42595) );
  IV U49166 ( .A(n36316), .Z(n36318) );
  NOR U49167 ( .A(n36318), .B(n36317), .Z(n42810) );
  NOR U49168 ( .A(n42595), .B(n42810), .Z(n39361) );
  XOR U49169 ( .A(n42596), .B(n39361), .Z(n36319) );
  IV U49170 ( .A(n36319), .Z(n39367) );
  XOR U49171 ( .A(n36320), .B(n39367), .Z(n39165) );
  NOR U49172 ( .A(n36321), .B(n39165), .Z(n36324) );
  IV U49173 ( .A(n36321), .Z(n36323) );
  XOR U49174 ( .A(n39364), .B(n39367), .Z(n36322) );
  NOR U49175 ( .A(n36323), .B(n36322), .Z(n42819) );
  NOR U49176 ( .A(n36324), .B(n42819), .Z(n36327) );
  NOR U49177 ( .A(n36325), .B(n39167), .Z(n36326) );
  XOR U49178 ( .A(n36327), .B(n36326), .Z(n36328) );
  IV U49179 ( .A(n36328), .Z(n39371) );
  XOR U49180 ( .A(n39370), .B(n39371), .Z(n39374) );
  XOR U49181 ( .A(n36329), .B(n39374), .Z(n36330) );
  IV U49182 ( .A(n36330), .Z(n39381) );
  IV U49183 ( .A(n36331), .Z(n36333) );
  NOR U49184 ( .A(n36333), .B(n36332), .Z(n39379) );
  XOR U49185 ( .A(n39381), .B(n39379), .Z(n39157) );
  XOR U49186 ( .A(n39158), .B(n39157), .Z(n39159) );
  IV U49187 ( .A(n36334), .Z(n36343) );
  IV U49188 ( .A(n36335), .Z(n36336) );
  NOR U49189 ( .A(n36343), .B(n36336), .Z(n39392) );
  IV U49190 ( .A(n36337), .Z(n36339) );
  NOR U49191 ( .A(n36339), .B(n36338), .Z(n39160) );
  NOR U49192 ( .A(n39392), .B(n39160), .Z(n36340) );
  XOR U49193 ( .A(n39159), .B(n36340), .Z(n39398) );
  IV U49194 ( .A(n36341), .Z(n36342) );
  NOR U49195 ( .A(n36343), .B(n36342), .Z(n39396) );
  XOR U49196 ( .A(n39398), .B(n39396), .Z(n39401) );
  XOR U49197 ( .A(n39399), .B(n39401), .Z(n39153) );
  XOR U49198 ( .A(n39152), .B(n39153), .Z(n39414) );
  XOR U49199 ( .A(n36344), .B(n39414), .Z(n39416) );
  XOR U49200 ( .A(n39417), .B(n39416), .Z(n39147) );
  IV U49201 ( .A(n36345), .Z(n36347) );
  NOR U49202 ( .A(n36347), .B(n36346), .Z(n39149) );
  IV U49203 ( .A(n36348), .Z(n36350) );
  NOR U49204 ( .A(n36350), .B(n36349), .Z(n39146) );
  NOR U49205 ( .A(n39149), .B(n39146), .Z(n36351) );
  XOR U49206 ( .A(n39147), .B(n36351), .Z(n39145) );
  XOR U49207 ( .A(n36352), .B(n39145), .Z(n39140) );
  IV U49208 ( .A(n36353), .Z(n36354) );
  NOR U49209 ( .A(n36354), .B(n36361), .Z(n36355) );
  NOR U49210 ( .A(n39140), .B(n36355), .Z(n36358) );
  IV U49211 ( .A(n36355), .Z(n39142) );
  XOR U49212 ( .A(n39143), .B(n39145), .Z(n36356) );
  NOR U49213 ( .A(n39142), .B(n36356), .Z(n36357) );
  NOR U49214 ( .A(n36358), .B(n36357), .Z(n36359) );
  IV U49215 ( .A(n36359), .Z(n39134) );
  IV U49216 ( .A(n36360), .Z(n36362) );
  NOR U49217 ( .A(n36362), .B(n36361), .Z(n39132) );
  XOR U49218 ( .A(n39134), .B(n39132), .Z(n39136) );
  XOR U49219 ( .A(n39135), .B(n39136), .Z(n39130) );
  XOR U49220 ( .A(n36363), .B(n39130), .Z(n39124) );
  XOR U49221 ( .A(n36364), .B(n39124), .Z(n42559) );
  XOR U49222 ( .A(n36365), .B(n42559), .Z(n39119) );
  IV U49223 ( .A(n36366), .Z(n36370) );
  NOR U49224 ( .A(n36368), .B(n36367), .Z(n36369) );
  IV U49225 ( .A(n36369), .Z(n36376) );
  NOR U49226 ( .A(n36370), .B(n36376), .Z(n36371) );
  IV U49227 ( .A(n36371), .Z(n39118) );
  XOR U49228 ( .A(n39119), .B(n39118), .Z(n39120) );
  IV U49229 ( .A(n36372), .Z(n36373) );
  NOR U49230 ( .A(n36374), .B(n36373), .Z(n39431) );
  IV U49231 ( .A(n36375), .Z(n36377) );
  NOR U49232 ( .A(n36377), .B(n36376), .Z(n39121) );
  NOR U49233 ( .A(n39431), .B(n39121), .Z(n36378) );
  XOR U49234 ( .A(n39120), .B(n36378), .Z(n39430) );
  XOR U49235 ( .A(n39428), .B(n39430), .Z(n36381) );
  NOR U49236 ( .A(n36379), .B(n36381), .Z(n42539) );
  NOR U49237 ( .A(n36380), .B(n36385), .Z(n36383) );
  IV U49238 ( .A(n36381), .Z(n36382) );
  NOR U49239 ( .A(n36383), .B(n36382), .Z(n36393) );
  IV U49240 ( .A(n36384), .Z(n36387) );
  NOR U49241 ( .A(n39430), .B(n36385), .Z(n36386) );
  IV U49242 ( .A(n36386), .Z(n36389) );
  NOR U49243 ( .A(n36387), .B(n36389), .Z(n42545) );
  IV U49244 ( .A(n36388), .Z(n36390) );
  NOR U49245 ( .A(n36390), .B(n36389), .Z(n42536) );
  NOR U49246 ( .A(n42545), .B(n42536), .Z(n36391) );
  IV U49247 ( .A(n36391), .Z(n36392) );
  NOR U49248 ( .A(n36393), .B(n36392), .Z(n36394) );
  NOR U49249 ( .A(n36395), .B(n36394), .Z(n36396) );
  NOR U49250 ( .A(n42539), .B(n36396), .Z(n36403) );
  IV U49251 ( .A(n36403), .Z(n39436) );
  NOR U49252 ( .A(n36404), .B(n39436), .Z(n42531) );
  IV U49253 ( .A(n36397), .Z(n36398) );
  NOR U49254 ( .A(n36399), .B(n36398), .Z(n39113) );
  IV U49255 ( .A(n36400), .Z(n36402) );
  NOR U49256 ( .A(n36402), .B(n36401), .Z(n39435) );
  XOR U49257 ( .A(n39435), .B(n36403), .Z(n39114) );
  XOR U49258 ( .A(n39113), .B(n39114), .Z(n36406) );
  NOR U49259 ( .A(n39114), .B(n36404), .Z(n36405) );
  NOR U49260 ( .A(n36406), .B(n36405), .Z(n36407) );
  NOR U49261 ( .A(n42531), .B(n36407), .Z(n39108) );
  XOR U49262 ( .A(n36408), .B(n39108), .Z(n39442) );
  XOR U49263 ( .A(n39440), .B(n39442), .Z(n39444) );
  XOR U49264 ( .A(n39443), .B(n39444), .Z(n39103) );
  XOR U49265 ( .A(n39102), .B(n39103), .Z(n42508) );
  IV U49266 ( .A(n36409), .Z(n36410) );
  NOR U49267 ( .A(n36411), .B(n36410), .Z(n42506) );
  IV U49268 ( .A(n36412), .Z(n36414) );
  NOR U49269 ( .A(n36414), .B(n36413), .Z(n42878) );
  NOR U49270 ( .A(n42506), .B(n42878), .Z(n39105) );
  XOR U49271 ( .A(n42508), .B(n39105), .Z(n39096) );
  XOR U49272 ( .A(n36415), .B(n39096), .Z(n39454) );
  IV U49273 ( .A(n36416), .Z(n36418) );
  NOR U49274 ( .A(n36418), .B(n36417), .Z(n39452) );
  XOR U49275 ( .A(n39454), .B(n39452), .Z(n39093) );
  IV U49276 ( .A(n36419), .Z(n36422) );
  IV U49277 ( .A(n36420), .Z(n36421) );
  NOR U49278 ( .A(n36422), .B(n36421), .Z(n39091) );
  XOR U49279 ( .A(n39093), .B(n39091), .Z(n39451) );
  IV U49280 ( .A(n36423), .Z(n36424) );
  NOR U49281 ( .A(n36427), .B(n36424), .Z(n39449) );
  XOR U49282 ( .A(n39451), .B(n39449), .Z(n39090) );
  IV U49283 ( .A(n36425), .Z(n36426) );
  NOR U49284 ( .A(n36427), .B(n36426), .Z(n39088) );
  XOR U49285 ( .A(n39090), .B(n39088), .Z(n39082) );
  XOR U49286 ( .A(n39081), .B(n39082), .Z(n39086) );
  IV U49287 ( .A(n36428), .Z(n36430) );
  NOR U49288 ( .A(n36430), .B(n36429), .Z(n39084) );
  XOR U49289 ( .A(n39086), .B(n39084), .Z(n39079) );
  XOR U49290 ( .A(n39080), .B(n39079), .Z(n39074) );
  IV U49291 ( .A(n36431), .Z(n36432) );
  NOR U49292 ( .A(n36433), .B(n36432), .Z(n39073) );
  NOR U49293 ( .A(n36435), .B(n36434), .Z(n39076) );
  NOR U49294 ( .A(n39073), .B(n39076), .Z(n36436) );
  XOR U49295 ( .A(n39074), .B(n36436), .Z(n39065) );
  XOR U49296 ( .A(n39064), .B(n39065), .Z(n39070) );
  XOR U49297 ( .A(n36437), .B(n39070), .Z(n39059) );
  IV U49298 ( .A(n36438), .Z(n36440) );
  NOR U49299 ( .A(n36440), .B(n36439), .Z(n39061) );
  IV U49300 ( .A(n36441), .Z(n36442) );
  NOR U49301 ( .A(n36443), .B(n36442), .Z(n39058) );
  NOR U49302 ( .A(n39061), .B(n39058), .Z(n36444) );
  XOR U49303 ( .A(n39059), .B(n36444), .Z(n39056) );
  XOR U49304 ( .A(n36445), .B(n39056), .Z(n39048) );
  XOR U49305 ( .A(n39046), .B(n39048), .Z(n39470) );
  IV U49306 ( .A(n36450), .Z(n36446) );
  NOR U49307 ( .A(n36446), .B(n36447), .Z(n39467) );
  XOR U49308 ( .A(n36448), .B(n36447), .Z(n36449) );
  NOR U49309 ( .A(n36450), .B(n36449), .Z(n36453) );
  IV U49310 ( .A(n36451), .Z(n36452) );
  NOR U49311 ( .A(n36453), .B(n36452), .Z(n39465) );
  NOR U49312 ( .A(n39467), .B(n39465), .Z(n36454) );
  XOR U49313 ( .A(n39470), .B(n36454), .Z(n39472) );
  IV U49314 ( .A(n36455), .Z(n36456) );
  NOR U49315 ( .A(n36457), .B(n36456), .Z(n42912) );
  IV U49316 ( .A(n36458), .Z(n36460) );
  NOR U49317 ( .A(n36460), .B(n36459), .Z(n42921) );
  NOR U49318 ( .A(n42912), .B(n42921), .Z(n39473) );
  XOR U49319 ( .A(n39472), .B(n39473), .Z(n39474) );
  XOR U49320 ( .A(n39475), .B(n39474), .Z(n36461) );
  NOR U49321 ( .A(n36466), .B(n36461), .Z(n36468) );
  IV U49322 ( .A(n36462), .Z(n36463) );
  NOR U49323 ( .A(n36464), .B(n36463), .Z(n36470) );
  IV U49324 ( .A(n36470), .Z(n36465) );
  NOR U49325 ( .A(n36468), .B(n36465), .Z(n42475) );
  IV U49326 ( .A(n36466), .Z(n36467) );
  NOR U49327 ( .A(n36467), .B(n39474), .Z(n49139) );
  NOR U49328 ( .A(n36468), .B(n49139), .Z(n36469) );
  NOR U49329 ( .A(n36470), .B(n36469), .Z(n36471) );
  NOR U49330 ( .A(n42475), .B(n36471), .Z(n39478) );
  XOR U49331 ( .A(n39479), .B(n39478), .Z(n39484) );
  XOR U49332 ( .A(n39482), .B(n39484), .Z(n39487) );
  XOR U49333 ( .A(n36472), .B(n39487), .Z(n39491) );
  XOR U49334 ( .A(n39489), .B(n39491), .Z(n39494) );
  IV U49335 ( .A(n36473), .Z(n36475) );
  NOR U49336 ( .A(n36475), .B(n36474), .Z(n39492) );
  XOR U49337 ( .A(n39494), .B(n39492), .Z(n42936) );
  IV U49338 ( .A(n36476), .Z(n36477) );
  NOR U49339 ( .A(n36478), .B(n36477), .Z(n42934) );
  IV U49340 ( .A(n36479), .Z(n36481) );
  NOR U49341 ( .A(n36481), .B(n36480), .Z(n42941) );
  NOR U49342 ( .A(n42934), .B(n42941), .Z(n39495) );
  XOR U49343 ( .A(n42936), .B(n39495), .Z(n39497) );
  XOR U49344 ( .A(n36482), .B(n39497), .Z(n42459) );
  XOR U49345 ( .A(n42457), .B(n42459), .Z(n42947) );
  IV U49346 ( .A(n36483), .Z(n36485) );
  NOR U49347 ( .A(n36485), .B(n36484), .Z(n39041) );
  NOR U49348 ( .A(n42945), .B(n39041), .Z(n36486) );
  XOR U49349 ( .A(n42947), .B(n36486), .Z(n39038) );
  IV U49350 ( .A(n36487), .Z(n36488) );
  NOR U49351 ( .A(n36489), .B(n36488), .Z(n39039) );
  IV U49352 ( .A(n36490), .Z(n36492) );
  NOR U49353 ( .A(n36492), .B(n36491), .Z(n39509) );
  NOR U49354 ( .A(n39039), .B(n39509), .Z(n36493) );
  XOR U49355 ( .A(n39038), .B(n36493), .Z(n39507) );
  XOR U49356 ( .A(n39506), .B(n39507), .Z(n39034) );
  IV U49357 ( .A(n36494), .Z(n36495) );
  NOR U49358 ( .A(n36496), .B(n36495), .Z(n39036) );
  IV U49359 ( .A(n36497), .Z(n36499) );
  NOR U49360 ( .A(n36499), .B(n36498), .Z(n39033) );
  NOR U49361 ( .A(n39036), .B(n39033), .Z(n36500) );
  XOR U49362 ( .A(n39034), .B(n36500), .Z(n39030) );
  IV U49363 ( .A(n36501), .Z(n36503) );
  NOR U49364 ( .A(n36503), .B(n36502), .Z(n39031) );
  IV U49365 ( .A(n36504), .Z(n36506) );
  NOR U49366 ( .A(n36506), .B(n36505), .Z(n39514) );
  NOR U49367 ( .A(n39031), .B(n39514), .Z(n36507) );
  XOR U49368 ( .A(n39030), .B(n36507), .Z(n39518) );
  XOR U49369 ( .A(n39517), .B(n39518), .Z(n42441) );
  XOR U49370 ( .A(n39029), .B(n42441), .Z(n39523) );
  XOR U49371 ( .A(n39524), .B(n39523), .Z(n39027) );
  XOR U49372 ( .A(n39026), .B(n39027), .Z(n39024) );
  XOR U49373 ( .A(n39023), .B(n39024), .Z(n39555) );
  XOR U49374 ( .A(n36508), .B(n39555), .Z(n39550) );
  XOR U49375 ( .A(n36509), .B(n39550), .Z(n39560) );
  XOR U49376 ( .A(n39558), .B(n39560), .Z(n42427) );
  XOR U49377 ( .A(n39568), .B(n42427), .Z(n39571) );
  XOR U49378 ( .A(n36510), .B(n39571), .Z(n39574) );
  IV U49379 ( .A(n36511), .Z(n36512) );
  NOR U49380 ( .A(n36513), .B(n36512), .Z(n43001) );
  NOR U49381 ( .A(n36515), .B(n36514), .Z(n42418) );
  NOR U49382 ( .A(n43001), .B(n42418), .Z(n39575) );
  XOR U49383 ( .A(n39574), .B(n39575), .Z(n39577) );
  XOR U49384 ( .A(n36516), .B(n39577), .Z(n39582) );
  XOR U49385 ( .A(n39581), .B(n39582), .Z(n42409) );
  XOR U49386 ( .A(n39584), .B(n42409), .Z(n36517) );
  IV U49387 ( .A(n36517), .Z(n39589) );
  XOR U49388 ( .A(n39587), .B(n39589), .Z(n39595) );
  XOR U49389 ( .A(n36518), .B(n39595), .Z(n39593) );
  XOR U49390 ( .A(n39592), .B(n39593), .Z(n36528) );
  IV U49391 ( .A(n36519), .Z(n36520) );
  NOR U49392 ( .A(n36521), .B(n36520), .Z(n36531) );
  IV U49393 ( .A(n36522), .Z(n36523) );
  NOR U49394 ( .A(n36524), .B(n36523), .Z(n36527) );
  NOR U49395 ( .A(n36531), .B(n36527), .Z(n36525) );
  IV U49396 ( .A(n36525), .Z(n36526) );
  NOR U49397 ( .A(n36528), .B(n36526), .Z(n36534) );
  IV U49398 ( .A(n36527), .Z(n36530) );
  IV U49399 ( .A(n36528), .Z(n36529) );
  NOR U49400 ( .A(n36530), .B(n36529), .Z(n43018) );
  IV U49401 ( .A(n36531), .Z(n36532) );
  NOR U49402 ( .A(n39593), .B(n36532), .Z(n42394) );
  NOR U49403 ( .A(n43018), .B(n42394), .Z(n36533) );
  IV U49404 ( .A(n36533), .Z(n39017) );
  NOR U49405 ( .A(n36534), .B(n39017), .Z(n39012) );
  XOR U49406 ( .A(n36535), .B(n39012), .Z(n39010) );
  XOR U49407 ( .A(n39008), .B(n39010), .Z(n39000) );
  XOR U49408 ( .A(n38999), .B(n39000), .Z(n39003) );
  XOR U49409 ( .A(n38994), .B(n39003), .Z(n43038) );
  XOR U49410 ( .A(n38992), .B(n43038), .Z(n36541) );
  IV U49411 ( .A(n36541), .Z(n38985) );
  NOR U49412 ( .A(n36537), .B(n38985), .Z(n36536) );
  IV U49413 ( .A(n36536), .Z(n42376) );
  NOR U49414 ( .A(n36538), .B(n42376), .Z(n39600) );
  NOR U49415 ( .A(n36538), .B(n36537), .Z(n36543) );
  NOR U49416 ( .A(n36539), .B(n38986), .Z(n36540) );
  XOR U49417 ( .A(n36541), .B(n36540), .Z(n36542) );
  NOR U49418 ( .A(n36543), .B(n36542), .Z(n36544) );
  NOR U49419 ( .A(n39600), .B(n36544), .Z(n38978) );
  IV U49420 ( .A(n36545), .Z(n38980) );
  XOR U49421 ( .A(n38978), .B(n38980), .Z(n38982) );
  XOR U49422 ( .A(n38981), .B(n38982), .Z(n43065) );
  XOR U49423 ( .A(n38973), .B(n43065), .Z(n38977) );
  XOR U49424 ( .A(n38975), .B(n38977), .Z(n36549) );
  NOR U49425 ( .A(n36546), .B(n36549), .Z(n43072) );
  NOR U49426 ( .A(n43068), .B(n36547), .Z(n36551) );
  IV U49427 ( .A(n36551), .Z(n36548) );
  NOR U49428 ( .A(n36548), .B(n43065), .Z(n42370) );
  IV U49429 ( .A(n36549), .Z(n36550) );
  NOR U49430 ( .A(n36551), .B(n36550), .Z(n36552) );
  NOR U49431 ( .A(n42370), .B(n36552), .Z(n36553) );
  NOR U49432 ( .A(n36554), .B(n36553), .Z(n36555) );
  NOR U49433 ( .A(n43072), .B(n36555), .Z(n39604) );
  XOR U49434 ( .A(n39605), .B(n39604), .Z(n39607) );
  XOR U49435 ( .A(n39606), .B(n39607), .Z(n38969) );
  NOR U49436 ( .A(n36567), .B(n38969), .Z(n42362) );
  IV U49437 ( .A(n36556), .Z(n38970) );
  NOR U49438 ( .A(n38970), .B(n36557), .Z(n36558) );
  XOR U49439 ( .A(n36558), .B(n38969), .Z(n39620) );
  IV U49440 ( .A(n36559), .Z(n36566) );
  NOR U49441 ( .A(n36561), .B(n36560), .Z(n36562) );
  IV U49442 ( .A(n36562), .Z(n36563) );
  NOR U49443 ( .A(n36564), .B(n36563), .Z(n36565) );
  IV U49444 ( .A(n36565), .Z(n36575) );
  NOR U49445 ( .A(n36566), .B(n36575), .Z(n36568) );
  IV U49446 ( .A(n36568), .Z(n39619) );
  XOR U49447 ( .A(n39620), .B(n39619), .Z(n36570) );
  NOR U49448 ( .A(n36568), .B(n36567), .Z(n36569) );
  NOR U49449 ( .A(n36570), .B(n36569), .Z(n36571) );
  NOR U49450 ( .A(n42362), .B(n36571), .Z(n38966) );
  IV U49451 ( .A(n36572), .Z(n36573) );
  NOR U49452 ( .A(n36573), .B(n36582), .Z(n38965) );
  IV U49453 ( .A(n36574), .Z(n36576) );
  NOR U49454 ( .A(n36576), .B(n36575), .Z(n39614) );
  NOR U49455 ( .A(n38965), .B(n39614), .Z(n36577) );
  XOR U49456 ( .A(n38966), .B(n36577), .Z(n39628) );
  IV U49457 ( .A(n36578), .Z(n36579) );
  NOR U49458 ( .A(n36580), .B(n36579), .Z(n39626) );
  IV U49459 ( .A(n36581), .Z(n36583) );
  NOR U49460 ( .A(n36583), .B(n36582), .Z(n38963) );
  NOR U49461 ( .A(n39626), .B(n38963), .Z(n36584) );
  XOR U49462 ( .A(n39628), .B(n36584), .Z(n39629) );
  XOR U49463 ( .A(n39631), .B(n39629), .Z(n43100) );
  XOR U49464 ( .A(n38962), .B(n43100), .Z(n38956) );
  XOR U49465 ( .A(n38957), .B(n38956), .Z(n38959) );
  IV U49466 ( .A(n36585), .Z(n36589) );
  NOR U49467 ( .A(n36587), .B(n36586), .Z(n36588) );
  IV U49468 ( .A(n36588), .Z(n36595) );
  NOR U49469 ( .A(n36589), .B(n36595), .Z(n36590) );
  IV U49470 ( .A(n36590), .Z(n36598) );
  NOR U49471 ( .A(n38959), .B(n36598), .Z(n43112) );
  IV U49472 ( .A(n36591), .Z(n36592) );
  NOR U49473 ( .A(n36593), .B(n36592), .Z(n38950) );
  IV U49474 ( .A(n36594), .Z(n36596) );
  NOR U49475 ( .A(n36596), .B(n36595), .Z(n36597) );
  IV U49476 ( .A(n36597), .Z(n38960) );
  XOR U49477 ( .A(n38960), .B(n38959), .Z(n38951) );
  XOR U49478 ( .A(n38950), .B(n38951), .Z(n36600) );
  NOR U49479 ( .A(n38951), .B(n36598), .Z(n36599) );
  NOR U49480 ( .A(n36600), .B(n36599), .Z(n36601) );
  NOR U49481 ( .A(n43112), .B(n36601), .Z(n38945) );
  IV U49482 ( .A(n36602), .Z(n36604) );
  NOR U49483 ( .A(n36604), .B(n36603), .Z(n38954) );
  IV U49484 ( .A(n36605), .Z(n36607) );
  NOR U49485 ( .A(n36607), .B(n36606), .Z(n39636) );
  NOR U49486 ( .A(n38954), .B(n39636), .Z(n36608) );
  XOR U49487 ( .A(n38945), .B(n36608), .Z(n38941) );
  IV U49488 ( .A(n36609), .Z(n36611) );
  NOR U49489 ( .A(n36611), .B(n36610), .Z(n38939) );
  XOR U49490 ( .A(n38941), .B(n38939), .Z(n39646) );
  XOR U49491 ( .A(n36612), .B(n39646), .Z(n39644) );
  XOR U49492 ( .A(n39642), .B(n39644), .Z(n45458) );
  XOR U49493 ( .A(n36613), .B(n45458), .Z(n39650) );
  NOR U49494 ( .A(n36618), .B(n39650), .Z(n39653) );
  IV U49495 ( .A(n36614), .Z(n36615) );
  NOR U49496 ( .A(n36616), .B(n36615), .Z(n36617) );
  IV U49497 ( .A(n36617), .Z(n39651) );
  XOR U49498 ( .A(n39651), .B(n39650), .Z(n38932) );
  XOR U49499 ( .A(n38931), .B(n38932), .Z(n36620) );
  NOR U49500 ( .A(n38932), .B(n36618), .Z(n36619) );
  NOR U49501 ( .A(n36620), .B(n36619), .Z(n36621) );
  NOR U49502 ( .A(n39653), .B(n36621), .Z(n42321) );
  XOR U49503 ( .A(n36622), .B(n42321), .Z(n39666) );
  IV U49504 ( .A(n36623), .Z(n36624) );
  NOR U49505 ( .A(n36625), .B(n36624), .Z(n36626) );
  NOR U49506 ( .A(n39667), .B(n36626), .Z(n36627) );
  XOR U49507 ( .A(n39666), .B(n36627), .Z(n39661) );
  XOR U49508 ( .A(n36628), .B(n39661), .Z(n39674) );
  XOR U49509 ( .A(n36629), .B(n39674), .Z(n36630) );
  IV U49510 ( .A(n36630), .Z(n38908) );
  XOR U49511 ( .A(n38907), .B(n38908), .Z(n43144) );
  XOR U49512 ( .A(n39679), .B(n43144), .Z(n36631) );
  IV U49513 ( .A(n36631), .Z(n39682) );
  IV U49514 ( .A(n36632), .Z(n36634) );
  NOR U49515 ( .A(n36634), .B(n36633), .Z(n39680) );
  XOR U49516 ( .A(n39682), .B(n39680), .Z(n38905) );
  XOR U49517 ( .A(n38906), .B(n38905), .Z(n38894) );
  NOR U49518 ( .A(n36635), .B(n38899), .Z(n36639) );
  IV U49519 ( .A(n36636), .Z(n36638) );
  IV U49520 ( .A(n36637), .Z(n36643) );
  NOR U49521 ( .A(n36638), .B(n36643), .Z(n38895) );
  NOR U49522 ( .A(n36639), .B(n38895), .Z(n36640) );
  XOR U49523 ( .A(n38894), .B(n36640), .Z(n38890) );
  IV U49524 ( .A(n36641), .Z(n36642) );
  NOR U49525 ( .A(n36643), .B(n36642), .Z(n38888) );
  XOR U49526 ( .A(n38890), .B(n38888), .Z(n38892) );
  XOR U49527 ( .A(n36644), .B(n38892), .Z(n38886) );
  XOR U49528 ( .A(n38887), .B(n38886), .Z(n39688) );
  IV U49529 ( .A(n36645), .Z(n36647) );
  NOR U49530 ( .A(n36647), .B(n36646), .Z(n45423) );
  NOR U49531 ( .A(n45431), .B(n45423), .Z(n39689) );
  XOR U49532 ( .A(n39688), .B(n39689), .Z(n39692) );
  XOR U49533 ( .A(n39690), .B(n39692), .Z(n39701) );
  XOR U49534 ( .A(n39700), .B(n39701), .Z(n39695) );
  XOR U49535 ( .A(n39694), .B(n39695), .Z(n39709) );
  IV U49536 ( .A(n36648), .Z(n36650) );
  NOR U49537 ( .A(n36650), .B(n36649), .Z(n39698) );
  IV U49538 ( .A(n36651), .Z(n36653) );
  NOR U49539 ( .A(n36653), .B(n36652), .Z(n39708) );
  NOR U49540 ( .A(n39698), .B(n39708), .Z(n36654) );
  XOR U49541 ( .A(n39709), .B(n36654), .Z(n36655) );
  NOR U49542 ( .A(n36656), .B(n36655), .Z(n36659) );
  IV U49543 ( .A(n36656), .Z(n36658) );
  XOR U49544 ( .A(n39698), .B(n39709), .Z(n36657) );
  NOR U49545 ( .A(n36658), .B(n36657), .Z(n42260) );
  NOR U49546 ( .A(n36659), .B(n42260), .Z(n38878) );
  IV U49547 ( .A(n36660), .Z(n36662) );
  NOR U49548 ( .A(n36662), .B(n36661), .Z(n38880) );
  IV U49549 ( .A(n36663), .Z(n36665) );
  NOR U49550 ( .A(n36665), .B(n36664), .Z(n38877) );
  NOR U49551 ( .A(n38880), .B(n38877), .Z(n36666) );
  XOR U49552 ( .A(n38878), .B(n36666), .Z(n38875) );
  XOR U49553 ( .A(n38873), .B(n38875), .Z(n39714) );
  XOR U49554 ( .A(n39712), .B(n39714), .Z(n39719) );
  XOR U49555 ( .A(n36667), .B(n39719), .Z(n43187) );
  XOR U49556 ( .A(n36668), .B(n43187), .Z(n38863) );
  XOR U49557 ( .A(n36669), .B(n38863), .Z(n36670) );
  IV U49558 ( .A(n36670), .Z(n38855) );
  XOR U49559 ( .A(n38854), .B(n38855), .Z(n38858) );
  XOR U49560 ( .A(n36671), .B(n38858), .Z(n36672) );
  IV U49561 ( .A(n36672), .Z(n38850) );
  IV U49562 ( .A(n36673), .Z(n36675) );
  NOR U49563 ( .A(n36675), .B(n36674), .Z(n38848) );
  XOR U49564 ( .A(n38850), .B(n38848), .Z(n39725) );
  XOR U49565 ( .A(n39724), .B(n39725), .Z(n38846) );
  XOR U49566 ( .A(n38845), .B(n38846), .Z(n42228) );
  IV U49567 ( .A(n36676), .Z(n36678) );
  NOR U49568 ( .A(n36678), .B(n36677), .Z(n42226) );
  NOR U49569 ( .A(n42231), .B(n42226), .Z(n38844) );
  XOR U49570 ( .A(n42228), .B(n38844), .Z(n38838) );
  XOR U49571 ( .A(n36679), .B(n38838), .Z(n39743) );
  XOR U49572 ( .A(n36680), .B(n39743), .Z(n38832) );
  XOR U49573 ( .A(n38830), .B(n38832), .Z(n42211) );
  IV U49574 ( .A(n36681), .Z(n36686) );
  IV U49575 ( .A(n36682), .Z(n36683) );
  NOR U49576 ( .A(n36686), .B(n36683), .Z(n42205) );
  IV U49577 ( .A(n36684), .Z(n36685) );
  NOR U49578 ( .A(n36686), .B(n36685), .Z(n42210) );
  NOR U49579 ( .A(n42205), .B(n42210), .Z(n38829) );
  XOR U49580 ( .A(n42211), .B(n38829), .Z(n39748) );
  XOR U49581 ( .A(n36687), .B(n39748), .Z(n43224) );
  XOR U49582 ( .A(n38825), .B(n43224), .Z(n36688) );
  NOR U49583 ( .A(n36689), .B(n36688), .Z(n36694) );
  IV U49584 ( .A(n36689), .Z(n36690) );
  NOR U49585 ( .A(n43224), .B(n36690), .Z(n46423) );
  NOR U49586 ( .A(n36694), .B(n46423), .Z(n36691) );
  NOR U49587 ( .A(n36692), .B(n36691), .Z(n36695) );
  IV U49588 ( .A(n36692), .Z(n36693) );
  NOR U49589 ( .A(n36694), .B(n36693), .Z(n46410) );
  NOR U49590 ( .A(n36695), .B(n46410), .Z(n36702) );
  IV U49591 ( .A(n36702), .Z(n38820) );
  NOR U49592 ( .A(n36703), .B(n38820), .Z(n43243) );
  IV U49593 ( .A(n36696), .Z(n36701) );
  IV U49594 ( .A(n36697), .Z(n36698) );
  NOR U49595 ( .A(n36701), .B(n36698), .Z(n38821) );
  IV U49596 ( .A(n36699), .Z(n36700) );
  NOR U49597 ( .A(n36701), .B(n36700), .Z(n38818) );
  XOR U49598 ( .A(n36702), .B(n38818), .Z(n38822) );
  XOR U49599 ( .A(n38821), .B(n38822), .Z(n36705) );
  NOR U49600 ( .A(n38822), .B(n36703), .Z(n36704) );
  NOR U49601 ( .A(n36705), .B(n36704), .Z(n36706) );
  NOR U49602 ( .A(n43243), .B(n36706), .Z(n39752) );
  IV U49603 ( .A(n36707), .Z(n36708) );
  NOR U49604 ( .A(n36709), .B(n36708), .Z(n36710) );
  IV U49605 ( .A(n36710), .Z(n39754) );
  XOR U49606 ( .A(n39752), .B(n39754), .Z(n39758) );
  XOR U49607 ( .A(n39756), .B(n39758), .Z(n39761) );
  XOR U49608 ( .A(n39759), .B(n39761), .Z(n38813) );
  XOR U49609 ( .A(n38812), .B(n38813), .Z(n38816) );
  XOR U49610 ( .A(n36711), .B(n38816), .Z(n36712) );
  IV U49611 ( .A(n36712), .Z(n38811) );
  IV U49612 ( .A(n36713), .Z(n36717) );
  XOR U49613 ( .A(n36715), .B(n36714), .Z(n36716) );
  NOR U49614 ( .A(n36717), .B(n36716), .Z(n38809) );
  XOR U49615 ( .A(n38811), .B(n38809), .Z(n39766) );
  IV U49616 ( .A(n36718), .Z(n36719) );
  NOR U49617 ( .A(n36720), .B(n36719), .Z(n38805) );
  IV U49618 ( .A(n36721), .Z(n36723) );
  NOR U49619 ( .A(n36723), .B(n36722), .Z(n39765) );
  NOR U49620 ( .A(n38805), .B(n39765), .Z(n36724) );
  XOR U49621 ( .A(n39766), .B(n36724), .Z(n38801) );
  IV U49622 ( .A(n36725), .Z(n36727) );
  NOR U49623 ( .A(n36727), .B(n36726), .Z(n38802) );
  IV U49624 ( .A(n36728), .Z(n36729) );
  NOR U49625 ( .A(n36732), .B(n36729), .Z(n39771) );
  NOR U49626 ( .A(n38802), .B(n39771), .Z(n36730) );
  XOR U49627 ( .A(n38801), .B(n36730), .Z(n39770) );
  IV U49628 ( .A(n36731), .Z(n36733) );
  NOR U49629 ( .A(n36733), .B(n36732), .Z(n39768) );
  XOR U49630 ( .A(n39770), .B(n39768), .Z(n38799) );
  IV U49631 ( .A(n36734), .Z(n36739) );
  IV U49632 ( .A(n36735), .Z(n36736) );
  NOR U49633 ( .A(n36739), .B(n36736), .Z(n38797) );
  XOR U49634 ( .A(n38799), .B(n38797), .Z(n39779) );
  IV U49635 ( .A(n36737), .Z(n36738) );
  NOR U49636 ( .A(n36739), .B(n36738), .Z(n39777) );
  XOR U49637 ( .A(n39779), .B(n39777), .Z(n39781) );
  XOR U49638 ( .A(n39780), .B(n39781), .Z(n39787) );
  IV U49639 ( .A(n36740), .Z(n36741) );
  NOR U49640 ( .A(n36741), .B(n36743), .Z(n39775) );
  IV U49641 ( .A(n36742), .Z(n36749) );
  NOR U49642 ( .A(n36744), .B(n36743), .Z(n36745) );
  IV U49643 ( .A(n36745), .Z(n36746) );
  NOR U49644 ( .A(n36747), .B(n36746), .Z(n36748) );
  IV U49645 ( .A(n36748), .Z(n36755) );
  NOR U49646 ( .A(n36749), .B(n36755), .Z(n39785) );
  NOR U49647 ( .A(n39775), .B(n39785), .Z(n36750) );
  XOR U49648 ( .A(n39787), .B(n36750), .Z(n38794) );
  IV U49649 ( .A(n36751), .Z(n36753) );
  NOR U49650 ( .A(n36753), .B(n36752), .Z(n39788) );
  IV U49651 ( .A(n36754), .Z(n36756) );
  NOR U49652 ( .A(n36756), .B(n36755), .Z(n38795) );
  NOR U49653 ( .A(n39788), .B(n38795), .Z(n36757) );
  XOR U49654 ( .A(n38794), .B(n36757), .Z(n39792) );
  XOR U49655 ( .A(n39791), .B(n39792), .Z(n42160) );
  XOR U49656 ( .A(n38790), .B(n42160), .Z(n36765) );
  NOR U49657 ( .A(n36759), .B(n36758), .Z(n42155) );
  IV U49658 ( .A(n36760), .Z(n36767) );
  IV U49659 ( .A(n36761), .Z(n36762) );
  NOR U49660 ( .A(n36767), .B(n36762), .Z(n42149) );
  NOR U49661 ( .A(n42155), .B(n42149), .Z(n38791) );
  XOR U49662 ( .A(n36765), .B(n38791), .Z(n36763) );
  NOR U49663 ( .A(n36764), .B(n36763), .Z(n42144) );
  IV U49664 ( .A(n36765), .Z(n42151) );
  IV U49665 ( .A(n36766), .Z(n36768) );
  NOR U49666 ( .A(n36768), .B(n36767), .Z(n38788) );
  IV U49667 ( .A(n38791), .Z(n36769) );
  NOR U49668 ( .A(n38788), .B(n36769), .Z(n36770) );
  XOR U49669 ( .A(n42151), .B(n36770), .Z(n36775) );
  NOR U49670 ( .A(n36771), .B(n36775), .Z(n36772) );
  NOR U49671 ( .A(n42144), .B(n36772), .Z(n36773) );
  NOR U49672 ( .A(n36774), .B(n36773), .Z(n36778) );
  IV U49673 ( .A(n36774), .Z(n36777) );
  IV U49674 ( .A(n36775), .Z(n36776) );
  NOR U49675 ( .A(n36777), .B(n36776), .Z(n42141) );
  NOR U49676 ( .A(n36778), .B(n42141), .Z(n36783) );
  IV U49677 ( .A(n36783), .Z(n38786) );
  NOR U49678 ( .A(n36792), .B(n38786), .Z(n43273) );
  IV U49679 ( .A(n36779), .Z(n36780) );
  NOR U49680 ( .A(n36781), .B(n36780), .Z(n36782) );
  IV U49681 ( .A(n36782), .Z(n38787) );
  XOR U49682 ( .A(n38787), .B(n36783), .Z(n38785) );
  IV U49683 ( .A(n36784), .Z(n36791) );
  NOR U49684 ( .A(n36786), .B(n36785), .Z(n36787) );
  IV U49685 ( .A(n36787), .Z(n36788) );
  NOR U49686 ( .A(n36789), .B(n36788), .Z(n36790) );
  IV U49687 ( .A(n36790), .Z(n36799) );
  NOR U49688 ( .A(n36791), .B(n36799), .Z(n36793) );
  IV U49689 ( .A(n36793), .Z(n38784) );
  XOR U49690 ( .A(n38785), .B(n38784), .Z(n36795) );
  NOR U49691 ( .A(n36793), .B(n36792), .Z(n36794) );
  NOR U49692 ( .A(n36795), .B(n36794), .Z(n36796) );
  NOR U49693 ( .A(n43273), .B(n36796), .Z(n38780) );
  NOR U49694 ( .A(n36797), .B(n38781), .Z(n36801) );
  IV U49695 ( .A(n36798), .Z(n36800) );
  NOR U49696 ( .A(n36800), .B(n36799), .Z(n39801) );
  NOR U49697 ( .A(n36801), .B(n39801), .Z(n36802) );
  XOR U49698 ( .A(n38780), .B(n36802), .Z(n39817) );
  XOR U49699 ( .A(n39815), .B(n39817), .Z(n39813) );
  XOR U49700 ( .A(n39812), .B(n39813), .Z(n38774) );
  XOR U49701 ( .A(n38773), .B(n38774), .Z(n38778) );
  XOR U49702 ( .A(n38776), .B(n38778), .Z(n43294) );
  XOR U49703 ( .A(n38771), .B(n43294), .Z(n38766) );
  XOR U49704 ( .A(n38765), .B(n38766), .Z(n38769) );
  XOR U49705 ( .A(n36803), .B(n38769), .Z(n38758) );
  IV U49706 ( .A(n36804), .Z(n36805) );
  NOR U49707 ( .A(n36806), .B(n36805), .Z(n38762) );
  IV U49708 ( .A(n36807), .Z(n36809) );
  NOR U49709 ( .A(n36809), .B(n36808), .Z(n38757) );
  NOR U49710 ( .A(n38762), .B(n38757), .Z(n36810) );
  XOR U49711 ( .A(n38758), .B(n36810), .Z(n38756) );
  IV U49712 ( .A(n38756), .Z(n36820) );
  IV U49713 ( .A(n36811), .Z(n36813) );
  NOR U49714 ( .A(n36813), .B(n36812), .Z(n38754) );
  IV U49715 ( .A(n36814), .Z(n36818) );
  NOR U49716 ( .A(n36816), .B(n36815), .Z(n36817) );
  IV U49717 ( .A(n36817), .Z(n36825) );
  NOR U49718 ( .A(n36818), .B(n36825), .Z(n38751) );
  NOR U49719 ( .A(n38754), .B(n38751), .Z(n36819) );
  XOR U49720 ( .A(n36820), .B(n36819), .Z(n39825) );
  IV U49721 ( .A(n36821), .Z(n36822) );
  NOR U49722 ( .A(n36823), .B(n36822), .Z(n36824) );
  IV U49723 ( .A(n36824), .Z(n36826) );
  NOR U49724 ( .A(n36826), .B(n36825), .Z(n36827) );
  IV U49725 ( .A(n36827), .Z(n39824) );
  XOR U49726 ( .A(n39825), .B(n39824), .Z(n38748) );
  IV U49727 ( .A(n36828), .Z(n36829) );
  NOR U49728 ( .A(n36830), .B(n36829), .Z(n39826) );
  IV U49729 ( .A(n36831), .Z(n36832) );
  NOR U49730 ( .A(n36832), .B(n36836), .Z(n38749) );
  NOR U49731 ( .A(n39826), .B(n38749), .Z(n36833) );
  XOR U49732 ( .A(n38748), .B(n36833), .Z(n38747) );
  IV U49733 ( .A(n36834), .Z(n36835) );
  NOR U49734 ( .A(n36836), .B(n36835), .Z(n38745) );
  XOR U49735 ( .A(n38747), .B(n38745), .Z(n38739) );
  XOR U49736 ( .A(n38738), .B(n38739), .Z(n38742) );
  XOR U49737 ( .A(n38741), .B(n38742), .Z(n38735) );
  XOR U49738 ( .A(n38734), .B(n38735), .Z(n39833) );
  XOR U49739 ( .A(n39831), .B(n39833), .Z(n43333) );
  IV U49740 ( .A(n36837), .Z(n39835) );
  NOR U49741 ( .A(n39835), .B(n36838), .Z(n36843) );
  NOR U49742 ( .A(n36840), .B(n36839), .Z(n43332) );
  NOR U49743 ( .A(n43332), .B(n36841), .Z(n38732) );
  IV U49744 ( .A(n38732), .Z(n36842) );
  NOR U49745 ( .A(n36843), .B(n36842), .Z(n36844) );
  XOR U49746 ( .A(n43333), .B(n36844), .Z(n38728) );
  XOR U49747 ( .A(n38729), .B(n38728), .Z(n38726) );
  IV U49748 ( .A(n36845), .Z(n36846) );
  NOR U49749 ( .A(n36846), .B(n36851), .Z(n39852) );
  IV U49750 ( .A(n36847), .Z(n36848) );
  NOR U49751 ( .A(n36849), .B(n36848), .Z(n39843) );
  IV U49752 ( .A(n36850), .Z(n36852) );
  NOR U49753 ( .A(n36852), .B(n36851), .Z(n38725) );
  NOR U49754 ( .A(n39843), .B(n38725), .Z(n36853) );
  IV U49755 ( .A(n36853), .Z(n36854) );
  NOR U49756 ( .A(n39852), .B(n36854), .Z(n36855) );
  XOR U49757 ( .A(n38726), .B(n36855), .Z(n42086) );
  IV U49758 ( .A(n36856), .Z(n36858) );
  NOR U49759 ( .A(n36858), .B(n36857), .Z(n38723) );
  NOR U49760 ( .A(n38724), .B(n38723), .Z(n36859) );
  XOR U49761 ( .A(n42086), .B(n36859), .Z(n36860) );
  NOR U49762 ( .A(n36861), .B(n36860), .Z(n36864) );
  IV U49763 ( .A(n36861), .Z(n36863) );
  XOR U49764 ( .A(n38724), .B(n42086), .Z(n36862) );
  NOR U49765 ( .A(n36863), .B(n36862), .Z(n42082) );
  NOR U49766 ( .A(n36864), .B(n42082), .Z(n38720) );
  XOR U49767 ( .A(n38721), .B(n38720), .Z(n39859) );
  XOR U49768 ( .A(n39858), .B(n39859), .Z(n38718) );
  IV U49769 ( .A(n36865), .Z(n36867) );
  NOR U49770 ( .A(n36867), .B(n36866), .Z(n38716) );
  XOR U49771 ( .A(n38718), .B(n38716), .Z(n39870) );
  IV U49772 ( .A(n36868), .Z(n36869) );
  NOR U49773 ( .A(n36870), .B(n36869), .Z(n39869) );
  IV U49774 ( .A(n36871), .Z(n36872) );
  NOR U49775 ( .A(n36873), .B(n36872), .Z(n39856) );
  NOR U49776 ( .A(n39869), .B(n39856), .Z(n36874) );
  XOR U49777 ( .A(n39870), .B(n36874), .Z(n38710) );
  IV U49778 ( .A(n36875), .Z(n36876) );
  NOR U49779 ( .A(n36877), .B(n36876), .Z(n39866) );
  IV U49780 ( .A(n36878), .Z(n36879) );
  NOR U49781 ( .A(n36880), .B(n36879), .Z(n38711) );
  NOR U49782 ( .A(n39866), .B(n38711), .Z(n36881) );
  XOR U49783 ( .A(n38710), .B(n36881), .Z(n38714) );
  XOR U49784 ( .A(n38713), .B(n38714), .Z(n38706) );
  XOR U49785 ( .A(n38705), .B(n38706), .Z(n38708) );
  XOR U49786 ( .A(n38709), .B(n38708), .Z(n39879) );
  XOR U49787 ( .A(n39878), .B(n39879), .Z(n39890) );
  IV U49788 ( .A(n36882), .Z(n36883) );
  NOR U49789 ( .A(n36884), .B(n36883), .Z(n39889) );
  IV U49790 ( .A(n36885), .Z(n36887) );
  NOR U49791 ( .A(n36887), .B(n36886), .Z(n38704) );
  NOR U49792 ( .A(n39889), .B(n38704), .Z(n36888) );
  XOR U49793 ( .A(n39890), .B(n36888), .Z(n36899) );
  IV U49794 ( .A(n36899), .Z(n38703) );
  IV U49795 ( .A(n36889), .Z(n36891) );
  NOR U49796 ( .A(n36891), .B(n36890), .Z(n36892) );
  IV U49797 ( .A(n36892), .Z(n36900) );
  NOR U49798 ( .A(n38703), .B(n36900), .Z(n42048) );
  IV U49799 ( .A(n36893), .Z(n36895) );
  NOR U49800 ( .A(n36895), .B(n36894), .Z(n39894) );
  IV U49801 ( .A(n36896), .Z(n36897) );
  NOR U49802 ( .A(n36898), .B(n36897), .Z(n38701) );
  XOR U49803 ( .A(n38701), .B(n36899), .Z(n39895) );
  XOR U49804 ( .A(n39894), .B(n39895), .Z(n36902) );
  NOR U49805 ( .A(n39895), .B(n36900), .Z(n36901) );
  NOR U49806 ( .A(n36902), .B(n36901), .Z(n36903) );
  NOR U49807 ( .A(n42048), .B(n36903), .Z(n39899) );
  XOR U49808 ( .A(n36904), .B(n39899), .Z(n46558) );
  XOR U49809 ( .A(n39907), .B(n46558), .Z(n36905) );
  IV U49810 ( .A(n36905), .Z(n38698) );
  XOR U49811 ( .A(n38697), .B(n38698), .Z(n39914) );
  XOR U49812 ( .A(n36906), .B(n39914), .Z(n38695) );
  XOR U49813 ( .A(n38694), .B(n38695), .Z(n38688) );
  XOR U49814 ( .A(n38689), .B(n38688), .Z(n38686) );
  IV U49815 ( .A(n36907), .Z(n36908) );
  NOR U49816 ( .A(n36909), .B(n36908), .Z(n38685) );
  IV U49817 ( .A(n36910), .Z(n36913) );
  IV U49818 ( .A(n36911), .Z(n36912) );
  NOR U49819 ( .A(n36913), .B(n36912), .Z(n38690) );
  NOR U49820 ( .A(n38685), .B(n38690), .Z(n36914) );
  XOR U49821 ( .A(n38686), .B(n36914), .Z(n39920) );
  XOR U49822 ( .A(n39918), .B(n39920), .Z(n39922) );
  XOR U49823 ( .A(n39921), .B(n39922), .Z(n38681) );
  XOR U49824 ( .A(n38679), .B(n38681), .Z(n38683) );
  XOR U49825 ( .A(n38682), .B(n38683), .Z(n38675) );
  XOR U49826 ( .A(n38673), .B(n38675), .Z(n38677) );
  XOR U49827 ( .A(n36915), .B(n38677), .Z(n39928) );
  IV U49828 ( .A(n36916), .Z(n36918) );
  NOR U49829 ( .A(n36918), .B(n36917), .Z(n43391) );
  NOR U49830 ( .A(n42023), .B(n43391), .Z(n39929) );
  XOR U49831 ( .A(n39928), .B(n39929), .Z(n39931) );
  XOR U49832 ( .A(n36919), .B(n39931), .Z(n39936) );
  XOR U49833 ( .A(n36920), .B(n39936), .Z(n39949) );
  XOR U49834 ( .A(n39948), .B(n39949), .Z(n39958) );
  XOR U49835 ( .A(n36921), .B(n39958), .Z(n39954) );
  XOR U49836 ( .A(n36922), .B(n39954), .Z(n39967) );
  XOR U49837 ( .A(n36923), .B(n39967), .Z(n42002) );
  XOR U49838 ( .A(n39964), .B(n42002), .Z(n39970) );
  XOR U49839 ( .A(n39971), .B(n39970), .Z(n36924) );
  IV U49840 ( .A(n36924), .Z(n39973) );
  XOR U49841 ( .A(n39972), .B(n39973), .Z(n39977) );
  XOR U49842 ( .A(n39976), .B(n39977), .Z(n39979) );
  NOR U49843 ( .A(n36925), .B(n39979), .Z(n36926) );
  IV U49844 ( .A(n36926), .Z(n36927) );
  NOR U49845 ( .A(n36928), .B(n36927), .Z(n41982) );
  NOR U49846 ( .A(n36928), .B(n36931), .Z(n36934) );
  IV U49847 ( .A(n36929), .Z(n36930) );
  NOR U49848 ( .A(n36931), .B(n36930), .Z(n36932) );
  IV U49849 ( .A(n36932), .Z(n39980) );
  XOR U49850 ( .A(n39980), .B(n39979), .Z(n36933) );
  NOR U49851 ( .A(n36934), .B(n36933), .Z(n36935) );
  NOR U49852 ( .A(n41982), .B(n36935), .Z(n39982) );
  XOR U49853 ( .A(n39984), .B(n39982), .Z(n41976) );
  IV U49854 ( .A(n36936), .Z(n36938) );
  NOR U49855 ( .A(n36938), .B(n36937), .Z(n41975) );
  IV U49856 ( .A(n36939), .Z(n36941) );
  NOR U49857 ( .A(n36941), .B(n36940), .Z(n43430) );
  NOR U49858 ( .A(n41975), .B(n43430), .Z(n39986) );
  XOR U49859 ( .A(n41976), .B(n39986), .Z(n39988) );
  XOR U49860 ( .A(n36942), .B(n39988), .Z(n40001) );
  XOR U49861 ( .A(n36943), .B(n40001), .Z(n36944) );
  IV U49862 ( .A(n36944), .Z(n40004) );
  XOR U49863 ( .A(n39997), .B(n40004), .Z(n36945) );
  NOR U49864 ( .A(n36946), .B(n36945), .Z(n41968) );
  IV U49865 ( .A(n36947), .Z(n36948) );
  NOR U49866 ( .A(n36949), .B(n36948), .Z(n40003) );
  NOR U49867 ( .A(n40003), .B(n39997), .Z(n36950) );
  XOR U49868 ( .A(n36950), .B(n40004), .Z(n36955) );
  NOR U49869 ( .A(n36951), .B(n36955), .Z(n36952) );
  NOR U49870 ( .A(n41968), .B(n36952), .Z(n36953) );
  NOR U49871 ( .A(n36954), .B(n36953), .Z(n36958) );
  IV U49872 ( .A(n36954), .Z(n36957) );
  IV U49873 ( .A(n36955), .Z(n36956) );
  NOR U49874 ( .A(n36957), .B(n36956), .Z(n46645) );
  NOR U49875 ( .A(n36958), .B(n46645), .Z(n40007) );
  IV U49876 ( .A(n36959), .Z(n36961) );
  NOR U49877 ( .A(n36961), .B(n36960), .Z(n36962) );
  IV U49878 ( .A(n36962), .Z(n40009) );
  XOR U49879 ( .A(n40007), .B(n40009), .Z(n38668) );
  XOR U49880 ( .A(n38666), .B(n38668), .Z(n40018) );
  XOR U49881 ( .A(n36963), .B(n40018), .Z(n38665) );
  XOR U49882 ( .A(n38663), .B(n38665), .Z(n41964) );
  XOR U49883 ( .A(n38660), .B(n41964), .Z(n38661) );
  XOR U49884 ( .A(n38662), .B(n38661), .Z(n40027) );
  XOR U49885 ( .A(n40029), .B(n40027), .Z(n36964) );
  IV U49886 ( .A(n36964), .Z(n40033) );
  XOR U49887 ( .A(n40032), .B(n40033), .Z(n40036) );
  XOR U49888 ( .A(n40035), .B(n40036), .Z(n36965) );
  NOR U49889 ( .A(n36966), .B(n36965), .Z(n41928) );
  IV U49890 ( .A(n36967), .Z(n36969) );
  NOR U49891 ( .A(n36969), .B(n36968), .Z(n38658) );
  XOR U49892 ( .A(n40032), .B(n40035), .Z(n36970) );
  NOR U49893 ( .A(n38658), .B(n36970), .Z(n36971) );
  XOR U49894 ( .A(n36971), .B(n40033), .Z(n36972) );
  NOR U49895 ( .A(n36973), .B(n36972), .Z(n36974) );
  NOR U49896 ( .A(n41928), .B(n36974), .Z(n38656) );
  NOR U49897 ( .A(n36976), .B(n36975), .Z(n45150) );
  IV U49898 ( .A(n36977), .Z(n36979) );
  NOR U49899 ( .A(n36979), .B(n36978), .Z(n45140) );
  NOR U49900 ( .A(n45150), .B(n45140), .Z(n38657) );
  XOR U49901 ( .A(n38656), .B(n38657), .Z(n38652) );
  XOR U49902 ( .A(n38650), .B(n38652), .Z(n38654) );
  XOR U49903 ( .A(n38653), .B(n38654), .Z(n38645) );
  XOR U49904 ( .A(n38644), .B(n38645), .Z(n38649) );
  XOR U49905 ( .A(n38647), .B(n38649), .Z(n38638) );
  XOR U49906 ( .A(n38637), .B(n38638), .Z(n38641) );
  XOR U49907 ( .A(n38640), .B(n38641), .Z(n38634) );
  XOR U49908 ( .A(n38633), .B(n38634), .Z(n40045) );
  XOR U49909 ( .A(n40047), .B(n40045), .Z(n38632) );
  IV U49910 ( .A(n36980), .Z(n41919) );
  NOR U49911 ( .A(n41919), .B(n36981), .Z(n40048) );
  IV U49912 ( .A(n36982), .Z(n36984) );
  NOR U49913 ( .A(n36984), .B(n36983), .Z(n38630) );
  NOR U49914 ( .A(n40048), .B(n38630), .Z(n36985) );
  XOR U49915 ( .A(n38632), .B(n36985), .Z(n38622) );
  XOR U49916 ( .A(n38623), .B(n38622), .Z(n38620) );
  IV U49917 ( .A(n36986), .Z(n36988) );
  NOR U49918 ( .A(n36988), .B(n36987), .Z(n38619) );
  NOR U49919 ( .A(n38626), .B(n38619), .Z(n36989) );
  XOR U49920 ( .A(n38620), .B(n36989), .Z(n40054) );
  XOR U49921 ( .A(n40053), .B(n40054), .Z(n40057) );
  XOR U49922 ( .A(n40056), .B(n40057), .Z(n40063) );
  XOR U49923 ( .A(n40062), .B(n40063), .Z(n40074) );
  XOR U49924 ( .A(n36990), .B(n40074), .Z(n43490) );
  XOR U49925 ( .A(n41900), .B(n43490), .Z(n40081) );
  IV U49926 ( .A(n36991), .Z(n36993) );
  NOR U49927 ( .A(n36993), .B(n36992), .Z(n43488) );
  IV U49928 ( .A(n36994), .Z(n36995) );
  NOR U49929 ( .A(n36996), .B(n36995), .Z(n40080) );
  NOR U49930 ( .A(n43488), .B(n40080), .Z(n36997) );
  XOR U49931 ( .A(n40081), .B(n36997), .Z(n40086) );
  NOR U49932 ( .A(n36999), .B(n36998), .Z(n40084) );
  XOR U49933 ( .A(n40086), .B(n40084), .Z(n40088) );
  XOR U49934 ( .A(n40087), .B(n40088), .Z(n40101) );
  XOR U49935 ( .A(n40099), .B(n40101), .Z(n40095) );
  XOR U49936 ( .A(n37000), .B(n40095), .Z(n40113) );
  XOR U49937 ( .A(n40111), .B(n40113), .Z(n40114) );
  XOR U49938 ( .A(n40115), .B(n40114), .Z(n38614) );
  IV U49939 ( .A(n37001), .Z(n37002) );
  NOR U49940 ( .A(n37002), .B(n37007), .Z(n40120) );
  IV U49941 ( .A(n37003), .Z(n37004) );
  NOR U49942 ( .A(n37005), .B(n37004), .Z(n45087) );
  IV U49943 ( .A(n37006), .Z(n37008) );
  NOR U49944 ( .A(n37008), .B(n37007), .Z(n45077) );
  NOR U49945 ( .A(n45087), .B(n45077), .Z(n38615) );
  IV U49946 ( .A(n38615), .Z(n37009) );
  NOR U49947 ( .A(n40120), .B(n37009), .Z(n37010) );
  XOR U49948 ( .A(n38614), .B(n37010), .Z(n40119) );
  IV U49949 ( .A(n37011), .Z(n37012) );
  NOR U49950 ( .A(n37013), .B(n37012), .Z(n40117) );
  XOR U49951 ( .A(n40119), .B(n40117), .Z(n38610) );
  XOR U49952 ( .A(n38608), .B(n38610), .Z(n38613) );
  XOR U49953 ( .A(n38611), .B(n38613), .Z(n41877) );
  XOR U49954 ( .A(n37014), .B(n41877), .Z(n38602) );
  XOR U49955 ( .A(n38601), .B(n38602), .Z(n38605) );
  XOR U49956 ( .A(n38604), .B(n38605), .Z(n38597) );
  IV U49957 ( .A(n37015), .Z(n37017) );
  NOR U49958 ( .A(n37017), .B(n37016), .Z(n38595) );
  XOR U49959 ( .A(n38597), .B(n38595), .Z(n40128) );
  IV U49960 ( .A(n37018), .Z(n37019) );
  NOR U49961 ( .A(n38589), .B(n37019), .Z(n37022) );
  IV U49962 ( .A(n37020), .Z(n37021) );
  NOR U49963 ( .A(n37025), .B(n37021), .Z(n40127) );
  NOR U49964 ( .A(n37022), .B(n40127), .Z(n37023) );
  XOR U49965 ( .A(n40128), .B(n37023), .Z(n38581) );
  IV U49966 ( .A(n37024), .Z(n37026) );
  NOR U49967 ( .A(n37026), .B(n37025), .Z(n38585) );
  IV U49968 ( .A(n37027), .Z(n37029) );
  NOR U49969 ( .A(n37029), .B(n37028), .Z(n38582) );
  NOR U49970 ( .A(n38585), .B(n38582), .Z(n37030) );
  XOR U49971 ( .A(n38581), .B(n37030), .Z(n40133) );
  IV U49972 ( .A(n37031), .Z(n37033) );
  NOR U49973 ( .A(n37033), .B(n37032), .Z(n40130) );
  NOR U49974 ( .A(n37034), .B(n40134), .Z(n37035) );
  NOR U49975 ( .A(n40130), .B(n37035), .Z(n37036) );
  XOR U49976 ( .A(n40133), .B(n37036), .Z(n37037) );
  IV U49977 ( .A(n37037), .Z(n38580) );
  IV U49978 ( .A(n37038), .Z(n37040) );
  NOR U49979 ( .A(n37040), .B(n37039), .Z(n38578) );
  XOR U49980 ( .A(n38580), .B(n38578), .Z(n38573) );
  XOR U49981 ( .A(n38572), .B(n38573), .Z(n38576) );
  NOR U49982 ( .A(n37048), .B(n38576), .Z(n41854) );
  IV U49983 ( .A(n37041), .Z(n37042) );
  NOR U49984 ( .A(n37043), .B(n37042), .Z(n38566) );
  IV U49985 ( .A(n37044), .Z(n37046) );
  NOR U49986 ( .A(n37046), .B(n37045), .Z(n38575) );
  NOR U49987 ( .A(n38575), .B(n38570), .Z(n37047) );
  XOR U49988 ( .A(n37047), .B(n38576), .Z(n38567) );
  XOR U49989 ( .A(n38566), .B(n38567), .Z(n37050) );
  NOR U49990 ( .A(n38567), .B(n37048), .Z(n37049) );
  NOR U49991 ( .A(n37050), .B(n37049), .Z(n37051) );
  NOR U49992 ( .A(n41854), .B(n37051), .Z(n38560) );
  IV U49993 ( .A(n37052), .Z(n37054) );
  NOR U49994 ( .A(n37054), .B(n37053), .Z(n37055) );
  IV U49995 ( .A(n37055), .Z(n38562) );
  XOR U49996 ( .A(n38560), .B(n38562), .Z(n43556) );
  XOR U49997 ( .A(n38563), .B(n43556), .Z(n38558) );
  XOR U49998 ( .A(n38559), .B(n38558), .Z(n43571) );
  XOR U49999 ( .A(n38553), .B(n43571), .Z(n38551) );
  IV U50000 ( .A(n37056), .Z(n37057) );
  NOR U50001 ( .A(n37058), .B(n37057), .Z(n38554) );
  IV U50002 ( .A(n37059), .Z(n37061) );
  NOR U50003 ( .A(n37061), .B(n37060), .Z(n38550) );
  NOR U50004 ( .A(n38554), .B(n38550), .Z(n37062) );
  XOR U50005 ( .A(n38551), .B(n37062), .Z(n38548) );
  NOR U50006 ( .A(n37064), .B(n37063), .Z(n38547) );
  IV U50007 ( .A(n37065), .Z(n38541) );
  NOR U50008 ( .A(n37066), .B(n38541), .Z(n37067) );
  NOR U50009 ( .A(n38547), .B(n37067), .Z(n37068) );
  XOR U50010 ( .A(n38548), .B(n37068), .Z(n40150) );
  XOR U50011 ( .A(n40151), .B(n40150), .Z(n38537) );
  XOR U50012 ( .A(n38536), .B(n38537), .Z(n40149) );
  XOR U50013 ( .A(n40147), .B(n40149), .Z(n40159) );
  XOR U50014 ( .A(n37069), .B(n40159), .Z(n38534) );
  IV U50015 ( .A(n37073), .Z(n37071) );
  IV U50016 ( .A(n37070), .Z(n37072) );
  NOR U50017 ( .A(n37071), .B(n37072), .Z(n38533) );
  XOR U50018 ( .A(n37073), .B(n37072), .Z(n37076) );
  IV U50019 ( .A(n37074), .Z(n37075) );
  NOR U50020 ( .A(n37076), .B(n37075), .Z(n40165) );
  NOR U50021 ( .A(n38533), .B(n40165), .Z(n37077) );
  XOR U50022 ( .A(n38534), .B(n37077), .Z(n40164) );
  XOR U50023 ( .A(n40162), .B(n40164), .Z(n38527) );
  XOR U50024 ( .A(n37078), .B(n38527), .Z(n38511) );
  XOR U50025 ( .A(n37079), .B(n38511), .Z(n38506) );
  XOR U50026 ( .A(n38504), .B(n38506), .Z(n38508) );
  XOR U50027 ( .A(n38507), .B(n38508), .Z(n40171) );
  IV U50028 ( .A(n37080), .Z(n37082) );
  NOR U50029 ( .A(n37082), .B(n37081), .Z(n40170) );
  IV U50030 ( .A(n37083), .Z(n37084) );
  NOR U50031 ( .A(n37085), .B(n37084), .Z(n38502) );
  NOR U50032 ( .A(n40170), .B(n38502), .Z(n37086) );
  XOR U50033 ( .A(n40171), .B(n37086), .Z(n38499) );
  XOR U50034 ( .A(n37087), .B(n38499), .Z(n40177) );
  XOR U50035 ( .A(n40176), .B(n40177), .Z(n37088) );
  NOR U50036 ( .A(n37089), .B(n37088), .Z(n41789) );
  IV U50037 ( .A(n37090), .Z(n37092) );
  NOR U50038 ( .A(n37092), .B(n37091), .Z(n38497) );
  NOR U50039 ( .A(n40176), .B(n38497), .Z(n37093) );
  XOR U50040 ( .A(n37093), .B(n40177), .Z(n37109) );
  NOR U50041 ( .A(n37094), .B(n37109), .Z(n37095) );
  NOR U50042 ( .A(n41789), .B(n37095), .Z(n37105) );
  IV U50043 ( .A(n37096), .Z(n37097) );
  NOR U50044 ( .A(n37098), .B(n37097), .Z(n37108) );
  IV U50045 ( .A(n37099), .Z(n37100) );
  NOR U50046 ( .A(n37101), .B(n37100), .Z(n37104) );
  NOR U50047 ( .A(n37108), .B(n37104), .Z(n37102) );
  IV U50048 ( .A(n37102), .Z(n37103) );
  NOR U50049 ( .A(n37105), .B(n37103), .Z(n37113) );
  IV U50050 ( .A(n37104), .Z(n37107) );
  IV U50051 ( .A(n37105), .Z(n37106) );
  NOR U50052 ( .A(n37107), .B(n37106), .Z(n41784) );
  IV U50053 ( .A(n37108), .Z(n37111) );
  IV U50054 ( .A(n37109), .Z(n37110) );
  NOR U50055 ( .A(n37111), .B(n37110), .Z(n41786) );
  NOR U50056 ( .A(n41784), .B(n41786), .Z(n37112) );
  IV U50057 ( .A(n37112), .Z(n38496) );
  NOR U50058 ( .A(n37113), .B(n38496), .Z(n38493) );
  IV U50059 ( .A(n37114), .Z(n37116) );
  NOR U50060 ( .A(n37116), .B(n37115), .Z(n37117) );
  IV U50061 ( .A(n37117), .Z(n38495) );
  XOR U50062 ( .A(n38493), .B(n38495), .Z(n38488) );
  XOR U50063 ( .A(n38487), .B(n38488), .Z(n38491) );
  XOR U50064 ( .A(n37118), .B(n38491), .Z(n38478) );
  IV U50065 ( .A(n37119), .Z(n37120) );
  NOR U50066 ( .A(n37121), .B(n37120), .Z(n38484) );
  IV U50067 ( .A(n37122), .Z(n37124) );
  NOR U50068 ( .A(n37124), .B(n37123), .Z(n38477) );
  NOR U50069 ( .A(n38484), .B(n38477), .Z(n37125) );
  XOR U50070 ( .A(n38478), .B(n37125), .Z(n40189) );
  XOR U50071 ( .A(n37126), .B(n40189), .Z(n38471) );
  XOR U50072 ( .A(n37127), .B(n38471), .Z(n38475) );
  XOR U50073 ( .A(n38474), .B(n38475), .Z(n38470) );
  NOR U50074 ( .A(n37134), .B(n38470), .Z(n41764) );
  IV U50075 ( .A(n37128), .Z(n37129) );
  NOR U50076 ( .A(n37130), .B(n37129), .Z(n38468) );
  XOR U50077 ( .A(n38470), .B(n38468), .Z(n38467) );
  IV U50078 ( .A(n37131), .Z(n37133) );
  NOR U50079 ( .A(n37133), .B(n37132), .Z(n37135) );
  IV U50080 ( .A(n37135), .Z(n38466) );
  XOR U50081 ( .A(n38467), .B(n38466), .Z(n37137) );
  NOR U50082 ( .A(n37135), .B(n37134), .Z(n37136) );
  NOR U50083 ( .A(n37137), .B(n37136), .Z(n37138) );
  NOR U50084 ( .A(n41764), .B(n37138), .Z(n38460) );
  XOR U50085 ( .A(n38462), .B(n38460), .Z(n38465) );
  IV U50086 ( .A(n37139), .Z(n37149) );
  IV U50087 ( .A(n37140), .Z(n37141) );
  NOR U50088 ( .A(n37149), .B(n37141), .Z(n38463) );
  XOR U50089 ( .A(n38465), .B(n38463), .Z(n40199) );
  IV U50090 ( .A(n40199), .Z(n37151) );
  IV U50091 ( .A(n37142), .Z(n37146) );
  NOR U50092 ( .A(n37144), .B(n37143), .Z(n37145) );
  IV U50093 ( .A(n37145), .Z(n37153) );
  NOR U50094 ( .A(n37146), .B(n37153), .Z(n40197) );
  IV U50095 ( .A(n37147), .Z(n37148) );
  NOR U50096 ( .A(n37149), .B(n37148), .Z(n40195) );
  NOR U50097 ( .A(n40197), .B(n40195), .Z(n37150) );
  XOR U50098 ( .A(n37151), .B(n37150), .Z(n38459) );
  IV U50099 ( .A(n37152), .Z(n37154) );
  NOR U50100 ( .A(n37154), .B(n37153), .Z(n38457) );
  XOR U50101 ( .A(n38459), .B(n38457), .Z(n37164) );
  NOR U50102 ( .A(n37162), .B(n37164), .Z(n37155) );
  IV U50103 ( .A(n37155), .Z(n37156) );
  NOR U50104 ( .A(n37157), .B(n37156), .Z(n43635) );
  IV U50105 ( .A(n37158), .Z(n37159) );
  NOR U50106 ( .A(n38459), .B(n37159), .Z(n37160) );
  IV U50107 ( .A(n37160), .Z(n37161) );
  NOR U50108 ( .A(n37162), .B(n37161), .Z(n38456) );
  NOR U50109 ( .A(n37163), .B(n37162), .Z(n37166) );
  IV U50110 ( .A(n37164), .Z(n37165) );
  NOR U50111 ( .A(n37166), .B(n37165), .Z(n37167) );
  NOR U50112 ( .A(n38456), .B(n37167), .Z(n37168) );
  IV U50113 ( .A(n37168), .Z(n37169) );
  NOR U50114 ( .A(n43635), .B(n37169), .Z(n38454) );
  XOR U50115 ( .A(n37170), .B(n38454), .Z(n38451) );
  IV U50116 ( .A(n37171), .Z(n37172) );
  NOR U50117 ( .A(n37173), .B(n37172), .Z(n38450) );
  IV U50118 ( .A(n37174), .Z(n37176) );
  NOR U50119 ( .A(n37176), .B(n37175), .Z(n38448) );
  NOR U50120 ( .A(n38450), .B(n38448), .Z(n37177) );
  XOR U50121 ( .A(n38451), .B(n37177), .Z(n40206) );
  XOR U50122 ( .A(n40207), .B(n40206), .Z(n38445) );
  XOR U50123 ( .A(n38444), .B(n38445), .Z(n40204) );
  XOR U50124 ( .A(n40205), .B(n40204), .Z(n38435) );
  IV U50125 ( .A(n37178), .Z(n38440) );
  NOR U50126 ( .A(n37179), .B(n38440), .Z(n40214) );
  IV U50127 ( .A(n37180), .Z(n37182) );
  NOR U50128 ( .A(n37182), .B(n37181), .Z(n38438) );
  NOR U50129 ( .A(n40214), .B(n38438), .Z(n37183) );
  XOR U50130 ( .A(n38435), .B(n37183), .Z(n40222) );
  XOR U50131 ( .A(n40220), .B(n40222), .Z(n43677) );
  XOR U50132 ( .A(n40223), .B(n43677), .Z(n40227) );
  IV U50133 ( .A(n37184), .Z(n37185) );
  NOR U50134 ( .A(n37186), .B(n37185), .Z(n40226) );
  IV U50135 ( .A(n37187), .Z(n37189) );
  NOR U50136 ( .A(n37189), .B(n37188), .Z(n40233) );
  NOR U50137 ( .A(n40226), .B(n40233), .Z(n37190) );
  XOR U50138 ( .A(n40227), .B(n37190), .Z(n38433) );
  IV U50139 ( .A(n37191), .Z(n37193) );
  NOR U50140 ( .A(n37193), .B(n37192), .Z(n38431) );
  XOR U50141 ( .A(n38433), .B(n38431), .Z(n40231) );
  XOR U50142 ( .A(n40230), .B(n40231), .Z(n38427) );
  XOR U50143 ( .A(n38425), .B(n38427), .Z(n38430) );
  XOR U50144 ( .A(n37194), .B(n38430), .Z(n38416) );
  IV U50145 ( .A(n37195), .Z(n37196) );
  NOR U50146 ( .A(n37197), .B(n37196), .Z(n38422) );
  IV U50147 ( .A(n37198), .Z(n37200) );
  NOR U50148 ( .A(n37200), .B(n37199), .Z(n38415) );
  NOR U50149 ( .A(n38422), .B(n38415), .Z(n37201) );
  XOR U50150 ( .A(n38416), .B(n37201), .Z(n38418) );
  NOR U50151 ( .A(n37209), .B(n38418), .Z(n43703) );
  IV U50152 ( .A(n37202), .Z(n37203) );
  NOR U50153 ( .A(n37204), .B(n37203), .Z(n38411) );
  IV U50154 ( .A(n37205), .Z(n37207) );
  NOR U50155 ( .A(n37207), .B(n37206), .Z(n37208) );
  IV U50156 ( .A(n37208), .Z(n38419) );
  XOR U50157 ( .A(n38419), .B(n38418), .Z(n38412) );
  XOR U50158 ( .A(n38411), .B(n38412), .Z(n37211) );
  NOR U50159 ( .A(n38412), .B(n37209), .Z(n37210) );
  NOR U50160 ( .A(n37211), .B(n37210), .Z(n37212) );
  NOR U50161 ( .A(n43703), .B(n37212), .Z(n38409) );
  IV U50162 ( .A(n37213), .Z(n37215) );
  NOR U50163 ( .A(n37215), .B(n37214), .Z(n38408) );
  IV U50164 ( .A(n37216), .Z(n37218) );
  NOR U50165 ( .A(n37218), .B(n37217), .Z(n40246) );
  NOR U50166 ( .A(n38408), .B(n40246), .Z(n37219) );
  XOR U50167 ( .A(n38409), .B(n37219), .Z(n40245) );
  IV U50168 ( .A(n37220), .Z(n37222) );
  NOR U50169 ( .A(n37222), .B(n37221), .Z(n40243) );
  XOR U50170 ( .A(n40245), .B(n40243), .Z(n40252) );
  XOR U50171 ( .A(n40251), .B(n40252), .Z(n40261) );
  XOR U50172 ( .A(n37223), .B(n40261), .Z(n40259) );
  XOR U50173 ( .A(n40257), .B(n40259), .Z(n41705) );
  IV U50174 ( .A(n37224), .Z(n37225) );
  NOR U50175 ( .A(n37226), .B(n37225), .Z(n41709) );
  IV U50176 ( .A(n37227), .Z(n37228) );
  NOR U50177 ( .A(n37229), .B(n37228), .Z(n41704) );
  NOR U50178 ( .A(n41709), .B(n41704), .Z(n38407) );
  XOR U50179 ( .A(n41705), .B(n38407), .Z(n38399) );
  XOR U50180 ( .A(n37230), .B(n38399), .Z(n40275) );
  XOR U50181 ( .A(n37231), .B(n40275), .Z(n37232) );
  IV U50182 ( .A(n37232), .Z(n40281) );
  XOR U50183 ( .A(n40280), .B(n40281), .Z(n40279) );
  XOR U50184 ( .A(n40277), .B(n40279), .Z(n38393) );
  XOR U50185 ( .A(n38391), .B(n38393), .Z(n38396) );
  XOR U50186 ( .A(n37233), .B(n38396), .Z(n37234) );
  IV U50187 ( .A(n37234), .Z(n38387) );
  IV U50188 ( .A(n37235), .Z(n37237) );
  NOR U50189 ( .A(n37237), .B(n37236), .Z(n38385) );
  XOR U50190 ( .A(n38387), .B(n38385), .Z(n40287) );
  XOR U50191 ( .A(n40288), .B(n40287), .Z(n38383) );
  NOR U50192 ( .A(n37239), .B(n37238), .Z(n38382) );
  IV U50193 ( .A(n37240), .Z(n37241) );
  NOR U50194 ( .A(n37242), .B(n37241), .Z(n40289) );
  NOR U50195 ( .A(n38382), .B(n40289), .Z(n37243) );
  XOR U50196 ( .A(n38383), .B(n37243), .Z(n38377) );
  XOR U50197 ( .A(n38376), .B(n38377), .Z(n38380) );
  XOR U50198 ( .A(n38379), .B(n38380), .Z(n40295) );
  XOR U50199 ( .A(n40294), .B(n40295), .Z(n40303) );
  XOR U50200 ( .A(n37244), .B(n40303), .Z(n40300) );
  XOR U50201 ( .A(n37245), .B(n40300), .Z(n40316) );
  IV U50202 ( .A(n37249), .Z(n37246) );
  NOR U50203 ( .A(n37246), .B(n37248), .Z(n40308) );
  IV U50204 ( .A(n37247), .Z(n37251) );
  XOR U50205 ( .A(n37249), .B(n37248), .Z(n37250) );
  NOR U50206 ( .A(n37251), .B(n37250), .Z(n40314) );
  NOR U50207 ( .A(n40308), .B(n40314), .Z(n37252) );
  XOR U50208 ( .A(n40316), .B(n37252), .Z(n38375) );
  XOR U50209 ( .A(n37253), .B(n38375), .Z(n40320) );
  XOR U50210 ( .A(n40318), .B(n40320), .Z(n38370) );
  XOR U50211 ( .A(n38368), .B(n38370), .Z(n38372) );
  XOR U50212 ( .A(n38371), .B(n38372), .Z(n38362) );
  XOR U50213 ( .A(n38360), .B(n38362), .Z(n38364) );
  IV U50214 ( .A(n37254), .Z(n37255) );
  NOR U50215 ( .A(n37256), .B(n37255), .Z(n38363) );
  IV U50216 ( .A(n37257), .Z(n37259) );
  NOR U50217 ( .A(n37259), .B(n37258), .Z(n38358) );
  NOR U50218 ( .A(n38363), .B(n38358), .Z(n37260) );
  XOR U50219 ( .A(n38364), .B(n37260), .Z(n37261) );
  NOR U50220 ( .A(n37262), .B(n37261), .Z(n37265) );
  IV U50221 ( .A(n37262), .Z(n37264) );
  XOR U50222 ( .A(n38358), .B(n38364), .Z(n37263) );
  NOR U50223 ( .A(n37264), .B(n37263), .Z(n41645) );
  NOR U50224 ( .A(n37265), .B(n41645), .Z(n37266) );
  IV U50225 ( .A(n37266), .Z(n40337) );
  NOR U50226 ( .A(n37268), .B(n37267), .Z(n40335) );
  XOR U50227 ( .A(n40337), .B(n40335), .Z(n40340) );
  XOR U50228 ( .A(n40339), .B(n40340), .Z(n40347) );
  IV U50229 ( .A(n37272), .Z(n37269) );
  NOR U50230 ( .A(n37271), .B(n37269), .Z(n40342) );
  IV U50231 ( .A(n37270), .Z(n37274) );
  XOR U50232 ( .A(n37272), .B(n37271), .Z(n37273) );
  NOR U50233 ( .A(n37274), .B(n37273), .Z(n40345) );
  NOR U50234 ( .A(n40342), .B(n40345), .Z(n37275) );
  XOR U50235 ( .A(n40347), .B(n37275), .Z(n38351) );
  IV U50236 ( .A(n37276), .Z(n40351) );
  NOR U50237 ( .A(n40351), .B(n40353), .Z(n37279) );
  NOR U50238 ( .A(n37277), .B(n38352), .Z(n37278) );
  NOR U50239 ( .A(n37279), .B(n37278), .Z(n37280) );
  XOR U50240 ( .A(n38351), .B(n37280), .Z(n38346) );
  NOR U50241 ( .A(n37282), .B(n37281), .Z(n37283) );
  IV U50242 ( .A(n37283), .Z(n37286) );
  NOR U50243 ( .A(n37284), .B(n37286), .Z(n38344) );
  XOR U50244 ( .A(n38346), .B(n38344), .Z(n38348) );
  IV U50245 ( .A(n37285), .Z(n37287) );
  NOR U50246 ( .A(n37287), .B(n37286), .Z(n37288) );
  IV U50247 ( .A(n37288), .Z(n38347) );
  XOR U50248 ( .A(n38348), .B(n38347), .Z(n38342) );
  IV U50249 ( .A(n37289), .Z(n37290) );
  NOR U50250 ( .A(n37291), .B(n37290), .Z(n38341) );
  IV U50251 ( .A(n37292), .Z(n37293) );
  NOR U50252 ( .A(n37294), .B(n37293), .Z(n40361) );
  NOR U50253 ( .A(n38341), .B(n40361), .Z(n37295) );
  XOR U50254 ( .A(n38342), .B(n37295), .Z(n40365) );
  XOR U50255 ( .A(n40364), .B(n40365), .Z(n40371) );
  XOR U50256 ( .A(n40370), .B(n40371), .Z(n38339) );
  XOR U50257 ( .A(n38338), .B(n38339), .Z(n40382) );
  XOR U50258 ( .A(n37296), .B(n40382), .Z(n37297) );
  IV U50259 ( .A(n37297), .Z(n40386) );
  IV U50260 ( .A(n37298), .Z(n37300) );
  NOR U50261 ( .A(n37300), .B(n37299), .Z(n40384) );
  XOR U50262 ( .A(n40386), .B(n40384), .Z(n38330) );
  XOR U50263 ( .A(n38331), .B(n38330), .Z(n38332) );
  IV U50264 ( .A(n37301), .Z(n37303) );
  NOR U50265 ( .A(n37303), .B(n37302), .Z(n43788) );
  IV U50266 ( .A(n37304), .Z(n37305) );
  NOR U50267 ( .A(n37306), .B(n37305), .Z(n41609) );
  NOR U50268 ( .A(n43788), .B(n41609), .Z(n38333) );
  XOR U50269 ( .A(n38332), .B(n38333), .Z(n38326) );
  XOR U50270 ( .A(n38324), .B(n38326), .Z(n38328) );
  XOR U50271 ( .A(n38327), .B(n38328), .Z(n38319) );
  XOR U50272 ( .A(n38318), .B(n38319), .Z(n38323) );
  XOR U50273 ( .A(n38321), .B(n38323), .Z(n38314) );
  XOR U50274 ( .A(n38313), .B(n38314), .Z(n41589) );
  XOR U50275 ( .A(n37307), .B(n41589), .Z(n40393) );
  XOR U50276 ( .A(n40392), .B(n40393), .Z(n40397) );
  IV U50277 ( .A(n37308), .Z(n37310) );
  NOR U50278 ( .A(n37310), .B(n37309), .Z(n40395) );
  XOR U50279 ( .A(n40397), .B(n40395), .Z(n38308) );
  XOR U50280 ( .A(n38307), .B(n38308), .Z(n38312) );
  IV U50281 ( .A(n37311), .Z(n37315) );
  NOR U50282 ( .A(n37313), .B(n37312), .Z(n37314) );
  IV U50283 ( .A(n37314), .Z(n37317) );
  NOR U50284 ( .A(n37315), .B(n37317), .Z(n38310) );
  XOR U50285 ( .A(n38312), .B(n38310), .Z(n38303) );
  IV U50286 ( .A(n37316), .Z(n37318) );
  NOR U50287 ( .A(n37318), .B(n37317), .Z(n37319) );
  IV U50288 ( .A(n37319), .Z(n38302) );
  XOR U50289 ( .A(n38303), .B(n38302), .Z(n38304) );
  IV U50290 ( .A(n37320), .Z(n37322) );
  NOR U50291 ( .A(n37322), .B(n37321), .Z(n41568) );
  IV U50292 ( .A(n37323), .Z(n37325) );
  NOR U50293 ( .A(n37325), .B(n37324), .Z(n43796) );
  NOR U50294 ( .A(n41568), .B(n43796), .Z(n38305) );
  XOR U50295 ( .A(n38304), .B(n38305), .Z(n38298) );
  XOR U50296 ( .A(n38296), .B(n38298), .Z(n38301) );
  XOR U50297 ( .A(n38299), .B(n38301), .Z(n40403) );
  XOR U50298 ( .A(n40401), .B(n40403), .Z(n43803) );
  XOR U50299 ( .A(n40404), .B(n43803), .Z(n38293) );
  IV U50300 ( .A(n37326), .Z(n37327) );
  NOR U50301 ( .A(n37328), .B(n37327), .Z(n40407) );
  IV U50302 ( .A(n37329), .Z(n37330) );
  NOR U50303 ( .A(n37334), .B(n37330), .Z(n38294) );
  NOR U50304 ( .A(n40407), .B(n38294), .Z(n37331) );
  XOR U50305 ( .A(n38293), .B(n37331), .Z(n38292) );
  IV U50306 ( .A(n37332), .Z(n37333) );
  NOR U50307 ( .A(n37334), .B(n37333), .Z(n38290) );
  XOR U50308 ( .A(n38292), .B(n38290), .Z(n38285) );
  XOR U50309 ( .A(n38284), .B(n38285), .Z(n38288) );
  XOR U50310 ( .A(n38287), .B(n38288), .Z(n38279) );
  XOR U50311 ( .A(n38278), .B(n38279), .Z(n41557) );
  XOR U50312 ( .A(n38281), .B(n41557), .Z(n38273) );
  IV U50313 ( .A(n37335), .Z(n37337) );
  NOR U50314 ( .A(n37337), .B(n37336), .Z(n41553) );
  IV U50315 ( .A(n37338), .Z(n37340) );
  NOR U50316 ( .A(n37340), .B(n37339), .Z(n41548) );
  NOR U50317 ( .A(n41553), .B(n41548), .Z(n38274) );
  XOR U50318 ( .A(n38273), .B(n38274), .Z(n40417) );
  XOR U50319 ( .A(n37341), .B(n40417), .Z(n38271) );
  XOR U50320 ( .A(n38272), .B(n38271), .Z(n38265) );
  IV U50321 ( .A(n37342), .Z(n37343) );
  NOR U50322 ( .A(n37343), .B(n37345), .Z(n41540) );
  IV U50323 ( .A(n37344), .Z(n37346) );
  NOR U50324 ( .A(n37346), .B(n37345), .Z(n43823) );
  NOR U50325 ( .A(n41540), .B(n43823), .Z(n38266) );
  XOR U50326 ( .A(n38265), .B(n38266), .Z(n38269) );
  XOR U50327 ( .A(n38267), .B(n38269), .Z(n38260) );
  XOR U50328 ( .A(n38259), .B(n38260), .Z(n38263) );
  XOR U50329 ( .A(n37347), .B(n38263), .Z(n38250) );
  XOR U50330 ( .A(n38248), .B(n38250), .Z(n40428) );
  XOR U50331 ( .A(n40429), .B(n40428), .Z(n40431) );
  IV U50332 ( .A(n37348), .Z(n37349) );
  NOR U50333 ( .A(n37350), .B(n37349), .Z(n40430) );
  IV U50334 ( .A(n37351), .Z(n37353) );
  NOR U50335 ( .A(n37353), .B(n37352), .Z(n40435) );
  NOR U50336 ( .A(n40430), .B(n40435), .Z(n37354) );
  XOR U50337 ( .A(n40431), .B(n37354), .Z(n38243) );
  XOR U50338 ( .A(n38241), .B(n38243), .Z(n38245) );
  XOR U50339 ( .A(n38244), .B(n38245), .Z(n40440) );
  XOR U50340 ( .A(n37355), .B(n40440), .Z(n40442) );
  XOR U50341 ( .A(n37356), .B(n40442), .Z(n40449) );
  XOR U50342 ( .A(n40448), .B(n40449), .Z(n40452) );
  XOR U50343 ( .A(n40451), .B(n40452), .Z(n40456) );
  XOR U50344 ( .A(n37357), .B(n40456), .Z(n40462) );
  IV U50345 ( .A(n37358), .Z(n37359) );
  NOR U50346 ( .A(n37360), .B(n37359), .Z(n41530) );
  IV U50347 ( .A(n37361), .Z(n37362) );
  NOR U50348 ( .A(n37363), .B(n37362), .Z(n43883) );
  NOR U50349 ( .A(n41530), .B(n43883), .Z(n40463) );
  XOR U50350 ( .A(n40462), .B(n40463), .Z(n40466) );
  XOR U50351 ( .A(n40464), .B(n40466), .Z(n40471) );
  XOR U50352 ( .A(n37364), .B(n40471), .Z(n38232) );
  XOR U50353 ( .A(n38230), .B(n38232), .Z(n41517) );
  IV U50354 ( .A(n37365), .Z(n37367) );
  NOR U50355 ( .A(n37367), .B(n37366), .Z(n41516) );
  IV U50356 ( .A(n37368), .Z(n37369) );
  NOR U50357 ( .A(n37369), .B(n37374), .Z(n43892) );
  NOR U50358 ( .A(n41516), .B(n43892), .Z(n38229) );
  XOR U50359 ( .A(n41517), .B(n38229), .Z(n37383) );
  IV U50360 ( .A(n37383), .Z(n37371) );
  NOR U50361 ( .A(n37371), .B(n37370), .Z(n37372) );
  IV U50362 ( .A(n37372), .Z(n37377) );
  NOR U50363 ( .A(n37374), .B(n37373), .Z(n37375) );
  IV U50364 ( .A(n37375), .Z(n37376) );
  NOR U50365 ( .A(n37377), .B(n37376), .Z(n37378) );
  IV U50366 ( .A(n37378), .Z(n37379) );
  NOR U50367 ( .A(n37380), .B(n37379), .Z(n41514) );
  NOR U50368 ( .A(n37381), .B(n37380), .Z(n37382) );
  NOR U50369 ( .A(n37383), .B(n37382), .Z(n37384) );
  NOR U50370 ( .A(n41514), .B(n37384), .Z(n38221) );
  XOR U50371 ( .A(n37385), .B(n38221), .Z(n38224) );
  XOR U50372 ( .A(n38223), .B(n38224), .Z(n38215) );
  XOR U50373 ( .A(n38216), .B(n38215), .Z(n38213) );
  IV U50374 ( .A(n37386), .Z(n37388) );
  NOR U50375 ( .A(n37388), .B(n37387), .Z(n38217) );
  IV U50376 ( .A(n37389), .Z(n37390) );
  NOR U50377 ( .A(n37390), .B(n37393), .Z(n38212) );
  NOR U50378 ( .A(n38217), .B(n38212), .Z(n37391) );
  XOR U50379 ( .A(n38213), .B(n37391), .Z(n38211) );
  IV U50380 ( .A(n37392), .Z(n37394) );
  NOR U50381 ( .A(n37394), .B(n37393), .Z(n38209) );
  XOR U50382 ( .A(n38211), .B(n38209), .Z(n41497) );
  XOR U50383 ( .A(n37395), .B(n41497), .Z(n41488) );
  XOR U50384 ( .A(n40479), .B(n41488), .Z(n43910) );
  XOR U50385 ( .A(n40487), .B(n43910), .Z(n37405) );
  IV U50386 ( .A(n37405), .Z(n40489) );
  IV U50387 ( .A(n37396), .Z(n37397) );
  NOR U50388 ( .A(n37397), .B(n37403), .Z(n37398) );
  IV U50389 ( .A(n37398), .Z(n37410) );
  NOR U50390 ( .A(n40489), .B(n37410), .Z(n40496) );
  IV U50391 ( .A(n37399), .Z(n37401) );
  NOR U50392 ( .A(n37401), .B(n37400), .Z(n40488) );
  IV U50393 ( .A(n37402), .Z(n37404) );
  NOR U50394 ( .A(n37404), .B(n37403), .Z(n40484) );
  NOR U50395 ( .A(n40488), .B(n40484), .Z(n37406) );
  XOR U50396 ( .A(n37406), .B(n37405), .Z(n38205) );
  IV U50397 ( .A(n37407), .Z(n37419) );
  IV U50398 ( .A(n37408), .Z(n37409) );
  NOR U50399 ( .A(n37419), .B(n37409), .Z(n37411) );
  IV U50400 ( .A(n37411), .Z(n38204) );
  XOR U50401 ( .A(n38205), .B(n38204), .Z(n37413) );
  NOR U50402 ( .A(n37411), .B(n37410), .Z(n37412) );
  NOR U50403 ( .A(n37413), .B(n37412), .Z(n37414) );
  NOR U50404 ( .A(n40496), .B(n37414), .Z(n38202) );
  IV U50405 ( .A(n37415), .Z(n37416) );
  NOR U50406 ( .A(n37416), .B(n37425), .Z(n38201) );
  IV U50407 ( .A(n37417), .Z(n37418) );
  NOR U50408 ( .A(n37419), .B(n37418), .Z(n38206) );
  NOR U50409 ( .A(n38201), .B(n38206), .Z(n37420) );
  XOR U50410 ( .A(n38202), .B(n37420), .Z(n38200) );
  IV U50411 ( .A(n37421), .Z(n37422) );
  NOR U50412 ( .A(n37423), .B(n37422), .Z(n38195) );
  IV U50413 ( .A(n37424), .Z(n37426) );
  NOR U50414 ( .A(n37426), .B(n37425), .Z(n38198) );
  NOR U50415 ( .A(n38195), .B(n38198), .Z(n37427) );
  XOR U50416 ( .A(n38200), .B(n37427), .Z(n40502) );
  NOR U50417 ( .A(n40508), .B(n40503), .Z(n37428) );
  IV U50418 ( .A(n37428), .Z(n37429) );
  NOR U50419 ( .A(n40506), .B(n37429), .Z(n37430) );
  XOR U50420 ( .A(n40502), .B(n37430), .Z(n40515) );
  NOR U50421 ( .A(n37432), .B(n37431), .Z(n40509) );
  IV U50422 ( .A(n37433), .Z(n40517) );
  NOR U50423 ( .A(n37434), .B(n40517), .Z(n37435) );
  NOR U50424 ( .A(n40509), .B(n37435), .Z(n37436) );
  XOR U50425 ( .A(n40515), .B(n37436), .Z(n40522) );
  XOR U50426 ( .A(n40520), .B(n40522), .Z(n37444) );
  IV U50427 ( .A(n37437), .Z(n37438) );
  NOR U50428 ( .A(n37453), .B(n37438), .Z(n37449) );
  IV U50429 ( .A(n37449), .Z(n37439) );
  NOR U50430 ( .A(n37444), .B(n37439), .Z(n41451) );
  IV U50431 ( .A(n37440), .Z(n37443) );
  NOR U50432 ( .A(n40522), .B(n37442), .Z(n37441) );
  IV U50433 ( .A(n37441), .Z(n47248) );
  NOR U50434 ( .A(n37443), .B(n47248), .Z(n38194) );
  NOR U50435 ( .A(n37443), .B(n37442), .Z(n37446) );
  IV U50436 ( .A(n37444), .Z(n37445) );
  NOR U50437 ( .A(n37446), .B(n37445), .Z(n37447) );
  NOR U50438 ( .A(n38194), .B(n37447), .Z(n37448) );
  NOR U50439 ( .A(n37449), .B(n37448), .Z(n37450) );
  NOR U50440 ( .A(n41451), .B(n37450), .Z(n40527) );
  IV U50441 ( .A(n37451), .Z(n37452) );
  NOR U50442 ( .A(n37453), .B(n37452), .Z(n37454) );
  IV U50443 ( .A(n37454), .Z(n40528) );
  XOR U50444 ( .A(n40527), .B(n40528), .Z(n38192) );
  NOR U50445 ( .A(n37456), .B(n37455), .Z(n38191) );
  IV U50446 ( .A(n37457), .Z(n38188) );
  NOR U50447 ( .A(n37458), .B(n38188), .Z(n37459) );
  NOR U50448 ( .A(n38191), .B(n37459), .Z(n37460) );
  XOR U50449 ( .A(n38192), .B(n37460), .Z(n40535) );
  XOR U50450 ( .A(n40536), .B(n40535), .Z(n40537) );
  XOR U50451 ( .A(n41442), .B(n40537), .Z(n40542) );
  IV U50452 ( .A(n37461), .Z(n37467) );
  IV U50453 ( .A(n37462), .Z(n37464) );
  NOR U50454 ( .A(n37464), .B(n37463), .Z(n37465) );
  IV U50455 ( .A(n37465), .Z(n37466) );
  NOR U50456 ( .A(n37467), .B(n37466), .Z(n44732) );
  NOR U50457 ( .A(n47271), .B(n44732), .Z(n40543) );
  XOR U50458 ( .A(n40542), .B(n40543), .Z(n40545) );
  XOR U50459 ( .A(n40544), .B(n40545), .Z(n40551) );
  XOR U50460 ( .A(n37468), .B(n40551), .Z(n40556) );
  XOR U50461 ( .A(n40554), .B(n40556), .Z(n40559) );
  IV U50462 ( .A(n37469), .Z(n37471) );
  NOR U50463 ( .A(n37471), .B(n37470), .Z(n40557) );
  XOR U50464 ( .A(n40559), .B(n40557), .Z(n38186) );
  IV U50465 ( .A(n37472), .Z(n37474) );
  NOR U50466 ( .A(n37474), .B(n37473), .Z(n38184) );
  XOR U50467 ( .A(n38186), .B(n38184), .Z(n38180) );
  XOR U50468 ( .A(n38179), .B(n38180), .Z(n38182) );
  XOR U50469 ( .A(n38183), .B(n38182), .Z(n38174) );
  IV U50470 ( .A(n37475), .Z(n37477) );
  NOR U50471 ( .A(n37477), .B(n37476), .Z(n41417) );
  IV U50472 ( .A(n37478), .Z(n37479) );
  NOR U50473 ( .A(n37480), .B(n37479), .Z(n41422) );
  NOR U50474 ( .A(n41417), .B(n41422), .Z(n38175) );
  XOR U50475 ( .A(n38174), .B(n38175), .Z(n38178) );
  XOR U50476 ( .A(n38176), .B(n38178), .Z(n38171) );
  XOR U50477 ( .A(n38168), .B(n38171), .Z(n38166) );
  XOR U50478 ( .A(n37481), .B(n38166), .Z(n38163) );
  XOR U50479 ( .A(n38161), .B(n38163), .Z(n40566) );
  IV U50480 ( .A(n37482), .Z(n37484) );
  NOR U50481 ( .A(n37484), .B(n37483), .Z(n40564) );
  XOR U50482 ( .A(n40566), .B(n40564), .Z(n41403) );
  IV U50483 ( .A(n37485), .Z(n37487) );
  NOR U50484 ( .A(n37487), .B(n37486), .Z(n43955) );
  IV U50485 ( .A(n37488), .Z(n37490) );
  NOR U50486 ( .A(n37490), .B(n37489), .Z(n41400) );
  NOR U50487 ( .A(n43955), .B(n41400), .Z(n40567) );
  XOR U50488 ( .A(n41403), .B(n40567), .Z(n40570) );
  XOR U50489 ( .A(n37491), .B(n40570), .Z(n40575) );
  XOR U50490 ( .A(n40576), .B(n40575), .Z(n40586) );
  IV U50491 ( .A(n37492), .Z(n40581) );
  NOR U50492 ( .A(n40581), .B(n37493), .Z(n37496) );
  IV U50493 ( .A(n37494), .Z(n37495) );
  NOR U50494 ( .A(n37499), .B(n37495), .Z(n40585) );
  NOR U50495 ( .A(n37496), .B(n40585), .Z(n37497) );
  XOR U50496 ( .A(n40586), .B(n37497), .Z(n40595) );
  IV U50497 ( .A(n37498), .Z(n37503) );
  NOR U50498 ( .A(n37500), .B(n37499), .Z(n37501) );
  IV U50499 ( .A(n37501), .Z(n37502) );
  NOR U50500 ( .A(n37503), .B(n37502), .Z(n40593) );
  XOR U50501 ( .A(n40595), .B(n40593), .Z(n40597) );
  XOR U50502 ( .A(n40596), .B(n40597), .Z(n38159) );
  XOR U50503 ( .A(n38158), .B(n38159), .Z(n38155) );
  XOR U50504 ( .A(n38153), .B(n38155), .Z(n38157) );
  NOR U50505 ( .A(n37504), .B(n38157), .Z(n43970) );
  IV U50506 ( .A(n37505), .Z(n37508) );
  IV U50507 ( .A(n37506), .Z(n37507) );
  NOR U50508 ( .A(n37508), .B(n37507), .Z(n37509) );
  IV U50509 ( .A(n37509), .Z(n38156) );
  XOR U50510 ( .A(n38157), .B(n38156), .Z(n37510) );
  NOR U50511 ( .A(n37511), .B(n37510), .Z(n38152) );
  IV U50512 ( .A(n37512), .Z(n37513) );
  NOR U50513 ( .A(n37514), .B(n37513), .Z(n38150) );
  XOR U50514 ( .A(n38152), .B(n38150), .Z(n37515) );
  NOR U50515 ( .A(n43970), .B(n37515), .Z(n38144) );
  XOR U50516 ( .A(n38146), .B(n38144), .Z(n38147) );
  XOR U50517 ( .A(n38148), .B(n38147), .Z(n38138) );
  IV U50518 ( .A(n37516), .Z(n37517) );
  NOR U50519 ( .A(n37518), .B(n37517), .Z(n38141) );
  IV U50520 ( .A(n37519), .Z(n37521) );
  NOR U50521 ( .A(n37521), .B(n37520), .Z(n38139) );
  NOR U50522 ( .A(n38141), .B(n38139), .Z(n37522) );
  XOR U50523 ( .A(n38138), .B(n37522), .Z(n40605) );
  XOR U50524 ( .A(n40603), .B(n40605), .Z(n40607) );
  XOR U50525 ( .A(n40606), .B(n40607), .Z(n38133) );
  XOR U50526 ( .A(n38132), .B(n38133), .Z(n38136) );
  XOR U50527 ( .A(n38135), .B(n38136), .Z(n41354) );
  XOR U50528 ( .A(n37523), .B(n41354), .Z(n40613) );
  XOR U50529 ( .A(n40612), .B(n40613), .Z(n40618) );
  XOR U50530 ( .A(n40617), .B(n40618), .Z(n40622) );
  IV U50531 ( .A(n37524), .Z(n37526) );
  IV U50532 ( .A(n37525), .Z(n37528) );
  NOR U50533 ( .A(n37526), .B(n37528), .Z(n40620) );
  XOR U50534 ( .A(n40622), .B(n40620), .Z(n40625) );
  IV U50535 ( .A(n37527), .Z(n37529) );
  NOR U50536 ( .A(n37529), .B(n37528), .Z(n37530) );
  IV U50537 ( .A(n37530), .Z(n40624) );
  XOR U50538 ( .A(n40625), .B(n40624), .Z(n38129) );
  IV U50539 ( .A(n37531), .Z(n37532) );
  NOR U50540 ( .A(n37533), .B(n37532), .Z(n40626) );
  IV U50541 ( .A(n37534), .Z(n37535) );
  NOR U50542 ( .A(n37536), .B(n37535), .Z(n38128) );
  NOR U50543 ( .A(n40626), .B(n38128), .Z(n37537) );
  XOR U50544 ( .A(n38129), .B(n37537), .Z(n38124) );
  XOR U50545 ( .A(n38123), .B(n38124), .Z(n44001) );
  XOR U50546 ( .A(n37538), .B(n44001), .Z(n44008) );
  XOR U50547 ( .A(n38119), .B(n44008), .Z(n44012) );
  XOR U50548 ( .A(n38121), .B(n44012), .Z(n38114) );
  XOR U50549 ( .A(n37539), .B(n38114), .Z(n38111) );
  IV U50550 ( .A(n37540), .Z(n37541) );
  NOR U50551 ( .A(n37542), .B(n37541), .Z(n38108) );
  IV U50552 ( .A(n37543), .Z(n37545) );
  NOR U50553 ( .A(n37545), .B(n37544), .Z(n38110) );
  NOR U50554 ( .A(n38108), .B(n38110), .Z(n37546) );
  XOR U50555 ( .A(n38111), .B(n37546), .Z(n38104) );
  XOR U50556 ( .A(n38105), .B(n38104), .Z(n40635) );
  IV U50557 ( .A(n37547), .Z(n37548) );
  NOR U50558 ( .A(n37549), .B(n37548), .Z(n40634) );
  IV U50559 ( .A(n37550), .Z(n37552) );
  NOR U50560 ( .A(n37552), .B(n37551), .Z(n38106) );
  NOR U50561 ( .A(n40634), .B(n38106), .Z(n37553) );
  XOR U50562 ( .A(n40635), .B(n37553), .Z(n38101) );
  IV U50563 ( .A(n37554), .Z(n37556) );
  NOR U50564 ( .A(n37556), .B(n37555), .Z(n38102) );
  IV U50565 ( .A(n37557), .Z(n37559) );
  NOR U50566 ( .A(n37559), .B(n37558), .Z(n40637) );
  NOR U50567 ( .A(n38102), .B(n40637), .Z(n37560) );
  XOR U50568 ( .A(n38101), .B(n37560), .Z(n38098) );
  XOR U50569 ( .A(n38097), .B(n38098), .Z(n40641) );
  XOR U50570 ( .A(n40640), .B(n40641), .Z(n40644) );
  XOR U50571 ( .A(n40643), .B(n40644), .Z(n51655) );
  XOR U50572 ( .A(n40658), .B(n51655), .Z(n40661) );
  IV U50573 ( .A(n37561), .Z(n51649) );
  NOR U50574 ( .A(n51649), .B(n51652), .Z(n40660) );
  IV U50575 ( .A(n37562), .Z(n37563) );
  NOR U50576 ( .A(n37564), .B(n37563), .Z(n38095) );
  NOR U50577 ( .A(n40660), .B(n38095), .Z(n37565) );
  XOR U50578 ( .A(n40661), .B(n37565), .Z(n37572) );
  IV U50579 ( .A(n37572), .Z(n40667) );
  NOR U50580 ( .A(n37573), .B(n40667), .Z(n44062) );
  IV U50581 ( .A(n37566), .Z(n37567) );
  NOR U50582 ( .A(n37568), .B(n37567), .Z(n40676) );
  IV U50583 ( .A(n37569), .Z(n37570) );
  NOR U50584 ( .A(n37571), .B(n37570), .Z(n40666) );
  XOR U50585 ( .A(n40666), .B(n37572), .Z(n40677) );
  XOR U50586 ( .A(n40676), .B(n40677), .Z(n37575) );
  NOR U50587 ( .A(n40677), .B(n37573), .Z(n37574) );
  NOR U50588 ( .A(n37575), .B(n37574), .Z(n37576) );
  NOR U50589 ( .A(n44062), .B(n37576), .Z(n37589) );
  IV U50590 ( .A(n37577), .Z(n37578) );
  NOR U50591 ( .A(n37579), .B(n37578), .Z(n40670) );
  IV U50592 ( .A(n37580), .Z(n37582) );
  NOR U50593 ( .A(n37582), .B(n37581), .Z(n40673) );
  NOR U50594 ( .A(n40670), .B(n40673), .Z(n37583) );
  XOR U50595 ( .A(n37589), .B(n37583), .Z(n37592) );
  NOR U50596 ( .A(n37596), .B(n37592), .Z(n40694) );
  IV U50597 ( .A(n37584), .Z(n37585) );
  NOR U50598 ( .A(n37601), .B(n37585), .Z(n40690) );
  IV U50599 ( .A(n37586), .Z(n37588) );
  NOR U50600 ( .A(n37588), .B(n37587), .Z(n37594) );
  IV U50601 ( .A(n37594), .Z(n37591) );
  IV U50602 ( .A(n37589), .Z(n40674) );
  XOR U50603 ( .A(n40670), .B(n40674), .Z(n37590) );
  NOR U50604 ( .A(n37591), .B(n37590), .Z(n41311) );
  IV U50605 ( .A(n37592), .Z(n37593) );
  NOR U50606 ( .A(n37594), .B(n37593), .Z(n37595) );
  NOR U50607 ( .A(n41311), .B(n37595), .Z(n40691) );
  XOR U50608 ( .A(n40690), .B(n40691), .Z(n37598) );
  NOR U50609 ( .A(n40691), .B(n37596), .Z(n37597) );
  NOR U50610 ( .A(n37598), .B(n37597), .Z(n37599) );
  NOR U50611 ( .A(n40694), .B(n37599), .Z(n40687) );
  IV U50612 ( .A(n37600), .Z(n37602) );
  NOR U50613 ( .A(n37602), .B(n37601), .Z(n40686) );
  IV U50614 ( .A(n37603), .Z(n37605) );
  NOR U50615 ( .A(n37605), .B(n37604), .Z(n40699) );
  NOR U50616 ( .A(n40686), .B(n40699), .Z(n37606) );
  XOR U50617 ( .A(n40687), .B(n37606), .Z(n38092) );
  XOR U50618 ( .A(n37607), .B(n38092), .Z(n40705) );
  IV U50619 ( .A(n37608), .Z(n37610) );
  NOR U50620 ( .A(n37610), .B(n37609), .Z(n40703) );
  XOR U50621 ( .A(n40705), .B(n40703), .Z(n38085) );
  XOR U50622 ( .A(n38084), .B(n38085), .Z(n38088) );
  XOR U50623 ( .A(n38087), .B(n38088), .Z(n38080) );
  XOR U50624 ( .A(n38078), .B(n38080), .Z(n38083) );
  XOR U50625 ( .A(n38081), .B(n38083), .Z(n38074) );
  XOR U50626 ( .A(n38072), .B(n38074), .Z(n38076) );
  XOR U50627 ( .A(n37611), .B(n38076), .Z(n38068) );
  XOR U50628 ( .A(n38069), .B(n38068), .Z(n40729) );
  XOR U50629 ( .A(n40728), .B(n40729), .Z(n40727) );
  XOR U50630 ( .A(n40725), .B(n40727), .Z(n40742) );
  XOR U50631 ( .A(n37612), .B(n40742), .Z(n38065) );
  IV U50632 ( .A(n37613), .Z(n37615) );
  NOR U50633 ( .A(n37615), .B(n37614), .Z(n40741) );
  IV U50634 ( .A(n37616), .Z(n37617) );
  NOR U50635 ( .A(n37618), .B(n37617), .Z(n38064) );
  NOR U50636 ( .A(n40741), .B(n38064), .Z(n37619) );
  XOR U50637 ( .A(n38065), .B(n37619), .Z(n38061) );
  IV U50638 ( .A(n37620), .Z(n37622) );
  NOR U50639 ( .A(n37622), .B(n37621), .Z(n38059) );
  IV U50640 ( .A(n37623), .Z(n37624) );
  NOR U50641 ( .A(n37625), .B(n37624), .Z(n38057) );
  NOR U50642 ( .A(n38059), .B(n38057), .Z(n37626) );
  XOR U50643 ( .A(n38061), .B(n37626), .Z(n37627) );
  NOR U50644 ( .A(n37628), .B(n37627), .Z(n37631) );
  IV U50645 ( .A(n37628), .Z(n37630) );
  XOR U50646 ( .A(n38059), .B(n38061), .Z(n37629) );
  NOR U50647 ( .A(n37630), .B(n37629), .Z(n44091) );
  NOR U50648 ( .A(n37631), .B(n44091), .Z(n37632) );
  IV U50649 ( .A(n37632), .Z(n38055) );
  XOR U50650 ( .A(n37633), .B(n38055), .Z(n38045) );
  NOR U50651 ( .A(n37634), .B(n38046), .Z(n37637) );
  NOR U50652 ( .A(n37636), .B(n37635), .Z(n40754) );
  NOR U50653 ( .A(n37637), .B(n40754), .Z(n37638) );
  XOR U50654 ( .A(n38045), .B(n37638), .Z(n38043) );
  XOR U50655 ( .A(n38041), .B(n38043), .Z(n40761) );
  XOR U50656 ( .A(n40760), .B(n40761), .Z(n40764) );
  XOR U50657 ( .A(n40763), .B(n40764), .Z(n40768) );
  XOR U50658 ( .A(n40767), .B(n40768), .Z(n40772) );
  XOR U50659 ( .A(n40770), .B(n40772), .Z(n40775) );
  XOR U50660 ( .A(n40774), .B(n40775), .Z(n40778) );
  XOR U50661 ( .A(n40777), .B(n40778), .Z(n40783) );
  XOR U50662 ( .A(n40781), .B(n40783), .Z(n40784) );
  NOR U50663 ( .A(n37646), .B(n40784), .Z(n41247) );
  IV U50664 ( .A(n37639), .Z(n37641) );
  NOR U50665 ( .A(n37641), .B(n37640), .Z(n38037) );
  IV U50666 ( .A(n37642), .Z(n37643) );
  NOR U50667 ( .A(n37644), .B(n37643), .Z(n37645) );
  IV U50668 ( .A(n37645), .Z(n40785) );
  XOR U50669 ( .A(n40785), .B(n40784), .Z(n38038) );
  XOR U50670 ( .A(n38037), .B(n38038), .Z(n37648) );
  NOR U50671 ( .A(n38038), .B(n37646), .Z(n37647) );
  NOR U50672 ( .A(n37648), .B(n37647), .Z(n37649) );
  NOR U50673 ( .A(n41247), .B(n37649), .Z(n37655) );
  IV U50674 ( .A(n37655), .Z(n40789) );
  NOR U50675 ( .A(n44600), .B(n40789), .Z(n40791) );
  IV U50676 ( .A(n37650), .Z(n37652) );
  NOR U50677 ( .A(n37652), .B(n37651), .Z(n41243) );
  NOR U50678 ( .A(n37654), .B(n37653), .Z(n40788) );
  XOR U50679 ( .A(n40788), .B(n37655), .Z(n40793) );
  XOR U50680 ( .A(n41243), .B(n40793), .Z(n37657) );
  NOR U50681 ( .A(n40793), .B(n44600), .Z(n37656) );
  NOR U50682 ( .A(n37657), .B(n37656), .Z(n37658) );
  NOR U50683 ( .A(n40791), .B(n37658), .Z(n40796) );
  IV U50684 ( .A(n37659), .Z(n37661) );
  NOR U50685 ( .A(n37661), .B(n37660), .Z(n40795) );
  IV U50686 ( .A(n37662), .Z(n37663) );
  NOR U50687 ( .A(n37663), .B(n37666), .Z(n40799) );
  NOR U50688 ( .A(n40795), .B(n40799), .Z(n37664) );
  XOR U50689 ( .A(n40796), .B(n37664), .Z(n40806) );
  XOR U50690 ( .A(n40802), .B(n40806), .Z(n40812) );
  IV U50691 ( .A(n37665), .Z(n37667) );
  NOR U50692 ( .A(n37667), .B(n37666), .Z(n40804) );
  IV U50693 ( .A(n37668), .Z(n37669) );
  NOR U50694 ( .A(n37670), .B(n37669), .Z(n40811) );
  NOR U50695 ( .A(n40804), .B(n40811), .Z(n37671) );
  XOR U50696 ( .A(n40812), .B(n37671), .Z(n40808) );
  XOR U50697 ( .A(n37672), .B(n40808), .Z(n40816) );
  XOR U50698 ( .A(n40815), .B(n40816), .Z(n38034) );
  XOR U50699 ( .A(n37673), .B(n38034), .Z(n40833) );
  XOR U50700 ( .A(n40832), .B(n40833), .Z(n40827) );
  XOR U50701 ( .A(n40828), .B(n40827), .Z(n40823) );
  IV U50702 ( .A(n37674), .Z(n37676) );
  NOR U50703 ( .A(n37676), .B(n37675), .Z(n40822) );
  NOR U50704 ( .A(n37678), .B(n37677), .Z(n37679) );
  IV U50705 ( .A(n37679), .Z(n37680) );
  NOR U50706 ( .A(n37681), .B(n37680), .Z(n40851) );
  NOR U50707 ( .A(n40822), .B(n40851), .Z(n37682) );
  XOR U50708 ( .A(n40823), .B(n37682), .Z(n41228) );
  XOR U50709 ( .A(n37683), .B(n41228), .Z(n38030) );
  XOR U50710 ( .A(n38029), .B(n38030), .Z(n40858) );
  XOR U50711 ( .A(n40857), .B(n40858), .Z(n40867) );
  IV U50712 ( .A(n37684), .Z(n37686) );
  NOR U50713 ( .A(n37686), .B(n37685), .Z(n40866) );
  NOR U50714 ( .A(n40860), .B(n40866), .Z(n37687) );
  XOR U50715 ( .A(n40867), .B(n37687), .Z(n38025) );
  IV U50716 ( .A(n37688), .Z(n37689) );
  NOR U50717 ( .A(n37690), .B(n37689), .Z(n40863) );
  IV U50718 ( .A(n37691), .Z(n37693) );
  NOR U50719 ( .A(n37693), .B(n37692), .Z(n38026) );
  NOR U50720 ( .A(n40863), .B(n38026), .Z(n37694) );
  XOR U50721 ( .A(n38025), .B(n37694), .Z(n40882) );
  IV U50722 ( .A(n40882), .Z(n37706) );
  IV U50723 ( .A(n37695), .Z(n37696) );
  NOR U50724 ( .A(n40871), .B(n37696), .Z(n37704) );
  IV U50725 ( .A(n37712), .Z(n37697) );
  NOR U50726 ( .A(n37708), .B(n37697), .Z(n37698) );
  IV U50727 ( .A(n37698), .Z(n37703) );
  NOR U50728 ( .A(n37700), .B(n37699), .Z(n37701) );
  IV U50729 ( .A(n37701), .Z(n37702) );
  NOR U50730 ( .A(n37703), .B(n37702), .Z(n40881) );
  NOR U50731 ( .A(n37704), .B(n40881), .Z(n37705) );
  XOR U50732 ( .A(n37706), .B(n37705), .Z(n40888) );
  IV U50733 ( .A(n37707), .Z(n37709) );
  NOR U50734 ( .A(n37709), .B(n37708), .Z(n37710) );
  IV U50735 ( .A(n37710), .Z(n37711) );
  NOR U50736 ( .A(n37712), .B(n37711), .Z(n40884) );
  XOR U50737 ( .A(n40888), .B(n40884), .Z(n40893) );
  IV U50738 ( .A(n37713), .Z(n37715) );
  NOR U50739 ( .A(n37715), .B(n37714), .Z(n40886) );
  IV U50740 ( .A(n37716), .Z(n37718) );
  NOR U50741 ( .A(n37718), .B(n37717), .Z(n40892) );
  NOR U50742 ( .A(n40886), .B(n40892), .Z(n37719) );
  XOR U50743 ( .A(n40893), .B(n37719), .Z(n40897) );
  XOR U50744 ( .A(n40898), .B(n40897), .Z(n38023) );
  XOR U50745 ( .A(n38022), .B(n38023), .Z(n38018) );
  XOR U50746 ( .A(n38017), .B(n38018), .Z(n38020) );
  XOR U50747 ( .A(n38021), .B(n38020), .Z(n38014) );
  IV U50748 ( .A(n37720), .Z(n37727) );
  NOR U50749 ( .A(n37722), .B(n37721), .Z(n37723) );
  IV U50750 ( .A(n37723), .Z(n37724) );
  NOR U50751 ( .A(n37725), .B(n37724), .Z(n37726) );
  IV U50752 ( .A(n37726), .Z(n37733) );
  NOR U50753 ( .A(n37727), .B(n37733), .Z(n40907) );
  IV U50754 ( .A(n37728), .Z(n37730) );
  NOR U50755 ( .A(n37730), .B(n37729), .Z(n38015) );
  NOR U50756 ( .A(n40907), .B(n38015), .Z(n37731) );
  XOR U50757 ( .A(n38014), .B(n37731), .Z(n40906) );
  IV U50758 ( .A(n37732), .Z(n37734) );
  NOR U50759 ( .A(n37734), .B(n37733), .Z(n40904) );
  XOR U50760 ( .A(n40906), .B(n40904), .Z(n37735) );
  NOR U50761 ( .A(n47611), .B(n37735), .Z(n44213) );
  IV U50762 ( .A(n37736), .Z(n37738) );
  NOR U50763 ( .A(n37738), .B(n37737), .Z(n38012) );
  NOR U50764 ( .A(n38012), .B(n40904), .Z(n37739) );
  XOR U50765 ( .A(n40906), .B(n37739), .Z(n47606) );
  NOR U50766 ( .A(n37740), .B(n47606), .Z(n37741) );
  NOR U50767 ( .A(n44213), .B(n37741), .Z(n38008) );
  IV U50768 ( .A(n37742), .Z(n37743) );
  NOR U50769 ( .A(n37744), .B(n37743), .Z(n41193) );
  IV U50770 ( .A(n37745), .Z(n37747) );
  NOR U50771 ( .A(n37747), .B(n37746), .Z(n44218) );
  NOR U50772 ( .A(n41193), .B(n44218), .Z(n38009) );
  XOR U50773 ( .A(n38008), .B(n38009), .Z(n40916) );
  XOR U50774 ( .A(n37748), .B(n40916), .Z(n40914) );
  IV U50775 ( .A(n37749), .Z(n37760) );
  NOR U50776 ( .A(n40914), .B(n37760), .Z(n37750) );
  IV U50777 ( .A(n37750), .Z(n37753) );
  NOR U50778 ( .A(n37751), .B(n37753), .Z(n44232) );
  IV U50779 ( .A(n37752), .Z(n37754) );
  NOR U50780 ( .A(n37754), .B(n37753), .Z(n41185) );
  IV U50781 ( .A(n37755), .Z(n37756) );
  NOR U50782 ( .A(n37756), .B(n37997), .Z(n37771) );
  NOR U50783 ( .A(n41185), .B(n37771), .Z(n37757) );
  IV U50784 ( .A(n37757), .Z(n37758) );
  NOR U50785 ( .A(n44232), .B(n37758), .Z(n37759) );
  IV U50786 ( .A(n37759), .Z(n37770) );
  NOR U50787 ( .A(n37761), .B(n37760), .Z(n37768) );
  IV U50788 ( .A(n37762), .Z(n37763) );
  NOR U50789 ( .A(n37767), .B(n37763), .Z(n37764) );
  IV U50790 ( .A(n37764), .Z(n38005) );
  IV U50791 ( .A(n37765), .Z(n37766) );
  NOR U50792 ( .A(n37767), .B(n37766), .Z(n40912) );
  XOR U50793 ( .A(n40912), .B(n40914), .Z(n38004) );
  XOR U50794 ( .A(n38005), .B(n38004), .Z(n37995) );
  NOR U50795 ( .A(n37768), .B(n37995), .Z(n37769) );
  NOR U50796 ( .A(n37770), .B(n37769), .Z(n37774) );
  IV U50797 ( .A(n37771), .Z(n37772) );
  NOR U50798 ( .A(n37995), .B(n37772), .Z(n37773) );
  NOR U50799 ( .A(n37774), .B(n37773), .Z(n40927) );
  XOR U50800 ( .A(n40920), .B(n40927), .Z(n37991) );
  IV U50801 ( .A(n37775), .Z(n37776) );
  NOR U50802 ( .A(n37777), .B(n37776), .Z(n40925) );
  IV U50803 ( .A(n37778), .Z(n37779) );
  NOR U50804 ( .A(n37780), .B(n37779), .Z(n37990) );
  NOR U50805 ( .A(n40925), .B(n37990), .Z(n37781) );
  XOR U50806 ( .A(n37991), .B(n37781), .Z(n37985) );
  IV U50807 ( .A(n37782), .Z(n37784) );
  NOR U50808 ( .A(n37784), .B(n37783), .Z(n37983) );
  XOR U50809 ( .A(n37985), .B(n37983), .Z(n37987) );
  XOR U50810 ( .A(n37986), .B(n37987), .Z(n37981) );
  XOR U50811 ( .A(n37979), .B(n37981), .Z(n40930) );
  XOR U50812 ( .A(n40929), .B(n40930), .Z(n40936) );
  XOR U50813 ( .A(n40932), .B(n40936), .Z(n37977) );
  XOR U50814 ( .A(n37785), .B(n37977), .Z(n40945) );
  XOR U50815 ( .A(n40938), .B(n40945), .Z(n40941) );
  IV U50816 ( .A(n37786), .Z(n37787) );
  NOR U50817 ( .A(n37788), .B(n37787), .Z(n37789) );
  IV U50818 ( .A(n37789), .Z(n40940) );
  XOR U50819 ( .A(n40941), .B(n40940), .Z(n40948) );
  NOR U50820 ( .A(n37791), .B(n37790), .Z(n40943) );
  NOR U50821 ( .A(n37793), .B(n37792), .Z(n40947) );
  NOR U50822 ( .A(n40943), .B(n40947), .Z(n37794) );
  XOR U50823 ( .A(n40948), .B(n37794), .Z(n40962) );
  XOR U50824 ( .A(n37974), .B(n40962), .Z(n40964) );
  XOR U50825 ( .A(n37795), .B(n40964), .Z(n37971) );
  NOR U50826 ( .A(n37797), .B(n37796), .Z(n40966) );
  IV U50827 ( .A(n40970), .Z(n37799) );
  IV U50828 ( .A(n37798), .Z(n40969) );
  NOR U50829 ( .A(n37799), .B(n40969), .Z(n37972) );
  NOR U50830 ( .A(n40966), .B(n37972), .Z(n37800) );
  XOR U50831 ( .A(n37971), .B(n37800), .Z(n40971) );
  IV U50832 ( .A(n37801), .Z(n40975) );
  NOR U50833 ( .A(n40975), .B(n40969), .Z(n37808) );
  IV U50834 ( .A(n37802), .Z(n37804) );
  NOR U50835 ( .A(n37804), .B(n37803), .Z(n37969) );
  NOR U50836 ( .A(n37808), .B(n37969), .Z(n37805) );
  XOR U50837 ( .A(n40971), .B(n37805), .Z(n37806) );
  NOR U50838 ( .A(n37807), .B(n37806), .Z(n37811) );
  IV U50839 ( .A(n37807), .Z(n37810) );
  XOR U50840 ( .A(n37808), .B(n40971), .Z(n37809) );
  NOR U50841 ( .A(n37810), .B(n37809), .Z(n41143) );
  NOR U50842 ( .A(n37811), .B(n41143), .Z(n40977) );
  XOR U50843 ( .A(n40976), .B(n40977), .Z(n40981) );
  IV U50844 ( .A(n37812), .Z(n37813) );
  NOR U50845 ( .A(n37814), .B(n37813), .Z(n40980) );
  NOR U50846 ( .A(n37816), .B(n37815), .Z(n40987) );
  NOR U50847 ( .A(n40980), .B(n40987), .Z(n37817) );
  XOR U50848 ( .A(n40981), .B(n37817), .Z(n40986) );
  IV U50849 ( .A(n37818), .Z(n37819) );
  NOR U50850 ( .A(n37820), .B(n37819), .Z(n40984) );
  XOR U50851 ( .A(n40986), .B(n40984), .Z(n40993) );
  XOR U50852 ( .A(n40991), .B(n40993), .Z(n40995) );
  XOR U50853 ( .A(n40994), .B(n40995), .Z(n44281) );
  XOR U50854 ( .A(n37821), .B(n44281), .Z(n37966) );
  XOR U50855 ( .A(n37965), .B(n37966), .Z(n37959) );
  XOR U50856 ( .A(n37958), .B(n37959), .Z(n37963) );
  IV U50857 ( .A(n37822), .Z(n37824) );
  NOR U50858 ( .A(n37824), .B(n37823), .Z(n37961) );
  XOR U50859 ( .A(n37963), .B(n37961), .Z(n37953) );
  XOR U50860 ( .A(n37952), .B(n37953), .Z(n37957) );
  NOR U50861 ( .A(n37826), .B(n37825), .Z(n37827) );
  IV U50862 ( .A(n37827), .Z(n37828) );
  NOR U50863 ( .A(n37829), .B(n37828), .Z(n37955) );
  XOR U50864 ( .A(n37957), .B(n37955), .Z(n41001) );
  IV U50865 ( .A(n37830), .Z(n37831) );
  NOR U50866 ( .A(n37832), .B(n37831), .Z(n37950) );
  IV U50867 ( .A(n37833), .Z(n37835) );
  NOR U50868 ( .A(n37835), .B(n37834), .Z(n41000) );
  NOR U50869 ( .A(n37950), .B(n41000), .Z(n37836) );
  XOR U50870 ( .A(n41001), .B(n37836), .Z(n37947) );
  IV U50871 ( .A(n37837), .Z(n37839) );
  NOR U50872 ( .A(n37839), .B(n37838), .Z(n37948) );
  IV U50873 ( .A(n37840), .Z(n37842) );
  NOR U50874 ( .A(n37842), .B(n37841), .Z(n41003) );
  NOR U50875 ( .A(n37948), .B(n41003), .Z(n37843) );
  XOR U50876 ( .A(n37947), .B(n37843), .Z(n47819) );
  IV U50877 ( .A(n37844), .Z(n37848) );
  NOR U50878 ( .A(n37846), .B(n37845), .Z(n37847) );
  IV U50879 ( .A(n37847), .Z(n37850) );
  NOR U50880 ( .A(n37848), .B(n37850), .Z(n41007) );
  IV U50881 ( .A(n37849), .Z(n37851) );
  NOR U50882 ( .A(n37851), .B(n37850), .Z(n47820) );
  NOR U50883 ( .A(n41007), .B(n47820), .Z(n37852) );
  XOR U50884 ( .A(n47819), .B(n37852), .Z(n41009) );
  XOR U50885 ( .A(n37853), .B(n41009), .Z(n41013) );
  XOR U50886 ( .A(n41012), .B(n41013), .Z(n41017) );
  XOR U50887 ( .A(n41016), .B(n41017), .Z(n44310) );
  IV U50888 ( .A(n37854), .Z(n37855) );
  NOR U50889 ( .A(n37855), .B(n37861), .Z(n37943) );
  IV U50890 ( .A(n37856), .Z(n37858) );
  NOR U50891 ( .A(n37858), .B(n37857), .Z(n44308) );
  IV U50892 ( .A(n37859), .Z(n37860) );
  NOR U50893 ( .A(n37861), .B(n37860), .Z(n44317) );
  NOR U50894 ( .A(n44308), .B(n44317), .Z(n37945) );
  IV U50895 ( .A(n37945), .Z(n37862) );
  NOR U50896 ( .A(n37943), .B(n37862), .Z(n37863) );
  XOR U50897 ( .A(n44310), .B(n37863), .Z(n37937) );
  NOR U50898 ( .A(n37869), .B(n37864), .Z(n37938) );
  IV U50899 ( .A(n37865), .Z(n37867) );
  NOR U50900 ( .A(n37867), .B(n37866), .Z(n37940) );
  NOR U50901 ( .A(n37938), .B(n37940), .Z(n37868) );
  XOR U50902 ( .A(n37937), .B(n37868), .Z(n37936) );
  NOR U50903 ( .A(n37870), .B(n37869), .Z(n37871) );
  IV U50904 ( .A(n37871), .Z(n37872) );
  NOR U50905 ( .A(n37873), .B(n37872), .Z(n37874) );
  IV U50906 ( .A(n37874), .Z(n37935) );
  XOR U50907 ( .A(n37936), .B(n37935), .Z(n37929) );
  NOR U50908 ( .A(n37876), .B(n37875), .Z(n44454) );
  IV U50909 ( .A(n37877), .Z(n37879) );
  NOR U50910 ( .A(n37879), .B(n37878), .Z(n44449) );
  NOR U50911 ( .A(n44454), .B(n44449), .Z(n41098) );
  XOR U50912 ( .A(n37929), .B(n41098), .Z(n37931) );
  XOR U50913 ( .A(n37930), .B(n37931), .Z(n41034) );
  XOR U50914 ( .A(n37880), .B(n41034), .Z(n41032) );
  XOR U50915 ( .A(n41030), .B(n41032), .Z(n41039) );
  IV U50916 ( .A(n37881), .Z(n37883) );
  NOR U50917 ( .A(n37883), .B(n37882), .Z(n41037) );
  XOR U50918 ( .A(n41039), .B(n41037), .Z(n41044) );
  IV U50919 ( .A(n37884), .Z(n37885) );
  NOR U50920 ( .A(n37886), .B(n37885), .Z(n41040) );
  IV U50921 ( .A(n37887), .Z(n37888) );
  NOR U50922 ( .A(n41073), .B(n37888), .Z(n41043) );
  NOR U50923 ( .A(n41040), .B(n41043), .Z(n37889) );
  XOR U50924 ( .A(n41044), .B(n37889), .Z(n37895) );
  IV U50925 ( .A(n37895), .Z(n41067) );
  NOR U50926 ( .A(n37890), .B(n41067), .Z(n44327) );
  IV U50927 ( .A(n37891), .Z(n37892) );
  NOR U50928 ( .A(n37893), .B(n37892), .Z(n37896) );
  IV U50929 ( .A(n37896), .Z(n37894) );
  XOR U50930 ( .A(n41040), .B(n41044), .Z(n47792) );
  NOR U50931 ( .A(n37894), .B(n47792), .Z(n41046) );
  NOR U50932 ( .A(n37896), .B(n37895), .Z(n37897) );
  NOR U50933 ( .A(n41046), .B(n37897), .Z(n37905) );
  NOR U50934 ( .A(n37898), .B(n37905), .Z(n37899) );
  NOR U50935 ( .A(n44327), .B(n37899), .Z(n37908) );
  IV U50936 ( .A(n37908), .Z(n37900) );
  NOR U50937 ( .A(n37901), .B(n37900), .Z(n41061) );
  IV U50938 ( .A(n37902), .Z(n37903) );
  NOR U50939 ( .A(n37904), .B(n37903), .Z(n37909) );
  IV U50940 ( .A(n37909), .Z(n37907) );
  IV U50941 ( .A(n37905), .Z(n37906) );
  NOR U50942 ( .A(n37907), .B(n37906), .Z(n37926) );
  NOR U50943 ( .A(n37909), .B(n37908), .Z(n37910) );
  NOR U50944 ( .A(n37926), .B(n37910), .Z(n37911) );
  NOR U50945 ( .A(n37912), .B(n37911), .Z(n37913) );
  NOR U50946 ( .A(n41061), .B(n37913), .Z(n37924) );
  IV U50947 ( .A(n37914), .Z(n37915) );
  NOR U50948 ( .A(n37916), .B(n37915), .Z(n41048) );
  IV U50949 ( .A(n37917), .Z(n37918) );
  NOR U50950 ( .A(n37919), .B(n37918), .Z(n37923) );
  NOR U50951 ( .A(n41048), .B(n37923), .Z(n37920) );
  XOR U50952 ( .A(n37924), .B(n37920), .Z(n44337) );
  XOR U50953 ( .A(n44336), .B(n44337), .Z(n44342) );
  IV U50954 ( .A(n44342), .Z(n37921) );
  NOR U50955 ( .A(n37922), .B(n37921), .Z(n44370) );
  IV U50956 ( .A(n44370), .Z(n41052) );
  IV U50957 ( .A(n37923), .Z(n37925) );
  IV U50958 ( .A(n37924), .Z(n41049) );
  NOR U50959 ( .A(n37925), .B(n41049), .Z(n44333) );
  IV U50960 ( .A(n37926), .Z(n44331) );
  IV U50961 ( .A(n37927), .Z(n37928) );
  NOR U50962 ( .A(n37928), .B(n37931), .Z(n41090) );
  IV U50963 ( .A(n37929), .Z(n41096) );
  NOR U50964 ( .A(n41098), .B(n41096), .Z(n37933) );
  IV U50965 ( .A(n37930), .Z(n37932) );
  NOR U50966 ( .A(n37932), .B(n37931), .Z(n41093) );
  NOR U50967 ( .A(n37933), .B(n41093), .Z(n37934) );
  IV U50968 ( .A(n37934), .Z(n41029) );
  NOR U50969 ( .A(n37936), .B(n37935), .Z(n41102) );
  IV U50970 ( .A(n37937), .Z(n37942) );
  IV U50971 ( .A(n37938), .Z(n37939) );
  NOR U50972 ( .A(n37942), .B(n37939), .Z(n41099) );
  IV U50973 ( .A(n37940), .Z(n37941) );
  NOR U50974 ( .A(n37942), .B(n37941), .Z(n41106) );
  IV U50975 ( .A(n37943), .Z(n37944) );
  NOR U50976 ( .A(n44310), .B(n37944), .Z(n44314) );
  NOR U50977 ( .A(n44310), .B(n37945), .Z(n41028) );
  IV U50978 ( .A(n47820), .Z(n37946) );
  NOR U50979 ( .A(n47819), .B(n37946), .Z(n41111) );
  IV U50980 ( .A(n41111), .Z(n41109) );
  IV U50981 ( .A(n37947), .Z(n41005) );
  IV U50982 ( .A(n37948), .Z(n37949) );
  NOR U50983 ( .A(n41005), .B(n37949), .Z(n44290) );
  IV U50984 ( .A(n37950), .Z(n37951) );
  NOR U50985 ( .A(n37951), .B(n41001), .Z(n41116) );
  IV U50986 ( .A(n37952), .Z(n37954) );
  NOR U50987 ( .A(n37954), .B(n37953), .Z(n41125) );
  IV U50988 ( .A(n37955), .Z(n37956) );
  NOR U50989 ( .A(n37957), .B(n37956), .Z(n41122) );
  NOR U50990 ( .A(n41125), .B(n41122), .Z(n40999) );
  IV U50991 ( .A(n37958), .Z(n37960) );
  NOR U50992 ( .A(n37960), .B(n37959), .Z(n41130) );
  IV U50993 ( .A(n37961), .Z(n37962) );
  NOR U50994 ( .A(n37963), .B(n37962), .Z(n41128) );
  NOR U50995 ( .A(n41130), .B(n41128), .Z(n40998) );
  NOR U50996 ( .A(n37964), .B(n44281), .Z(n37968) );
  IV U50997 ( .A(n37965), .Z(n37967) );
  NOR U50998 ( .A(n37967), .B(n37966), .Z(n41133) );
  NOR U50999 ( .A(n37968), .B(n41133), .Z(n40997) );
  IV U51000 ( .A(n37969), .Z(n37970) );
  NOR U51001 ( .A(n37970), .B(n40971), .Z(n41148) );
  IV U51002 ( .A(n37971), .Z(n40968) );
  IV U51003 ( .A(n37972), .Z(n37973) );
  NOR U51004 ( .A(n40968), .B(n37973), .Z(n44262) );
  IV U51005 ( .A(n37974), .Z(n37975) );
  NOR U51006 ( .A(n40962), .B(n37975), .Z(n40955) );
  IV U51007 ( .A(n37976), .Z(n37978) );
  NOR U51008 ( .A(n37978), .B(n37977), .Z(n41163) );
  IV U51009 ( .A(n37979), .Z(n37980) );
  NOR U51010 ( .A(n37981), .B(n37980), .Z(n37982) );
  IV U51011 ( .A(n37982), .Z(n41172) );
  IV U51012 ( .A(n37983), .Z(n37984) );
  NOR U51013 ( .A(n37985), .B(n37984), .Z(n44243) );
  IV U51014 ( .A(n37986), .Z(n37988) );
  NOR U51015 ( .A(n37988), .B(n37987), .Z(n41174) );
  NOR U51016 ( .A(n44243), .B(n41174), .Z(n37989) );
  IV U51017 ( .A(n37989), .Z(n40928) );
  IV U51018 ( .A(n37990), .Z(n37993) );
  IV U51019 ( .A(n37991), .Z(n37992) );
  NOR U51020 ( .A(n37993), .B(n37992), .Z(n44240) );
  IV U51021 ( .A(n37994), .Z(n38002) );
  IV U51022 ( .A(n37995), .Z(n37996) );
  NOR U51023 ( .A(n37997), .B(n37996), .Z(n37998) );
  IV U51024 ( .A(n37998), .Z(n37999) );
  NOR U51025 ( .A(n38000), .B(n37999), .Z(n38001) );
  IV U51026 ( .A(n38001), .Z(n40922) );
  NOR U51027 ( .A(n38002), .B(n40922), .Z(n38003) );
  IV U51028 ( .A(n38003), .Z(n41183) );
  NOR U51029 ( .A(n38005), .B(n38004), .Z(n44224) );
  NOR U51030 ( .A(n44224), .B(n41185), .Z(n40919) );
  IV U51031 ( .A(n38006), .Z(n38007) );
  NOR U51032 ( .A(n38007), .B(n40916), .Z(n41190) );
  IV U51033 ( .A(n38008), .Z(n41195) );
  NOR U51034 ( .A(n38009), .B(n41195), .Z(n38010) );
  NOR U51035 ( .A(n44213), .B(n38010), .Z(n38011) );
  IV U51036 ( .A(n38011), .Z(n40911) );
  IV U51037 ( .A(n38012), .Z(n38013) );
  NOR U51038 ( .A(n40906), .B(n38013), .Z(n44211) );
  IV U51039 ( .A(n38014), .Z(n40909) );
  IV U51040 ( .A(n38015), .Z(n38016) );
  NOR U51041 ( .A(n40909), .B(n38016), .Z(n41198) );
  IV U51042 ( .A(n38017), .Z(n38019) );
  NOR U51043 ( .A(n38019), .B(n38018), .Z(n44201) );
  NOR U51044 ( .A(n38021), .B(n38020), .Z(n41204) );
  NOR U51045 ( .A(n44201), .B(n41204), .Z(n40903) );
  IV U51046 ( .A(n38022), .Z(n38024) );
  NOR U51047 ( .A(n38024), .B(n38023), .Z(n40901) );
  IV U51048 ( .A(n40901), .Z(n40896) );
  IV U51049 ( .A(n38025), .Z(n40865) );
  IV U51050 ( .A(n38026), .Z(n38027) );
  NOR U51051 ( .A(n40865), .B(n38027), .Z(n41208) );
  NOR U51052 ( .A(n38028), .B(n41228), .Z(n41221) );
  IV U51053 ( .A(n38029), .Z(n38031) );
  NOR U51054 ( .A(n38031), .B(n38030), .Z(n41224) );
  NOR U51055 ( .A(n41221), .B(n41224), .Z(n40855) );
  IV U51056 ( .A(n40833), .Z(n44152) );
  NOR U51057 ( .A(n40832), .B(n44152), .Z(n40836) );
  IV U51058 ( .A(n38032), .Z(n38033) );
  NOR U51059 ( .A(n38034), .B(n38033), .Z(n44157) );
  IV U51060 ( .A(n38035), .Z(n38036) );
  NOR U51061 ( .A(n38036), .B(n40816), .Z(n41234) );
  IV U51062 ( .A(n38037), .Z(n38040) );
  IV U51063 ( .A(n38038), .Z(n38039) );
  NOR U51064 ( .A(n38040), .B(n38039), .Z(n44118) );
  IV U51065 ( .A(n38041), .Z(n38042) );
  NOR U51066 ( .A(n38043), .B(n38042), .Z(n40758) );
  IV U51067 ( .A(n40758), .Z(n40753) );
  IV U51068 ( .A(n38044), .Z(n38048) );
  IV U51069 ( .A(n38045), .Z(n40756) );
  NOR U51070 ( .A(n40756), .B(n38046), .Z(n38047) );
  IV U51071 ( .A(n38047), .Z(n38050) );
  NOR U51072 ( .A(n38048), .B(n38050), .Z(n41261) );
  IV U51073 ( .A(n38049), .Z(n38051) );
  NOR U51074 ( .A(n38051), .B(n38050), .Z(n41259) );
  IV U51075 ( .A(n38052), .Z(n38053) );
  NOR U51076 ( .A(n38053), .B(n38055), .Z(n41264) );
  NOR U51077 ( .A(n41259), .B(n41264), .Z(n40750) );
  IV U51078 ( .A(n38054), .Z(n38056) );
  NOR U51079 ( .A(n38056), .B(n38055), .Z(n44095) );
  NOR U51080 ( .A(n44091), .B(n44095), .Z(n40749) );
  IV U51081 ( .A(n38057), .Z(n38058) );
  NOR U51082 ( .A(n38061), .B(n38058), .Z(n44088) );
  IV U51083 ( .A(n38059), .Z(n38060) );
  NOR U51084 ( .A(n38061), .B(n38060), .Z(n41267) );
  NOR U51085 ( .A(n44088), .B(n41267), .Z(n40748) );
  IV U51086 ( .A(n38062), .Z(n38063) );
  NOR U51087 ( .A(n38063), .B(n40742), .Z(n44082) );
  IV U51088 ( .A(n38064), .Z(n38067) );
  IV U51089 ( .A(n38065), .Z(n38066) );
  NOR U51090 ( .A(n38067), .B(n38066), .Z(n41273) );
  NOR U51091 ( .A(n44082), .B(n41273), .Z(n40747) );
  IV U51092 ( .A(n38068), .Z(n40716) );
  NOR U51093 ( .A(n38069), .B(n40716), .Z(n40714) );
  IV U51094 ( .A(n38070), .Z(n38071) );
  NOR U51095 ( .A(n38071), .B(n38076), .Z(n41278) );
  IV U51096 ( .A(n38072), .Z(n38073) );
  NOR U51097 ( .A(n38074), .B(n38073), .Z(n41284) );
  IV U51098 ( .A(n38075), .Z(n38077) );
  NOR U51099 ( .A(n38077), .B(n38076), .Z(n44074) );
  NOR U51100 ( .A(n41284), .B(n44074), .Z(n40712) );
  IV U51101 ( .A(n38078), .Z(n38079) );
  NOR U51102 ( .A(n38080), .B(n38079), .Z(n41286) );
  IV U51103 ( .A(n38081), .Z(n38082) );
  NOR U51104 ( .A(n38083), .B(n38082), .Z(n41281) );
  NOR U51105 ( .A(n41286), .B(n41281), .Z(n40711) );
  IV U51106 ( .A(n38084), .Z(n38086) );
  NOR U51107 ( .A(n38086), .B(n38085), .Z(n41292) );
  IV U51108 ( .A(n38087), .Z(n38089) );
  NOR U51109 ( .A(n38089), .B(n38088), .Z(n41290) );
  NOR U51110 ( .A(n41292), .B(n41290), .Z(n40710) );
  IV U51111 ( .A(n38090), .Z(n38094) );
  NOR U51112 ( .A(n38092), .B(n38091), .Z(n38093) );
  IV U51113 ( .A(n38093), .Z(n40707) );
  NOR U51114 ( .A(n38094), .B(n40707), .Z(n44069) );
  IV U51115 ( .A(n38095), .Z(n38096) );
  NOR U51116 ( .A(n38096), .B(n40661), .Z(n40664) );
  IV U51117 ( .A(n40664), .Z(n40657) );
  IV U51118 ( .A(n38097), .Z(n38099) );
  NOR U51119 ( .A(n38099), .B(n38098), .Z(n38100) );
  IV U51120 ( .A(n38100), .Z(n44042) );
  IV U51121 ( .A(n38101), .Z(n40639) );
  IV U51122 ( .A(n38102), .Z(n38103) );
  NOR U51123 ( .A(n40639), .B(n38103), .Z(n44043) );
  IV U51124 ( .A(n38104), .Z(n41327) );
  NOR U51125 ( .A(n38105), .B(n41327), .Z(n41321) );
  IV U51126 ( .A(n38106), .Z(n38107) );
  NOR U51127 ( .A(n40635), .B(n38107), .Z(n44030) );
  NOR U51128 ( .A(n41321), .B(n44030), .Z(n40632) );
  IV U51129 ( .A(n38108), .Z(n38109) );
  NOR U51130 ( .A(n38109), .B(n38111), .Z(n41334) );
  IV U51131 ( .A(n38110), .Z(n38112) );
  NOR U51132 ( .A(n38112), .B(n38111), .Z(n41331) );
  IV U51133 ( .A(n38113), .Z(n38115) );
  IV U51134 ( .A(n38114), .Z(n38117) );
  NOR U51135 ( .A(n38115), .B(n38117), .Z(n44027) );
  IV U51136 ( .A(n38116), .Z(n38118) );
  NOR U51137 ( .A(n38118), .B(n38117), .Z(n44024) );
  IV U51138 ( .A(n38119), .Z(n38120) );
  NOR U51139 ( .A(n38120), .B(n44008), .Z(n41338) );
  NOR U51140 ( .A(n38121), .B(n44012), .Z(n38122) );
  NOR U51141 ( .A(n41338), .B(n38122), .Z(n40631) );
  IV U51142 ( .A(n38123), .Z(n38125) );
  NOR U51143 ( .A(n38125), .B(n38124), .Z(n41340) );
  NOR U51144 ( .A(n38126), .B(n44001), .Z(n38127) );
  NOR U51145 ( .A(n41340), .B(n38127), .Z(n40630) );
  IV U51146 ( .A(n38128), .Z(n38130) );
  IV U51147 ( .A(n38129), .Z(n40627) );
  NOR U51148 ( .A(n38130), .B(n40627), .Z(n41343) );
  IV U51149 ( .A(n41355), .Z(n38131) );
  NOR U51150 ( .A(n41354), .B(n38131), .Z(n43987) );
  IV U51151 ( .A(n38132), .Z(n38134) );
  NOR U51152 ( .A(n38134), .B(n38133), .Z(n41365) );
  IV U51153 ( .A(n38135), .Z(n38137) );
  NOR U51154 ( .A(n38137), .B(n38136), .Z(n41360) );
  NOR U51155 ( .A(n41365), .B(n41360), .Z(n40610) );
  IV U51156 ( .A(n38138), .Z(n38143) );
  IV U51157 ( .A(n38139), .Z(n38140) );
  NOR U51158 ( .A(n38143), .B(n38140), .Z(n41368) );
  IV U51159 ( .A(n38141), .Z(n38142) );
  NOR U51160 ( .A(n38143), .B(n38142), .Z(n43977) );
  IV U51161 ( .A(n38144), .Z(n38145) );
  NOR U51162 ( .A(n38146), .B(n38145), .Z(n43974) );
  NOR U51163 ( .A(n38148), .B(n38147), .Z(n43980) );
  NOR U51164 ( .A(n43974), .B(n43980), .Z(n38149) );
  IV U51165 ( .A(n38149), .Z(n40602) );
  IV U51166 ( .A(n38150), .Z(n38151) );
  NOR U51167 ( .A(n38152), .B(n38151), .Z(n43972) );
  NOR U51168 ( .A(n43970), .B(n43972), .Z(n40601) );
  IV U51169 ( .A(n38153), .Z(n38154) );
  NOR U51170 ( .A(n38155), .B(n38154), .Z(n43961) );
  NOR U51171 ( .A(n38157), .B(n38156), .Z(n41374) );
  NOR U51172 ( .A(n43961), .B(n41374), .Z(n40600) );
  IV U51173 ( .A(n38158), .Z(n38160) );
  NOR U51174 ( .A(n38160), .B(n38159), .Z(n41378) );
  IV U51175 ( .A(n38161), .Z(n38162) );
  NOR U51176 ( .A(n38163), .B(n38162), .Z(n38164) );
  IV U51177 ( .A(n38164), .Z(n43951) );
  IV U51178 ( .A(n38165), .Z(n38167) );
  NOR U51179 ( .A(n38167), .B(n38166), .Z(n43947) );
  IV U51180 ( .A(n38168), .Z(n38169) );
  NOR U51181 ( .A(n38169), .B(n38171), .Z(n41413) );
  IV U51182 ( .A(n38170), .Z(n38172) );
  NOR U51183 ( .A(n38172), .B(n38171), .Z(n41406) );
  NOR U51184 ( .A(n41413), .B(n41406), .Z(n38173) );
  IV U51185 ( .A(n38173), .Z(n40563) );
  IV U51186 ( .A(n38174), .Z(n41418) );
  NOR U51187 ( .A(n38175), .B(n41418), .Z(n41412) );
  IV U51188 ( .A(n38176), .Z(n38177) );
  NOR U51189 ( .A(n38178), .B(n38177), .Z(n41410) );
  NOR U51190 ( .A(n41412), .B(n41410), .Z(n40562) );
  IV U51191 ( .A(n38179), .Z(n38181) );
  NOR U51192 ( .A(n38181), .B(n38180), .Z(n41428) );
  NOR U51193 ( .A(n38183), .B(n38182), .Z(n41425) );
  NOR U51194 ( .A(n41428), .B(n41425), .Z(n40561) );
  IV U51195 ( .A(n38184), .Z(n38185) );
  NOR U51196 ( .A(n38186), .B(n38185), .Z(n43938) );
  IV U51197 ( .A(n38187), .Z(n38190) );
  NOR U51198 ( .A(n38188), .B(n38192), .Z(n38189) );
  IV U51199 ( .A(n38189), .Z(n40533) );
  NOR U51200 ( .A(n38190), .B(n40533), .Z(n43927) );
  IV U51201 ( .A(n38191), .Z(n38193) );
  NOR U51202 ( .A(n38193), .B(n38192), .Z(n41444) );
  NOR U51203 ( .A(n43927), .B(n41444), .Z(n40531) );
  IV U51204 ( .A(n38194), .Z(n41450) );
  IV U51205 ( .A(n38195), .Z(n38196) );
  NOR U51206 ( .A(n38200), .B(n38196), .Z(n38197) );
  IV U51207 ( .A(n38197), .Z(n41477) );
  IV U51208 ( .A(n38198), .Z(n38199) );
  NOR U51209 ( .A(n38200), .B(n38199), .Z(n41473) );
  IV U51210 ( .A(n38201), .Z(n38203) );
  IV U51211 ( .A(n38202), .Z(n38207) );
  NOR U51212 ( .A(n38203), .B(n38207), .Z(n41478) );
  NOR U51213 ( .A(n38205), .B(n38204), .Z(n41484) );
  IV U51214 ( .A(n38206), .Z(n38208) );
  NOR U51215 ( .A(n38208), .B(n38207), .Z(n41482) );
  NOR U51216 ( .A(n41484), .B(n41482), .Z(n40501) );
  IV U51217 ( .A(n38209), .Z(n38210) );
  NOR U51218 ( .A(n38211), .B(n38210), .Z(n41500) );
  IV U51219 ( .A(n38212), .Z(n38214) );
  IV U51220 ( .A(n38213), .Z(n38218) );
  NOR U51221 ( .A(n38214), .B(n38218), .Z(n41506) );
  NOR U51222 ( .A(n41500), .B(n41506), .Z(n40477) );
  NOR U51223 ( .A(n38216), .B(n38215), .Z(n43899) );
  IV U51224 ( .A(n38217), .Z(n38219) );
  NOR U51225 ( .A(n38219), .B(n38218), .Z(n41509) );
  NOR U51226 ( .A(n43899), .B(n41509), .Z(n40476) );
  IV U51227 ( .A(n38220), .Z(n38222) );
  IV U51228 ( .A(n38221), .Z(n38228) );
  NOR U51229 ( .A(n38222), .B(n38228), .Z(n43895) );
  IV U51230 ( .A(n38223), .Z(n38225) );
  NOR U51231 ( .A(n38225), .B(n38224), .Z(n43902) );
  NOR U51232 ( .A(n43895), .B(n43902), .Z(n40475) );
  IV U51233 ( .A(n38226), .Z(n38227) );
  NOR U51234 ( .A(n38228), .B(n38227), .Z(n41511) );
  NOR U51235 ( .A(n41514), .B(n41511), .Z(n40474) );
  NOR U51236 ( .A(n38229), .B(n41517), .Z(n40473) );
  IV U51237 ( .A(n38230), .Z(n38231) );
  NOR U51238 ( .A(n38232), .B(n38231), .Z(n43889) );
  IV U51239 ( .A(n38233), .Z(n38234) );
  NOR U51240 ( .A(n40471), .B(n38234), .Z(n41524) );
  NOR U51241 ( .A(n43889), .B(n41524), .Z(n38235) );
  IV U51242 ( .A(n38235), .Z(n40472) );
  IV U51243 ( .A(n38236), .Z(n38237) );
  NOR U51244 ( .A(n38237), .B(n40456), .Z(n38238) );
  IV U51245 ( .A(n38238), .Z(n43882) );
  IV U51246 ( .A(n38239), .Z(n38240) );
  NOR U51247 ( .A(n38240), .B(n38245), .Z(n43854) );
  IV U51248 ( .A(n38241), .Z(n38242) );
  NOR U51249 ( .A(n38243), .B(n38242), .Z(n43848) );
  IV U51250 ( .A(n38244), .Z(n38246) );
  NOR U51251 ( .A(n38246), .B(n38245), .Z(n43851) );
  NOR U51252 ( .A(n43848), .B(n43851), .Z(n38247) );
  IV U51253 ( .A(n38247), .Z(n40438) );
  IV U51254 ( .A(n38248), .Z(n38249) );
  NOR U51255 ( .A(n38250), .B(n38249), .Z(n41534) );
  IV U51256 ( .A(n38251), .Z(n38254) );
  NOR U51257 ( .A(n38252), .B(n38263), .Z(n38253) );
  IV U51258 ( .A(n38253), .Z(n38256) );
  NOR U51259 ( .A(n38254), .B(n38256), .Z(n43835) );
  IV U51260 ( .A(n38255), .Z(n38257) );
  NOR U51261 ( .A(n38257), .B(n38256), .Z(n43833) );
  XOR U51262 ( .A(n43835), .B(n43833), .Z(n38258) );
  NOR U51263 ( .A(n41534), .B(n38258), .Z(n40427) );
  IV U51264 ( .A(n38259), .Z(n38261) );
  NOR U51265 ( .A(n38261), .B(n38260), .Z(n41538) );
  IV U51266 ( .A(n38262), .Z(n38264) );
  NOR U51267 ( .A(n38264), .B(n38263), .Z(n43830) );
  NOR U51268 ( .A(n41538), .B(n43830), .Z(n40426) );
  IV U51269 ( .A(n38265), .Z(n41543) );
  NOR U51270 ( .A(n38266), .B(n41543), .Z(n38270) );
  IV U51271 ( .A(n38267), .Z(n38268) );
  NOR U51272 ( .A(n38269), .B(n38268), .Z(n43826) );
  NOR U51273 ( .A(n38270), .B(n43826), .Z(n40425) );
  NOR U51274 ( .A(n38272), .B(n38271), .Z(n40423) );
  IV U51275 ( .A(n40423), .Z(n40415) );
  IV U51276 ( .A(n38273), .Z(n41549) );
  NOR U51277 ( .A(n38274), .B(n41549), .Z(n38277) );
  IV U51278 ( .A(n38275), .Z(n38276) );
  NOR U51279 ( .A(n38276), .B(n40417), .Z(n41546) );
  NOR U51280 ( .A(n38277), .B(n41546), .Z(n40413) );
  IV U51281 ( .A(n38278), .Z(n38280) );
  NOR U51282 ( .A(n38280), .B(n38279), .Z(n43819) );
  NOR U51283 ( .A(n38281), .B(n41557), .Z(n38282) );
  NOR U51284 ( .A(n43819), .B(n38282), .Z(n38283) );
  IV U51285 ( .A(n38283), .Z(n40412) );
  IV U51286 ( .A(n38284), .Z(n38286) );
  NOR U51287 ( .A(n38286), .B(n38285), .Z(n50537) );
  IV U51288 ( .A(n38287), .Z(n38289) );
  NOR U51289 ( .A(n38289), .B(n38288), .Z(n48254) );
  NOR U51290 ( .A(n50537), .B(n48254), .Z(n47127) );
  IV U51291 ( .A(n38290), .Z(n38291) );
  NOR U51292 ( .A(n38292), .B(n38291), .Z(n43814) );
  IV U51293 ( .A(n38293), .Z(n40408) );
  IV U51294 ( .A(n38294), .Z(n38295) );
  NOR U51295 ( .A(n40408), .B(n38295), .Z(n41563) );
  NOR U51296 ( .A(n43814), .B(n41563), .Z(n40411) );
  IV U51297 ( .A(n38296), .Z(n38297) );
  NOR U51298 ( .A(n38298), .B(n38297), .Z(n44868) );
  IV U51299 ( .A(n38299), .Z(n38300) );
  NOR U51300 ( .A(n38301), .B(n38300), .Z(n44861) );
  NOR U51301 ( .A(n44868), .B(n44861), .Z(n43795) );
  NOR U51302 ( .A(n38303), .B(n38302), .Z(n41575) );
  IV U51303 ( .A(n38304), .Z(n41570) );
  NOR U51304 ( .A(n38305), .B(n41570), .Z(n38306) );
  NOR U51305 ( .A(n41575), .B(n38306), .Z(n40400) );
  IV U51306 ( .A(n38307), .Z(n38309) );
  NOR U51307 ( .A(n38309), .B(n38308), .Z(n41579) );
  IV U51308 ( .A(n38310), .Z(n38311) );
  NOR U51309 ( .A(n38312), .B(n38311), .Z(n41573) );
  NOR U51310 ( .A(n41579), .B(n41573), .Z(n40399) );
  IV U51311 ( .A(n38313), .Z(n38315) );
  NOR U51312 ( .A(n38315), .B(n38314), .Z(n41595) );
  NOR U51313 ( .A(n38316), .B(n41589), .Z(n38317) );
  NOR U51314 ( .A(n41595), .B(n38317), .Z(n40391) );
  IV U51315 ( .A(n38318), .Z(n38320) );
  NOR U51316 ( .A(n38320), .B(n38319), .Z(n41603) );
  IV U51317 ( .A(n38321), .Z(n38322) );
  NOR U51318 ( .A(n38323), .B(n38322), .Z(n41598) );
  NOR U51319 ( .A(n41603), .B(n41598), .Z(n40390) );
  IV U51320 ( .A(n38324), .Z(n38325) );
  NOR U51321 ( .A(n38326), .B(n38325), .Z(n41606) );
  IV U51322 ( .A(n38327), .Z(n38329) );
  NOR U51323 ( .A(n38329), .B(n38328), .Z(n41601) );
  NOR U51324 ( .A(n41606), .B(n41601), .Z(n40389) );
  NOR U51325 ( .A(n38331), .B(n38330), .Z(n43784) );
  IV U51326 ( .A(n38332), .Z(n41611) );
  NOR U51327 ( .A(n38333), .B(n41611), .Z(n38334) );
  NOR U51328 ( .A(n43784), .B(n38334), .Z(n40388) );
  IV U51329 ( .A(n38335), .Z(n38336) );
  NOR U51330 ( .A(n38336), .B(n40382), .Z(n38337) );
  IV U51331 ( .A(n38337), .Z(n43778) );
  IV U51332 ( .A(n38338), .Z(n38340) );
  NOR U51333 ( .A(n38340), .B(n38339), .Z(n40379) );
  IV U51334 ( .A(n40379), .Z(n40369) );
  IV U51335 ( .A(n38341), .Z(n38343) );
  IV U51336 ( .A(n38342), .Z(n40362) );
  NOR U51337 ( .A(n38343), .B(n40362), .Z(n41619) );
  IV U51338 ( .A(n38344), .Z(n38345) );
  NOR U51339 ( .A(n38346), .B(n38345), .Z(n41624) );
  NOR U51340 ( .A(n38348), .B(n38347), .Z(n41622) );
  NOR U51341 ( .A(n41624), .B(n41622), .Z(n38349) );
  IV U51342 ( .A(n38349), .Z(n40360) );
  IV U51343 ( .A(n38350), .Z(n38354) );
  IV U51344 ( .A(n38351), .Z(n40350) );
  NOR U51345 ( .A(n40350), .B(n38352), .Z(n38353) );
  IV U51346 ( .A(n38353), .Z(n38356) );
  NOR U51347 ( .A(n38354), .B(n38356), .Z(n43771) );
  IV U51348 ( .A(n38355), .Z(n38357) );
  NOR U51349 ( .A(n38357), .B(n38356), .Z(n40357) );
  IV U51350 ( .A(n40357), .Z(n40349) );
  IV U51351 ( .A(n38358), .Z(n38359) );
  NOR U51352 ( .A(n38364), .B(n38359), .Z(n41650) );
  IV U51353 ( .A(n38360), .Z(n38361) );
  NOR U51354 ( .A(n38362), .B(n38361), .Z(n41657) );
  IV U51355 ( .A(n38363), .Z(n38365) );
  NOR U51356 ( .A(n38365), .B(n38364), .Z(n41649) );
  NOR U51357 ( .A(n41657), .B(n41649), .Z(n38366) );
  IV U51358 ( .A(n38366), .Z(n38367) );
  NOR U51359 ( .A(n41650), .B(n38367), .Z(n40334) );
  IV U51360 ( .A(n38368), .Z(n38369) );
  NOR U51361 ( .A(n38370), .B(n38369), .Z(n41662) );
  IV U51362 ( .A(n38371), .Z(n38373) );
  NOR U51363 ( .A(n38373), .B(n38372), .Z(n41660) );
  NOR U51364 ( .A(n41662), .B(n41660), .Z(n40333) );
  IV U51365 ( .A(n38374), .Z(n40328) );
  IV U51366 ( .A(n38375), .Z(n40324) );
  IV U51367 ( .A(n38376), .Z(n38378) );
  NOR U51368 ( .A(n38378), .B(n38377), .Z(n41687) );
  IV U51369 ( .A(n38379), .Z(n38381) );
  NOR U51370 ( .A(n38381), .B(n38380), .Z(n43755) );
  NOR U51371 ( .A(n41687), .B(n43755), .Z(n40293) );
  IV U51372 ( .A(n38382), .Z(n38384) );
  IV U51373 ( .A(n38383), .Z(n40291) );
  NOR U51374 ( .A(n38384), .B(n40291), .Z(n41684) );
  IV U51375 ( .A(n38385), .Z(n38386) );
  NOR U51376 ( .A(n38387), .B(n38386), .Z(n38388) );
  IV U51377 ( .A(n38388), .Z(n43739) );
  IV U51378 ( .A(n38389), .Z(n38390) );
  NOR U51379 ( .A(n38390), .B(n38396), .Z(n43742) );
  IV U51380 ( .A(n38391), .Z(n38392) );
  NOR U51381 ( .A(n38393), .B(n38392), .Z(n44925) );
  IV U51382 ( .A(n38394), .Z(n38395) );
  NOR U51383 ( .A(n38396), .B(n38395), .Z(n46992) );
  NOR U51384 ( .A(n44925), .B(n46992), .Z(n43732) );
  IV U51385 ( .A(n38397), .Z(n38398) );
  NOR U51386 ( .A(n40275), .B(n38398), .Z(n43719) );
  IV U51387 ( .A(n38399), .Z(n38403) );
  IV U51388 ( .A(n38400), .Z(n38401) );
  NOR U51389 ( .A(n38403), .B(n38401), .Z(n41695) );
  NOR U51390 ( .A(n43719), .B(n41695), .Z(n40268) );
  IV U51391 ( .A(n38402), .Z(n38406) );
  NOR U51392 ( .A(n38404), .B(n38403), .Z(n38405) );
  IV U51393 ( .A(n38405), .Z(n40266) );
  NOR U51394 ( .A(n38406), .B(n40266), .Z(n41700) );
  NOR U51395 ( .A(n38407), .B(n41705), .Z(n40264) );
  IV U51396 ( .A(n38408), .Z(n38410) );
  IV U51397 ( .A(n38409), .Z(n40247) );
  NOR U51398 ( .A(n38410), .B(n40247), .Z(n43709) );
  IV U51399 ( .A(n38411), .Z(n38414) );
  IV U51400 ( .A(n38412), .Z(n38413) );
  NOR U51401 ( .A(n38414), .B(n38413), .Z(n41723) );
  IV U51402 ( .A(n38415), .Z(n38417) );
  IV U51403 ( .A(n38416), .Z(n38423) );
  NOR U51404 ( .A(n38417), .B(n38423), .Z(n43694) );
  NOR U51405 ( .A(n38419), .B(n38418), .Z(n43698) );
  NOR U51406 ( .A(n43694), .B(n43698), .Z(n40242) );
  IV U51407 ( .A(n38420), .Z(n38421) );
  NOR U51408 ( .A(n38421), .B(n38430), .Z(n46923) );
  IV U51409 ( .A(n38422), .Z(n38424) );
  NOR U51410 ( .A(n38424), .B(n38423), .Z(n46941) );
  NOR U51411 ( .A(n46923), .B(n46941), .Z(n43693) );
  IV U51412 ( .A(n38425), .Z(n38426) );
  NOR U51413 ( .A(n38427), .B(n38426), .Z(n41726) );
  IV U51414 ( .A(n38428), .Z(n38429) );
  NOR U51415 ( .A(n38430), .B(n38429), .Z(n43689) );
  NOR U51416 ( .A(n41726), .B(n43689), .Z(n40241) );
  IV U51417 ( .A(n38431), .Z(n38432) );
  NOR U51418 ( .A(n38433), .B(n38432), .Z(n38434) );
  IV U51419 ( .A(n38434), .Z(n40237) );
  IV U51420 ( .A(n38435), .Z(n40215) );
  IV U51421 ( .A(n38438), .Z(n38436) );
  NOR U51422 ( .A(n40215), .B(n38436), .Z(n43669) );
  IV U51423 ( .A(n38437), .Z(n38443) );
  XOR U51424 ( .A(n38438), .B(n40215), .Z(n38439) );
  NOR U51425 ( .A(n38440), .B(n38439), .Z(n38441) );
  IV U51426 ( .A(n38441), .Z(n38442) );
  NOR U51427 ( .A(n38443), .B(n38442), .Z(n43666) );
  NOR U51428 ( .A(n43669), .B(n43666), .Z(n41742) );
  IV U51429 ( .A(n38444), .Z(n38446) );
  NOR U51430 ( .A(n38446), .B(n38445), .Z(n38447) );
  IV U51431 ( .A(n38447), .Z(n40209) );
  IV U51432 ( .A(n38448), .Z(n38449) );
  NOR U51433 ( .A(n38449), .B(n38451), .Z(n43651) );
  IV U51434 ( .A(n43651), .Z(n43649) );
  IV U51435 ( .A(n38450), .Z(n38452) );
  NOR U51436 ( .A(n38452), .B(n38451), .Z(n43644) );
  IV U51437 ( .A(n38453), .Z(n38455) );
  IV U51438 ( .A(n38454), .Z(n40201) );
  NOR U51439 ( .A(n38455), .B(n40201), .Z(n43641) );
  IV U51440 ( .A(n38456), .Z(n41751) );
  IV U51441 ( .A(n38457), .Z(n38458) );
  NOR U51442 ( .A(n38459), .B(n38458), .Z(n41748) );
  IV U51443 ( .A(n38460), .Z(n38461) );
  NOR U51444 ( .A(n38462), .B(n38461), .Z(n44973) );
  IV U51445 ( .A(n38463), .Z(n38464) );
  NOR U51446 ( .A(n38465), .B(n38464), .Z(n46868) );
  NOR U51447 ( .A(n44973), .B(n46868), .Z(n41762) );
  NOR U51448 ( .A(n38467), .B(n38466), .Z(n41759) );
  IV U51449 ( .A(n38468), .Z(n38469) );
  NOR U51450 ( .A(n38470), .B(n38469), .Z(n43627) );
  NOR U51451 ( .A(n43627), .B(n41764), .Z(n40192) );
  IV U51452 ( .A(n38471), .Z(n40186) );
  IV U51453 ( .A(n38472), .Z(n38473) );
  NOR U51454 ( .A(n40186), .B(n38473), .Z(n41768) );
  IV U51455 ( .A(n38474), .Z(n38476) );
  NOR U51456 ( .A(n38476), .B(n38475), .Z(n43630) );
  NOR U51457 ( .A(n41768), .B(n43630), .Z(n40191) );
  IV U51458 ( .A(n38477), .Z(n38479) );
  IV U51459 ( .A(n38478), .Z(n38485) );
  NOR U51460 ( .A(n38479), .B(n38485), .Z(n43619) );
  IV U51461 ( .A(n38480), .Z(n38481) );
  NOR U51462 ( .A(n38481), .B(n40189), .Z(n43624) );
  NOR U51463 ( .A(n43619), .B(n43624), .Z(n40183) );
  IV U51464 ( .A(n38482), .Z(n38483) );
  NOR U51465 ( .A(n38483), .B(n38491), .Z(n44988) );
  IV U51466 ( .A(n38484), .Z(n38486) );
  NOR U51467 ( .A(n38486), .B(n38485), .Z(n44984) );
  NOR U51468 ( .A(n44988), .B(n44984), .Z(n43618) );
  IV U51469 ( .A(n38487), .Z(n38489) );
  NOR U51470 ( .A(n38489), .B(n38488), .Z(n41778) );
  IV U51471 ( .A(n38490), .Z(n38492) );
  NOR U51472 ( .A(n38492), .B(n38491), .Z(n41774) );
  NOR U51473 ( .A(n41778), .B(n41774), .Z(n40182) );
  IV U51474 ( .A(n38493), .Z(n38494) );
  NOR U51475 ( .A(n38495), .B(n38494), .Z(n41781) );
  NOR U51476 ( .A(n38496), .B(n41781), .Z(n40181) );
  IV U51477 ( .A(n38497), .Z(n38498) );
  NOR U51478 ( .A(n38498), .B(n40177), .Z(n41794) );
  NOR U51479 ( .A(n41794), .B(n41789), .Z(n40180) );
  IV U51480 ( .A(n38499), .Z(n40175) );
  IV U51481 ( .A(n38500), .Z(n38501) );
  NOR U51482 ( .A(n40175), .B(n38501), .Z(n43605) );
  IV U51483 ( .A(n38502), .Z(n38503) );
  NOR U51484 ( .A(n40171), .B(n38503), .Z(n43608) );
  IV U51485 ( .A(n38504), .Z(n38505) );
  NOR U51486 ( .A(n38506), .B(n38505), .Z(n43602) );
  IV U51487 ( .A(n38507), .Z(n38509) );
  NOR U51488 ( .A(n38509), .B(n38508), .Z(n41805) );
  NOR U51489 ( .A(n43602), .B(n41805), .Z(n38510) );
  IV U51490 ( .A(n38510), .Z(n40169) );
  IV U51491 ( .A(n38511), .Z(n38522) );
  IV U51492 ( .A(n38512), .Z(n38513) );
  NOR U51493 ( .A(n38522), .B(n38513), .Z(n43598) );
  IV U51494 ( .A(n38514), .Z(n38515) );
  NOR U51495 ( .A(n38522), .B(n38515), .Z(n43595) );
  IV U51496 ( .A(n38516), .Z(n38517) );
  NOR U51497 ( .A(n38522), .B(n38517), .Z(n38518) );
  IV U51498 ( .A(n38518), .Z(n38519) );
  NOR U51499 ( .A(n38520), .B(n38519), .Z(n41807) );
  IV U51500 ( .A(n38520), .Z(n38525) );
  NOR U51501 ( .A(n38522), .B(n38521), .Z(n38523) );
  IV U51502 ( .A(n38523), .Z(n38524) );
  NOR U51503 ( .A(n38525), .B(n38524), .Z(n43591) );
  IV U51504 ( .A(n38526), .Z(n38528) );
  NOR U51505 ( .A(n38528), .B(n38527), .Z(n43588) );
  IV U51506 ( .A(n38529), .Z(n38530) );
  NOR U51507 ( .A(n40164), .B(n38530), .Z(n43584) );
  IV U51508 ( .A(n38531), .Z(n38532) );
  NOR U51509 ( .A(n38532), .B(n40159), .Z(n41819) );
  IV U51510 ( .A(n38533), .Z(n38535) );
  IV U51511 ( .A(n38534), .Z(n40166) );
  NOR U51512 ( .A(n38535), .B(n40166), .Z(n41814) );
  NOR U51513 ( .A(n41819), .B(n41814), .Z(n40161) );
  IV U51514 ( .A(n38536), .Z(n38538) );
  NOR U51515 ( .A(n38538), .B(n38537), .Z(n38539) );
  IV U51516 ( .A(n38539), .Z(n40153) );
  IV U51517 ( .A(n38540), .Z(n38543) );
  NOR U51518 ( .A(n38541), .B(n38548), .Z(n38542) );
  IV U51519 ( .A(n38542), .Z(n38545) );
  NOR U51520 ( .A(n38543), .B(n38545), .Z(n41832) );
  IV U51521 ( .A(n38544), .Z(n38546) );
  NOR U51522 ( .A(n38546), .B(n38545), .Z(n41844) );
  IV U51523 ( .A(n38547), .Z(n38549) );
  NOR U51524 ( .A(n38549), .B(n38548), .Z(n41841) );
  IV U51525 ( .A(n38550), .Z(n38552) );
  IV U51526 ( .A(n38551), .Z(n38555) );
  NOR U51527 ( .A(n38552), .B(n38555), .Z(n41847) );
  NOR U51528 ( .A(n38553), .B(n43571), .Z(n38557) );
  IV U51529 ( .A(n38554), .Z(n38556) );
  NOR U51530 ( .A(n38556), .B(n38555), .Z(n41850) );
  NOR U51531 ( .A(n38557), .B(n41850), .Z(n40145) );
  IV U51532 ( .A(n38558), .Z(n43563) );
  NOR U51533 ( .A(n38559), .B(n43563), .Z(n40144) );
  IV U51534 ( .A(n38560), .Z(n38561) );
  NOR U51535 ( .A(n38562), .B(n38561), .Z(n43552) );
  NOR U51536 ( .A(n38563), .B(n43556), .Z(n38564) );
  NOR U51537 ( .A(n43552), .B(n38564), .Z(n38565) );
  IV U51538 ( .A(n38565), .Z(n40143) );
  IV U51539 ( .A(n38566), .Z(n38569) );
  IV U51540 ( .A(n38567), .Z(n38568) );
  NOR U51541 ( .A(n38569), .B(n38568), .Z(n41856) );
  IV U51542 ( .A(n38570), .Z(n38571) );
  NOR U51543 ( .A(n38571), .B(n38576), .Z(n43545) );
  NOR U51544 ( .A(n43545), .B(n41854), .Z(n40142) );
  IV U51545 ( .A(n38572), .Z(n38574) );
  NOR U51546 ( .A(n38574), .B(n38573), .Z(n43543) );
  IV U51547 ( .A(n38575), .Z(n38577) );
  NOR U51548 ( .A(n38577), .B(n38576), .Z(n43548) );
  NOR U51549 ( .A(n43543), .B(n43548), .Z(n40141) );
  IV U51550 ( .A(n38578), .Z(n38579) );
  NOR U51551 ( .A(n38580), .B(n38579), .Z(n41862) );
  IV U51552 ( .A(n38581), .Z(n38587) );
  IV U51553 ( .A(n38582), .Z(n38583) );
  NOR U51554 ( .A(n38587), .B(n38583), .Z(n38584) );
  IV U51555 ( .A(n38584), .Z(n43534) );
  IV U51556 ( .A(n38585), .Z(n38586) );
  NOR U51557 ( .A(n38587), .B(n38586), .Z(n41865) );
  IV U51558 ( .A(n38588), .Z(n38594) );
  NOR U51559 ( .A(n38589), .B(n38605), .Z(n38590) );
  IV U51560 ( .A(n38590), .Z(n38591) );
  NOR U51561 ( .A(n38592), .B(n38591), .Z(n38593) );
  IV U51562 ( .A(n38593), .Z(n38599) );
  NOR U51563 ( .A(n38594), .B(n38599), .Z(n41869) );
  IV U51564 ( .A(n38595), .Z(n38596) );
  NOR U51565 ( .A(n38597), .B(n38596), .Z(n43522) );
  IV U51566 ( .A(n38598), .Z(n38600) );
  NOR U51567 ( .A(n38600), .B(n38599), .Z(n43529) );
  NOR U51568 ( .A(n43522), .B(n43529), .Z(n40126) );
  IV U51569 ( .A(n38601), .Z(n38603) );
  NOR U51570 ( .A(n38603), .B(n38602), .Z(n43518) );
  IV U51571 ( .A(n38604), .Z(n38606) );
  NOR U51572 ( .A(n38606), .B(n38605), .Z(n43525) );
  NOR U51573 ( .A(n43518), .B(n43525), .Z(n40125) );
  NOR U51574 ( .A(n38607), .B(n41877), .Z(n40124) );
  IV U51575 ( .A(n38608), .Z(n38609) );
  NOR U51576 ( .A(n38610), .B(n38609), .Z(n43506) );
  IV U51577 ( .A(n38611), .Z(n38612) );
  NOR U51578 ( .A(n38613), .B(n38612), .Z(n43511) );
  NOR U51579 ( .A(n43506), .B(n43511), .Z(n40123) );
  IV U51580 ( .A(n38614), .Z(n45081) );
  NOR U51581 ( .A(n38615), .B(n45081), .Z(n38616) );
  IV U51582 ( .A(n38616), .Z(n41883) );
  IV U51583 ( .A(n38617), .Z(n38618) );
  NOR U51584 ( .A(n38618), .B(n40074), .Z(n40071) );
  IV U51585 ( .A(n40071), .Z(n40061) );
  IV U51586 ( .A(n38619), .Z(n38621) );
  IV U51587 ( .A(n38620), .Z(n38627) );
  NOR U51588 ( .A(n38621), .B(n38627), .Z(n41911) );
  IV U51589 ( .A(n38622), .Z(n38625) );
  IV U51590 ( .A(n38623), .Z(n38624) );
  NOR U51591 ( .A(n38625), .B(n38624), .Z(n43474) );
  IV U51592 ( .A(n38626), .Z(n38628) );
  NOR U51593 ( .A(n38628), .B(n38627), .Z(n41909) );
  NOR U51594 ( .A(n43474), .B(n41909), .Z(n38629) );
  IV U51595 ( .A(n38629), .Z(n40052) );
  IV U51596 ( .A(n38630), .Z(n38631) );
  NOR U51597 ( .A(n38632), .B(n38631), .Z(n43471) );
  IV U51598 ( .A(n38633), .Z(n38635) );
  NOR U51599 ( .A(n38635), .B(n38634), .Z(n38636) );
  IV U51600 ( .A(n38636), .Z(n41920) );
  IV U51601 ( .A(n38637), .Z(n38639) );
  NOR U51602 ( .A(n38639), .B(n38638), .Z(n41923) );
  IV U51603 ( .A(n38640), .Z(n38642) );
  NOR U51604 ( .A(n38642), .B(n38641), .Z(n41921) );
  NOR U51605 ( .A(n41923), .B(n41921), .Z(n38643) );
  IV U51606 ( .A(n38643), .Z(n40043) );
  IV U51607 ( .A(n38644), .Z(n38646) );
  NOR U51608 ( .A(n38646), .B(n38645), .Z(n43463) );
  IV U51609 ( .A(n38647), .Z(n38648) );
  NOR U51610 ( .A(n38649), .B(n38648), .Z(n43465) );
  NOR U51611 ( .A(n43463), .B(n43465), .Z(n40042) );
  IV U51612 ( .A(n38650), .Z(n38651) );
  NOR U51613 ( .A(n38652), .B(n38651), .Z(n41926) );
  IV U51614 ( .A(n38653), .Z(n38655) );
  NOR U51615 ( .A(n38655), .B(n38654), .Z(n43459) );
  NOR U51616 ( .A(n41926), .B(n43459), .Z(n40041) );
  IV U51617 ( .A(n38656), .Z(n45145) );
  NOR U51618 ( .A(n38657), .B(n45145), .Z(n41931) );
  IV U51619 ( .A(n38658), .Z(n38659) );
  NOR U51620 ( .A(n38659), .B(n40033), .Z(n41933) );
  NOR U51621 ( .A(n41928), .B(n41933), .Z(n40039) );
  NOR U51622 ( .A(n40029), .B(n40027), .Z(n40024) );
  NOR U51623 ( .A(n38660), .B(n41964), .Z(n40025) );
  IV U51624 ( .A(n38661), .Z(n41957) );
  NOR U51625 ( .A(n38662), .B(n41957), .Z(n41950) );
  NOR U51626 ( .A(n40025), .B(n41950), .Z(n40023) );
  IV U51627 ( .A(n38663), .Z(n38664) );
  NOR U51628 ( .A(n38665), .B(n38664), .Z(n40020) );
  IV U51629 ( .A(n40020), .Z(n40011) );
  IV U51630 ( .A(n38666), .Z(n38667) );
  NOR U51631 ( .A(n38668), .B(n38667), .Z(n43442) );
  IV U51632 ( .A(n38669), .Z(n38670) );
  NOR U51633 ( .A(n38670), .B(n39967), .Z(n43414) );
  IV U51634 ( .A(n38671), .Z(n38672) );
  NOR U51635 ( .A(n38672), .B(n38677), .Z(n42021) );
  IV U51636 ( .A(n38673), .Z(n38674) );
  NOR U51637 ( .A(n38675), .B(n38674), .Z(n48710) );
  IV U51638 ( .A(n38676), .Z(n38678) );
  NOR U51639 ( .A(n38678), .B(n38677), .Z(n50035) );
  NOR U51640 ( .A(n48710), .B(n50035), .Z(n42031) );
  IV U51641 ( .A(n38679), .Z(n38680) );
  NOR U51642 ( .A(n38681), .B(n38680), .Z(n42032) );
  IV U51643 ( .A(n38682), .Z(n38684) );
  NOR U51644 ( .A(n38684), .B(n38683), .Z(n42028) );
  NOR U51645 ( .A(n42032), .B(n42028), .Z(n39924) );
  IV U51646 ( .A(n38685), .Z(n38687) );
  IV U51647 ( .A(n38686), .Z(n38692) );
  NOR U51648 ( .A(n38687), .B(n38692), .Z(n43383) );
  NOR U51649 ( .A(n38689), .B(n38688), .Z(n43376) );
  IV U51650 ( .A(n38690), .Z(n38691) );
  NOR U51651 ( .A(n38692), .B(n38691), .Z(n43379) );
  NOR U51652 ( .A(n43376), .B(n43379), .Z(n38693) );
  IV U51653 ( .A(n38693), .Z(n39917) );
  IV U51654 ( .A(n38694), .Z(n38696) );
  NOR U51655 ( .A(n38696), .B(n38695), .Z(n42038) );
  IV U51656 ( .A(n38697), .Z(n38699) );
  NOR U51657 ( .A(n38699), .B(n38698), .Z(n38700) );
  IV U51658 ( .A(n38700), .Z(n39909) );
  IV U51659 ( .A(n38701), .Z(n38702) );
  NOR U51660 ( .A(n38703), .B(n38702), .Z(n42054) );
  NOR U51661 ( .A(n42054), .B(n42048), .Z(n39893) );
  IV U51662 ( .A(n39879), .Z(n39877) );
  IV U51663 ( .A(n38704), .Z(n39885) );
  IV U51664 ( .A(n38705), .Z(n38707) );
  NOR U51665 ( .A(n38707), .B(n38706), .Z(n43361) );
  NOR U51666 ( .A(n38709), .B(n38708), .Z(n42060) );
  NOR U51667 ( .A(n43361), .B(n42060), .Z(n39874) );
  IV U51668 ( .A(n38710), .Z(n39868) );
  IV U51669 ( .A(n38711), .Z(n38712) );
  NOR U51670 ( .A(n39868), .B(n38712), .Z(n43356) );
  IV U51671 ( .A(n38713), .Z(n38715) );
  NOR U51672 ( .A(n38715), .B(n38714), .Z(n43358) );
  NOR U51673 ( .A(n43356), .B(n43358), .Z(n39873) );
  IV U51674 ( .A(n38716), .Z(n38717) );
  NOR U51675 ( .A(n38718), .B(n38717), .Z(n38719) );
  IV U51676 ( .A(n38719), .Z(n39862) );
  IV U51677 ( .A(n38720), .Z(n42076) );
  NOR U51678 ( .A(n38721), .B(n42076), .Z(n38722) );
  NOR U51679 ( .A(n42082), .B(n38722), .Z(n39855) );
  IV U51680 ( .A(n38723), .Z(n43353) );
  IV U51681 ( .A(n38725), .Z(n38727) );
  IV U51682 ( .A(n38726), .Z(n39853) );
  NOR U51683 ( .A(n38727), .B(n39853), .Z(n39847) );
  IV U51684 ( .A(n38728), .Z(n38731) );
  IV U51685 ( .A(n38729), .Z(n38730) );
  NOR U51686 ( .A(n38731), .B(n38730), .Z(n43337) );
  NOR U51687 ( .A(n38732), .B(n43333), .Z(n42092) );
  NOR U51688 ( .A(n43337), .B(n42092), .Z(n38733) );
  IV U51689 ( .A(n38733), .Z(n39842) );
  IV U51690 ( .A(n38734), .Z(n38736) );
  NOR U51691 ( .A(n38736), .B(n38735), .Z(n38737) );
  IV U51692 ( .A(n38737), .Z(n42108) );
  IV U51693 ( .A(n38738), .Z(n38740) );
  NOR U51694 ( .A(n38740), .B(n38739), .Z(n42117) );
  IV U51695 ( .A(n38741), .Z(n38743) );
  NOR U51696 ( .A(n38743), .B(n38742), .Z(n42114) );
  NOR U51697 ( .A(n42117), .B(n42114), .Z(n38744) );
  IV U51698 ( .A(n38744), .Z(n39830) );
  IV U51699 ( .A(n38745), .Z(n38746) );
  NOR U51700 ( .A(n38747), .B(n38746), .Z(n42119) );
  IV U51701 ( .A(n38748), .Z(n39827) );
  IV U51702 ( .A(n38749), .Z(n38750) );
  NOR U51703 ( .A(n39827), .B(n38750), .Z(n43326) );
  IV U51704 ( .A(n38751), .Z(n38752) );
  NOR U51705 ( .A(n38756), .B(n38752), .Z(n38753) );
  IV U51706 ( .A(n38753), .Z(n43318) );
  IV U51707 ( .A(n38754), .Z(n38755) );
  NOR U51708 ( .A(n38756), .B(n38755), .Z(n43313) );
  IV U51709 ( .A(n38757), .Z(n38759) );
  IV U51710 ( .A(n38758), .Z(n38763) );
  NOR U51711 ( .A(n38759), .B(n38763), .Z(n43310) );
  IV U51712 ( .A(n38760), .Z(n38761) );
  NOR U51713 ( .A(n38761), .B(n38769), .Z(n42123) );
  IV U51714 ( .A(n38762), .Z(n38764) );
  NOR U51715 ( .A(n38764), .B(n38763), .Z(n43307) );
  NOR U51716 ( .A(n42123), .B(n43307), .Z(n39823) );
  IV U51717 ( .A(n38765), .Z(n38767) );
  NOR U51718 ( .A(n38767), .B(n38766), .Z(n48818) );
  IV U51719 ( .A(n38768), .Z(n38770) );
  NOR U51720 ( .A(n38770), .B(n38769), .Z(n48805) );
  NOR U51721 ( .A(n48818), .B(n48805), .Z(n42122) );
  IV U51722 ( .A(n38771), .Z(n38772) );
  NOR U51723 ( .A(n43294), .B(n38772), .Z(n42128) );
  IV U51724 ( .A(n38773), .Z(n38775) );
  NOR U51725 ( .A(n38775), .B(n38774), .Z(n43290) );
  IV U51726 ( .A(n38776), .Z(n38777) );
  NOR U51727 ( .A(n38778), .B(n38777), .Z(n43303) );
  NOR U51728 ( .A(n43290), .B(n43303), .Z(n39822) );
  IV U51729 ( .A(n38779), .Z(n38783) );
  IV U51730 ( .A(n38780), .Z(n39802) );
  NOR U51731 ( .A(n38781), .B(n39802), .Z(n38782) );
  IV U51732 ( .A(n38782), .Z(n39799) );
  NOR U51733 ( .A(n38783), .B(n39799), .Z(n43281) );
  NOR U51734 ( .A(n38785), .B(n38784), .Z(n42135) );
  NOR U51735 ( .A(n38787), .B(n38786), .Z(n43276) );
  NOR U51736 ( .A(n42141), .B(n43276), .Z(n39797) );
  IV U51737 ( .A(n38788), .Z(n38789) );
  NOR U51738 ( .A(n38789), .B(n42151), .Z(n42146) );
  NOR U51739 ( .A(n42146), .B(n42144), .Z(n39796) );
  NOR U51740 ( .A(n38790), .B(n42160), .Z(n38793) );
  NOR U51741 ( .A(n38791), .B(n42151), .Z(n38792) );
  NOR U51742 ( .A(n38793), .B(n38792), .Z(n39795) );
  IV U51743 ( .A(n38794), .Z(n39790) );
  IV U51744 ( .A(n38795), .Z(n38796) );
  NOR U51745 ( .A(n39790), .B(n38796), .Z(n43268) );
  IV U51746 ( .A(n38797), .Z(n38798) );
  NOR U51747 ( .A(n38799), .B(n38798), .Z(n38800) );
  IV U51748 ( .A(n38800), .Z(n42180) );
  IV U51749 ( .A(n38801), .Z(n39773) );
  IV U51750 ( .A(n38802), .Z(n38803) );
  NOR U51751 ( .A(n39773), .B(n38803), .Z(n38804) );
  IV U51752 ( .A(n38804), .Z(n43262) );
  IV U51753 ( .A(n38805), .Z(n38806) );
  NOR U51754 ( .A(n38806), .B(n39766), .Z(n42185) );
  IV U51755 ( .A(n38807), .Z(n38808) );
  NOR U51756 ( .A(n38808), .B(n38816), .Z(n43252) );
  IV U51757 ( .A(n38809), .Z(n38810) );
  NOR U51758 ( .A(n38811), .B(n38810), .Z(n43255) );
  NOR U51759 ( .A(n43252), .B(n43255), .Z(n39764) );
  IV U51760 ( .A(n38812), .Z(n38814) );
  NOR U51761 ( .A(n38814), .B(n38813), .Z(n42189) );
  IV U51762 ( .A(n38815), .Z(n38817) );
  NOR U51763 ( .A(n38817), .B(n38816), .Z(n43249) );
  NOR U51764 ( .A(n42189), .B(n43249), .Z(n39763) );
  IV U51765 ( .A(n38818), .Z(n38819) );
  NOR U51766 ( .A(n38820), .B(n38819), .Z(n43235) );
  IV U51767 ( .A(n38821), .Z(n38824) );
  IV U51768 ( .A(n38822), .Z(n38823) );
  NOR U51769 ( .A(n38824), .B(n38823), .Z(n43240) );
  NOR U51770 ( .A(n43235), .B(n43240), .Z(n39751) );
  NOR U51771 ( .A(n43224), .B(n38825), .Z(n42200) );
  IV U51772 ( .A(n38826), .Z(n38828) );
  XOR U51773 ( .A(n42210), .B(n42211), .Z(n38827) );
  NOR U51774 ( .A(n38828), .B(n38827), .Z(n43216) );
  NOR U51775 ( .A(n38829), .B(n38832), .Z(n39746) );
  IV U51776 ( .A(n38830), .Z(n38831) );
  NOR U51777 ( .A(n38832), .B(n38831), .Z(n42216) );
  IV U51778 ( .A(n38833), .Z(n38834) );
  NOR U51779 ( .A(n39743), .B(n38834), .Z(n43213) );
  NOR U51780 ( .A(n42216), .B(n43213), .Z(n38835) );
  IV U51781 ( .A(n38835), .Z(n39745) );
  IV U51782 ( .A(n38836), .Z(n38837) );
  NOR U51783 ( .A(n38837), .B(n39743), .Z(n42218) );
  IV U51784 ( .A(n38840), .Z(n38839) );
  IV U51785 ( .A(n38838), .Z(n39740) );
  NOR U51786 ( .A(n38839), .B(n39740), .Z(n46399) );
  XOR U51787 ( .A(n38840), .B(n39740), .Z(n38843) );
  IV U51788 ( .A(n38841), .Z(n38842) );
  NOR U51789 ( .A(n38843), .B(n38842), .Z(n46405) );
  NOR U51790 ( .A(n46399), .B(n46405), .Z(n42221) );
  NOR U51791 ( .A(n38844), .B(n42228), .Z(n39738) );
  IV U51792 ( .A(n38845), .Z(n38847) );
  NOR U51793 ( .A(n38847), .B(n38846), .Z(n39728) );
  IV U51794 ( .A(n38848), .Z(n38849) );
  NOR U51795 ( .A(n38850), .B(n38849), .Z(n38851) );
  IV U51796 ( .A(n38851), .Z(n43205) );
  IV U51797 ( .A(n38852), .Z(n38853) );
  NOR U51798 ( .A(n38858), .B(n38853), .Z(n43201) );
  IV U51799 ( .A(n38854), .Z(n38856) );
  NOR U51800 ( .A(n38856), .B(n38855), .Z(n42240) );
  IV U51801 ( .A(n38857), .Z(n38859) );
  NOR U51802 ( .A(n38859), .B(n38858), .Z(n42235) );
  NOR U51803 ( .A(n42240), .B(n42235), .Z(n38860) );
  IV U51804 ( .A(n38860), .Z(n39722) );
  IV U51805 ( .A(n38861), .Z(n38862) );
  NOR U51806 ( .A(n38863), .B(n38862), .Z(n42237) );
  IV U51807 ( .A(n38864), .Z(n38865) );
  NOR U51808 ( .A(n43187), .B(n38865), .Z(n42246) );
  IV U51809 ( .A(n38866), .Z(n38869) );
  NOR U51810 ( .A(n43187), .B(n38867), .Z(n38868) );
  IV U51811 ( .A(n38868), .Z(n38871) );
  NOR U51812 ( .A(n38869), .B(n38871), .Z(n42243) );
  IV U51813 ( .A(n38870), .Z(n38872) );
  NOR U51814 ( .A(n38872), .B(n38871), .Z(n39721) );
  IV U51815 ( .A(n38873), .Z(n38874) );
  NOR U51816 ( .A(n38875), .B(n38874), .Z(n38876) );
  IV U51817 ( .A(n38876), .Z(n43174) );
  IV U51818 ( .A(n38877), .Z(n38879) );
  IV U51819 ( .A(n38878), .Z(n38881) );
  NOR U51820 ( .A(n38879), .B(n38881), .Z(n43175) );
  IV U51821 ( .A(n38880), .Z(n38882) );
  NOR U51822 ( .A(n38882), .B(n38881), .Z(n42254) );
  NOR U51823 ( .A(n42260), .B(n42254), .Z(n38883) );
  IV U51824 ( .A(n38883), .Z(n39711) );
  IV U51825 ( .A(n38884), .Z(n38885) );
  NOR U51826 ( .A(n38885), .B(n38892), .Z(n42277) );
  NOR U51827 ( .A(n38887), .B(n38886), .Z(n42275) );
  NOR U51828 ( .A(n42277), .B(n42275), .Z(n39687) );
  IV U51829 ( .A(n38888), .Z(n38889) );
  NOR U51830 ( .A(n38890), .B(n38889), .Z(n43162) );
  IV U51831 ( .A(n38891), .Z(n38893) );
  NOR U51832 ( .A(n38893), .B(n38892), .Z(n42281) );
  NOR U51833 ( .A(n43162), .B(n42281), .Z(n39686) );
  IV U51834 ( .A(n38894), .Z(n38897) );
  IV U51835 ( .A(n38895), .Z(n38896) );
  NOR U51836 ( .A(n38897), .B(n38896), .Z(n43165) );
  IV U51837 ( .A(n38898), .Z(n38901) );
  NOR U51838 ( .A(n38899), .B(n38905), .Z(n38900) );
  IV U51839 ( .A(n38900), .Z(n38903) );
  NOR U51840 ( .A(n38901), .B(n38903), .Z(n43160) );
  NOR U51841 ( .A(n43165), .B(n43160), .Z(n39685) );
  IV U51842 ( .A(n38902), .Z(n38904) );
  NOR U51843 ( .A(n38904), .B(n38903), .Z(n42283) );
  NOR U51844 ( .A(n38906), .B(n38905), .Z(n43153) );
  IV U51845 ( .A(n38907), .Z(n38909) );
  NOR U51846 ( .A(n38909), .B(n38908), .Z(n38910) );
  IV U51847 ( .A(n38910), .Z(n43141) );
  IV U51848 ( .A(n38911), .Z(n38912) );
  NOR U51849 ( .A(n39674), .B(n38912), .Z(n42290) );
  IV U51850 ( .A(n38913), .Z(n38916) );
  NOR U51851 ( .A(n38914), .B(n39666), .Z(n38915) );
  IV U51852 ( .A(n38915), .Z(n38928) );
  NOR U51853 ( .A(n38916), .B(n38928), .Z(n45444) );
  NOR U51854 ( .A(n39667), .B(n39666), .Z(n38917) );
  IV U51855 ( .A(n38917), .Z(n38918) );
  NOR U51856 ( .A(n38919), .B(n38918), .Z(n38920) );
  IV U51857 ( .A(n38920), .Z(n38921) );
  NOR U51858 ( .A(n38922), .B(n38921), .Z(n38923) );
  IV U51859 ( .A(n38923), .Z(n39658) );
  NOR U51860 ( .A(n38924), .B(n39658), .Z(n46302) );
  NOR U51861 ( .A(n45444), .B(n46302), .Z(n42311) );
  IV U51862 ( .A(n38925), .Z(n38926) );
  IV U51863 ( .A(n42321), .Z(n42315) );
  NOR U51864 ( .A(n38926), .B(n42315), .Z(n38930) );
  IV U51865 ( .A(n38927), .Z(n38929) );
  NOR U51866 ( .A(n38929), .B(n38928), .Z(n42312) );
  NOR U51867 ( .A(n38930), .B(n42312), .Z(n39656) );
  IV U51868 ( .A(n38931), .Z(n38934) );
  IV U51869 ( .A(n38932), .Z(n38933) );
  NOR U51870 ( .A(n38934), .B(n38933), .Z(n42335) );
  IV U51871 ( .A(n42322), .Z(n38935) );
  NOR U51872 ( .A(n38935), .B(n42315), .Z(n43134) );
  NOR U51873 ( .A(n42335), .B(n43134), .Z(n39655) );
  IV U51874 ( .A(n39653), .Z(n39648) );
  IV U51875 ( .A(n38936), .Z(n38937) );
  NOR U51876 ( .A(n38941), .B(n38937), .Z(n38938) );
  IV U51877 ( .A(n38938), .Z(n42346) );
  IV U51878 ( .A(n38939), .Z(n38940) );
  NOR U51879 ( .A(n38941), .B(n38940), .Z(n42342) );
  IV U51880 ( .A(n39641), .Z(n38942) );
  NOR U51881 ( .A(n38943), .B(n38942), .Z(n38944) );
  IV U51882 ( .A(n38944), .Z(n38949) );
  IV U51883 ( .A(n38945), .Z(n39637) );
  NOR U51884 ( .A(n39637), .B(n38946), .Z(n38947) );
  IV U51885 ( .A(n38947), .Z(n38948) );
  NOR U51886 ( .A(n38949), .B(n38948), .Z(n43118) );
  IV U51887 ( .A(n38950), .Z(n38953) );
  IV U51888 ( .A(n38951), .Z(n38952) );
  NOR U51889 ( .A(n38953), .B(n38952), .Z(n45486) );
  IV U51890 ( .A(n38954), .Z(n38955) );
  NOR U51891 ( .A(n38955), .B(n39637), .Z(n45481) );
  NOR U51892 ( .A(n45486), .B(n45481), .Z(n42347) );
  IV U51893 ( .A(n42347), .Z(n39635) );
  IV U51894 ( .A(n38956), .Z(n38958) );
  NOR U51895 ( .A(n38958), .B(n38957), .Z(n42349) );
  NOR U51896 ( .A(n38960), .B(n38959), .Z(n43109) );
  NOR U51897 ( .A(n42349), .B(n43109), .Z(n43114) );
  IV U51898 ( .A(n43114), .Z(n38961) );
  NOR U51899 ( .A(n43112), .B(n38961), .Z(n39634) );
  NOR U51900 ( .A(n38962), .B(n43100), .Z(n39633) );
  IV U51901 ( .A(n38963), .Z(n38964) );
  NOR U51902 ( .A(n39628), .B(n38964), .Z(n42351) );
  IV U51903 ( .A(n38965), .Z(n38967) );
  IV U51904 ( .A(n38966), .Z(n39615) );
  NOR U51905 ( .A(n38967), .B(n39615), .Z(n42356) );
  IV U51906 ( .A(n38968), .Z(n38972) );
  NOR U51907 ( .A(n38970), .B(n38969), .Z(n38971) );
  IV U51908 ( .A(n38971), .Z(n39612) );
  NOR U51909 ( .A(n38972), .B(n39612), .Z(n43086) );
  NOR U51910 ( .A(n43072), .B(n42370), .Z(n39603) );
  IV U51911 ( .A(n38973), .Z(n38974) );
  NOR U51912 ( .A(n38974), .B(n43065), .Z(n43055) );
  IV U51913 ( .A(n38975), .Z(n38976) );
  NOR U51914 ( .A(n38977), .B(n38976), .Z(n43061) );
  NOR U51915 ( .A(n43055), .B(n43061), .Z(n39602) );
  IV U51916 ( .A(n38978), .Z(n38979) );
  NOR U51917 ( .A(n38980), .B(n38979), .Z(n43051) );
  IV U51918 ( .A(n38981), .Z(n38983) );
  NOR U51919 ( .A(n38983), .B(n38982), .Z(n43057) );
  NOR U51920 ( .A(n43051), .B(n43057), .Z(n39601) );
  IV U51921 ( .A(n38984), .Z(n38988) );
  NOR U51922 ( .A(n38986), .B(n38985), .Z(n38987) );
  IV U51923 ( .A(n38987), .Z(n38990) );
  NOR U51924 ( .A(n38988), .B(n38990), .Z(n42385) );
  IV U51925 ( .A(n38989), .Z(n38991) );
  NOR U51926 ( .A(n38991), .B(n38990), .Z(n42382) );
  NOR U51927 ( .A(n38992), .B(n43038), .Z(n42388) );
  IV U51928 ( .A(n38993), .Z(n38998) );
  IV U51929 ( .A(n38994), .Z(n38995) );
  NOR U51930 ( .A(n38995), .B(n39003), .Z(n38996) );
  IV U51931 ( .A(n38996), .Z(n38997) );
  NOR U51932 ( .A(n38998), .B(n38997), .Z(n42390) );
  IV U51933 ( .A(n38999), .Z(n39001) );
  NOR U51934 ( .A(n39001), .B(n39000), .Z(n46231) );
  IV U51935 ( .A(n39002), .Z(n39007) );
  NOR U51936 ( .A(n39004), .B(n39003), .Z(n39005) );
  IV U51937 ( .A(n39005), .Z(n39006) );
  NOR U51938 ( .A(n39007), .B(n39006), .Z(n45551) );
  NOR U51939 ( .A(n46231), .B(n45551), .Z(n43031) );
  IV U51940 ( .A(n39008), .Z(n39009) );
  NOR U51941 ( .A(n39010), .B(n39009), .Z(n43028) );
  IV U51942 ( .A(n39011), .Z(n39013) );
  IV U51943 ( .A(n39012), .Z(n39015) );
  NOR U51944 ( .A(n39013), .B(n39015), .Z(n43021) );
  IV U51945 ( .A(n39014), .Z(n39016) );
  NOR U51946 ( .A(n39016), .B(n39015), .Z(n43024) );
  NOR U51947 ( .A(n39017), .B(n43024), .Z(n39598) );
  IV U51948 ( .A(n39018), .Z(n39019) );
  NOR U51949 ( .A(n39019), .B(n39577), .Z(n39020) );
  IV U51950 ( .A(n39020), .Z(n43005) );
  IV U51951 ( .A(n39021), .Z(n39022) );
  NOR U51952 ( .A(n39022), .B(n39571), .Z(n42997) );
  IV U51953 ( .A(n39023), .Z(n39025) );
  NOR U51954 ( .A(n39025), .B(n39024), .Z(n39541) );
  IV U51955 ( .A(n39026), .Z(n39028) );
  NOR U51956 ( .A(n39028), .B(n39027), .Z(n39538) );
  IV U51957 ( .A(n39538), .Z(n39522) );
  NOR U51958 ( .A(n39029), .B(n42441), .Z(n39521) );
  IV U51959 ( .A(n39030), .Z(n39516) );
  IV U51960 ( .A(n39031), .Z(n39032) );
  NOR U51961 ( .A(n39516), .B(n39032), .Z(n42972) );
  IV U51962 ( .A(n39033), .Z(n39035) );
  NOR U51963 ( .A(n39035), .B(n39034), .Z(n42962) );
  NOR U51964 ( .A(n42972), .B(n42962), .Z(n39513) );
  IV U51965 ( .A(n39036), .Z(n39037) );
  NOR U51966 ( .A(n39037), .B(n39507), .Z(n42958) );
  IV U51967 ( .A(n39038), .Z(n39511) );
  IV U51968 ( .A(n39039), .Z(n39040) );
  NOR U51969 ( .A(n39511), .B(n39040), .Z(n42951) );
  IV U51970 ( .A(n39041), .Z(n39042) );
  NOR U51971 ( .A(n42459), .B(n39042), .Z(n42452) );
  NOR U51972 ( .A(n42951), .B(n42452), .Z(n39505) );
  NOR U51973 ( .A(n39043), .B(n42459), .Z(n39504) );
  IV U51974 ( .A(n39044), .Z(n39045) );
  NOR U51975 ( .A(n39045), .B(n39487), .Z(n42465) );
  IV U51976 ( .A(n39046), .Z(n39047) );
  NOR U51977 ( .A(n39048), .B(n39047), .Z(n42908) );
  IV U51978 ( .A(n39467), .Z(n39049) );
  NOR U51979 ( .A(n39470), .B(n39049), .Z(n42477) );
  NOR U51980 ( .A(n42908), .B(n42477), .Z(n39050) );
  IV U51981 ( .A(n39050), .Z(n39464) );
  IV U51982 ( .A(n39051), .Z(n39052) );
  NOR U51983 ( .A(n39052), .B(n39056), .Z(n42905) );
  IV U51984 ( .A(n39053), .Z(n39054) );
  NOR U51985 ( .A(n39054), .B(n39056), .Z(n42901) );
  IV U51986 ( .A(n39055), .Z(n39057) );
  NOR U51987 ( .A(n39057), .B(n39056), .Z(n42898) );
  IV U51988 ( .A(n39058), .Z(n39060) );
  IV U51989 ( .A(n39059), .Z(n39062) );
  NOR U51990 ( .A(n39060), .B(n39062), .Z(n42482) );
  IV U51991 ( .A(n39061), .Z(n39063) );
  NOR U51992 ( .A(n39063), .B(n39062), .Z(n42479) );
  IV U51993 ( .A(n39064), .Z(n39066) );
  NOR U51994 ( .A(n39066), .B(n39065), .Z(n42491) );
  IV U51995 ( .A(n39067), .Z(n39068) );
  NOR U51996 ( .A(n39068), .B(n39070), .Z(n42486) );
  NOR U51997 ( .A(n42491), .B(n42486), .Z(n39463) );
  IV U51998 ( .A(n39069), .Z(n39071) );
  NOR U51999 ( .A(n39071), .B(n39070), .Z(n39072) );
  IV U52000 ( .A(n39072), .Z(n42485) );
  IV U52001 ( .A(n39073), .Z(n39075) );
  IV U52002 ( .A(n39074), .Z(n39078) );
  NOR U52003 ( .A(n39075), .B(n39078), .Z(n42488) );
  IV U52004 ( .A(n39076), .Z(n39077) );
  NOR U52005 ( .A(n39078), .B(n39077), .Z(n42497) );
  NOR U52006 ( .A(n39080), .B(n39079), .Z(n42494) );
  IV U52007 ( .A(n39081), .Z(n39083) );
  NOR U52008 ( .A(n39083), .B(n39082), .Z(n42503) );
  IV U52009 ( .A(n39084), .Z(n39085) );
  NOR U52010 ( .A(n39086), .B(n39085), .Z(n42500) );
  NOR U52011 ( .A(n42503), .B(n42500), .Z(n39087) );
  IV U52012 ( .A(n39087), .Z(n39461) );
  IV U52013 ( .A(n39088), .Z(n39089) );
  NOR U52014 ( .A(n39090), .B(n39089), .Z(n42890) );
  IV U52015 ( .A(n39091), .Z(n39092) );
  NOR U52016 ( .A(n39093), .B(n39092), .Z(n39094) );
  IV U52017 ( .A(n39094), .Z(n39456) );
  IV U52018 ( .A(n39095), .Z(n39097) );
  IV U52019 ( .A(n39096), .Z(n39100) );
  NOR U52020 ( .A(n39097), .B(n39100), .Z(n42882) );
  IV U52021 ( .A(n39098), .Z(n39099) );
  NOR U52022 ( .A(n39100), .B(n39099), .Z(n49185) );
  NOR U52023 ( .A(n42882), .B(n49185), .Z(n39101) );
  IV U52024 ( .A(n39101), .Z(n39448) );
  IV U52025 ( .A(n39102), .Z(n39104) );
  NOR U52026 ( .A(n39104), .B(n39103), .Z(n42517) );
  NOR U52027 ( .A(n39105), .B(n42508), .Z(n39106) );
  NOR U52028 ( .A(n42517), .B(n39106), .Z(n39447) );
  IV U52029 ( .A(n39107), .Z(n39109) );
  IV U52030 ( .A(n39108), .Z(n39111) );
  NOR U52031 ( .A(n39109), .B(n39111), .Z(n42525) );
  IV U52032 ( .A(n39110), .Z(n39112) );
  NOR U52033 ( .A(n39112), .B(n39111), .Z(n42522) );
  IV U52034 ( .A(n39113), .Z(n39116) );
  IV U52035 ( .A(n39114), .Z(n39115) );
  NOR U52036 ( .A(n39116), .B(n39115), .Z(n42529) );
  XOR U52037 ( .A(n42531), .B(n42529), .Z(n39117) );
  NOR U52038 ( .A(n42522), .B(n39117), .Z(n39439) );
  NOR U52039 ( .A(n39119), .B(n39118), .Z(n42554) );
  IV U52040 ( .A(n39120), .Z(n39432) );
  IV U52041 ( .A(n39121), .Z(n39122) );
  NOR U52042 ( .A(n39432), .B(n39122), .Z(n42551) );
  NOR U52043 ( .A(n42554), .B(n42551), .Z(n39427) );
  NOR U52044 ( .A(n39123), .B(n42559), .Z(n39426) );
  IV U52045 ( .A(n39124), .Z(n39425) );
  IV U52046 ( .A(n39125), .Z(n39126) );
  NOR U52047 ( .A(n39425), .B(n39126), .Z(n42861) );
  IV U52048 ( .A(n39127), .Z(n39128) );
  NOR U52049 ( .A(n39128), .B(n39130), .Z(n42855) );
  NOR U52050 ( .A(n42861), .B(n42855), .Z(n39421) );
  IV U52051 ( .A(n39129), .Z(n39131) );
  NOR U52052 ( .A(n39131), .B(n39130), .Z(n42852) );
  IV U52053 ( .A(n39132), .Z(n39133) );
  NOR U52054 ( .A(n39134), .B(n39133), .Z(n42569) );
  IV U52055 ( .A(n39135), .Z(n39137) );
  NOR U52056 ( .A(n39137), .B(n39136), .Z(n42567) );
  NOR U52057 ( .A(n42569), .B(n42567), .Z(n39420) );
  IV U52058 ( .A(n39138), .Z(n39139) );
  NOR U52059 ( .A(n39145), .B(n39139), .Z(n42845) );
  IV U52060 ( .A(n39140), .Z(n39141) );
  NOR U52061 ( .A(n39142), .B(n39141), .Z(n42849) );
  NOR U52062 ( .A(n42845), .B(n42849), .Z(n39419) );
  IV U52063 ( .A(n39143), .Z(n39144) );
  NOR U52064 ( .A(n39145), .B(n39144), .Z(n42843) );
  IV U52065 ( .A(n39146), .Z(n39148) );
  IV U52066 ( .A(n39147), .Z(n39150) );
  NOR U52067 ( .A(n39148), .B(n39150), .Z(n42839) );
  IV U52068 ( .A(n39149), .Z(n39151) );
  NOR U52069 ( .A(n39151), .B(n39150), .Z(n42836) );
  IV U52070 ( .A(n39152), .Z(n39154) );
  NOR U52071 ( .A(n39154), .B(n39153), .Z(n45964) );
  IV U52072 ( .A(n39155), .Z(n39156) );
  NOR U52073 ( .A(n39156), .B(n39414), .Z(n45970) );
  NOR U52074 ( .A(n45964), .B(n45970), .Z(n42578) );
  NOR U52075 ( .A(n39158), .B(n39157), .Z(n42587) );
  IV U52076 ( .A(n39159), .Z(n39394) );
  IV U52077 ( .A(n39160), .Z(n39161) );
  NOR U52078 ( .A(n39394), .B(n39161), .Z(n42585) );
  NOR U52079 ( .A(n42587), .B(n42585), .Z(n39391) );
  IV U52080 ( .A(n39162), .Z(n39163) );
  NOR U52081 ( .A(n39163), .B(n39374), .Z(n39383) );
  IV U52082 ( .A(n39164), .Z(n39169) );
  IV U52083 ( .A(n39165), .Z(n39166) );
  NOR U52084 ( .A(n39167), .B(n39166), .Z(n39168) );
  IV U52085 ( .A(n39168), .Z(n39171) );
  NOR U52086 ( .A(n39169), .B(n39171), .Z(n42826) );
  IV U52087 ( .A(n39170), .Z(n39172) );
  NOR U52088 ( .A(n39172), .B(n39171), .Z(n42823) );
  IV U52089 ( .A(n42608), .Z(n42806) );
  NOR U52090 ( .A(n42806), .B(n42607), .Z(n39346) );
  IV U52091 ( .A(n39173), .Z(n39175) );
  IV U52092 ( .A(n39174), .Z(n42799) );
  NOR U52093 ( .A(n39175), .B(n42799), .Z(n42618) );
  IV U52094 ( .A(n42800), .Z(n39176) );
  NOR U52095 ( .A(n39176), .B(n42799), .Z(n42616) );
  NOR U52096 ( .A(n42786), .B(n42616), .Z(n39177) );
  IV U52097 ( .A(n39177), .Z(n39178) );
  NOR U52098 ( .A(n42618), .B(n39178), .Z(n39345) );
  IV U52099 ( .A(n39179), .Z(n39180) );
  NOR U52100 ( .A(n39181), .B(n39180), .Z(n39337) );
  IV U52101 ( .A(n39337), .Z(n39328) );
  IV U52102 ( .A(n39182), .Z(n39185) );
  IV U52103 ( .A(n39183), .Z(n39184) );
  NOR U52104 ( .A(n39185), .B(n39184), .Z(n42628) );
  NOR U52105 ( .A(n39187), .B(n39186), .Z(n42634) );
  IV U52106 ( .A(n39188), .Z(n39189) );
  NOR U52107 ( .A(n39190), .B(n39189), .Z(n42632) );
  NOR U52108 ( .A(n42634), .B(n42632), .Z(n39326) );
  IV U52109 ( .A(n39191), .Z(n39194) );
  NOR U52110 ( .A(n39197), .B(n39192), .Z(n39193) );
  IV U52111 ( .A(n39193), .Z(n39199) );
  NOR U52112 ( .A(n39194), .B(n39199), .Z(n42774) );
  NOR U52113 ( .A(n42637), .B(n42774), .Z(n39325) );
  IV U52114 ( .A(n39195), .Z(n39196) );
  NOR U52115 ( .A(n39197), .B(n39196), .Z(n49406) );
  IV U52116 ( .A(n39198), .Z(n39200) );
  NOR U52117 ( .A(n39200), .B(n39199), .Z(n49415) );
  NOR U52118 ( .A(n49406), .B(n49415), .Z(n42765) );
  IV U52119 ( .A(n39201), .Z(n39202) );
  NOR U52120 ( .A(n39202), .B(n39323), .Z(n42640) );
  IV U52121 ( .A(n39203), .Z(n39204) );
  NOR U52122 ( .A(n39204), .B(n39206), .Z(n42757) );
  IV U52123 ( .A(n39205), .Z(n39207) );
  NOR U52124 ( .A(n39207), .B(n39206), .Z(n42753) );
  NOR U52125 ( .A(n42751), .B(n42753), .Z(n39208) );
  IV U52126 ( .A(n39208), .Z(n39312) );
  IV U52127 ( .A(n39209), .Z(n39210) );
  NOR U52128 ( .A(n39213), .B(n39210), .Z(n42746) );
  IV U52129 ( .A(n39211), .Z(n39212) );
  NOR U52130 ( .A(n39213), .B(n39212), .Z(n42656) );
  NOR U52131 ( .A(n42661), .B(n39214), .Z(n42740) );
  NOR U52132 ( .A(n42661), .B(n39215), .Z(n39311) );
  IV U52133 ( .A(n39216), .Z(n39218) );
  NOR U52134 ( .A(n39218), .B(n39217), .Z(n39222) );
  IV U52135 ( .A(n39219), .Z(n39221) );
  NOR U52136 ( .A(n39221), .B(n39220), .Z(n42667) );
  NOR U52137 ( .A(n39222), .B(n42667), .Z(n39223) );
  IV U52138 ( .A(n39223), .Z(n39310) );
  IV U52139 ( .A(n39224), .Z(n39226) );
  NOR U52140 ( .A(n39226), .B(n39225), .Z(n42681) );
  IV U52141 ( .A(n39227), .Z(n39228) );
  NOR U52142 ( .A(n39228), .B(n42669), .Z(n42677) );
  NOR U52143 ( .A(n42681), .B(n42677), .Z(n39309) );
  IV U52144 ( .A(n39229), .Z(n39231) );
  NOR U52145 ( .A(n39231), .B(n39230), .Z(n39268) );
  IV U52146 ( .A(n39232), .Z(n39234) );
  NOR U52147 ( .A(n39234), .B(n39233), .Z(n42704) );
  NOR U52148 ( .A(n39236), .B(n39235), .Z(n39237) );
  NOR U52149 ( .A(n39238), .B(n39237), .Z(n42714) );
  NOR U52150 ( .A(n39240), .B(n39239), .Z(n39245) );
  IV U52151 ( .A(n39241), .Z(n39242) );
  NOR U52152 ( .A(n39243), .B(n39242), .Z(n39244) );
  NOR U52153 ( .A(n39245), .B(n39244), .Z(n42713) );
  NOR U52154 ( .A(n39247), .B(n39246), .Z(n39257) );
  IV U52155 ( .A(n39248), .Z(n39253) );
  NOR U52156 ( .A(n39250), .B(n39249), .Z(n39251) );
  IV U52157 ( .A(n39251), .Z(n39252) );
  NOR U52158 ( .A(n39253), .B(n39252), .Z(n39255) );
  NOR U52159 ( .A(n39255), .B(n39254), .Z(n39256) );
  NOR U52160 ( .A(n39257), .B(n39256), .Z(n42712) );
  XOR U52161 ( .A(n42713), .B(n42712), .Z(n39258) );
  XOR U52162 ( .A(n42714), .B(n39258), .Z(n39259) );
  IV U52163 ( .A(n39259), .Z(n42706) );
  XOR U52164 ( .A(n42704), .B(n42706), .Z(n42708) );
  IV U52165 ( .A(n39260), .Z(n39261) );
  NOR U52166 ( .A(n39262), .B(n39261), .Z(n42707) );
  IV U52167 ( .A(n39263), .Z(n39264) );
  NOR U52168 ( .A(n39265), .B(n39264), .Z(n42702) );
  NOR U52169 ( .A(n42707), .B(n42702), .Z(n39266) );
  XOR U52170 ( .A(n42708), .B(n39266), .Z(n39267) );
  NOR U52171 ( .A(n39268), .B(n39267), .Z(n39271) );
  IV U52172 ( .A(n39268), .Z(n39270) );
  XOR U52173 ( .A(n42707), .B(n42708), .Z(n39269) );
  NOR U52174 ( .A(n39270), .B(n39269), .Z(n42718) );
  NOR U52175 ( .A(n39271), .B(n42718), .Z(n39272) );
  IV U52176 ( .A(n39272), .Z(n42721) );
  IV U52177 ( .A(n39273), .Z(n39274) );
  NOR U52178 ( .A(n39275), .B(n39274), .Z(n42715) );
  IV U52179 ( .A(n39276), .Z(n39278) );
  NOR U52180 ( .A(n39278), .B(n39277), .Z(n42720) );
  NOR U52181 ( .A(n42715), .B(n42720), .Z(n39279) );
  XOR U52182 ( .A(n42721), .B(n39279), .Z(n42692) );
  IV U52183 ( .A(n39280), .Z(n39282) );
  NOR U52184 ( .A(n39282), .B(n39281), .Z(n42699) );
  IV U52185 ( .A(n39283), .Z(n39284) );
  NOR U52186 ( .A(n39284), .B(n39287), .Z(n42693) );
  NOR U52187 ( .A(n42699), .B(n42693), .Z(n39285) );
  XOR U52188 ( .A(n42692), .B(n39285), .Z(n42697) );
  IV U52189 ( .A(n39286), .Z(n39288) );
  NOR U52190 ( .A(n39288), .B(n39287), .Z(n42695) );
  XOR U52191 ( .A(n42697), .B(n42695), .Z(n42732) );
  IV U52192 ( .A(n39289), .Z(n42689) );
  NOR U52193 ( .A(n42689), .B(n39290), .Z(n39293) );
  IV U52194 ( .A(n39291), .Z(n39292) );
  NOR U52195 ( .A(n39292), .B(n39297), .Z(n42730) );
  NOR U52196 ( .A(n39293), .B(n42730), .Z(n39294) );
  XOR U52197 ( .A(n42732), .B(n39294), .Z(n42685) );
  IV U52198 ( .A(n39295), .Z(n39296) );
  NOR U52199 ( .A(n39297), .B(n39296), .Z(n42728) );
  IV U52200 ( .A(n39298), .Z(n39299) );
  NOR U52201 ( .A(n39302), .B(n39299), .Z(n42734) );
  IV U52202 ( .A(n39300), .Z(n39301) );
  NOR U52203 ( .A(n39302), .B(n39301), .Z(n42686) );
  NOR U52204 ( .A(n42734), .B(n42686), .Z(n39303) );
  IV U52205 ( .A(n39303), .Z(n39304) );
  NOR U52206 ( .A(n42728), .B(n39304), .Z(n39305) );
  XOR U52207 ( .A(n42685), .B(n39305), .Z(n45788) );
  IV U52208 ( .A(n39306), .Z(n39307) );
  NOR U52209 ( .A(n39308), .B(n39307), .Z(n45836) );
  NOR U52210 ( .A(n45787), .B(n45836), .Z(n42680) );
  XOR U52211 ( .A(n45788), .B(n42680), .Z(n42678) );
  XOR U52212 ( .A(n39309), .B(n42678), .Z(n42670) );
  XOR U52213 ( .A(n39310), .B(n42670), .Z(n42660) );
  XOR U52214 ( .A(n39311), .B(n42660), .Z(n42741) );
  XOR U52215 ( .A(n42740), .B(n42741), .Z(n42657) );
  XOR U52216 ( .A(n42656), .B(n42657), .Z(n42747) );
  XOR U52217 ( .A(n42746), .B(n42747), .Z(n42754) );
  XOR U52218 ( .A(n39312), .B(n42754), .Z(n42761) );
  XOR U52219 ( .A(n42757), .B(n42761), .Z(n42654) );
  IV U52220 ( .A(n39313), .Z(n39315) );
  NOR U52221 ( .A(n39315), .B(n39314), .Z(n42653) );
  NOR U52222 ( .A(n42759), .B(n42653), .Z(n39316) );
  XOR U52223 ( .A(n42654), .B(n39316), .Z(n42645) );
  IV U52224 ( .A(n39317), .Z(n42646) );
  NOR U52225 ( .A(n39318), .B(n42646), .Z(n39320) );
  NOR U52226 ( .A(n39320), .B(n39319), .Z(n39321) );
  XOR U52227 ( .A(n42645), .B(n39321), .Z(n42768) );
  IV U52228 ( .A(n39322), .Z(n39324) );
  NOR U52229 ( .A(n39324), .B(n39323), .Z(n42766) );
  XOR U52230 ( .A(n42768), .B(n42766), .Z(n42641) );
  XOR U52231 ( .A(n42640), .B(n42641), .Z(n49411) );
  XOR U52232 ( .A(n42765), .B(n49411), .Z(n42638) );
  XOR U52233 ( .A(n39325), .B(n42638), .Z(n42636) );
  XOR U52234 ( .A(n39326), .B(n42636), .Z(n39327) );
  IV U52235 ( .A(n39327), .Z(n42626) );
  XOR U52236 ( .A(n42625), .B(n42626), .Z(n42629) );
  XOR U52237 ( .A(n42628), .B(n42629), .Z(n39332) );
  NOR U52238 ( .A(n39328), .B(n39332), .Z(n45906) );
  IV U52239 ( .A(n39329), .Z(n39330) );
  NOR U52240 ( .A(n39331), .B(n39330), .Z(n39334) );
  IV U52241 ( .A(n39332), .Z(n39333) );
  NOR U52242 ( .A(n39334), .B(n39333), .Z(n39336) );
  IV U52243 ( .A(n39334), .Z(n39335) );
  NOR U52244 ( .A(n39335), .B(n42626), .Z(n45903) );
  NOR U52245 ( .A(n39336), .B(n45903), .Z(n42622) );
  NOR U52246 ( .A(n39337), .B(n42622), .Z(n39338) );
  NOR U52247 ( .A(n45906), .B(n39338), .Z(n42780) );
  IV U52248 ( .A(n39339), .Z(n39340) );
  NOR U52249 ( .A(n39340), .B(n39342), .Z(n42779) );
  IV U52250 ( .A(n39341), .Z(n39343) );
  NOR U52251 ( .A(n39343), .B(n39342), .Z(n42621) );
  NOR U52252 ( .A(n42779), .B(n42621), .Z(n39344) );
  XOR U52253 ( .A(n42780), .B(n39344), .Z(n42785) );
  XOR U52254 ( .A(n42783), .B(n42785), .Z(n42787) );
  XOR U52255 ( .A(n39345), .B(n42787), .Z(n42801) );
  NOR U52256 ( .A(n39346), .B(n42801), .Z(n39350) );
  XOR U52257 ( .A(n42786), .B(n42787), .Z(n39348) );
  IV U52258 ( .A(n39346), .Z(n39347) );
  NOR U52259 ( .A(n39348), .B(n39347), .Z(n39349) );
  NOR U52260 ( .A(n39350), .B(n39349), .Z(n42600) );
  IV U52261 ( .A(n39351), .Z(n39352) );
  NOR U52262 ( .A(n39352), .B(n42607), .Z(n42610) );
  IV U52263 ( .A(n39353), .Z(n39355) );
  IV U52264 ( .A(n39354), .Z(n39359) );
  NOR U52265 ( .A(n39355), .B(n39359), .Z(n39356) );
  NOR U52266 ( .A(n42610), .B(n39356), .Z(n39357) );
  XOR U52267 ( .A(n42600), .B(n39357), .Z(n42597) );
  IV U52268 ( .A(n39358), .Z(n39360) );
  NOR U52269 ( .A(n39360), .B(n39359), .Z(n42593) );
  NOR U52270 ( .A(n39361), .B(n42596), .Z(n39362) );
  NOR U52271 ( .A(n42593), .B(n39362), .Z(n39363) );
  XOR U52272 ( .A(n42597), .B(n39363), .Z(n42591) );
  IV U52273 ( .A(n39364), .Z(n39365) );
  NOR U52274 ( .A(n39365), .B(n39367), .Z(n42590) );
  IV U52275 ( .A(n39366), .Z(n39368) );
  NOR U52276 ( .A(n39368), .B(n39367), .Z(n42816) );
  NOR U52277 ( .A(n42590), .B(n42816), .Z(n39369) );
  XOR U52278 ( .A(n42591), .B(n39369), .Z(n42820) );
  XOR U52279 ( .A(n42819), .B(n42820), .Z(n42825) );
  XOR U52280 ( .A(n42823), .B(n42825), .Z(n42827) );
  XOR U52281 ( .A(n42826), .B(n42827), .Z(n42833) );
  IV U52282 ( .A(n39370), .Z(n39372) );
  NOR U52283 ( .A(n39372), .B(n39371), .Z(n42830) );
  IV U52284 ( .A(n39373), .Z(n39375) );
  NOR U52285 ( .A(n39375), .B(n39374), .Z(n42832) );
  NOR U52286 ( .A(n42830), .B(n42832), .Z(n39376) );
  XOR U52287 ( .A(n42833), .B(n39376), .Z(n39377) );
  NOR U52288 ( .A(n39383), .B(n39377), .Z(n39378) );
  IV U52289 ( .A(n39378), .Z(n39382) );
  IV U52290 ( .A(n39379), .Z(n39380) );
  NOR U52291 ( .A(n39381), .B(n39380), .Z(n39385) );
  NOR U52292 ( .A(n39382), .B(n39385), .Z(n39390) );
  IV U52293 ( .A(n39383), .Z(n39384) );
  NOR U52294 ( .A(n39384), .B(n42833), .Z(n45736) );
  IV U52295 ( .A(n39385), .Z(n39387) );
  XOR U52296 ( .A(n42830), .B(n42833), .Z(n39386) );
  NOR U52297 ( .A(n39387), .B(n39386), .Z(n45956) );
  NOR U52298 ( .A(n45736), .B(n45956), .Z(n39388) );
  IV U52299 ( .A(n39388), .Z(n39389) );
  NOR U52300 ( .A(n39390), .B(n39389), .Z(n42584) );
  XOR U52301 ( .A(n39391), .B(n42584), .Z(n42583) );
  IV U52302 ( .A(n39392), .Z(n39393) );
  NOR U52303 ( .A(n39394), .B(n39393), .Z(n39395) );
  IV U52304 ( .A(n39395), .Z(n42582) );
  XOR U52305 ( .A(n42583), .B(n42582), .Z(n39405) );
  IV U52306 ( .A(n39396), .Z(n39397) );
  NOR U52307 ( .A(n39398), .B(n39397), .Z(n39408) );
  IV U52308 ( .A(n39399), .Z(n39400) );
  NOR U52309 ( .A(n39401), .B(n39400), .Z(n39404) );
  NOR U52310 ( .A(n39408), .B(n39404), .Z(n39402) );
  IV U52311 ( .A(n39402), .Z(n39403) );
  NOR U52312 ( .A(n39405), .B(n39403), .Z(n39411) );
  IV U52313 ( .A(n39404), .Z(n39407) );
  IV U52314 ( .A(n39405), .Z(n39406) );
  NOR U52315 ( .A(n39407), .B(n39406), .Z(n45724) );
  IV U52316 ( .A(n39408), .Z(n39409) );
  NOR U52317 ( .A(n39409), .B(n42583), .Z(n45729) );
  NOR U52318 ( .A(n45724), .B(n45729), .Z(n39410) );
  IV U52319 ( .A(n39410), .Z(n42580) );
  NOR U52320 ( .A(n39411), .B(n42580), .Z(n39412) );
  IV U52321 ( .A(n39412), .Z(n45966) );
  XOR U52322 ( .A(n42578), .B(n45966), .Z(n42573) );
  IV U52323 ( .A(n39413), .Z(n39415) );
  NOR U52324 ( .A(n39415), .B(n39414), .Z(n42575) );
  NOR U52325 ( .A(n39417), .B(n39416), .Z(n42572) );
  NOR U52326 ( .A(n42575), .B(n42572), .Z(n39418) );
  XOR U52327 ( .A(n42573), .B(n39418), .Z(n42837) );
  XOR U52328 ( .A(n42836), .B(n42837), .Z(n42840) );
  XOR U52329 ( .A(n42839), .B(n42840), .Z(n42846) );
  XOR U52330 ( .A(n42843), .B(n42846), .Z(n42851) );
  XOR U52331 ( .A(n39419), .B(n42851), .Z(n42566) );
  XOR U52332 ( .A(n39420), .B(n42566), .Z(n42853) );
  XOR U52333 ( .A(n42852), .B(n42853), .Z(n42863) );
  XOR U52334 ( .A(n39421), .B(n42863), .Z(n39422) );
  IV U52335 ( .A(n39422), .Z(n42564) );
  IV U52336 ( .A(n39423), .Z(n39424) );
  NOR U52337 ( .A(n39425), .B(n39424), .Z(n42562) );
  XOR U52338 ( .A(n42564), .B(n42562), .Z(n42555) );
  XOR U52339 ( .A(n39426), .B(n42555), .Z(n42552) );
  XOR U52340 ( .A(n39427), .B(n42552), .Z(n42542) );
  IV U52341 ( .A(n39428), .Z(n39429) );
  NOR U52342 ( .A(n39430), .B(n39429), .Z(n42543) );
  IV U52343 ( .A(n39431), .Z(n39433) );
  NOR U52344 ( .A(n39433), .B(n39432), .Z(n42548) );
  NOR U52345 ( .A(n42543), .B(n42548), .Z(n39434) );
  XOR U52346 ( .A(n42542), .B(n39434), .Z(n42546) );
  XOR U52347 ( .A(n42545), .B(n42546), .Z(n42537) );
  XOR U52348 ( .A(n42536), .B(n42537), .Z(n42540) );
  IV U52349 ( .A(n39435), .Z(n39437) );
  NOR U52350 ( .A(n39437), .B(n39436), .Z(n42534) );
  NOR U52351 ( .A(n42539), .B(n42534), .Z(n39438) );
  XOR U52352 ( .A(n42540), .B(n39438), .Z(n42523) );
  XOR U52353 ( .A(n39439), .B(n42523), .Z(n42526) );
  XOR U52354 ( .A(n42525), .B(n42526), .Z(n42514) );
  IV U52355 ( .A(n39440), .Z(n39441) );
  NOR U52356 ( .A(n39442), .B(n39441), .Z(n42513) );
  IV U52357 ( .A(n39443), .Z(n39445) );
  NOR U52358 ( .A(n39445), .B(n39444), .Z(n42511) );
  NOR U52359 ( .A(n42513), .B(n42511), .Z(n39446) );
  XOR U52360 ( .A(n42514), .B(n39446), .Z(n42507) );
  XOR U52361 ( .A(n39447), .B(n42507), .Z(n49184) );
  XOR U52362 ( .A(n39448), .B(n49184), .Z(n42883) );
  NOR U52363 ( .A(n39456), .B(n42883), .Z(n42505) );
  IV U52364 ( .A(n39449), .Z(n39450) );
  NOR U52365 ( .A(n39451), .B(n39450), .Z(n42886) );
  IV U52366 ( .A(n39452), .Z(n39453) );
  NOR U52367 ( .A(n39454), .B(n39453), .Z(n39455) );
  IV U52368 ( .A(n39455), .Z(n42884) );
  XOR U52369 ( .A(n42884), .B(n42883), .Z(n42887) );
  XOR U52370 ( .A(n42886), .B(n42887), .Z(n39458) );
  NOR U52371 ( .A(n42887), .B(n39456), .Z(n39457) );
  NOR U52372 ( .A(n39458), .B(n39457), .Z(n39459) );
  NOR U52373 ( .A(n42505), .B(n39459), .Z(n39460) );
  IV U52374 ( .A(n39460), .Z(n42891) );
  XOR U52375 ( .A(n42890), .B(n42891), .Z(n42501) );
  XOR U52376 ( .A(n39461), .B(n42501), .Z(n42496) );
  XOR U52377 ( .A(n42494), .B(n42496), .Z(n42498) );
  XOR U52378 ( .A(n42497), .B(n42498), .Z(n42489) );
  XOR U52379 ( .A(n42488), .B(n42489), .Z(n42492) );
  XOR U52380 ( .A(n42485), .B(n42492), .Z(n39462) );
  XOR U52381 ( .A(n39463), .B(n39462), .Z(n42481) );
  XOR U52382 ( .A(n42479), .B(n42481), .Z(n42483) );
  XOR U52383 ( .A(n42482), .B(n42483), .Z(n42900) );
  XOR U52384 ( .A(n42898), .B(n42900), .Z(n42903) );
  XOR U52385 ( .A(n42901), .B(n42903), .Z(n42907) );
  XOR U52386 ( .A(n42905), .B(n42907), .Z(n42909) );
  XOR U52387 ( .A(n39464), .B(n42909), .Z(n42913) );
  IV U52388 ( .A(n39465), .Z(n39466) );
  NOR U52389 ( .A(n39467), .B(n39466), .Z(n39468) );
  IV U52390 ( .A(n39468), .Z(n39469) );
  NOR U52391 ( .A(n39470), .B(n39469), .Z(n39471) );
  IV U52392 ( .A(n39471), .Z(n42911) );
  XOR U52393 ( .A(n42913), .B(n42911), .Z(n42919) );
  IV U52394 ( .A(n39472), .Z(n42914) );
  NOR U52395 ( .A(n42914), .B(n39473), .Z(n39476) );
  NOR U52396 ( .A(n39475), .B(n39474), .Z(n42918) );
  NOR U52397 ( .A(n39476), .B(n42918), .Z(n39477) );
  XOR U52398 ( .A(n42919), .B(n39477), .Z(n49138) );
  XOR U52399 ( .A(n49139), .B(n49138), .Z(n42476) );
  IV U52400 ( .A(n39478), .Z(n42472) );
  NOR U52401 ( .A(n39479), .B(n42472), .Z(n39480) );
  NOR U52402 ( .A(n42475), .B(n39480), .Z(n39481) );
  XOR U52403 ( .A(n42476), .B(n39481), .Z(n42466) );
  IV U52404 ( .A(n39482), .Z(n39483) );
  NOR U52405 ( .A(n39484), .B(n39483), .Z(n42469) );
  IV U52406 ( .A(n39485), .Z(n39486) );
  NOR U52407 ( .A(n39487), .B(n39486), .Z(n42930) );
  NOR U52408 ( .A(n42469), .B(n42930), .Z(n39488) );
  XOR U52409 ( .A(n42466), .B(n39488), .Z(n45631) );
  XOR U52410 ( .A(n42465), .B(n45631), .Z(n46121) );
  IV U52411 ( .A(n39489), .Z(n39490) );
  NOR U52412 ( .A(n39491), .B(n39490), .Z(n45629) );
  IV U52413 ( .A(n39492), .Z(n39493) );
  NOR U52414 ( .A(n39494), .B(n39493), .Z(n46120) );
  NOR U52415 ( .A(n45629), .B(n46120), .Z(n42933) );
  XOR U52416 ( .A(n46121), .B(n42933), .Z(n42462) );
  NOR U52417 ( .A(n39495), .B(n42936), .Z(n39499) );
  IV U52418 ( .A(n39496), .Z(n39498) );
  IV U52419 ( .A(n39497), .Z(n39502) );
  NOR U52420 ( .A(n39498), .B(n39502), .Z(n42463) );
  NOR U52421 ( .A(n39499), .B(n42463), .Z(n39500) );
  XOR U52422 ( .A(n42462), .B(n39500), .Z(n42456) );
  IV U52423 ( .A(n39501), .Z(n39503) );
  NOR U52424 ( .A(n39503), .B(n39502), .Z(n42454) );
  XOR U52425 ( .A(n42456), .B(n42454), .Z(n42946) );
  XOR U52426 ( .A(n39504), .B(n42946), .Z(n42953) );
  XOR U52427 ( .A(n39505), .B(n42953), .Z(n42954) );
  IV U52428 ( .A(n39506), .Z(n39508) );
  NOR U52429 ( .A(n39508), .B(n39507), .Z(n42964) );
  IV U52430 ( .A(n39509), .Z(n39510) );
  NOR U52431 ( .A(n39511), .B(n39510), .Z(n42955) );
  NOR U52432 ( .A(n42964), .B(n42955), .Z(n39512) );
  XOR U52433 ( .A(n42954), .B(n39512), .Z(n42959) );
  XOR U52434 ( .A(n42958), .B(n42959), .Z(n42973) );
  XOR U52435 ( .A(n39513), .B(n42973), .Z(n42450) );
  IV U52436 ( .A(n39514), .Z(n39515) );
  NOR U52437 ( .A(n39516), .B(n39515), .Z(n42975) );
  IV U52438 ( .A(n39517), .Z(n39519) );
  NOR U52439 ( .A(n39519), .B(n39518), .Z(n42449) );
  NOR U52440 ( .A(n42975), .B(n42449), .Z(n39520) );
  XOR U52441 ( .A(n42450), .B(n39520), .Z(n42440) );
  XOR U52442 ( .A(n39521), .B(n42440), .Z(n39525) );
  NOR U52443 ( .A(n39522), .B(n39525), .Z(n42438) );
  IV U52444 ( .A(n39523), .Z(n39529) );
  NOR U52445 ( .A(n39524), .B(n39529), .Z(n39527) );
  IV U52446 ( .A(n39525), .Z(n39526) );
  NOR U52447 ( .A(n39527), .B(n39526), .Z(n39537) );
  IV U52448 ( .A(n39528), .Z(n39531) );
  NOR U52449 ( .A(n39529), .B(n42440), .Z(n39530) );
  IV U52450 ( .A(n39530), .Z(n39533) );
  NOR U52451 ( .A(n39531), .B(n39533), .Z(n46168) );
  IV U52452 ( .A(n39532), .Z(n39534) );
  NOR U52453 ( .A(n39534), .B(n39533), .Z(n46154) );
  NOR U52454 ( .A(n46168), .B(n46154), .Z(n39535) );
  IV U52455 ( .A(n39535), .Z(n39536) );
  NOR U52456 ( .A(n39537), .B(n39536), .Z(n39542) );
  NOR U52457 ( .A(n39538), .B(n39542), .Z(n39539) );
  NOR U52458 ( .A(n42438), .B(n39539), .Z(n39540) );
  NOR U52459 ( .A(n39541), .B(n39540), .Z(n39545) );
  IV U52460 ( .A(n39541), .Z(n39544) );
  IV U52461 ( .A(n39542), .Z(n39543) );
  NOR U52462 ( .A(n39544), .B(n39543), .Z(n46174) );
  NOR U52463 ( .A(n39545), .B(n46174), .Z(n39546) );
  IV U52464 ( .A(n39546), .Z(n42985) );
  IV U52465 ( .A(n39547), .Z(n39548) );
  NOR U52466 ( .A(n39548), .B(n39555), .Z(n42980) );
  XOR U52467 ( .A(n42985), .B(n42980), .Z(n42437) );
  IV U52468 ( .A(n39549), .Z(n39553) );
  NOR U52469 ( .A(n39551), .B(n39550), .Z(n39552) );
  IV U52470 ( .A(n39552), .Z(n39563) );
  NOR U52471 ( .A(n39553), .B(n39563), .Z(n42435) );
  IV U52472 ( .A(n39554), .Z(n39556) );
  NOR U52473 ( .A(n39556), .B(n39555), .Z(n42983) );
  NOR U52474 ( .A(n42435), .B(n42983), .Z(n39557) );
  XOR U52475 ( .A(n42437), .B(n39557), .Z(n39565) );
  IV U52476 ( .A(n39565), .Z(n42433) );
  IV U52477 ( .A(n39558), .Z(n39559) );
  NOR U52478 ( .A(n39560), .B(n39559), .Z(n39566) );
  IV U52479 ( .A(n39566), .Z(n39561) );
  NOR U52480 ( .A(n42433), .B(n39561), .Z(n45590) );
  IV U52481 ( .A(n39562), .Z(n39564) );
  NOR U52482 ( .A(n39564), .B(n39563), .Z(n42431) );
  XOR U52483 ( .A(n42431), .B(n39565), .Z(n42425) );
  NOR U52484 ( .A(n39566), .B(n42425), .Z(n39567) );
  NOR U52485 ( .A(n45590), .B(n39567), .Z(n42419) );
  IV U52486 ( .A(n39568), .Z(n39569) );
  NOR U52487 ( .A(n39569), .B(n42427), .Z(n42988) );
  IV U52488 ( .A(n39570), .Z(n39572) );
  NOR U52489 ( .A(n39572), .B(n39571), .Z(n42994) );
  NOR U52490 ( .A(n42988), .B(n42994), .Z(n39573) );
  XOR U52491 ( .A(n42419), .B(n39573), .Z(n42998) );
  XOR U52492 ( .A(n42997), .B(n42998), .Z(n43008) );
  IV U52493 ( .A(n39574), .Z(n42421) );
  NOR U52494 ( .A(n39575), .B(n42421), .Z(n39579) );
  IV U52495 ( .A(n39576), .Z(n39578) );
  NOR U52496 ( .A(n39578), .B(n39577), .Z(n43007) );
  NOR U52497 ( .A(n39579), .B(n43007), .Z(n39580) );
  XOR U52498 ( .A(n43008), .B(n39580), .Z(n43004) );
  XOR U52499 ( .A(n43005), .B(n43004), .Z(n42416) );
  IV U52500 ( .A(n39581), .Z(n39583) );
  NOR U52501 ( .A(n39583), .B(n39582), .Z(n42415) );
  NOR U52502 ( .A(n39584), .B(n42409), .Z(n39585) );
  NOR U52503 ( .A(n42415), .B(n39585), .Z(n39586) );
  XOR U52504 ( .A(n42416), .B(n39586), .Z(n42402) );
  IV U52505 ( .A(n39587), .Z(n39588) );
  NOR U52506 ( .A(n39589), .B(n39588), .Z(n45561) );
  IV U52507 ( .A(n39590), .Z(n39591) );
  NOR U52508 ( .A(n39595), .B(n39591), .Z(n46194) );
  NOR U52509 ( .A(n45561), .B(n46194), .Z(n42403) );
  XOR U52510 ( .A(n42402), .B(n42403), .Z(n42400) );
  NOR U52511 ( .A(n39593), .B(n39592), .Z(n42399) );
  IV U52512 ( .A(n39594), .Z(n39596) );
  NOR U52513 ( .A(n39596), .B(n39595), .Z(n42397) );
  NOR U52514 ( .A(n42399), .B(n42397), .Z(n39597) );
  XOR U52515 ( .A(n42400), .B(n39597), .Z(n43019) );
  XOR U52516 ( .A(n39598), .B(n43019), .Z(n43023) );
  XOR U52517 ( .A(n43021), .B(n43023), .Z(n46235) );
  XOR U52518 ( .A(n43028), .B(n46235), .Z(n43030) );
  XOR U52519 ( .A(n43031), .B(n43030), .Z(n39599) );
  IV U52520 ( .A(n39599), .Z(n42391) );
  XOR U52521 ( .A(n42390), .B(n42391), .Z(n43035) );
  XOR U52522 ( .A(n42388), .B(n43035), .Z(n42383) );
  XOR U52523 ( .A(n42382), .B(n42383), .Z(n42386) );
  XOR U52524 ( .A(n42385), .B(n42386), .Z(n43052) );
  XOR U52525 ( .A(n39600), .B(n43052), .Z(n43058) );
  XOR U52526 ( .A(n39601), .B(n43058), .Z(n43054) );
  XOR U52527 ( .A(n39602), .B(n43054), .Z(n43073) );
  XOR U52528 ( .A(n39603), .B(n43073), .Z(n42366) );
  IV U52529 ( .A(n39604), .Z(n42372) );
  NOR U52530 ( .A(n39605), .B(n42372), .Z(n39609) );
  IV U52531 ( .A(n39606), .Z(n39608) );
  NOR U52532 ( .A(n39608), .B(n39607), .Z(n42365) );
  NOR U52533 ( .A(n39609), .B(n42365), .Z(n39610) );
  XOR U52534 ( .A(n42366), .B(n39610), .Z(n43085) );
  IV U52535 ( .A(n39611), .Z(n39613) );
  NOR U52536 ( .A(n39613), .B(n39612), .Z(n43083) );
  XOR U52537 ( .A(n43085), .B(n43083), .Z(n43088) );
  XOR U52538 ( .A(n43086), .B(n43088), .Z(n42363) );
  XOR U52539 ( .A(n42362), .B(n42363), .Z(n39618) );
  IV U52540 ( .A(n39614), .Z(n39616) );
  NOR U52541 ( .A(n39616), .B(n39615), .Z(n39623) );
  IV U52542 ( .A(n39623), .Z(n39617) );
  NOR U52543 ( .A(n39618), .B(n39617), .Z(n49023) );
  NOR U52544 ( .A(n39620), .B(n39619), .Z(n42359) );
  NOR U52545 ( .A(n42359), .B(n42362), .Z(n39621) );
  XOR U52546 ( .A(n42363), .B(n39621), .Z(n39622) );
  NOR U52547 ( .A(n39623), .B(n39622), .Z(n39624) );
  NOR U52548 ( .A(n49023), .B(n39624), .Z(n39625) );
  IV U52549 ( .A(n39625), .Z(n42357) );
  XOR U52550 ( .A(n42356), .B(n42357), .Z(n42352) );
  XOR U52551 ( .A(n42351), .B(n42352), .Z(n43097) );
  IV U52552 ( .A(n39626), .Z(n39627) );
  NOR U52553 ( .A(n39628), .B(n39627), .Z(n42354) );
  IV U52554 ( .A(n39629), .Z(n39630) );
  NOR U52555 ( .A(n39631), .B(n39630), .Z(n43096) );
  NOR U52556 ( .A(n42354), .B(n43096), .Z(n39632) );
  XOR U52557 ( .A(n43097), .B(n39632), .Z(n42348) );
  XOR U52558 ( .A(n39633), .B(n42348), .Z(n43113) );
  XOR U52559 ( .A(n39634), .B(n43113), .Z(n45483) );
  XOR U52560 ( .A(n39635), .B(n45483), .Z(n43119) );
  XOR U52561 ( .A(n43118), .B(n43119), .Z(n43123) );
  IV U52562 ( .A(n39636), .Z(n39638) );
  NOR U52563 ( .A(n39638), .B(n39637), .Z(n39639) );
  IV U52564 ( .A(n39639), .Z(n39640) );
  NOR U52565 ( .A(n39641), .B(n39640), .Z(n43121) );
  XOR U52566 ( .A(n43123), .B(n43121), .Z(n42343) );
  XOR U52567 ( .A(n42342), .B(n42343), .Z(n42345) );
  XOR U52568 ( .A(n42346), .B(n42345), .Z(n42340) );
  IV U52569 ( .A(n39642), .Z(n39643) );
  NOR U52570 ( .A(n39644), .B(n39643), .Z(n45464) );
  IV U52571 ( .A(n39645), .Z(n39647) );
  NOR U52572 ( .A(n39647), .B(n39646), .Z(n45470) );
  NOR U52573 ( .A(n45464), .B(n45470), .Z(n42341) );
  XOR U52574 ( .A(n42340), .B(n42341), .Z(n45455) );
  NOR U52575 ( .A(n39648), .B(n45455), .Z(n45451) );
  NOR U52576 ( .A(n39649), .B(n45458), .Z(n42339) );
  NOR U52577 ( .A(n39651), .B(n39650), .Z(n42337) );
  NOR U52578 ( .A(n42339), .B(n42337), .Z(n39652) );
  XOR U52579 ( .A(n39652), .B(n45455), .Z(n42336) );
  NOR U52580 ( .A(n39653), .B(n42336), .Z(n39654) );
  NOR U52581 ( .A(n45451), .B(n39654), .Z(n43129) );
  XOR U52582 ( .A(n39655), .B(n43129), .Z(n42325) );
  XOR U52583 ( .A(n39656), .B(n42325), .Z(n42310) );
  XOR U52584 ( .A(n42311), .B(n42310), .Z(n42309) );
  IV U52585 ( .A(n39657), .Z(n39659) );
  NOR U52586 ( .A(n39659), .B(n39658), .Z(n42307) );
  XOR U52587 ( .A(n42309), .B(n42307), .Z(n42300) );
  IV U52588 ( .A(n39660), .Z(n39665) );
  IV U52589 ( .A(n39661), .Z(n39662) );
  NOR U52590 ( .A(n39663), .B(n39662), .Z(n39664) );
  IV U52591 ( .A(n39664), .Z(n39676) );
  NOR U52592 ( .A(n39665), .B(n39676), .Z(n42299) );
  XOR U52593 ( .A(n39667), .B(n39666), .Z(n39670) );
  IV U52594 ( .A(n39668), .Z(n39669) );
  NOR U52595 ( .A(n39670), .B(n39669), .Z(n42297) );
  NOR U52596 ( .A(n42299), .B(n42297), .Z(n39671) );
  XOR U52597 ( .A(n42300), .B(n39671), .Z(n42294) );
  IV U52598 ( .A(n39672), .Z(n39673) );
  NOR U52599 ( .A(n39674), .B(n39673), .Z(n42295) );
  IV U52600 ( .A(n39675), .Z(n39677) );
  NOR U52601 ( .A(n39677), .B(n39676), .Z(n42303) );
  NOR U52602 ( .A(n42295), .B(n42303), .Z(n39678) );
  XOR U52603 ( .A(n42294), .B(n39678), .Z(n42292) );
  XOR U52604 ( .A(n42290), .B(n42292), .Z(n43143) );
  XOR U52605 ( .A(n43141), .B(n43143), .Z(n42287) );
  NOR U52606 ( .A(n39679), .B(n43144), .Z(n39683) );
  IV U52607 ( .A(n39680), .Z(n39681) );
  NOR U52608 ( .A(n39682), .B(n39681), .Z(n42286) );
  NOR U52609 ( .A(n39683), .B(n42286), .Z(n39684) );
  XOR U52610 ( .A(n42287), .B(n39684), .Z(n43155) );
  XOR U52611 ( .A(n43153), .B(n43155), .Z(n42284) );
  XOR U52612 ( .A(n42283), .B(n42284), .Z(n43167) );
  XOR U52613 ( .A(n39685), .B(n43167), .Z(n42280) );
  XOR U52614 ( .A(n39686), .B(n42280), .Z(n42278) );
  XOR U52615 ( .A(n39687), .B(n42278), .Z(n42270) );
  IV U52616 ( .A(n39688), .Z(n45428) );
  NOR U52617 ( .A(n39689), .B(n45428), .Z(n42273) );
  IV U52618 ( .A(n39690), .Z(n39691) );
  NOR U52619 ( .A(n39692), .B(n39691), .Z(n42269) );
  NOR U52620 ( .A(n42273), .B(n42269), .Z(n39693) );
  XOR U52621 ( .A(n42270), .B(n39693), .Z(n42268) );
  IV U52622 ( .A(n39694), .Z(n39696) );
  NOR U52623 ( .A(n39696), .B(n39695), .Z(n39697) );
  IV U52624 ( .A(n39697), .Z(n39704) );
  NOR U52625 ( .A(n42268), .B(n39704), .Z(n46354) );
  IV U52626 ( .A(n39698), .Z(n39699) );
  NOR U52627 ( .A(n39699), .B(n39709), .Z(n42263) );
  IV U52628 ( .A(n39700), .Z(n39702) );
  NOR U52629 ( .A(n39702), .B(n39701), .Z(n39703) );
  IV U52630 ( .A(n39703), .Z(n42267) );
  XOR U52631 ( .A(n42267), .B(n42268), .Z(n42264) );
  XOR U52632 ( .A(n42263), .B(n42264), .Z(n39706) );
  NOR U52633 ( .A(n42264), .B(n39704), .Z(n39705) );
  NOR U52634 ( .A(n39706), .B(n39705), .Z(n39707) );
  NOR U52635 ( .A(n46354), .B(n39707), .Z(n42257) );
  IV U52636 ( .A(n39708), .Z(n39710) );
  NOR U52637 ( .A(n39710), .B(n39709), .Z(n42256) );
  IV U52638 ( .A(n42256), .Z(n42259) );
  XOR U52639 ( .A(n42257), .B(n42259), .Z(n45413) );
  XOR U52640 ( .A(n39711), .B(n45413), .Z(n43177) );
  XOR U52641 ( .A(n43175), .B(n43177), .Z(n43173) );
  XOR U52642 ( .A(n43174), .B(n43173), .Z(n42249) );
  IV U52643 ( .A(n39712), .Z(n39713) );
  NOR U52644 ( .A(n39714), .B(n39713), .Z(n43170) );
  IV U52645 ( .A(n39715), .Z(n39716) );
  NOR U52646 ( .A(n39719), .B(n39716), .Z(n42250) );
  NOR U52647 ( .A(n43170), .B(n42250), .Z(n39717) );
  XOR U52648 ( .A(n42249), .B(n39717), .Z(n43185) );
  IV U52649 ( .A(n39718), .Z(n39720) );
  NOR U52650 ( .A(n39720), .B(n39719), .Z(n43183) );
  XOR U52651 ( .A(n43185), .B(n43183), .Z(n43190) );
  XOR U52652 ( .A(n39721), .B(n43190), .Z(n42245) );
  XOR U52653 ( .A(n42243), .B(n42245), .Z(n42248) );
  XOR U52654 ( .A(n42246), .B(n42248), .Z(n42239) );
  XOR U52655 ( .A(n42237), .B(n42239), .Z(n42241) );
  XOR U52656 ( .A(n39722), .B(n42241), .Z(n43202) );
  XOR U52657 ( .A(n43201), .B(n43202), .Z(n43204) );
  XOR U52658 ( .A(n43205), .B(n43204), .Z(n39729) );
  NOR U52659 ( .A(n39728), .B(n39729), .Z(n39723) );
  IV U52660 ( .A(n39723), .Z(n39727) );
  IV U52661 ( .A(n39724), .Z(n39726) );
  NOR U52662 ( .A(n39726), .B(n39725), .Z(n39732) );
  NOR U52663 ( .A(n39727), .B(n39732), .Z(n39736) );
  IV U52664 ( .A(n39728), .Z(n39731) );
  IV U52665 ( .A(n39729), .Z(n39730) );
  NOR U52666 ( .A(n39731), .B(n39730), .Z(n46388) );
  IV U52667 ( .A(n39732), .Z(n39733) );
  NOR U52668 ( .A(n39733), .B(n43204), .Z(n42234) );
  NOR U52669 ( .A(n46388), .B(n42234), .Z(n39734) );
  IV U52670 ( .A(n39734), .Z(n39735) );
  NOR U52671 ( .A(n39736), .B(n39735), .Z(n39737) );
  IV U52672 ( .A(n39737), .Z(n42227) );
  XOR U52673 ( .A(n39738), .B(n42227), .Z(n46401) );
  XOR U52674 ( .A(n42221), .B(n46401), .Z(n42222) );
  IV U52675 ( .A(n39739), .Z(n39741) );
  NOR U52676 ( .A(n39741), .B(n39740), .Z(n48896) );
  IV U52677 ( .A(n39742), .Z(n39744) );
  NOR U52678 ( .A(n39744), .B(n39743), .Z(n49797) );
  NOR U52679 ( .A(n48896), .B(n49797), .Z(n45383) );
  XOR U52680 ( .A(n42222), .B(n45383), .Z(n42220) );
  XOR U52681 ( .A(n42218), .B(n42220), .Z(n43215) );
  XOR U52682 ( .A(n39745), .B(n43215), .Z(n42215) );
  XOR U52683 ( .A(n39746), .B(n42215), .Z(n43218) );
  XOR U52684 ( .A(n43216), .B(n43218), .Z(n43221) );
  IV U52685 ( .A(n39747), .Z(n39750) );
  IV U52686 ( .A(n39748), .Z(n39749) );
  NOR U52687 ( .A(n39750), .B(n39749), .Z(n43219) );
  XOR U52688 ( .A(n43221), .B(n43219), .Z(n43223) );
  XOR U52689 ( .A(n42200), .B(n43223), .Z(n46411) );
  NOR U52690 ( .A(n46423), .B(n46410), .Z(n43234) );
  XOR U52691 ( .A(n46411), .B(n43234), .Z(n43236) );
  XOR U52692 ( .A(n39751), .B(n43236), .Z(n43244) );
  IV U52693 ( .A(n39752), .Z(n39753) );
  NOR U52694 ( .A(n39754), .B(n39753), .Z(n42197) );
  NOR U52695 ( .A(n43243), .B(n42197), .Z(n39755) );
  XOR U52696 ( .A(n43244), .B(n39755), .Z(n42192) );
  IV U52697 ( .A(n39756), .Z(n39757) );
  NOR U52698 ( .A(n39758), .B(n39757), .Z(n42194) );
  IV U52699 ( .A(n39759), .Z(n39760) );
  NOR U52700 ( .A(n39761), .B(n39760), .Z(n42191) );
  NOR U52701 ( .A(n42194), .B(n42191), .Z(n39762) );
  XOR U52702 ( .A(n42192), .B(n39762), .Z(n43251) );
  XOR U52703 ( .A(n39763), .B(n43251), .Z(n43253) );
  XOR U52704 ( .A(n39764), .B(n43253), .Z(n42187) );
  XOR U52705 ( .A(n42185), .B(n42187), .Z(n43260) );
  IV U52706 ( .A(n39765), .Z(n39767) );
  NOR U52707 ( .A(n39767), .B(n39766), .Z(n43258) );
  XOR U52708 ( .A(n43260), .B(n43258), .Z(n43261) );
  XOR U52709 ( .A(n43262), .B(n43261), .Z(n42177) );
  IV U52710 ( .A(n39768), .Z(n39769) );
  NOR U52711 ( .A(n39770), .B(n39769), .Z(n42176) );
  IV U52712 ( .A(n39771), .Z(n39772) );
  NOR U52713 ( .A(n39773), .B(n39772), .Z(n42182) );
  NOR U52714 ( .A(n42176), .B(n42182), .Z(n39774) );
  XOR U52715 ( .A(n42177), .B(n39774), .Z(n42179) );
  XOR U52716 ( .A(n42180), .B(n42179), .Z(n42171) );
  IV U52717 ( .A(n39775), .Z(n39776) );
  NOR U52718 ( .A(n39781), .B(n39776), .Z(n42172) );
  IV U52719 ( .A(n39777), .Z(n39778) );
  NOR U52720 ( .A(n39779), .B(n39778), .Z(n48852) );
  IV U52721 ( .A(n39780), .Z(n39782) );
  NOR U52722 ( .A(n39782), .B(n39781), .Z(n49865) );
  NOR U52723 ( .A(n48852), .B(n49865), .Z(n42175) );
  IV U52724 ( .A(n42175), .Z(n39783) );
  NOR U52725 ( .A(n42172), .B(n39783), .Z(n39784) );
  XOR U52726 ( .A(n42171), .B(n39784), .Z(n43267) );
  IV U52727 ( .A(n39785), .Z(n39786) );
  NOR U52728 ( .A(n39787), .B(n39786), .Z(n43265) );
  XOR U52729 ( .A(n43267), .B(n43265), .Z(n43269) );
  XOR U52730 ( .A(n43268), .B(n43269), .Z(n42169) );
  IV U52731 ( .A(n39788), .Z(n39789) );
  NOR U52732 ( .A(n39790), .B(n39789), .Z(n42168) );
  IV U52733 ( .A(n39791), .Z(n39793) );
  NOR U52734 ( .A(n39793), .B(n39792), .Z(n42166) );
  NOR U52735 ( .A(n42168), .B(n42166), .Z(n39794) );
  XOR U52736 ( .A(n42169), .B(n39794), .Z(n42150) );
  XOR U52737 ( .A(n39795), .B(n42150), .Z(n42148) );
  XOR U52738 ( .A(n39796), .B(n42148), .Z(n42142) );
  XOR U52739 ( .A(n39797), .B(n42142), .Z(n43275) );
  XOR U52740 ( .A(n43273), .B(n43275), .Z(n42136) );
  XOR U52741 ( .A(n42135), .B(n42136), .Z(n42140) );
  IV U52742 ( .A(n42140), .Z(n39805) );
  IV U52743 ( .A(n39798), .Z(n39800) );
  NOR U52744 ( .A(n39800), .B(n39799), .Z(n42133) );
  IV U52745 ( .A(n39801), .Z(n39803) );
  NOR U52746 ( .A(n39803), .B(n39802), .Z(n42138) );
  NOR U52747 ( .A(n42133), .B(n42138), .Z(n39804) );
  XOR U52748 ( .A(n39805), .B(n39804), .Z(n43283) );
  XOR U52749 ( .A(n43281), .B(n43283), .Z(n43284) );
  NOR U52750 ( .A(n39817), .B(n43284), .Z(n39806) );
  IV U52751 ( .A(n39806), .Z(n39811) );
  NOR U52752 ( .A(n39808), .B(n39807), .Z(n39809) );
  IV U52753 ( .A(n39809), .Z(n39810) );
  NOR U52754 ( .A(n39811), .B(n39810), .Z(n45291) );
  IV U52755 ( .A(n39812), .Z(n39814) );
  NOR U52756 ( .A(n39814), .B(n39813), .Z(n39820) );
  IV U52757 ( .A(n39815), .Z(n39816) );
  NOR U52758 ( .A(n39817), .B(n39816), .Z(n39818) );
  IV U52759 ( .A(n39818), .Z(n43285) );
  XOR U52760 ( .A(n43285), .B(n43284), .Z(n39819) );
  NOR U52761 ( .A(n39820), .B(n39819), .Z(n39821) );
  NOR U52762 ( .A(n45291), .B(n39821), .Z(n43291) );
  XOR U52763 ( .A(n39822), .B(n43291), .Z(n43295) );
  XOR U52764 ( .A(n42128), .B(n43295), .Z(n48815) );
  XOR U52765 ( .A(n42122), .B(n48815), .Z(n42124) );
  XOR U52766 ( .A(n39823), .B(n42124), .Z(n43312) );
  XOR U52767 ( .A(n43310), .B(n43312), .Z(n43314) );
  XOR U52768 ( .A(n43313), .B(n43314), .Z(n43317) );
  XOR U52769 ( .A(n43318), .B(n43317), .Z(n43320) );
  NOR U52770 ( .A(n39825), .B(n39824), .Z(n43319) );
  IV U52771 ( .A(n39826), .Z(n39828) );
  NOR U52772 ( .A(n39828), .B(n39827), .Z(n43323) );
  NOR U52773 ( .A(n43319), .B(n43323), .Z(n39829) );
  XOR U52774 ( .A(n43320), .B(n39829), .Z(n43328) );
  XOR U52775 ( .A(n43326), .B(n43328), .Z(n42120) );
  XOR U52776 ( .A(n42119), .B(n42120), .Z(n42115) );
  XOR U52777 ( .A(n39830), .B(n42115), .Z(n42109) );
  XOR U52778 ( .A(n42108), .B(n42109), .Z(n42101) );
  IV U52779 ( .A(n39831), .Z(n39832) );
  NOR U52780 ( .A(n39833), .B(n39832), .Z(n42110) );
  IV U52781 ( .A(n39834), .Z(n42102) );
  NOR U52782 ( .A(n39835), .B(n43333), .Z(n39836) );
  IV U52783 ( .A(n39836), .Z(n39840) );
  NOR U52784 ( .A(n42102), .B(n39840), .Z(n39837) );
  NOR U52785 ( .A(n42110), .B(n39837), .Z(n39838) );
  XOR U52786 ( .A(n42101), .B(n39838), .Z(n42100) );
  IV U52787 ( .A(n39839), .Z(n39841) );
  NOR U52788 ( .A(n39841), .B(n39840), .Z(n42098) );
  XOR U52789 ( .A(n42100), .B(n42098), .Z(n43338) );
  XOR U52790 ( .A(n39842), .B(n43338), .Z(n43341) );
  IV U52791 ( .A(n39843), .Z(n39844) );
  NOR U52792 ( .A(n39844), .B(n39853), .Z(n39845) );
  IV U52793 ( .A(n39845), .Z(n43340) );
  XOR U52794 ( .A(n43341), .B(n43340), .Z(n39846) );
  NOR U52795 ( .A(n39847), .B(n39846), .Z(n39850) );
  IV U52796 ( .A(n39847), .Z(n39849) );
  XOR U52797 ( .A(n42092), .B(n43338), .Z(n39848) );
  NOR U52798 ( .A(n39849), .B(n39848), .Z(n46528) );
  NOR U52799 ( .A(n39850), .B(n46528), .Z(n39851) );
  IV U52800 ( .A(n39851), .Z(n43345) );
  IV U52801 ( .A(n39852), .Z(n39854) );
  NOR U52802 ( .A(n39854), .B(n39853), .Z(n43343) );
  XOR U52803 ( .A(n39855), .B(n42075), .Z(n42072) );
  NOR U52804 ( .A(n39862), .B(n42072), .Z(n48770) );
  IV U52805 ( .A(n39856), .Z(n39857) );
  NOR U52806 ( .A(n39870), .B(n39857), .Z(n42068) );
  IV U52807 ( .A(n39858), .Z(n39860) );
  NOR U52808 ( .A(n39860), .B(n39859), .Z(n39861) );
  IV U52809 ( .A(n39861), .Z(n42073) );
  XOR U52810 ( .A(n42073), .B(n42072), .Z(n42069) );
  XOR U52811 ( .A(n42068), .B(n42069), .Z(n39864) );
  NOR U52812 ( .A(n42069), .B(n39862), .Z(n39863) );
  NOR U52813 ( .A(n39864), .B(n39863), .Z(n39865) );
  NOR U52814 ( .A(n48770), .B(n39865), .Z(n42063) );
  IV U52815 ( .A(n39866), .Z(n39867) );
  NOR U52816 ( .A(n39868), .B(n39867), .Z(n42062) );
  IV U52817 ( .A(n39869), .Z(n39871) );
  NOR U52818 ( .A(n39871), .B(n39870), .Z(n42065) );
  NOR U52819 ( .A(n42062), .B(n42065), .Z(n39872) );
  XOR U52820 ( .A(n42063), .B(n39872), .Z(n43359) );
  XOR U52821 ( .A(n39873), .B(n43359), .Z(n42059) );
  XOR U52822 ( .A(n39874), .B(n42059), .Z(n42057) );
  NOR U52823 ( .A(n39885), .B(n42057), .Z(n39875) );
  IV U52824 ( .A(n39875), .Z(n39876) );
  NOR U52825 ( .A(n39877), .B(n39876), .Z(n52508) );
  NOR U52826 ( .A(n39878), .B(n39877), .Z(n39882) );
  IV U52827 ( .A(n39882), .Z(n42058) );
  XOR U52828 ( .A(n42058), .B(n42057), .Z(n39887) );
  NOR U52829 ( .A(n39880), .B(n39879), .Z(n39881) );
  NOR U52830 ( .A(n39882), .B(n39881), .Z(n39883) );
  IV U52831 ( .A(n39883), .Z(n39884) );
  NOR U52832 ( .A(n39885), .B(n39884), .Z(n39886) );
  NOR U52833 ( .A(n39887), .B(n39886), .Z(n39888) );
  NOR U52834 ( .A(n52508), .B(n39888), .Z(n43364) );
  IV U52835 ( .A(n39889), .Z(n39891) );
  NOR U52836 ( .A(n39891), .B(n39890), .Z(n39892) );
  IV U52837 ( .A(n39892), .Z(n43365) );
  XOR U52838 ( .A(n43364), .B(n43365), .Z(n42055) );
  XOR U52839 ( .A(n39893), .B(n42055), .Z(n42045) );
  IV U52840 ( .A(n39894), .Z(n39897) );
  IV U52841 ( .A(n39895), .Z(n39896) );
  NOR U52842 ( .A(n39897), .B(n39896), .Z(n42050) );
  IV U52843 ( .A(n39898), .Z(n39900) );
  IV U52844 ( .A(n39899), .Z(n39903) );
  NOR U52845 ( .A(n39900), .B(n39903), .Z(n42044) );
  NOR U52846 ( .A(n42050), .B(n42044), .Z(n39901) );
  XOR U52847 ( .A(n42045), .B(n39901), .Z(n43371) );
  IV U52848 ( .A(n39902), .Z(n39904) );
  NOR U52849 ( .A(n39904), .B(n39903), .Z(n43369) );
  XOR U52850 ( .A(n43371), .B(n43369), .Z(n46555) );
  NOR U52851 ( .A(n39909), .B(n46555), .Z(n45223) );
  IV U52852 ( .A(n39905), .Z(n39906) );
  NOR U52853 ( .A(n39914), .B(n39906), .Z(n42040) );
  NOR U52854 ( .A(n46558), .B(n39907), .Z(n39908) );
  IV U52855 ( .A(n39908), .Z(n43372) );
  XOR U52856 ( .A(n43372), .B(n46555), .Z(n42041) );
  XOR U52857 ( .A(n42040), .B(n42041), .Z(n39911) );
  NOR U52858 ( .A(n42041), .B(n39909), .Z(n39910) );
  NOR U52859 ( .A(n39911), .B(n39910), .Z(n39912) );
  NOR U52860 ( .A(n45223), .B(n39912), .Z(n42035) );
  IV U52861 ( .A(n39913), .Z(n39915) );
  NOR U52862 ( .A(n39915), .B(n39914), .Z(n39916) );
  IV U52863 ( .A(n39916), .Z(n42037) );
  XOR U52864 ( .A(n42035), .B(n42037), .Z(n43377) );
  XOR U52865 ( .A(n42038), .B(n43377), .Z(n43380) );
  XOR U52866 ( .A(n39917), .B(n43380), .Z(n43385) );
  XOR U52867 ( .A(n43383), .B(n43385), .Z(n46587) );
  IV U52868 ( .A(n39918), .Z(n39919) );
  NOR U52869 ( .A(n39920), .B(n39919), .Z(n46585) );
  IV U52870 ( .A(n39921), .Z(n39923) );
  NOR U52871 ( .A(n39923), .B(n39922), .Z(n46593) );
  NOR U52872 ( .A(n46585), .B(n46593), .Z(n43386) );
  XOR U52873 ( .A(n46587), .B(n43386), .Z(n42029) );
  XOR U52874 ( .A(n39924), .B(n42029), .Z(n48713) );
  XOR U52875 ( .A(n42031), .B(n48713), .Z(n39925) );
  IV U52876 ( .A(n39925), .Z(n42024) );
  XOR U52877 ( .A(n42021), .B(n42024), .Z(n42020) );
  IV U52878 ( .A(n39926), .Z(n48709) );
  NOR U52879 ( .A(n48709), .B(n39931), .Z(n39927) );
  IV U52880 ( .A(n39927), .Z(n39939) );
  NOR U52881 ( .A(n42020), .B(n39939), .Z(n43397) );
  IV U52882 ( .A(n39928), .Z(n42025) );
  NOR U52883 ( .A(n39929), .B(n42025), .Z(n39933) );
  IV U52884 ( .A(n39930), .Z(n39932) );
  NOR U52885 ( .A(n39932), .B(n39931), .Z(n42018) );
  NOR U52886 ( .A(n39933), .B(n42018), .Z(n39934) );
  IV U52887 ( .A(n39934), .Z(n39935) );
  XOR U52888 ( .A(n39935), .B(n42020), .Z(n43403) );
  IV U52889 ( .A(n39936), .Z(n39947) );
  IV U52890 ( .A(n39937), .Z(n39938) );
  NOR U52891 ( .A(n39947), .B(n39938), .Z(n39940) );
  IV U52892 ( .A(n39940), .Z(n43402) );
  XOR U52893 ( .A(n43403), .B(n43402), .Z(n39942) );
  NOR U52894 ( .A(n39940), .B(n39939), .Z(n39941) );
  NOR U52895 ( .A(n39942), .B(n39941), .Z(n39943) );
  NOR U52896 ( .A(n43397), .B(n39943), .Z(n39944) );
  IV U52897 ( .A(n39944), .Z(n43407) );
  IV U52898 ( .A(n39945), .Z(n39946) );
  NOR U52899 ( .A(n39947), .B(n39946), .Z(n43405) );
  XOR U52900 ( .A(n43407), .B(n43405), .Z(n43413) );
  IV U52901 ( .A(n39948), .Z(n39950) );
  NOR U52902 ( .A(n39950), .B(n39949), .Z(n43408) );
  IV U52903 ( .A(n39951), .Z(n39952) );
  NOR U52904 ( .A(n39952), .B(n39958), .Z(n43411) );
  NOR U52905 ( .A(n43408), .B(n43411), .Z(n39953) );
  XOR U52906 ( .A(n43413), .B(n39953), .Z(n42015) );
  IV U52907 ( .A(n39954), .Z(n39963) );
  IV U52908 ( .A(n39955), .Z(n39956) );
  NOR U52909 ( .A(n39963), .B(n39956), .Z(n43417) );
  IV U52910 ( .A(n39957), .Z(n39959) );
  NOR U52911 ( .A(n39959), .B(n39958), .Z(n42016) );
  NOR U52912 ( .A(n43417), .B(n42016), .Z(n39960) );
  XOR U52913 ( .A(n42015), .B(n39960), .Z(n42013) );
  IV U52914 ( .A(n39961), .Z(n39962) );
  NOR U52915 ( .A(n39963), .B(n39962), .Z(n42011) );
  XOR U52916 ( .A(n42013), .B(n42011), .Z(n43415) );
  XOR U52917 ( .A(n43414), .B(n43415), .Z(n42010) );
  IV U52918 ( .A(n39964), .Z(n39965) );
  NOR U52919 ( .A(n42002), .B(n39965), .Z(n42006) );
  IV U52920 ( .A(n39966), .Z(n39968) );
  NOR U52921 ( .A(n39968), .B(n39967), .Z(n42008) );
  NOR U52922 ( .A(n42006), .B(n42008), .Z(n39969) );
  XOR U52923 ( .A(n42010), .B(n39969), .Z(n41989) );
  NOR U52924 ( .A(n39971), .B(n39970), .Z(n41995) );
  IV U52925 ( .A(n39972), .Z(n39974) );
  NOR U52926 ( .A(n39974), .B(n39973), .Z(n41992) );
  NOR U52927 ( .A(n41995), .B(n41992), .Z(n39975) );
  XOR U52928 ( .A(n41989), .B(n39975), .Z(n41986) );
  IV U52929 ( .A(n39976), .Z(n39978) );
  NOR U52930 ( .A(n39978), .B(n39977), .Z(n41988) );
  NOR U52931 ( .A(n39980), .B(n39979), .Z(n41985) );
  NOR U52932 ( .A(n41988), .B(n41985), .Z(n39981) );
  XOR U52933 ( .A(n41986), .B(n39981), .Z(n41979) );
  IV U52934 ( .A(n39982), .Z(n39983) );
  NOR U52935 ( .A(n39984), .B(n39983), .Z(n41980) );
  NOR U52936 ( .A(n41982), .B(n41980), .Z(n39985) );
  XOR U52937 ( .A(n41979), .B(n39985), .Z(n43428) );
  NOR U52938 ( .A(n39986), .B(n41976), .Z(n39990) );
  IV U52939 ( .A(n39987), .Z(n39989) );
  IV U52940 ( .A(n39988), .Z(n39995) );
  NOR U52941 ( .A(n39989), .B(n39995), .Z(n43427) );
  NOR U52942 ( .A(n39990), .B(n43427), .Z(n39991) );
  XOR U52943 ( .A(n43428), .B(n39991), .Z(n43434) );
  IV U52944 ( .A(n39992), .Z(n39993) );
  NOR U52945 ( .A(n40001), .B(n39993), .Z(n50093) );
  IV U52946 ( .A(n39994), .Z(n39996) );
  NOR U52947 ( .A(n39996), .B(n39995), .Z(n48664) );
  NOR U52948 ( .A(n50093), .B(n48664), .Z(n43435) );
  XOR U52949 ( .A(n43434), .B(n43435), .Z(n43438) );
  IV U52950 ( .A(n39997), .Z(n39998) );
  NOR U52951 ( .A(n40004), .B(n39998), .Z(n41970) );
  IV U52952 ( .A(n39999), .Z(n40000) );
  NOR U52953 ( .A(n40001), .B(n40000), .Z(n43436) );
  NOR U52954 ( .A(n41970), .B(n43436), .Z(n40002) );
  XOR U52955 ( .A(n43438), .B(n40002), .Z(n41967) );
  IV U52956 ( .A(n40003), .Z(n40005) );
  NOR U52957 ( .A(n40005), .B(n40004), .Z(n41972) );
  NOR U52958 ( .A(n41968), .B(n41972), .Z(n40006) );
  XOR U52959 ( .A(n41967), .B(n40006), .Z(n45160) );
  IV U52960 ( .A(n40007), .Z(n40008) );
  NOR U52961 ( .A(n40009), .B(n40008), .Z(n45159) );
  NOR U52962 ( .A(n46645), .B(n45159), .Z(n43441) );
  XOR U52963 ( .A(n45160), .B(n43441), .Z(n40014) );
  IV U52964 ( .A(n40014), .Z(n43447) );
  XOR U52965 ( .A(n43442), .B(n43447), .Z(n40010) );
  NOR U52966 ( .A(n40011), .B(n40010), .Z(n45154) );
  IV U52967 ( .A(n40012), .Z(n40013) );
  NOR U52968 ( .A(n40018), .B(n40013), .Z(n43446) );
  NOR U52969 ( .A(n43442), .B(n43446), .Z(n40015) );
  XOR U52970 ( .A(n40015), .B(n40014), .Z(n43450) );
  IV U52971 ( .A(n40016), .Z(n40017) );
  NOR U52972 ( .A(n40018), .B(n40017), .Z(n40019) );
  IV U52973 ( .A(n40019), .Z(n43449) );
  XOR U52974 ( .A(n43450), .B(n43449), .Z(n41962) );
  NOR U52975 ( .A(n40020), .B(n41962), .Z(n40021) );
  NOR U52976 ( .A(n45154), .B(n40021), .Z(n40022) );
  IV U52977 ( .A(n40022), .Z(n41956) );
  XOR U52978 ( .A(n40023), .B(n41956), .Z(n41941) );
  NOR U52979 ( .A(n40024), .B(n41941), .Z(n40031) );
  XOR U52980 ( .A(n40025), .B(n41956), .Z(n40026) );
  NOR U52981 ( .A(n40027), .B(n40026), .Z(n40028) );
  IV U52982 ( .A(n40028), .Z(n41947) );
  NOR U52983 ( .A(n41947), .B(n40029), .Z(n40030) );
  NOR U52984 ( .A(n40031), .B(n40030), .Z(n41937) );
  IV U52985 ( .A(n40032), .Z(n40034) );
  NOR U52986 ( .A(n40034), .B(n40033), .Z(n41940) );
  IV U52987 ( .A(n40035), .Z(n40037) );
  NOR U52988 ( .A(n40037), .B(n40036), .Z(n41936) );
  NOR U52989 ( .A(n41940), .B(n41936), .Z(n40038) );
  XOR U52990 ( .A(n41937), .B(n40038), .Z(n41935) );
  XOR U52991 ( .A(n40039), .B(n41935), .Z(n40040) );
  IV U52992 ( .A(n40040), .Z(n45142) );
  XOR U52993 ( .A(n41931), .B(n45142), .Z(n43460) );
  XOR U52994 ( .A(n40041), .B(n43460), .Z(n43462) );
  XOR U52995 ( .A(n40042), .B(n43462), .Z(n41924) );
  XOR U52996 ( .A(n40043), .B(n41924), .Z(n43469) );
  XOR U52997 ( .A(n41920), .B(n43469), .Z(n41914) );
  IV U52998 ( .A(n40047), .Z(n40044) );
  NOR U52999 ( .A(n40044), .B(n40045), .Z(n43468) );
  IV U53000 ( .A(n40045), .Z(n40046) );
  NOR U53001 ( .A(n40047), .B(n40046), .Z(n40050) );
  IV U53002 ( .A(n40048), .Z(n40049) );
  NOR U53003 ( .A(n40050), .B(n40049), .Z(n40051) );
  NOR U53004 ( .A(n43468), .B(n40051), .Z(n41916) );
  XOR U53005 ( .A(n41914), .B(n41916), .Z(n43473) );
  XOR U53006 ( .A(n43471), .B(n43473), .Z(n43475) );
  XOR U53007 ( .A(n40052), .B(n43475), .Z(n41912) );
  XOR U53008 ( .A(n41911), .B(n41912), .Z(n43481) );
  IV U53009 ( .A(n40053), .Z(n40055) );
  NOR U53010 ( .A(n40055), .B(n40054), .Z(n43480) );
  IV U53011 ( .A(n40056), .Z(n40058) );
  NOR U53012 ( .A(n40058), .B(n40057), .Z(n43478) );
  NOR U53013 ( .A(n43480), .B(n43478), .Z(n40059) );
  XOR U53014 ( .A(n43481), .B(n40059), .Z(n40065) );
  IV U53015 ( .A(n40065), .Z(n40060) );
  NOR U53016 ( .A(n40061), .B(n40060), .Z(n45113) );
  IV U53017 ( .A(n40062), .Z(n40064) );
  NOR U53018 ( .A(n40064), .B(n40063), .Z(n40066) );
  NOR U53019 ( .A(n40066), .B(n40065), .Z(n40069) );
  IV U53020 ( .A(n40066), .Z(n40068) );
  XOR U53021 ( .A(n43480), .B(n43481), .Z(n40067) );
  NOR U53022 ( .A(n40068), .B(n40067), .Z(n45110) );
  NOR U53023 ( .A(n40069), .B(n45110), .Z(n40070) );
  NOR U53024 ( .A(n40071), .B(n40070), .Z(n40072) );
  NOR U53025 ( .A(n45113), .B(n40072), .Z(n41902) );
  IV U53026 ( .A(n40073), .Z(n40075) );
  NOR U53027 ( .A(n40075), .B(n40074), .Z(n41906) );
  NOR U53028 ( .A(n40076), .B(n43488), .Z(n40077) );
  NOR U53029 ( .A(n43490), .B(n40077), .Z(n40078) );
  NOR U53030 ( .A(n41906), .B(n40078), .Z(n40079) );
  XOR U53031 ( .A(n41902), .B(n40079), .Z(n43487) );
  IV U53032 ( .A(n40080), .Z(n40083) );
  IV U53033 ( .A(n40081), .Z(n40082) );
  NOR U53034 ( .A(n40083), .B(n40082), .Z(n43485) );
  XOR U53035 ( .A(n43487), .B(n43485), .Z(n41898) );
  IV U53036 ( .A(n40084), .Z(n40085) );
  NOR U53037 ( .A(n40086), .B(n40085), .Z(n41897) );
  IV U53038 ( .A(n40087), .Z(n40089) );
  NOR U53039 ( .A(n40089), .B(n40088), .Z(n41892) );
  NOR U53040 ( .A(n41897), .B(n41892), .Z(n40090) );
  XOR U53041 ( .A(n41898), .B(n40090), .Z(n40102) );
  IV U53042 ( .A(n40102), .Z(n41895) );
  IV U53043 ( .A(n40091), .Z(n40092) );
  NOR U53044 ( .A(n40092), .B(n40101), .Z(n40093) );
  IV U53045 ( .A(n40093), .Z(n40103) );
  NOR U53046 ( .A(n41895), .B(n40103), .Z(n46714) );
  IV U53047 ( .A(n40094), .Z(n40098) );
  NOR U53048 ( .A(n40096), .B(n40095), .Z(n40097) );
  IV U53049 ( .A(n40097), .Z(n40108) );
  NOR U53050 ( .A(n40098), .B(n40108), .Z(n41887) );
  IV U53051 ( .A(n40099), .Z(n40100) );
  NOR U53052 ( .A(n40101), .B(n40100), .Z(n41894) );
  XOR U53053 ( .A(n41894), .B(n40102), .Z(n41888) );
  XOR U53054 ( .A(n41887), .B(n41888), .Z(n40105) );
  NOR U53055 ( .A(n41888), .B(n40103), .Z(n40104) );
  NOR U53056 ( .A(n40105), .B(n40104), .Z(n40106) );
  NOR U53057 ( .A(n46714), .B(n40106), .Z(n43496) );
  IV U53058 ( .A(n40107), .Z(n40109) );
  NOR U53059 ( .A(n40109), .B(n40108), .Z(n40110) );
  IV U53060 ( .A(n40110), .Z(n43497) );
  XOR U53061 ( .A(n43496), .B(n43497), .Z(n43503) );
  IV U53062 ( .A(n40111), .Z(n40112) );
  NOR U53063 ( .A(n40113), .B(n40112), .Z(n43499) );
  NOR U53064 ( .A(n40115), .B(n40114), .Z(n43502) );
  NOR U53065 ( .A(n43499), .B(n43502), .Z(n40116) );
  XOR U53066 ( .A(n43503), .B(n40116), .Z(n41882) );
  XOR U53067 ( .A(n41883), .B(n41882), .Z(n43507) );
  IV U53068 ( .A(n40117), .Z(n40118) );
  NOR U53069 ( .A(n40119), .B(n40118), .Z(n41880) );
  IV U53070 ( .A(n40120), .Z(n40121) );
  NOR U53071 ( .A(n45081), .B(n40121), .Z(n43508) );
  NOR U53072 ( .A(n41880), .B(n43508), .Z(n40122) );
  XOR U53073 ( .A(n43507), .B(n40122), .Z(n43512) );
  XOR U53074 ( .A(n40123), .B(n43512), .Z(n43520) );
  XOR U53075 ( .A(n40124), .B(n43520), .Z(n43527) );
  XOR U53076 ( .A(n40125), .B(n43527), .Z(n43523) );
  XOR U53077 ( .A(n40126), .B(n43523), .Z(n41871) );
  XOR U53078 ( .A(n41869), .B(n41871), .Z(n41874) );
  IV U53079 ( .A(n40127), .Z(n40129) );
  NOR U53080 ( .A(n40129), .B(n40128), .Z(n41872) );
  XOR U53081 ( .A(n41874), .B(n41872), .Z(n41866) );
  XOR U53082 ( .A(n41865), .B(n41866), .Z(n43533) );
  XOR U53083 ( .A(n43534), .B(n43533), .Z(n43535) );
  IV U53084 ( .A(n40130), .Z(n40131) );
  NOR U53085 ( .A(n40131), .B(n40133), .Z(n43536) );
  IV U53086 ( .A(n40132), .Z(n40136) );
  NOR U53087 ( .A(n40134), .B(n40133), .Z(n40135) );
  IV U53088 ( .A(n40135), .Z(n40139) );
  NOR U53089 ( .A(n40136), .B(n40139), .Z(n43539) );
  NOR U53090 ( .A(n43536), .B(n43539), .Z(n40137) );
  XOR U53091 ( .A(n43535), .B(n40137), .Z(n41861) );
  IV U53092 ( .A(n40138), .Z(n40140) );
  NOR U53093 ( .A(n40140), .B(n40139), .Z(n41859) );
  XOR U53094 ( .A(n41861), .B(n41859), .Z(n41863) );
  XOR U53095 ( .A(n41862), .B(n41863), .Z(n43549) );
  XOR U53096 ( .A(n40141), .B(n43549), .Z(n41853) );
  XOR U53097 ( .A(n40142), .B(n41853), .Z(n41857) );
  XOR U53098 ( .A(n41856), .B(n41857), .Z(n43555) );
  XOR U53099 ( .A(n40143), .B(n43555), .Z(n43572) );
  XOR U53100 ( .A(n40144), .B(n43572), .Z(n41852) );
  XOR U53101 ( .A(n40145), .B(n41852), .Z(n40146) );
  IV U53102 ( .A(n40146), .Z(n41848) );
  XOR U53103 ( .A(n41847), .B(n41848), .Z(n41843) );
  XOR U53104 ( .A(n41841), .B(n41843), .Z(n41845) );
  XOR U53105 ( .A(n41844), .B(n41845), .Z(n41833) );
  XOR U53106 ( .A(n41832), .B(n41833), .Z(n41836) );
  NOR U53107 ( .A(n40153), .B(n41836), .Z(n45041) );
  IV U53108 ( .A(n40147), .Z(n40148) );
  NOR U53109 ( .A(n40149), .B(n40148), .Z(n41823) );
  IV U53110 ( .A(n40150), .Z(n41837) );
  NOR U53111 ( .A(n41837), .B(n40151), .Z(n40152) );
  IV U53112 ( .A(n40152), .Z(n41828) );
  XOR U53113 ( .A(n41828), .B(n41836), .Z(n41824) );
  XOR U53114 ( .A(n41823), .B(n41824), .Z(n40155) );
  NOR U53115 ( .A(n41824), .B(n40153), .Z(n40154) );
  NOR U53116 ( .A(n40155), .B(n40154), .Z(n40156) );
  NOR U53117 ( .A(n45041), .B(n40156), .Z(n41816) );
  IV U53118 ( .A(n40157), .Z(n40158) );
  NOR U53119 ( .A(n40159), .B(n40158), .Z(n40160) );
  IV U53120 ( .A(n40160), .Z(n41818) );
  XOR U53121 ( .A(n41816), .B(n41818), .Z(n41820) );
  XOR U53122 ( .A(n40161), .B(n41820), .Z(n41811) );
  IV U53123 ( .A(n40162), .Z(n40163) );
  NOR U53124 ( .A(n40164), .B(n40163), .Z(n43581) );
  IV U53125 ( .A(n40165), .Z(n40167) );
  NOR U53126 ( .A(n40167), .B(n40166), .Z(n41812) );
  NOR U53127 ( .A(n43581), .B(n41812), .Z(n40168) );
  XOR U53128 ( .A(n41811), .B(n40168), .Z(n43585) );
  XOR U53129 ( .A(n43584), .B(n43585), .Z(n43590) );
  XOR U53130 ( .A(n43588), .B(n43590), .Z(n43593) );
  XOR U53131 ( .A(n43591), .B(n43593), .Z(n41809) );
  XOR U53132 ( .A(n41807), .B(n41809), .Z(n43597) );
  XOR U53133 ( .A(n43595), .B(n43597), .Z(n43600) );
  XOR U53134 ( .A(n43598), .B(n43600), .Z(n43603) );
  XOR U53135 ( .A(n40169), .B(n43603), .Z(n43610) );
  XOR U53136 ( .A(n43608), .B(n43610), .Z(n41803) );
  IV U53137 ( .A(n40170), .Z(n40172) );
  NOR U53138 ( .A(n40172), .B(n40171), .Z(n41801) );
  XOR U53139 ( .A(n41803), .B(n41801), .Z(n43606) );
  XOR U53140 ( .A(n43605), .B(n43606), .Z(n41798) );
  IV U53141 ( .A(n40173), .Z(n40174) );
  NOR U53142 ( .A(n40175), .B(n40174), .Z(n41797) );
  IV U53143 ( .A(n40176), .Z(n40178) );
  NOR U53144 ( .A(n40178), .B(n40177), .Z(n41792) );
  NOR U53145 ( .A(n41797), .B(n41792), .Z(n40179) );
  XOR U53146 ( .A(n41798), .B(n40179), .Z(n41790) );
  XOR U53147 ( .A(n40180), .B(n41790), .Z(n41788) );
  XOR U53148 ( .A(n40181), .B(n41788), .Z(n41775) );
  XOR U53149 ( .A(n40182), .B(n41775), .Z(n44985) );
  XOR U53150 ( .A(n43618), .B(n44985), .Z(n43620) );
  XOR U53151 ( .A(n40183), .B(n43620), .Z(n41773) );
  IV U53152 ( .A(n40184), .Z(n40185) );
  NOR U53153 ( .A(n40186), .B(n40185), .Z(n41766) );
  IV U53154 ( .A(n40187), .Z(n40188) );
  NOR U53155 ( .A(n40189), .B(n40188), .Z(n41771) );
  NOR U53156 ( .A(n41766), .B(n41771), .Z(n40190) );
  XOR U53157 ( .A(n41773), .B(n40190), .Z(n41769) );
  XOR U53158 ( .A(n40191), .B(n41769), .Z(n43629) );
  XOR U53159 ( .A(n40192), .B(n43629), .Z(n40193) );
  IV U53160 ( .A(n40193), .Z(n41760) );
  XOR U53161 ( .A(n41759), .B(n41760), .Z(n44974) );
  XOR U53162 ( .A(n41762), .B(n44974), .Z(n40194) );
  IV U53163 ( .A(n40194), .Z(n41755) );
  IV U53164 ( .A(n40195), .Z(n40196) );
  NOR U53165 ( .A(n40199), .B(n40196), .Z(n41753) );
  XOR U53166 ( .A(n41755), .B(n41753), .Z(n41758) );
  IV U53167 ( .A(n40197), .Z(n40198) );
  NOR U53168 ( .A(n40199), .B(n40198), .Z(n41756) );
  XOR U53169 ( .A(n41758), .B(n41756), .Z(n41749) );
  XOR U53170 ( .A(n41748), .B(n41749), .Z(n54159) );
  XOR U53171 ( .A(n41751), .B(n54159), .Z(n43636) );
  IV U53172 ( .A(n40200), .Z(n40202) );
  NOR U53173 ( .A(n40202), .B(n40201), .Z(n43639) );
  NOR U53174 ( .A(n43635), .B(n43639), .Z(n40203) );
  XOR U53175 ( .A(n43636), .B(n40203), .Z(n43643) );
  XOR U53176 ( .A(n43641), .B(n43643), .Z(n43645) );
  XOR U53177 ( .A(n43644), .B(n43645), .Z(n43648) );
  IV U53178 ( .A(n43648), .Z(n43650) );
  XOR U53179 ( .A(n43649), .B(n43650), .Z(n43659) );
  NOR U53180 ( .A(n40209), .B(n43659), .Z(n46880) );
  NOR U53181 ( .A(n40205), .B(n40204), .Z(n41743) );
  IV U53182 ( .A(n40206), .Z(n43653) );
  NOR U53183 ( .A(n40207), .B(n43653), .Z(n40208) );
  IV U53184 ( .A(n40208), .Z(n43660) );
  XOR U53185 ( .A(n43660), .B(n43659), .Z(n41744) );
  XOR U53186 ( .A(n41743), .B(n41744), .Z(n40211) );
  NOR U53187 ( .A(n41744), .B(n40209), .Z(n40210) );
  NOR U53188 ( .A(n40211), .B(n40210), .Z(n40212) );
  NOR U53189 ( .A(n46880), .B(n40212), .Z(n41741) );
  XOR U53190 ( .A(n41742), .B(n41741), .Z(n41738) );
  IV U53191 ( .A(n40213), .Z(n40219) );
  IV U53192 ( .A(n40214), .Z(n40216) );
  NOR U53193 ( .A(n40216), .B(n40215), .Z(n40217) );
  IV U53194 ( .A(n40217), .Z(n40218) );
  NOR U53195 ( .A(n40219), .B(n40218), .Z(n41736) );
  XOR U53196 ( .A(n41738), .B(n41736), .Z(n43676) );
  IV U53197 ( .A(n40220), .Z(n40221) );
  NOR U53198 ( .A(n40222), .B(n40221), .Z(n41739) );
  NOR U53199 ( .A(n40223), .B(n43677), .Z(n40224) );
  NOR U53200 ( .A(n41739), .B(n40224), .Z(n40225) );
  XOR U53201 ( .A(n43676), .B(n40225), .Z(n43681) );
  IV U53202 ( .A(n40226), .Z(n40228) );
  IV U53203 ( .A(n40227), .Z(n40234) );
  NOR U53204 ( .A(n40228), .B(n40234), .Z(n40229) );
  IV U53205 ( .A(n40229), .Z(n43682) );
  XOR U53206 ( .A(n43681), .B(n43682), .Z(n41729) );
  NOR U53207 ( .A(n40237), .B(n41729), .Z(n46916) );
  IV U53208 ( .A(n40230), .Z(n40232) );
  NOR U53209 ( .A(n40232), .B(n40231), .Z(n41731) );
  IV U53210 ( .A(n40233), .Z(n40235) );
  NOR U53211 ( .A(n40235), .B(n40234), .Z(n40236) );
  IV U53212 ( .A(n40236), .Z(n41730) );
  XOR U53213 ( .A(n41730), .B(n41729), .Z(n41732) );
  XOR U53214 ( .A(n41731), .B(n41732), .Z(n40239) );
  NOR U53215 ( .A(n41732), .B(n40237), .Z(n40238) );
  NOR U53216 ( .A(n40239), .B(n40238), .Z(n40240) );
  NOR U53217 ( .A(n46916), .B(n40240), .Z(n41727) );
  XOR U53218 ( .A(n40241), .B(n41727), .Z(n46925) );
  XOR U53219 ( .A(n43693), .B(n46925), .Z(n43695) );
  XOR U53220 ( .A(n40242), .B(n43695), .Z(n43705) );
  XOR U53221 ( .A(n43703), .B(n43705), .Z(n41724) );
  XOR U53222 ( .A(n41723), .B(n41724), .Z(n43716) );
  XOR U53223 ( .A(n43709), .B(n43716), .Z(n43713) );
  IV U53224 ( .A(n40243), .Z(n40244) );
  NOR U53225 ( .A(n40245), .B(n40244), .Z(n43715) );
  IV U53226 ( .A(n40246), .Z(n40248) );
  NOR U53227 ( .A(n40248), .B(n40247), .Z(n43711) );
  NOR U53228 ( .A(n43715), .B(n43711), .Z(n40249) );
  XOR U53229 ( .A(n43713), .B(n40249), .Z(n40250) );
  IV U53230 ( .A(n40250), .Z(n41722) );
  IV U53231 ( .A(n40251), .Z(n40253) );
  NOR U53232 ( .A(n40253), .B(n40252), .Z(n41720) );
  IV U53233 ( .A(n40254), .Z(n40255) );
  NOR U53234 ( .A(n40255), .B(n40261), .Z(n41718) );
  NOR U53235 ( .A(n41720), .B(n41718), .Z(n40256) );
  XOR U53236 ( .A(n41722), .B(n40256), .Z(n41713) );
  IV U53237 ( .A(n40257), .Z(n40258) );
  NOR U53238 ( .A(n40259), .B(n40258), .Z(n41712) );
  IV U53239 ( .A(n40260), .Z(n40262) );
  NOR U53240 ( .A(n40262), .B(n40261), .Z(n41715) );
  NOR U53241 ( .A(n41712), .B(n41715), .Z(n40263) );
  XOR U53242 ( .A(n41713), .B(n40263), .Z(n41706) );
  XOR U53243 ( .A(n40264), .B(n41706), .Z(n41699) );
  IV U53244 ( .A(n40265), .Z(n40267) );
  NOR U53245 ( .A(n40267), .B(n40266), .Z(n41697) );
  XOR U53246 ( .A(n41699), .B(n41697), .Z(n41701) );
  XOR U53247 ( .A(n41700), .B(n41701), .Z(n43721) );
  XOR U53248 ( .A(n40268), .B(n43721), .Z(n43723) );
  IV U53249 ( .A(n40285), .Z(n40272) );
  NOR U53250 ( .A(n40269), .B(n40281), .Z(n40270) );
  IV U53251 ( .A(n40270), .Z(n40271) );
  NOR U53252 ( .A(n40272), .B(n40271), .Z(n43726) );
  IV U53253 ( .A(n40273), .Z(n40274) );
  NOR U53254 ( .A(n40275), .B(n40274), .Z(n43722) );
  NOR U53255 ( .A(n43726), .B(n43722), .Z(n40276) );
  XOR U53256 ( .A(n43723), .B(n40276), .Z(n43735) );
  IV U53257 ( .A(n40277), .Z(n40278) );
  NOR U53258 ( .A(n40279), .B(n40278), .Z(n43733) );
  IV U53259 ( .A(n40280), .Z(n40282) );
  NOR U53260 ( .A(n40282), .B(n40281), .Z(n40283) );
  IV U53261 ( .A(n40283), .Z(n40284) );
  NOR U53262 ( .A(n40285), .B(n40284), .Z(n43729) );
  NOR U53263 ( .A(n43733), .B(n43729), .Z(n40286) );
  XOR U53264 ( .A(n43735), .B(n40286), .Z(n43731) );
  XOR U53265 ( .A(n43732), .B(n43731), .Z(n43743) );
  XOR U53266 ( .A(n43742), .B(n43743), .Z(n43738) );
  XOR U53267 ( .A(n43739), .B(n43738), .Z(n41690) );
  NOR U53268 ( .A(n40288), .B(n40287), .Z(n41693) );
  IV U53269 ( .A(n40289), .Z(n40290) );
  NOR U53270 ( .A(n40291), .B(n40290), .Z(n41689) );
  NOR U53271 ( .A(n41693), .B(n41689), .Z(n40292) );
  XOR U53272 ( .A(n41690), .B(n40292), .Z(n41686) );
  XOR U53273 ( .A(n41684), .B(n41686), .Z(n43756) );
  XOR U53274 ( .A(n40293), .B(n43756), .Z(n43759) );
  IV U53275 ( .A(n40294), .Z(n40296) );
  NOR U53276 ( .A(n40296), .B(n40295), .Z(n43758) );
  IV U53277 ( .A(n40297), .Z(n40298) );
  NOR U53278 ( .A(n40298), .B(n40303), .Z(n43762) );
  NOR U53279 ( .A(n43758), .B(n43762), .Z(n40299) );
  XOR U53280 ( .A(n43759), .B(n40299), .Z(n41683) );
  IV U53281 ( .A(n40300), .Z(n40309) );
  IV U53282 ( .A(n40310), .Z(n40301) );
  NOR U53283 ( .A(n40309), .B(n40301), .Z(n41679) );
  IV U53284 ( .A(n40302), .Z(n40304) );
  NOR U53285 ( .A(n40304), .B(n40303), .Z(n41681) );
  NOR U53286 ( .A(n41679), .B(n41681), .Z(n40305) );
  XOR U53287 ( .A(n41683), .B(n40305), .Z(n41674) );
  IV U53288 ( .A(n40306), .Z(n40307) );
  NOR U53289 ( .A(n40309), .B(n40307), .Z(n41676) );
  IV U53290 ( .A(n40308), .Z(n40312) );
  XOR U53291 ( .A(n40310), .B(n40309), .Z(n40311) );
  NOR U53292 ( .A(n40312), .B(n40311), .Z(n41673) );
  NOR U53293 ( .A(n41676), .B(n41673), .Z(n40313) );
  XOR U53294 ( .A(n41674), .B(n40313), .Z(n41669) );
  IV U53295 ( .A(n40314), .Z(n40315) );
  NOR U53296 ( .A(n40316), .B(n40315), .Z(n41667) );
  XOR U53297 ( .A(n41669), .B(n41667), .Z(n40323) );
  NOR U53298 ( .A(n40324), .B(n40323), .Z(n40317) );
  IV U53299 ( .A(n40317), .Z(n41670) );
  NOR U53300 ( .A(n40328), .B(n41670), .Z(n44899) );
  IV U53301 ( .A(n40318), .Z(n40319) );
  NOR U53302 ( .A(n40320), .B(n40319), .Z(n40325) );
  IV U53303 ( .A(n40325), .Z(n41666) );
  IV U53304 ( .A(n40321), .Z(n41671) );
  NOR U53305 ( .A(n40324), .B(n41671), .Z(n40322) );
  XOR U53306 ( .A(n40323), .B(n40322), .Z(n41665) );
  XOR U53307 ( .A(n41666), .B(n41665), .Z(n40330) );
  NOR U53308 ( .A(n40325), .B(n40324), .Z(n40326) );
  IV U53309 ( .A(n40326), .Z(n40327) );
  NOR U53310 ( .A(n40328), .B(n40327), .Z(n40329) );
  NOR U53311 ( .A(n40330), .B(n40329), .Z(n40331) );
  NOR U53312 ( .A(n44899), .B(n40331), .Z(n40332) );
  IV U53313 ( .A(n40332), .Z(n41663) );
  XOR U53314 ( .A(n40333), .B(n41663), .Z(n41651) );
  XOR U53315 ( .A(n40334), .B(n41651), .Z(n41647) );
  IV U53316 ( .A(n40335), .Z(n40336) );
  NOR U53317 ( .A(n40337), .B(n40336), .Z(n41643) );
  NOR U53318 ( .A(n41645), .B(n41643), .Z(n40338) );
  XOR U53319 ( .A(n41647), .B(n40338), .Z(n41636) );
  IV U53320 ( .A(n40339), .Z(n40341) );
  NOR U53321 ( .A(n40341), .B(n40340), .Z(n41635) );
  IV U53322 ( .A(n40342), .Z(n40343) );
  NOR U53323 ( .A(n40343), .B(n40347), .Z(n41638) );
  NOR U53324 ( .A(n41635), .B(n41638), .Z(n40344) );
  XOR U53325 ( .A(n41636), .B(n40344), .Z(n41634) );
  IV U53326 ( .A(n40345), .Z(n40346) );
  NOR U53327 ( .A(n40347), .B(n40346), .Z(n41632) );
  XOR U53328 ( .A(n41634), .B(n41632), .Z(n40348) );
  NOR U53329 ( .A(n40349), .B(n40348), .Z(n44880) );
  NOR U53330 ( .A(n40351), .B(n40350), .Z(n40352) );
  IV U53331 ( .A(n40352), .Z(n41628) );
  NOR U53332 ( .A(n40353), .B(n41628), .Z(n40354) );
  NOR U53333 ( .A(n41632), .B(n40354), .Z(n40355) );
  XOR U53334 ( .A(n41634), .B(n40355), .Z(n40356) );
  NOR U53335 ( .A(n40357), .B(n40356), .Z(n40358) );
  NOR U53336 ( .A(n44880), .B(n40358), .Z(n40359) );
  IV U53337 ( .A(n40359), .Z(n43772) );
  XOR U53338 ( .A(n43771), .B(n43772), .Z(n41625) );
  XOR U53339 ( .A(n40360), .B(n41625), .Z(n41620) );
  XOR U53340 ( .A(n41619), .B(n41620), .Z(n41617) );
  IV U53341 ( .A(n40361), .Z(n40363) );
  NOR U53342 ( .A(n40363), .B(n40362), .Z(n41616) );
  IV U53343 ( .A(n40364), .Z(n40366) );
  NOR U53344 ( .A(n40366), .B(n40365), .Z(n41614) );
  NOR U53345 ( .A(n41616), .B(n41614), .Z(n40367) );
  XOR U53346 ( .A(n41617), .B(n40367), .Z(n40375) );
  IV U53347 ( .A(n40375), .Z(n40368) );
  NOR U53348 ( .A(n40369), .B(n40368), .Z(n47056) );
  IV U53349 ( .A(n40370), .Z(n40372) );
  NOR U53350 ( .A(n40372), .B(n40371), .Z(n40376) );
  IV U53351 ( .A(n40376), .Z(n40374) );
  XOR U53352 ( .A(n41616), .B(n41617), .Z(n40373) );
  NOR U53353 ( .A(n40374), .B(n40373), .Z(n47053) );
  NOR U53354 ( .A(n40376), .B(n40375), .Z(n40377) );
  NOR U53355 ( .A(n47053), .B(n40377), .Z(n40378) );
  NOR U53356 ( .A(n40379), .B(n40378), .Z(n40380) );
  NOR U53357 ( .A(n47056), .B(n40380), .Z(n43776) );
  XOR U53358 ( .A(n43778), .B(n43776), .Z(n43782) );
  IV U53359 ( .A(n40381), .Z(n40383) );
  NOR U53360 ( .A(n40383), .B(n40382), .Z(n43779) );
  IV U53361 ( .A(n40384), .Z(n40385) );
  NOR U53362 ( .A(n40386), .B(n40385), .Z(n43781) );
  NOR U53363 ( .A(n43779), .B(n43781), .Z(n40387) );
  XOR U53364 ( .A(n43782), .B(n40387), .Z(n41610) );
  XOR U53365 ( .A(n40388), .B(n41610), .Z(n41608) );
  XOR U53366 ( .A(n40389), .B(n41608), .Z(n41599) );
  XOR U53367 ( .A(n40390), .B(n41599), .Z(n41597) );
  XOR U53368 ( .A(n40391), .B(n41597), .Z(n41583) );
  IV U53369 ( .A(n40392), .Z(n40394) );
  NOR U53370 ( .A(n40394), .B(n40393), .Z(n41585) );
  IV U53371 ( .A(n40395), .Z(n40396) );
  NOR U53372 ( .A(n40397), .B(n40396), .Z(n41582) );
  NOR U53373 ( .A(n41585), .B(n41582), .Z(n40398) );
  XOR U53374 ( .A(n41583), .B(n40398), .Z(n41581) );
  XOR U53375 ( .A(n40399), .B(n41581), .Z(n41569) );
  XOR U53376 ( .A(n40400), .B(n41569), .Z(n44862) );
  XOR U53377 ( .A(n43795), .B(n44862), .Z(n43802) );
  IV U53378 ( .A(n40401), .Z(n40402) );
  NOR U53379 ( .A(n40403), .B(n40402), .Z(n43806) );
  NOR U53380 ( .A(n40404), .B(n43803), .Z(n40405) );
  NOR U53381 ( .A(n43806), .B(n40405), .Z(n40406) );
  XOR U53382 ( .A(n43802), .B(n40406), .Z(n43816) );
  IV U53383 ( .A(n40407), .Z(n40409) );
  NOR U53384 ( .A(n40409), .B(n40408), .Z(n41566) );
  XOR U53385 ( .A(n43816), .B(n41566), .Z(n40410) );
  XOR U53386 ( .A(n40411), .B(n40410), .Z(n43813) );
  XOR U53387 ( .A(n47127), .B(n43813), .Z(n43820) );
  XOR U53388 ( .A(n40412), .B(n43820), .Z(n41550) );
  XOR U53389 ( .A(n40413), .B(n41550), .Z(n40420) );
  IV U53390 ( .A(n40420), .Z(n40414) );
  NOR U53391 ( .A(n40415), .B(n40414), .Z(n48239) );
  IV U53392 ( .A(n40416), .Z(n40418) );
  NOR U53393 ( .A(n40418), .B(n40417), .Z(n40421) );
  IV U53394 ( .A(n40421), .Z(n40419) );
  NOR U53395 ( .A(n41550), .B(n40419), .Z(n47137) );
  NOR U53396 ( .A(n40421), .B(n40420), .Z(n40422) );
  NOR U53397 ( .A(n47137), .B(n40422), .Z(n41541) );
  NOR U53398 ( .A(n40423), .B(n41541), .Z(n40424) );
  NOR U53399 ( .A(n48239), .B(n40424), .Z(n43827) );
  XOR U53400 ( .A(n40425), .B(n43827), .Z(n43832) );
  XOR U53401 ( .A(n40426), .B(n43832), .Z(n43836) );
  XOR U53402 ( .A(n40427), .B(n43836), .Z(n43844) );
  IV U53403 ( .A(n43844), .Z(n40434) );
  NOR U53404 ( .A(n40429), .B(n40428), .Z(n41536) );
  IV U53405 ( .A(n40430), .Z(n40432) );
  IV U53406 ( .A(n40431), .Z(n40436) );
  NOR U53407 ( .A(n40432), .B(n40436), .Z(n43842) );
  NOR U53408 ( .A(n41536), .B(n43842), .Z(n40433) );
  XOR U53409 ( .A(n40434), .B(n40433), .Z(n43847) );
  IV U53410 ( .A(n40435), .Z(n40437) );
  NOR U53411 ( .A(n40437), .B(n40436), .Z(n43845) );
  XOR U53412 ( .A(n43847), .B(n43845), .Z(n43852) );
  XOR U53413 ( .A(n40438), .B(n43852), .Z(n43855) );
  XOR U53414 ( .A(n43854), .B(n43855), .Z(n43860) );
  IV U53415 ( .A(n40439), .Z(n40441) );
  NOR U53416 ( .A(n40441), .B(n40440), .Z(n43858) );
  XOR U53417 ( .A(n43860), .B(n43858), .Z(n43863) );
  IV U53418 ( .A(n40442), .Z(n40447) );
  IV U53419 ( .A(n40443), .Z(n40444) );
  NOR U53420 ( .A(n40447), .B(n40444), .Z(n43861) );
  XOR U53421 ( .A(n43863), .B(n43861), .Z(n43867) );
  IV U53422 ( .A(n40445), .Z(n40446) );
  NOR U53423 ( .A(n40447), .B(n40446), .Z(n43865) );
  XOR U53424 ( .A(n43867), .B(n43865), .Z(n43872) );
  IV U53425 ( .A(n40448), .Z(n40450) );
  NOR U53426 ( .A(n40450), .B(n40449), .Z(n43868) );
  IV U53427 ( .A(n40451), .Z(n40453) );
  NOR U53428 ( .A(n40453), .B(n40452), .Z(n43871) );
  NOR U53429 ( .A(n43868), .B(n43871), .Z(n40454) );
  XOR U53430 ( .A(n43872), .B(n40454), .Z(n43874) );
  IV U53431 ( .A(n40457), .Z(n40455) );
  NOR U53432 ( .A(n40456), .B(n40455), .Z(n43875) );
  XOR U53433 ( .A(n40457), .B(n40456), .Z(n40460) );
  IV U53434 ( .A(n40458), .Z(n40459) );
  NOR U53435 ( .A(n40460), .B(n40459), .Z(n43877) );
  NOR U53436 ( .A(n43875), .B(n43877), .Z(n40461) );
  XOR U53437 ( .A(n43874), .B(n40461), .Z(n43881) );
  XOR U53438 ( .A(n43882), .B(n43881), .Z(n41527) );
  IV U53439 ( .A(n40462), .Z(n41531) );
  NOR U53440 ( .A(n40463), .B(n41531), .Z(n40467) );
  IV U53441 ( .A(n40464), .Z(n40465) );
  NOR U53442 ( .A(n40466), .B(n40465), .Z(n41526) );
  NOR U53443 ( .A(n40467), .B(n41526), .Z(n40468) );
  XOR U53444 ( .A(n41527), .B(n40468), .Z(n41523) );
  IV U53445 ( .A(n40469), .Z(n40470) );
  NOR U53446 ( .A(n40471), .B(n40470), .Z(n41521) );
  XOR U53447 ( .A(n41523), .B(n41521), .Z(n43890) );
  XOR U53448 ( .A(n40472), .B(n43890), .Z(n41518) );
  XOR U53449 ( .A(n40473), .B(n41518), .Z(n41513) );
  XOR U53450 ( .A(n40474), .B(n41513), .Z(n43896) );
  XOR U53451 ( .A(n40475), .B(n43896), .Z(n43901) );
  XOR U53452 ( .A(n40476), .B(n43901), .Z(n41501) );
  XOR U53453 ( .A(n40477), .B(n41501), .Z(n41496) );
  IV U53454 ( .A(n41496), .Z(n40483) );
  NOR U53455 ( .A(n40478), .B(n41497), .Z(n40481) );
  IV U53456 ( .A(n40479), .Z(n40480) );
  NOR U53457 ( .A(n40480), .B(n41488), .Z(n41493) );
  NOR U53458 ( .A(n40481), .B(n41493), .Z(n40482) );
  XOR U53459 ( .A(n40483), .B(n40482), .Z(n43911) );
  IV U53460 ( .A(n40484), .Z(n40485) );
  NOR U53461 ( .A(n40489), .B(n40485), .Z(n40493) );
  IV U53462 ( .A(n40493), .Z(n40486) );
  NOR U53463 ( .A(n43911), .B(n40486), .Z(n47204) );
  NOR U53464 ( .A(n40487), .B(n43910), .Z(n40491) );
  IV U53465 ( .A(n40488), .Z(n40490) );
  NOR U53466 ( .A(n40490), .B(n40489), .Z(n43907) );
  NOR U53467 ( .A(n40491), .B(n43907), .Z(n40492) );
  XOR U53468 ( .A(n43911), .B(n40492), .Z(n40497) );
  NOR U53469 ( .A(n40493), .B(n40497), .Z(n40494) );
  NOR U53470 ( .A(n47204), .B(n40494), .Z(n40495) );
  NOR U53471 ( .A(n40496), .B(n40495), .Z(n40500) );
  IV U53472 ( .A(n40496), .Z(n40499) );
  IV U53473 ( .A(n40497), .Z(n40498) );
  NOR U53474 ( .A(n40499), .B(n40498), .Z(n47200) );
  NOR U53475 ( .A(n40500), .B(n47200), .Z(n41481) );
  XOR U53476 ( .A(n40501), .B(n41481), .Z(n41480) );
  XOR U53477 ( .A(n41478), .B(n41480), .Z(n41474) );
  XOR U53478 ( .A(n41473), .B(n41474), .Z(n41476) );
  XOR U53479 ( .A(n41477), .B(n41476), .Z(n41463) );
  IV U53480 ( .A(n40502), .Z(n40510) );
  NOR U53481 ( .A(n40503), .B(n40510), .Z(n40504) );
  IV U53482 ( .A(n40504), .Z(n40505) );
  NOR U53483 ( .A(n40506), .B(n40505), .Z(n40507) );
  IV U53484 ( .A(n40507), .Z(n41467) );
  NOR U53485 ( .A(n40508), .B(n41467), .Z(n40512) );
  IV U53486 ( .A(n40509), .Z(n40511) );
  NOR U53487 ( .A(n40511), .B(n40510), .Z(n41464) );
  NOR U53488 ( .A(n40512), .B(n41464), .Z(n40513) );
  XOR U53489 ( .A(n41463), .B(n40513), .Z(n41459) );
  IV U53490 ( .A(n40514), .Z(n40519) );
  IV U53491 ( .A(n40515), .Z(n40516) );
  NOR U53492 ( .A(n40517), .B(n40516), .Z(n40518) );
  IV U53493 ( .A(n40518), .Z(n40524) );
  NOR U53494 ( .A(n40519), .B(n40524), .Z(n41457) );
  XOR U53495 ( .A(n41459), .B(n41457), .Z(n41462) );
  IV U53496 ( .A(n40520), .Z(n40521) );
  NOR U53497 ( .A(n40522), .B(n40521), .Z(n41455) );
  IV U53498 ( .A(n40523), .Z(n40525) );
  NOR U53499 ( .A(n40525), .B(n40524), .Z(n41460) );
  NOR U53500 ( .A(n41455), .B(n41460), .Z(n40526) );
  XOR U53501 ( .A(n41462), .B(n40526), .Z(n41449) );
  XOR U53502 ( .A(n41450), .B(n41449), .Z(n41452) );
  IV U53503 ( .A(n40527), .Z(n40529) );
  NOR U53504 ( .A(n40529), .B(n40528), .Z(n41447) );
  NOR U53505 ( .A(n41451), .B(n41447), .Z(n40530) );
  XOR U53506 ( .A(n41452), .B(n40530), .Z(n41443) );
  XOR U53507 ( .A(n40531), .B(n41443), .Z(n43932) );
  IV U53508 ( .A(n40532), .Z(n40534) );
  NOR U53509 ( .A(n40534), .B(n40533), .Z(n43930) );
  XOR U53510 ( .A(n43932), .B(n43930), .Z(n43935) );
  IV U53511 ( .A(n40535), .Z(n41439) );
  NOR U53512 ( .A(n41439), .B(n40536), .Z(n43934) );
  NOR U53513 ( .A(n41442), .B(n40537), .Z(n40538) );
  NOR U53514 ( .A(n43934), .B(n40538), .Z(n40539) );
  XOR U53515 ( .A(n43935), .B(n40539), .Z(n41435) );
  IV U53516 ( .A(n40540), .Z(n40541) );
  NOR U53517 ( .A(n40545), .B(n40541), .Z(n41436) );
  IV U53518 ( .A(n40542), .Z(n44736) );
  NOR U53519 ( .A(n40543), .B(n44736), .Z(n40547) );
  IV U53520 ( .A(n40544), .Z(n40546) );
  NOR U53521 ( .A(n40546), .B(n40545), .Z(n47277) );
  NOR U53522 ( .A(n40547), .B(n47277), .Z(n41438) );
  IV U53523 ( .A(n41438), .Z(n40548) );
  NOR U53524 ( .A(n41436), .B(n40548), .Z(n40549) );
  XOR U53525 ( .A(n41435), .B(n40549), .Z(n41431) );
  IV U53526 ( .A(n40550), .Z(n40552) );
  NOR U53527 ( .A(n40552), .B(n40551), .Z(n40553) );
  IV U53528 ( .A(n40553), .Z(n41430) );
  XOR U53529 ( .A(n41431), .B(n41430), .Z(n41433) );
  IV U53530 ( .A(n40554), .Z(n40555) );
  NOR U53531 ( .A(n40556), .B(n40555), .Z(n41432) );
  IV U53532 ( .A(n40557), .Z(n40558) );
  NOR U53533 ( .A(n40559), .B(n40558), .Z(n43941) );
  NOR U53534 ( .A(n41432), .B(n43941), .Z(n40560) );
  XOR U53535 ( .A(n41433), .B(n40560), .Z(n43940) );
  XOR U53536 ( .A(n43938), .B(n43940), .Z(n41426) );
  XOR U53537 ( .A(n40561), .B(n41426), .Z(n41409) );
  XOR U53538 ( .A(n40562), .B(n41409), .Z(n41407) );
  XOR U53539 ( .A(n40563), .B(n41407), .Z(n43949) );
  XOR U53540 ( .A(n43947), .B(n43949), .Z(n43950) );
  XOR U53541 ( .A(n43951), .B(n43950), .Z(n41401) );
  IV U53542 ( .A(n40564), .Z(n40565) );
  NOR U53543 ( .A(n40566), .B(n40565), .Z(n43945) );
  NOR U53544 ( .A(n40567), .B(n41403), .Z(n40568) );
  NOR U53545 ( .A(n43945), .B(n40568), .Z(n40569) );
  XOR U53546 ( .A(n41401), .B(n40569), .Z(n41399) );
  IV U53547 ( .A(n40570), .Z(n40578) );
  IV U53548 ( .A(n40571), .Z(n40572) );
  NOR U53549 ( .A(n40578), .B(n40572), .Z(n41395) );
  IV U53550 ( .A(n40579), .Z(n40573) );
  NOR U53551 ( .A(n40573), .B(n40578), .Z(n41397) );
  NOR U53552 ( .A(n41395), .B(n41397), .Z(n40574) );
  XOR U53553 ( .A(n41399), .B(n40574), .Z(n41388) );
  NOR U53554 ( .A(n40576), .B(n40575), .Z(n41392) );
  IV U53555 ( .A(n40577), .Z(n40583) );
  XOR U53556 ( .A(n40579), .B(n40578), .Z(n40580) );
  NOR U53557 ( .A(n40581), .B(n40580), .Z(n40582) );
  IV U53558 ( .A(n40582), .Z(n40590) );
  NOR U53559 ( .A(n40583), .B(n40590), .Z(n41390) );
  NOR U53560 ( .A(n41392), .B(n41390), .Z(n40584) );
  XOR U53561 ( .A(n41388), .B(n40584), .Z(n41386) );
  IV U53562 ( .A(n40585), .Z(n40588) );
  IV U53563 ( .A(n40586), .Z(n40587) );
  NOR U53564 ( .A(n40588), .B(n40587), .Z(n41384) );
  IV U53565 ( .A(n40589), .Z(n40591) );
  NOR U53566 ( .A(n40591), .B(n40590), .Z(n41387) );
  NOR U53567 ( .A(n41384), .B(n41387), .Z(n40592) );
  XOR U53568 ( .A(n41386), .B(n40592), .Z(n41382) );
  IV U53569 ( .A(n40593), .Z(n40594) );
  NOR U53570 ( .A(n40595), .B(n40594), .Z(n41381) );
  IV U53571 ( .A(n40596), .Z(n40598) );
  NOR U53572 ( .A(n40598), .B(n40597), .Z(n43958) );
  NOR U53573 ( .A(n41381), .B(n43958), .Z(n40599) );
  XOR U53574 ( .A(n41382), .B(n40599), .Z(n43963) );
  XOR U53575 ( .A(n41378), .B(n43963), .Z(n41375) );
  XOR U53576 ( .A(n40600), .B(n41375), .Z(n43969) );
  XOR U53577 ( .A(n40601), .B(n43969), .Z(n43981) );
  XOR U53578 ( .A(n40602), .B(n43981), .Z(n43979) );
  XOR U53579 ( .A(n43977), .B(n43979), .Z(n41369) );
  XOR U53580 ( .A(n41368), .B(n41369), .Z(n41372) );
  IV U53581 ( .A(n40603), .Z(n40604) );
  NOR U53582 ( .A(n40605), .B(n40604), .Z(n41371) );
  IV U53583 ( .A(n40606), .Z(n40608) );
  NOR U53584 ( .A(n40608), .B(n40607), .Z(n41363) );
  NOR U53585 ( .A(n41371), .B(n41363), .Z(n40609) );
  XOR U53586 ( .A(n41372), .B(n40609), .Z(n41361) );
  XOR U53587 ( .A(n40610), .B(n41361), .Z(n43989) );
  XOR U53588 ( .A(n43987), .B(n43989), .Z(n43995) );
  IV U53589 ( .A(n40611), .Z(n41359) );
  NOR U53590 ( .A(n41354), .B(n41359), .Z(n40615) );
  IV U53591 ( .A(n40612), .Z(n40614) );
  NOR U53592 ( .A(n40614), .B(n40613), .Z(n43994) );
  NOR U53593 ( .A(n40615), .B(n43994), .Z(n40616) );
  XOR U53594 ( .A(n43995), .B(n40616), .Z(n41348) );
  IV U53595 ( .A(n40617), .Z(n40619) );
  NOR U53596 ( .A(n40619), .B(n40618), .Z(n41351) );
  IV U53597 ( .A(n40620), .Z(n40621) );
  NOR U53598 ( .A(n40622), .B(n40621), .Z(n41349) );
  NOR U53599 ( .A(n41351), .B(n41349), .Z(n40623) );
  XOR U53600 ( .A(n41348), .B(n40623), .Z(n44677) );
  NOR U53601 ( .A(n40625), .B(n40624), .Z(n47354) );
  IV U53602 ( .A(n40626), .Z(n40628) );
  NOR U53603 ( .A(n40628), .B(n40627), .Z(n44676) );
  NOR U53604 ( .A(n47354), .B(n44676), .Z(n41342) );
  XOR U53605 ( .A(n44677), .B(n41342), .Z(n40629) );
  IV U53606 ( .A(n40629), .Z(n41344) );
  XOR U53607 ( .A(n41343), .B(n41344), .Z(n44000) );
  XOR U53608 ( .A(n40630), .B(n44000), .Z(n41337) );
  XOR U53609 ( .A(n40631), .B(n41337), .Z(n44025) );
  XOR U53610 ( .A(n44024), .B(n44025), .Z(n44028) );
  XOR U53611 ( .A(n44027), .B(n44028), .Z(n41332) );
  XOR U53612 ( .A(n41331), .B(n41332), .Z(n41336) );
  XOR U53613 ( .A(n41334), .B(n41336), .Z(n44031) );
  XOR U53614 ( .A(n40632), .B(n44031), .Z(n40633) );
  IV U53615 ( .A(n40633), .Z(n44035) );
  IV U53616 ( .A(n40634), .Z(n40636) );
  NOR U53617 ( .A(n40636), .B(n40635), .Z(n44033) );
  XOR U53618 ( .A(n44035), .B(n44033), .Z(n44044) );
  XOR U53619 ( .A(n44043), .B(n44044), .Z(n44039) );
  IV U53620 ( .A(n40637), .Z(n40638) );
  NOR U53621 ( .A(n40639), .B(n40638), .Z(n44037) );
  XOR U53622 ( .A(n44039), .B(n44037), .Z(n44041) );
  XOR U53623 ( .A(n44042), .B(n44041), .Z(n40649) );
  IV U53624 ( .A(n40640), .Z(n40642) );
  NOR U53625 ( .A(n40642), .B(n40641), .Z(n40652) );
  IV U53626 ( .A(n40643), .Z(n40645) );
  NOR U53627 ( .A(n40645), .B(n40644), .Z(n40648) );
  NOR U53628 ( .A(n40652), .B(n40648), .Z(n40646) );
  IV U53629 ( .A(n40646), .Z(n40647) );
  NOR U53630 ( .A(n40649), .B(n40647), .Z(n40655) );
  IV U53631 ( .A(n40648), .Z(n40651) );
  IV U53632 ( .A(n40649), .Z(n40650) );
  NOR U53633 ( .A(n40651), .B(n40650), .Z(n47386) );
  IV U53634 ( .A(n40652), .Z(n40653) );
  NOR U53635 ( .A(n40653), .B(n44041), .Z(n44652) );
  NOR U53636 ( .A(n47386), .B(n44652), .Z(n40654) );
  IV U53637 ( .A(n40654), .Z(n44055) );
  NOR U53638 ( .A(n40655), .B(n44055), .Z(n40656) );
  IV U53639 ( .A(n40656), .Z(n51650) );
  NOR U53640 ( .A(n40657), .B(n51650), .Z(n41317) );
  IV U53641 ( .A(n40658), .Z(n40659) );
  NOR U53642 ( .A(n40659), .B(n51655), .Z(n44053) );
  IV U53643 ( .A(n40660), .Z(n40662) );
  NOR U53644 ( .A(n40662), .B(n40661), .Z(n41318) );
  NOR U53645 ( .A(n44053), .B(n41318), .Z(n40663) );
  XOR U53646 ( .A(n40663), .B(n51650), .Z(n44059) );
  NOR U53647 ( .A(n40664), .B(n44059), .Z(n40665) );
  NOR U53648 ( .A(n41317), .B(n40665), .Z(n44063) );
  IV U53649 ( .A(n40666), .Z(n40668) );
  NOR U53650 ( .A(n40668), .B(n40667), .Z(n44058) );
  NOR U53651 ( .A(n44058), .B(n44062), .Z(n40669) );
  XOR U53652 ( .A(n44063), .B(n40669), .Z(n41315) );
  IV U53653 ( .A(n40670), .Z(n40671) );
  NOR U53654 ( .A(n40671), .B(n40674), .Z(n40672) );
  IV U53655 ( .A(n40672), .Z(n40681) );
  NOR U53656 ( .A(n41315), .B(n40681), .Z(n50838) );
  IV U53657 ( .A(n40673), .Z(n40675) );
  NOR U53658 ( .A(n40675), .B(n40674), .Z(n41307) );
  IV U53659 ( .A(n40676), .Z(n40679) );
  IV U53660 ( .A(n40677), .Z(n40678) );
  NOR U53661 ( .A(n40679), .B(n40678), .Z(n40680) );
  IV U53662 ( .A(n40680), .Z(n41314) );
  XOR U53663 ( .A(n41314), .B(n41315), .Z(n41308) );
  XOR U53664 ( .A(n41307), .B(n41308), .Z(n40683) );
  NOR U53665 ( .A(n41308), .B(n40681), .Z(n40682) );
  NOR U53666 ( .A(n40683), .B(n40682), .Z(n40684) );
  NOR U53667 ( .A(n50838), .B(n40684), .Z(n40685) );
  IV U53668 ( .A(n40685), .Z(n41312) );
  XOR U53669 ( .A(n41312), .B(n41311), .Z(n41301) );
  IV U53670 ( .A(n40686), .Z(n40688) );
  IV U53671 ( .A(n40687), .Z(n40700) );
  NOR U53672 ( .A(n40688), .B(n40700), .Z(n40689) );
  IV U53673 ( .A(n40689), .Z(n40695) );
  NOR U53674 ( .A(n41301), .B(n40695), .Z(n41300) );
  IV U53675 ( .A(n40690), .Z(n40693) );
  IV U53676 ( .A(n40691), .Z(n40692) );
  NOR U53677 ( .A(n40693), .B(n40692), .Z(n41303) );
  IV U53678 ( .A(n40694), .Z(n41302) );
  XOR U53679 ( .A(n41302), .B(n41301), .Z(n41304) );
  XOR U53680 ( .A(n41303), .B(n41304), .Z(n40697) );
  NOR U53681 ( .A(n41304), .B(n40695), .Z(n40696) );
  NOR U53682 ( .A(n40697), .B(n40696), .Z(n40698) );
  NOR U53683 ( .A(n41300), .B(n40698), .Z(n44066) );
  IV U53684 ( .A(n40699), .Z(n40701) );
  NOR U53685 ( .A(n40701), .B(n40700), .Z(n40702) );
  IV U53686 ( .A(n40702), .Z(n44067) );
  XOR U53687 ( .A(n44066), .B(n44067), .Z(n44070) );
  XOR U53688 ( .A(n44069), .B(n44070), .Z(n41296) );
  IV U53689 ( .A(n40703), .Z(n40704) );
  NOR U53690 ( .A(n40705), .B(n40704), .Z(n41295) );
  IV U53691 ( .A(n40706), .Z(n40708) );
  NOR U53692 ( .A(n40708), .B(n40707), .Z(n41298) );
  NOR U53693 ( .A(n41295), .B(n41298), .Z(n40709) );
  XOR U53694 ( .A(n41296), .B(n40709), .Z(n41289) );
  XOR U53695 ( .A(n40710), .B(n41289), .Z(n41287) );
  XOR U53696 ( .A(n40711), .B(n41287), .Z(n41283) );
  XOR U53697 ( .A(n40712), .B(n41283), .Z(n41280) );
  XOR U53698 ( .A(n41278), .B(n41280), .Z(n40731) );
  IV U53699 ( .A(n40731), .Z(n40713) );
  NOR U53700 ( .A(n40714), .B(n40713), .Z(n40724) );
  IV U53701 ( .A(n40715), .Z(n40718) );
  NOR U53702 ( .A(n40716), .B(n41280), .Z(n40717) );
  IV U53703 ( .A(n40717), .Z(n40720) );
  NOR U53704 ( .A(n40718), .B(n40720), .Z(n47434) );
  IV U53705 ( .A(n40719), .Z(n40721) );
  NOR U53706 ( .A(n40721), .B(n40720), .Z(n44626) );
  NOR U53707 ( .A(n47434), .B(n44626), .Z(n40722) );
  IV U53708 ( .A(n40722), .Z(n40723) );
  NOR U53709 ( .A(n40724), .B(n40723), .Z(n44077) );
  IV U53710 ( .A(n40725), .Z(n40726) );
  NOR U53711 ( .A(n40727), .B(n40726), .Z(n40737) );
  IV U53712 ( .A(n40737), .Z(n44079) );
  NOR U53713 ( .A(n44077), .B(n44079), .Z(n40739) );
  IV U53714 ( .A(n40728), .Z(n40730) );
  NOR U53715 ( .A(n40730), .B(n40729), .Z(n40733) );
  IV U53716 ( .A(n40733), .Z(n40732) );
  NOR U53717 ( .A(n40732), .B(n40731), .Z(n41277) );
  NOR U53718 ( .A(n44077), .B(n40733), .Z(n40734) );
  NOR U53719 ( .A(n41277), .B(n40734), .Z(n40735) );
  IV U53720 ( .A(n40735), .Z(n40736) );
  NOR U53721 ( .A(n40737), .B(n40736), .Z(n40738) );
  NOR U53722 ( .A(n40739), .B(n40738), .Z(n44083) );
  IV U53723 ( .A(n40743), .Z(n40740) );
  NOR U53724 ( .A(n40740), .B(n40742), .Z(n44084) );
  IV U53725 ( .A(n40741), .Z(n40745) );
  XOR U53726 ( .A(n40743), .B(n40742), .Z(n40744) );
  NOR U53727 ( .A(n40745), .B(n40744), .Z(n41270) );
  NOR U53728 ( .A(n44084), .B(n41270), .Z(n40746) );
  XOR U53729 ( .A(n44083), .B(n40746), .Z(n41272) );
  XOR U53730 ( .A(n40747), .B(n41272), .Z(n44090) );
  XOR U53731 ( .A(n40748), .B(n44090), .Z(n44092) );
  XOR U53732 ( .A(n40749), .B(n44092), .Z(n41266) );
  XOR U53733 ( .A(n40750), .B(n41266), .Z(n40751) );
  IV U53734 ( .A(n40751), .Z(n41262) );
  XOR U53735 ( .A(n41261), .B(n41262), .Z(n40752) );
  NOR U53736 ( .A(n40753), .B(n40752), .Z(n47466) );
  IV U53737 ( .A(n40754), .Z(n40755) );
  NOR U53738 ( .A(n40756), .B(n40755), .Z(n41257) );
  NOR U53739 ( .A(n41261), .B(n41257), .Z(n40757) );
  XOR U53740 ( .A(n40757), .B(n41262), .Z(n41254) );
  NOR U53741 ( .A(n40758), .B(n41254), .Z(n40759) );
  NOR U53742 ( .A(n47466), .B(n40759), .Z(n44100) );
  IV U53743 ( .A(n40760), .Z(n40762) );
  NOR U53744 ( .A(n40762), .B(n40761), .Z(n41253) );
  IV U53745 ( .A(n40763), .Z(n40765) );
  NOR U53746 ( .A(n40765), .B(n40764), .Z(n44099) );
  NOR U53747 ( .A(n41253), .B(n44099), .Z(n40766) );
  XOR U53748 ( .A(n44100), .B(n40766), .Z(n44111) );
  IV U53749 ( .A(n40767), .Z(n40769) );
  NOR U53750 ( .A(n40769), .B(n40768), .Z(n44107) );
  IV U53751 ( .A(n40770), .Z(n40771) );
  NOR U53752 ( .A(n40772), .B(n40771), .Z(n44109) );
  NOR U53753 ( .A(n44107), .B(n44109), .Z(n40773) );
  XOR U53754 ( .A(n44111), .B(n40773), .Z(n44105) );
  IV U53755 ( .A(n40774), .Z(n40776) );
  NOR U53756 ( .A(n40776), .B(n40775), .Z(n44104) );
  IV U53757 ( .A(n40777), .Z(n40779) );
  NOR U53758 ( .A(n40779), .B(n40778), .Z(n44115) );
  NOR U53759 ( .A(n44104), .B(n44115), .Z(n40780) );
  XOR U53760 ( .A(n44105), .B(n40780), .Z(n44123) );
  IV U53761 ( .A(n44123), .Z(n40787) );
  IV U53762 ( .A(n40781), .Z(n40782) );
  NOR U53763 ( .A(n40783), .B(n40782), .Z(n41251) );
  NOR U53764 ( .A(n40785), .B(n40784), .Z(n44121) );
  NOR U53765 ( .A(n41251), .B(n44121), .Z(n40786) );
  XOR U53766 ( .A(n40787), .B(n40786), .Z(n41248) );
  XOR U53767 ( .A(n41247), .B(n41248), .Z(n44119) );
  XOR U53768 ( .A(n44118), .B(n44119), .Z(n44130) );
  IV U53769 ( .A(n40788), .Z(n40790) );
  NOR U53770 ( .A(n40790), .B(n40789), .Z(n44129) );
  NOR U53771 ( .A(n44129), .B(n40791), .Z(n40792) );
  XOR U53772 ( .A(n44130), .B(n40792), .Z(n44135) );
  IV U53773 ( .A(n41243), .Z(n40794) );
  IV U53774 ( .A(n40793), .Z(n41244) );
  NOR U53775 ( .A(n40794), .B(n41244), .Z(n47492) );
  IV U53776 ( .A(n40795), .Z(n40797) );
  IV U53777 ( .A(n40796), .Z(n40800) );
  NOR U53778 ( .A(n40797), .B(n40800), .Z(n44136) );
  NOR U53779 ( .A(n47492), .B(n44136), .Z(n40798) );
  XOR U53780 ( .A(n44135), .B(n40798), .Z(n44139) );
  IV U53781 ( .A(n40799), .Z(n40801) );
  NOR U53782 ( .A(n40801), .B(n40800), .Z(n41240) );
  XOR U53783 ( .A(n44139), .B(n41240), .Z(n41239) );
  IV U53784 ( .A(n40802), .Z(n40803) );
  NOR U53785 ( .A(n40806), .B(n40803), .Z(n44138) );
  IV U53786 ( .A(n40804), .Z(n40805) );
  NOR U53787 ( .A(n40806), .B(n40805), .Z(n41237) );
  NOR U53788 ( .A(n44138), .B(n41237), .Z(n40807) );
  XOR U53789 ( .A(n41239), .B(n40807), .Z(n44141) );
  IV U53790 ( .A(n40808), .Z(n40820) );
  IV U53791 ( .A(n40809), .Z(n40810) );
  NOR U53792 ( .A(n40820), .B(n40810), .Z(n44146) );
  IV U53793 ( .A(n40811), .Z(n40813) );
  NOR U53794 ( .A(n40813), .B(n40812), .Z(n44142) );
  NOR U53795 ( .A(n44146), .B(n44142), .Z(n40814) );
  XOR U53796 ( .A(n44141), .B(n40814), .Z(n47520) );
  IV U53797 ( .A(n40815), .Z(n40817) );
  NOR U53798 ( .A(n40817), .B(n40816), .Z(n47527) );
  IV U53799 ( .A(n40818), .Z(n40819) );
  NOR U53800 ( .A(n40820), .B(n40819), .Z(n47518) );
  NOR U53801 ( .A(n47527), .B(n47518), .Z(n44145) );
  XOR U53802 ( .A(n47520), .B(n44145), .Z(n40821) );
  IV U53803 ( .A(n40821), .Z(n41236) );
  XOR U53804 ( .A(n41234), .B(n41236), .Z(n44159) );
  XOR U53805 ( .A(n44157), .B(n44159), .Z(n40835) );
  XOR U53806 ( .A(n40836), .B(n40835), .Z(n40826) );
  IV U53807 ( .A(n40822), .Z(n40824) );
  IV U53808 ( .A(n40823), .Z(n40852) );
  NOR U53809 ( .A(n40824), .B(n40852), .Z(n40849) );
  IV U53810 ( .A(n40849), .Z(n40825) );
  NOR U53811 ( .A(n40826), .B(n40825), .Z(n47550) );
  IV U53812 ( .A(n40826), .Z(n40830) );
  NOR U53813 ( .A(n40828), .B(n40827), .Z(n40829) );
  NOR U53814 ( .A(n40830), .B(n40829), .Z(n40847) );
  IV U53815 ( .A(n40831), .Z(n40841) );
  IV U53816 ( .A(n40832), .Z(n40834) );
  NOR U53817 ( .A(n40834), .B(n40833), .Z(n40839) );
  NOR U53818 ( .A(n40836), .B(n40835), .Z(n40837) );
  IV U53819 ( .A(n40837), .Z(n40838) );
  NOR U53820 ( .A(n40839), .B(n40838), .Z(n40840) );
  IV U53821 ( .A(n40840), .Z(n40843) );
  NOR U53822 ( .A(n40841), .B(n40843), .Z(n47547) );
  IV U53823 ( .A(n40842), .Z(n40844) );
  NOR U53824 ( .A(n40844), .B(n40843), .Z(n47541) );
  NOR U53825 ( .A(n47547), .B(n47541), .Z(n40845) );
  IV U53826 ( .A(n40845), .Z(n40846) );
  NOR U53827 ( .A(n40847), .B(n40846), .Z(n40848) );
  NOR U53828 ( .A(n40849), .B(n40848), .Z(n40850) );
  NOR U53829 ( .A(n47550), .B(n40850), .Z(n41231) );
  IV U53830 ( .A(n40851), .Z(n40853) );
  NOR U53831 ( .A(n40853), .B(n40852), .Z(n40854) );
  IV U53832 ( .A(n40854), .Z(n41233) );
  XOR U53833 ( .A(n41231), .B(n41233), .Z(n41227) );
  XOR U53834 ( .A(n40855), .B(n41227), .Z(n40856) );
  IV U53835 ( .A(n40856), .Z(n41219) );
  IV U53836 ( .A(n40857), .Z(n40859) );
  NOR U53837 ( .A(n40859), .B(n40858), .Z(n41220) );
  IV U53838 ( .A(n40860), .Z(n40861) );
  NOR U53839 ( .A(n40861), .B(n40867), .Z(n41217) );
  NOR U53840 ( .A(n41220), .B(n41217), .Z(n40862) );
  XOR U53841 ( .A(n41219), .B(n40862), .Z(n41211) );
  IV U53842 ( .A(n40863), .Z(n40864) );
  NOR U53843 ( .A(n40865), .B(n40864), .Z(n41212) );
  IV U53844 ( .A(n40866), .Z(n40868) );
  NOR U53845 ( .A(n40868), .B(n40867), .Z(n41214) );
  NOR U53846 ( .A(n41212), .B(n41214), .Z(n40869) );
  XOR U53847 ( .A(n41211), .B(n40869), .Z(n41209) );
  XOR U53848 ( .A(n41208), .B(n41209), .Z(n44176) );
  IV U53849 ( .A(n40870), .Z(n40876) );
  NOR U53850 ( .A(n40871), .B(n40882), .Z(n40872) );
  IV U53851 ( .A(n40872), .Z(n40878) );
  NOR U53852 ( .A(n40873), .B(n40878), .Z(n40874) );
  IV U53853 ( .A(n40874), .Z(n40875) );
  NOR U53854 ( .A(n40876), .B(n40875), .Z(n44174) );
  XOR U53855 ( .A(n44176), .B(n44174), .Z(n44178) );
  IV U53856 ( .A(n40877), .Z(n40879) );
  NOR U53857 ( .A(n40879), .B(n40878), .Z(n40880) );
  IV U53858 ( .A(n40880), .Z(n44177) );
  XOR U53859 ( .A(n44178), .B(n44177), .Z(n44182) );
  IV U53860 ( .A(n40881), .Z(n40883) );
  NOR U53861 ( .A(n40883), .B(n40882), .Z(n44184) );
  IV U53862 ( .A(n40884), .Z(n40885) );
  NOR U53863 ( .A(n40888), .B(n40885), .Z(n44181) );
  IV U53864 ( .A(n40886), .Z(n40887) );
  NOR U53865 ( .A(n40888), .B(n40887), .Z(n44190) );
  NOR U53866 ( .A(n44181), .B(n44190), .Z(n40889) );
  IV U53867 ( .A(n40889), .Z(n40890) );
  NOR U53868 ( .A(n44184), .B(n40890), .Z(n40891) );
  XOR U53869 ( .A(n44182), .B(n40891), .Z(n44197) );
  IV U53870 ( .A(n40892), .Z(n40894) );
  NOR U53871 ( .A(n40894), .B(n40893), .Z(n44195) );
  XOR U53872 ( .A(n44197), .B(n44195), .Z(n40895) );
  NOR U53873 ( .A(n40896), .B(n40895), .Z(n44576) );
  IV U53874 ( .A(n40897), .Z(n40899) );
  NOR U53875 ( .A(n40899), .B(n40898), .Z(n44193) );
  NOR U53876 ( .A(n44193), .B(n44195), .Z(n40900) );
  XOR U53877 ( .A(n44197), .B(n40900), .Z(n44202) );
  NOR U53878 ( .A(n40901), .B(n44202), .Z(n40902) );
  NOR U53879 ( .A(n44576), .B(n40902), .Z(n41205) );
  XOR U53880 ( .A(n40903), .B(n41205), .Z(n41200) );
  XOR U53881 ( .A(n41198), .B(n41200), .Z(n44208) );
  IV U53882 ( .A(n40904), .Z(n40905) );
  NOR U53883 ( .A(n40906), .B(n40905), .Z(n44207) );
  IV U53884 ( .A(n40907), .Z(n40908) );
  NOR U53885 ( .A(n40909), .B(n40908), .Z(n41201) );
  NOR U53886 ( .A(n44207), .B(n41201), .Z(n40910) );
  XOR U53887 ( .A(n44208), .B(n40910), .Z(n44210) );
  IV U53888 ( .A(n44210), .Z(n47602) );
  XOR U53889 ( .A(n44211), .B(n47602), .Z(n41194) );
  XOR U53890 ( .A(n40911), .B(n41194), .Z(n41192) );
  XOR U53891 ( .A(n41190), .B(n41192), .Z(n44222) );
  IV U53892 ( .A(n40912), .Z(n40913) );
  NOR U53893 ( .A(n40914), .B(n40913), .Z(n44221) );
  IV U53894 ( .A(n40915), .Z(n40917) );
  NOR U53895 ( .A(n40917), .B(n40916), .Z(n41188) );
  NOR U53896 ( .A(n44221), .B(n41188), .Z(n40918) );
  XOR U53897 ( .A(n44222), .B(n40918), .Z(n41186) );
  XOR U53898 ( .A(n40919), .B(n41186), .Z(n44234) );
  XOR U53899 ( .A(n44232), .B(n44234), .Z(n41182) );
  XOR U53900 ( .A(n41183), .B(n41182), .Z(n41180) );
  NOR U53901 ( .A(n40927), .B(n40920), .Z(n41179) );
  IV U53902 ( .A(n40921), .Z(n40923) );
  NOR U53903 ( .A(n40923), .B(n40922), .Z(n44229) );
  NOR U53904 ( .A(n41179), .B(n44229), .Z(n40924) );
  XOR U53905 ( .A(n41180), .B(n40924), .Z(n41178) );
  IV U53906 ( .A(n40925), .Z(n40926) );
  NOR U53907 ( .A(n40927), .B(n40926), .Z(n41176) );
  XOR U53908 ( .A(n41178), .B(n41176), .Z(n44242) );
  XOR U53909 ( .A(n44240), .B(n44242), .Z(n44244) );
  XOR U53910 ( .A(n40928), .B(n44244), .Z(n41173) );
  XOR U53911 ( .A(n41172), .B(n41173), .Z(n41167) );
  IV U53912 ( .A(n40929), .Z(n40931) );
  NOR U53913 ( .A(n40931), .B(n40930), .Z(n41170) );
  IV U53914 ( .A(n40932), .Z(n40933) );
  NOR U53915 ( .A(n40933), .B(n40936), .Z(n41166) );
  NOR U53916 ( .A(n41170), .B(n41166), .Z(n40934) );
  XOR U53917 ( .A(n41167), .B(n40934), .Z(n41162) );
  IV U53918 ( .A(n40935), .Z(n40937) );
  NOR U53919 ( .A(n40937), .B(n40936), .Z(n41160) );
  XOR U53920 ( .A(n41162), .B(n41160), .Z(n41165) );
  XOR U53921 ( .A(n41163), .B(n41165), .Z(n44253) );
  IV U53922 ( .A(n40938), .Z(n40939) );
  NOR U53923 ( .A(n40945), .B(n40939), .Z(n44250) );
  NOR U53924 ( .A(n40941), .B(n40940), .Z(n44252) );
  NOR U53925 ( .A(n44250), .B(n44252), .Z(n40942) );
  XOR U53926 ( .A(n44253), .B(n40942), .Z(n40951) );
  IV U53927 ( .A(n40951), .Z(n40957) );
  IV U53928 ( .A(n40943), .Z(n40944) );
  NOR U53929 ( .A(n40945), .B(n40944), .Z(n40952) );
  IV U53930 ( .A(n40952), .Z(n40946) );
  NOR U53931 ( .A(n40957), .B(n40946), .Z(n44524) );
  IV U53932 ( .A(n40947), .Z(n40950) );
  IV U53933 ( .A(n40948), .Z(n40949) );
  NOR U53934 ( .A(n40950), .B(n40949), .Z(n44255) );
  NOR U53935 ( .A(n40952), .B(n40951), .Z(n44257) );
  XOR U53936 ( .A(n44255), .B(n44257), .Z(n40953) );
  NOR U53937 ( .A(n44524), .B(n40953), .Z(n40954) );
  NOR U53938 ( .A(n40955), .B(n40954), .Z(n40958) );
  IV U53939 ( .A(n40955), .Z(n40956) );
  NOR U53940 ( .A(n40957), .B(n40956), .Z(n47651) );
  NOR U53941 ( .A(n40958), .B(n47651), .Z(n40959) );
  IV U53942 ( .A(n40959), .Z(n41159) );
  IV U53943 ( .A(n40960), .Z(n40961) );
  NOR U53944 ( .A(n40962), .B(n40961), .Z(n41157) );
  XOR U53945 ( .A(n41159), .B(n41157), .Z(n41153) );
  IV U53946 ( .A(n40963), .Z(n40965) );
  NOR U53947 ( .A(n40965), .B(n40964), .Z(n41151) );
  XOR U53948 ( .A(n41153), .B(n41151), .Z(n41156) );
  IV U53949 ( .A(n40966), .Z(n40967) );
  NOR U53950 ( .A(n40968), .B(n40967), .Z(n41154) );
  XOR U53951 ( .A(n41156), .B(n41154), .Z(n44263) );
  XOR U53952 ( .A(n44262), .B(n44263), .Z(n44267) );
  XOR U53953 ( .A(n40970), .B(n40969), .Z(n40972) );
  NOR U53954 ( .A(n40972), .B(n40971), .Z(n40973) );
  IV U53955 ( .A(n40973), .Z(n40974) );
  NOR U53956 ( .A(n40975), .B(n40974), .Z(n44265) );
  XOR U53957 ( .A(n44267), .B(n44265), .Z(n41149) );
  XOR U53958 ( .A(n41148), .B(n41149), .Z(n41146) );
  XOR U53959 ( .A(n41143), .B(n41146), .Z(n41142) );
  IV U53960 ( .A(n40976), .Z(n40979) );
  IV U53961 ( .A(n40977), .Z(n40978) );
  NOR U53962 ( .A(n40979), .B(n40978), .Z(n41145) );
  IV U53963 ( .A(n40980), .Z(n40982) );
  IV U53964 ( .A(n40981), .Z(n40988) );
  NOR U53965 ( .A(n40982), .B(n40988), .Z(n41140) );
  NOR U53966 ( .A(n41145), .B(n41140), .Z(n40983) );
  XOR U53967 ( .A(n41142), .B(n40983), .Z(n41136) );
  IV U53968 ( .A(n40984), .Z(n40985) );
  NOR U53969 ( .A(n40986), .B(n40985), .Z(n41137) );
  IV U53970 ( .A(n40987), .Z(n40989) );
  NOR U53971 ( .A(n40989), .B(n40988), .Z(n44275) );
  NOR U53972 ( .A(n41137), .B(n44275), .Z(n40990) );
  XOR U53973 ( .A(n41136), .B(n40990), .Z(n44505) );
  IV U53974 ( .A(n40991), .Z(n40992) );
  NOR U53975 ( .A(n40993), .B(n40992), .Z(n47672) );
  IV U53976 ( .A(n40994), .Z(n40996) );
  NOR U53977 ( .A(n40996), .B(n40995), .Z(n44504) );
  NOR U53978 ( .A(n47672), .B(n44504), .Z(n44278) );
  XOR U53979 ( .A(n44505), .B(n44278), .Z(n41134) );
  XOR U53980 ( .A(n40997), .B(n41134), .Z(n41132) );
  XOR U53981 ( .A(n40998), .B(n41132), .Z(n41123) );
  XOR U53982 ( .A(n40999), .B(n41123), .Z(n41118) );
  XOR U53983 ( .A(n41116), .B(n41118), .Z(n41121) );
  IV U53984 ( .A(n41000), .Z(n41002) );
  NOR U53985 ( .A(n41002), .B(n41001), .Z(n41119) );
  XOR U53986 ( .A(n41121), .B(n41119), .Z(n44291) );
  XOR U53987 ( .A(n44290), .B(n44291), .Z(n44294) );
  IV U53988 ( .A(n41003), .Z(n41004) );
  NOR U53989 ( .A(n41005), .B(n41004), .Z(n41006) );
  IV U53990 ( .A(n41006), .Z(n44293) );
  XOR U53991 ( .A(n44294), .B(n44293), .Z(n41110) );
  XOR U53992 ( .A(n41109), .B(n41110), .Z(n44298) );
  IV U53993 ( .A(n41007), .Z(n47817) );
  NOR U53994 ( .A(n47819), .B(n47817), .Z(n41112) );
  IV U53995 ( .A(n41008), .Z(n41010) );
  IV U53996 ( .A(n41009), .Z(n41021) );
  NOR U53997 ( .A(n41010), .B(n41021), .Z(n44297) );
  NOR U53998 ( .A(n41112), .B(n44297), .Z(n41011) );
  XOR U53999 ( .A(n44298), .B(n41011), .Z(n41022) );
  IV U54000 ( .A(n41022), .Z(n44302) );
  IV U54001 ( .A(n41012), .Z(n41014) );
  NOR U54002 ( .A(n41014), .B(n41013), .Z(n41015) );
  IV U54003 ( .A(n41015), .Z(n41023) );
  NOR U54004 ( .A(n44302), .B(n41023), .Z(n47687) );
  IV U54005 ( .A(n41016), .Z(n41018) );
  NOR U54006 ( .A(n41018), .B(n41017), .Z(n44304) );
  IV U54007 ( .A(n41019), .Z(n41020) );
  NOR U54008 ( .A(n41021), .B(n41020), .Z(n44300) );
  XOR U54009 ( .A(n44300), .B(n41022), .Z(n44305) );
  XOR U54010 ( .A(n44304), .B(n44305), .Z(n41025) );
  NOR U54011 ( .A(n44305), .B(n41023), .Z(n41024) );
  NOR U54012 ( .A(n41025), .B(n41024), .Z(n41026) );
  NOR U54013 ( .A(n47687), .B(n41026), .Z(n41027) );
  IV U54014 ( .A(n41027), .Z(n44309) );
  XOR U54015 ( .A(n41028), .B(n44309), .Z(n44316) );
  XOR U54016 ( .A(n44314), .B(n44316), .Z(n41107) );
  XOR U54017 ( .A(n41106), .B(n41107), .Z(n41100) );
  XOR U54018 ( .A(n41099), .B(n41100), .Z(n41103) );
  XOR U54019 ( .A(n41102), .B(n41103), .Z(n41094) );
  XOR U54020 ( .A(n41029), .B(n41094), .Z(n41092) );
  XOR U54021 ( .A(n41090), .B(n41092), .Z(n41089) );
  IV U54022 ( .A(n41030), .Z(n41031) );
  NOR U54023 ( .A(n41032), .B(n41031), .Z(n41085) );
  IV U54024 ( .A(n41033), .Z(n41035) );
  NOR U54025 ( .A(n41035), .B(n41034), .Z(n41087) );
  NOR U54026 ( .A(n41085), .B(n41087), .Z(n41036) );
  XOR U54027 ( .A(n41089), .B(n41036), .Z(n41078) );
  IV U54028 ( .A(n41037), .Z(n41038) );
  NOR U54029 ( .A(n41039), .B(n41038), .Z(n41082) );
  IV U54030 ( .A(n41040), .Z(n41041) );
  NOR U54031 ( .A(n41041), .B(n41044), .Z(n41079) );
  NOR U54032 ( .A(n41082), .B(n41079), .Z(n41042) );
  XOR U54033 ( .A(n41078), .B(n41042), .Z(n41076) );
  IV U54034 ( .A(n41043), .Z(n41045) );
  NOR U54035 ( .A(n41045), .B(n41044), .Z(n41075) );
  XOR U54036 ( .A(n41075), .B(n41046), .Z(n41047) );
  XOR U54037 ( .A(n41076), .B(n41047), .Z(n44328) );
  XOR U54038 ( .A(n44327), .B(n44328), .Z(n44330) );
  XOR U54039 ( .A(n44331), .B(n44330), .Z(n41058) );
  IV U54040 ( .A(n41048), .Z(n41050) );
  NOR U54041 ( .A(n41050), .B(n41049), .Z(n41059) );
  NOR U54042 ( .A(n41061), .B(n41059), .Z(n41051) );
  XOR U54043 ( .A(n41058), .B(n41051), .Z(n44335) );
  XOR U54044 ( .A(n44333), .B(n44335), .Z(n44365) );
  NOR U54045 ( .A(n41052), .B(n44365), .Z(n44417) );
  NOR U54046 ( .A(n41054), .B(n41053), .Z(n41055) );
  IV U54047 ( .A(n41055), .Z(n44341) );
  NOR U54048 ( .A(n44337), .B(n44341), .Z(n44363) );
  IV U54049 ( .A(n44363), .Z(n41056) );
  NOR U54050 ( .A(n41056), .B(n44365), .Z(n41057) );
  IV U54051 ( .A(n41057), .Z(n44424) );
  IV U54052 ( .A(n41058), .Z(n41062) );
  IV U54053 ( .A(n41059), .Z(n41060) );
  NOR U54054 ( .A(n41062), .B(n41060), .Z(n47722) );
  IV U54055 ( .A(n41061), .Z(n41063) );
  NOR U54056 ( .A(n41063), .B(n41062), .Z(n44431) );
  NOR U54057 ( .A(n41076), .B(n41064), .Z(n41065) );
  IV U54058 ( .A(n41065), .Z(n41070) );
  NOR U54059 ( .A(n41067), .B(n41066), .Z(n41068) );
  IV U54060 ( .A(n41068), .Z(n41069) );
  NOR U54061 ( .A(n41070), .B(n41069), .Z(n41071) );
  IV U54062 ( .A(n41071), .Z(n41072) );
  NOR U54063 ( .A(n41073), .B(n41072), .Z(n41074) );
  IV U54064 ( .A(n41074), .Z(n44438) );
  IV U54065 ( .A(n41075), .Z(n41077) );
  NOR U54066 ( .A(n41077), .B(n41076), .Z(n41081) );
  IV U54067 ( .A(n41078), .Z(n41084) );
  IV U54068 ( .A(n41079), .Z(n41080) );
  NOR U54069 ( .A(n41084), .B(n41080), .Z(n51168) );
  NOR U54070 ( .A(n41081), .B(n51168), .Z(n44445) );
  IV U54071 ( .A(n44445), .Z(n44326) );
  IV U54072 ( .A(n41082), .Z(n41083) );
  NOR U54073 ( .A(n41084), .B(n41083), .Z(n44442) );
  IV U54074 ( .A(n41085), .Z(n41086) );
  NOR U54075 ( .A(n41086), .B(n41089), .Z(n44446) );
  IV U54076 ( .A(n41087), .Z(n41088) );
  NOR U54077 ( .A(n41089), .B(n41088), .Z(n47708) );
  IV U54078 ( .A(n41090), .Z(n41091) );
  NOR U54079 ( .A(n41092), .B(n41091), .Z(n47705) );
  IV U54080 ( .A(n41093), .Z(n41095) );
  NOR U54081 ( .A(n41095), .B(n41094), .Z(n47701) );
  NOR U54082 ( .A(n47705), .B(n47701), .Z(n44324) );
  NOR U54083 ( .A(n41096), .B(n41103), .Z(n41097) );
  IV U54084 ( .A(n41097), .Z(n44450) );
  NOR U54085 ( .A(n44450), .B(n41098), .Z(n44323) );
  IV U54086 ( .A(n41099), .Z(n41101) );
  NOR U54087 ( .A(n41101), .B(n41100), .Z(n44459) );
  IV U54088 ( .A(n41102), .Z(n41104) );
  NOR U54089 ( .A(n41104), .B(n41103), .Z(n44457) );
  NOR U54090 ( .A(n44459), .B(n44457), .Z(n41105) );
  IV U54091 ( .A(n41105), .Z(n44322) );
  IV U54092 ( .A(n41106), .Z(n41108) );
  NOR U54093 ( .A(n41108), .B(n41107), .Z(n47690) );
  IV U54094 ( .A(n41110), .Z(n47822) );
  NOR U54095 ( .A(n41109), .B(n47822), .Z(n51139) );
  NOR U54096 ( .A(n41111), .B(n41110), .Z(n41114) );
  IV U54097 ( .A(n41112), .Z(n41113) );
  NOR U54098 ( .A(n41114), .B(n41113), .Z(n41115) );
  NOR U54099 ( .A(n51139), .B(n41115), .Z(n44476) );
  IV U54100 ( .A(n44476), .Z(n44296) );
  IV U54101 ( .A(n41116), .Z(n41117) );
  NOR U54102 ( .A(n41118), .B(n41117), .Z(n44488) );
  IV U54103 ( .A(n41119), .Z(n41120) );
  NOR U54104 ( .A(n41121), .B(n41120), .Z(n44483) );
  NOR U54105 ( .A(n44488), .B(n44483), .Z(n44289) );
  IV U54106 ( .A(n41122), .Z(n41124) );
  IV U54107 ( .A(n41123), .Z(n41126) );
  NOR U54108 ( .A(n41124), .B(n41126), .Z(n44485) );
  IV U54109 ( .A(n41125), .Z(n41127) );
  NOR U54110 ( .A(n41127), .B(n41126), .Z(n44494) );
  IV U54111 ( .A(n41128), .Z(n41129) );
  NOR U54112 ( .A(n41132), .B(n41129), .Z(n44491) );
  IV U54113 ( .A(n41130), .Z(n41131) );
  NOR U54114 ( .A(n41132), .B(n41131), .Z(n44497) );
  IV U54115 ( .A(n41133), .Z(n41135) );
  IV U54116 ( .A(n41134), .Z(n44280) );
  NOR U54117 ( .A(n41135), .B(n44280), .Z(n47679) );
  IV U54118 ( .A(n41136), .Z(n44277) );
  IV U54119 ( .A(n41137), .Z(n41138) );
  NOR U54120 ( .A(n44277), .B(n41138), .Z(n41139) );
  IV U54121 ( .A(n41139), .Z(n47671) );
  IV U54122 ( .A(n41140), .Z(n41141) );
  NOR U54123 ( .A(n41142), .B(n41141), .Z(n44514) );
  IV U54124 ( .A(n41143), .Z(n41144) );
  NOR U54125 ( .A(n41144), .B(n41146), .Z(n47667) );
  IV U54126 ( .A(n41145), .Z(n41147) );
  NOR U54127 ( .A(n41147), .B(n41146), .Z(n44512) );
  NOR U54128 ( .A(n47667), .B(n44512), .Z(n44274) );
  IV U54129 ( .A(n41148), .Z(n41150) );
  NOR U54130 ( .A(n41150), .B(n41149), .Z(n44270) );
  IV U54131 ( .A(n41151), .Z(n41152) );
  NOR U54132 ( .A(n41153), .B(n41152), .Z(n47654) );
  IV U54133 ( .A(n41154), .Z(n41155) );
  NOR U54134 ( .A(n41156), .B(n41155), .Z(n47660) );
  NOR U54135 ( .A(n47654), .B(n47660), .Z(n44260) );
  IV U54136 ( .A(n41157), .Z(n41158) );
  NOR U54137 ( .A(n41159), .B(n41158), .Z(n47656) );
  NOR U54138 ( .A(n47651), .B(n47656), .Z(n44259) );
  IV U54139 ( .A(n41160), .Z(n41161) );
  NOR U54140 ( .A(n41162), .B(n41161), .Z(n47638) );
  IV U54141 ( .A(n41163), .Z(n41164) );
  NOR U54142 ( .A(n41165), .B(n41164), .Z(n44534) );
  NOR U54143 ( .A(n47638), .B(n44534), .Z(n44248) );
  IV U54144 ( .A(n41166), .Z(n41169) );
  IV U54145 ( .A(n41167), .Z(n41168) );
  NOR U54146 ( .A(n41169), .B(n41168), .Z(n44536) );
  IV U54147 ( .A(n41170), .Z(n41171) );
  NOR U54148 ( .A(n41173), .B(n41171), .Z(n47641) );
  NOR U54149 ( .A(n41173), .B(n41172), .Z(n44541) );
  IV U54150 ( .A(n41174), .Z(n41175) );
  NOR U54151 ( .A(n41175), .B(n44244), .Z(n44543) );
  NOR U54152 ( .A(n44541), .B(n44543), .Z(n44247) );
  IV U54153 ( .A(n41176), .Z(n41177) );
  NOR U54154 ( .A(n41178), .B(n41177), .Z(n47883) );
  IV U54155 ( .A(n41179), .Z(n41181) );
  IV U54156 ( .A(n41180), .Z(n44231) );
  NOR U54157 ( .A(n41181), .B(n44231), .Z(n47879) );
  NOR U54158 ( .A(n47883), .B(n47879), .Z(n44549) );
  NOR U54159 ( .A(n41183), .B(n41182), .Z(n41184) );
  IV U54160 ( .A(n41184), .Z(n44236) );
  IV U54161 ( .A(n41185), .Z(n41187) );
  IV U54162 ( .A(n41186), .Z(n44225) );
  NOR U54163 ( .A(n41187), .B(n44225), .Z(n44558) );
  IV U54164 ( .A(n41188), .Z(n41189) );
  NOR U54165 ( .A(n44222), .B(n41189), .Z(n47624) );
  IV U54166 ( .A(n41190), .Z(n41191) );
  NOR U54167 ( .A(n41192), .B(n41191), .Z(n47613) );
  IV U54168 ( .A(n41193), .Z(n41197) );
  NOR U54169 ( .A(n41195), .B(n41194), .Z(n41196) );
  IV U54170 ( .A(n41196), .Z(n44219) );
  NOR U54171 ( .A(n41197), .B(n44219), .Z(n47616) );
  IV U54172 ( .A(n41198), .Z(n41199) );
  NOR U54173 ( .A(n41200), .B(n41199), .Z(n44567) );
  IV U54174 ( .A(n41201), .Z(n41202) );
  NOR U54175 ( .A(n44208), .B(n41202), .Z(n47596) );
  NOR U54176 ( .A(n44567), .B(n47596), .Z(n41203) );
  IV U54177 ( .A(n41203), .Z(n44206) );
  IV U54178 ( .A(n41204), .Z(n41207) );
  IV U54179 ( .A(n41205), .Z(n41206) );
  NOR U54180 ( .A(n41207), .B(n41206), .Z(n44573) );
  IV U54181 ( .A(n41208), .Z(n41210) );
  NOR U54182 ( .A(n41210), .B(n41209), .Z(n44586) );
  IV U54183 ( .A(n41211), .Z(n41216) );
  IV U54184 ( .A(n41212), .Z(n41213) );
  NOR U54185 ( .A(n41216), .B(n41213), .Z(n44588) );
  NOR U54186 ( .A(n44586), .B(n44588), .Z(n44173) );
  IV U54187 ( .A(n41214), .Z(n41215) );
  NOR U54188 ( .A(n41216), .B(n41215), .Z(n47566) );
  IV U54189 ( .A(n41217), .Z(n41218) );
  NOR U54190 ( .A(n41219), .B(n41218), .Z(n47562) );
  IV U54191 ( .A(n41220), .Z(n41223) );
  XOR U54192 ( .A(n41221), .B(n41227), .Z(n41222) );
  NOR U54193 ( .A(n41223), .B(n41222), .Z(n47569) );
  IV U54194 ( .A(n41224), .Z(n41225) );
  NOR U54195 ( .A(n41225), .B(n41227), .Z(n51009) );
  IV U54196 ( .A(n41226), .Z(n41230) );
  NOR U54197 ( .A(n41228), .B(n41227), .Z(n41229) );
  IV U54198 ( .A(n41229), .Z(n44170) );
  NOR U54199 ( .A(n41230), .B(n44170), .Z(n47937) );
  NOR U54200 ( .A(n51009), .B(n47937), .Z(n47559) );
  IV U54201 ( .A(n41231), .Z(n41232) );
  NOR U54202 ( .A(n41233), .B(n41232), .Z(n47551) );
  NOR U54203 ( .A(n47550), .B(n47551), .Z(n50997) );
  IV U54204 ( .A(n41234), .Z(n41235) );
  NOR U54205 ( .A(n41236), .B(n41235), .Z(n47524) );
  IV U54206 ( .A(n41237), .Z(n41238) );
  NOR U54207 ( .A(n41239), .B(n41238), .Z(n44592) );
  IV U54208 ( .A(n41240), .Z(n41241) );
  NOR U54209 ( .A(n44139), .B(n41241), .Z(n47501) );
  NOR U54210 ( .A(n41243), .B(n41242), .Z(n41246) );
  NOR U54211 ( .A(n41244), .B(n44130), .Z(n41245) );
  IV U54212 ( .A(n41245), .Z(n44597) );
  NOR U54213 ( .A(n41246), .B(n44597), .Z(n44133) );
  IV U54214 ( .A(n41247), .Z(n41249) );
  NOR U54215 ( .A(n41249), .B(n41248), .Z(n41250) );
  IV U54216 ( .A(n41250), .Z(n44125) );
  IV U54217 ( .A(n41251), .Z(n41252) );
  NOR U54218 ( .A(n44123), .B(n41252), .Z(n47485) );
  IV U54219 ( .A(n41253), .Z(n41256) );
  IV U54220 ( .A(n41254), .Z(n41255) );
  NOR U54221 ( .A(n41256), .B(n41255), .Z(n47470) );
  IV U54222 ( .A(n41257), .Z(n41258) );
  NOR U54223 ( .A(n41262), .B(n41258), .Z(n47463) );
  IV U54224 ( .A(n41259), .Z(n41260) );
  NOR U54225 ( .A(n41266), .B(n41260), .Z(n47977) );
  IV U54226 ( .A(n41261), .Z(n41263) );
  NOR U54227 ( .A(n41263), .B(n41262), .Z(n50911) );
  NOR U54228 ( .A(n47977), .B(n50911), .Z(n47460) );
  IV U54229 ( .A(n47460), .Z(n44098) );
  IV U54230 ( .A(n41264), .Z(n41265) );
  NOR U54231 ( .A(n41266), .B(n41265), .Z(n47457) );
  IV U54232 ( .A(n41267), .Z(n41268) );
  NOR U54233 ( .A(n44090), .B(n41268), .Z(n41269) );
  IV U54234 ( .A(n41269), .Z(n47444) );
  IV U54235 ( .A(n41270), .Z(n41271) );
  NOR U54236 ( .A(n41271), .B(n44083), .Z(n44619) );
  IV U54237 ( .A(n41272), .Z(n41275) );
  IV U54238 ( .A(n41273), .Z(n41274) );
  NOR U54239 ( .A(n41275), .B(n41274), .Z(n44613) );
  NOR U54240 ( .A(n44619), .B(n44613), .Z(n41276) );
  IV U54241 ( .A(n41276), .Z(n44087) );
  IV U54242 ( .A(n41277), .Z(n47438) );
  IV U54243 ( .A(n41278), .Z(n41279) );
  NOR U54244 ( .A(n41280), .B(n41279), .Z(n47424) );
  IV U54245 ( .A(n41281), .Z(n41282) );
  NOR U54246 ( .A(n41282), .B(n41287), .Z(n50870) );
  IV U54247 ( .A(n41283), .Z(n44076) );
  IV U54248 ( .A(n41284), .Z(n41285) );
  NOR U54249 ( .A(n44076), .B(n41285), .Z(n47999) );
  NOR U54250 ( .A(n50870), .B(n47999), .Z(n47427) );
  IV U54251 ( .A(n41286), .Z(n41288) );
  NOR U54252 ( .A(n41288), .B(n41287), .Z(n47420) );
  IV U54253 ( .A(n41289), .Z(n41294) );
  IV U54254 ( .A(n41290), .Z(n41291) );
  NOR U54255 ( .A(n41294), .B(n41291), .Z(n47417) );
  IV U54256 ( .A(n41292), .Z(n41293) );
  NOR U54257 ( .A(n41294), .B(n41293), .Z(n44636) );
  IV U54258 ( .A(n41295), .Z(n41297) );
  NOR U54259 ( .A(n41297), .B(n41296), .Z(n44633) );
  IV U54260 ( .A(n41298), .Z(n41299) );
  NOR U54261 ( .A(n44070), .B(n41299), .Z(n47413) );
  IV U54262 ( .A(n41300), .Z(n47405) );
  NOR U54263 ( .A(n41302), .B(n41301), .Z(n48022) );
  IV U54264 ( .A(n41303), .Z(n41306) );
  IV U54265 ( .A(n41304), .Z(n41305) );
  NOR U54266 ( .A(n41306), .B(n41305), .Z(n50851) );
  NOR U54267 ( .A(n48022), .B(n50851), .Z(n44640) );
  IV U54268 ( .A(n41307), .Z(n41310) );
  IV U54269 ( .A(n41308), .Z(n41309) );
  NOR U54270 ( .A(n41310), .B(n41309), .Z(n50836) );
  IV U54271 ( .A(n41311), .Z(n41313) );
  NOR U54272 ( .A(n41313), .B(n41312), .Z(n50829) );
  NOR U54273 ( .A(n50836), .B(n50829), .Z(n47399) );
  IV U54274 ( .A(n50838), .Z(n47398) );
  NOR U54275 ( .A(n41315), .B(n41314), .Z(n41316) );
  IV U54276 ( .A(n41316), .Z(n44645) );
  IV U54277 ( .A(n41317), .Z(n47393) );
  IV U54278 ( .A(n41318), .Z(n41319) );
  NOR U54279 ( .A(n41319), .B(n51650), .Z(n47388) );
  IV U54280 ( .A(n47388), .Z(n44052) );
  IV U54281 ( .A(n41320), .Z(n41325) );
  IV U54282 ( .A(n41321), .Z(n41322) );
  NOR U54283 ( .A(n41322), .B(n44031), .Z(n41323) );
  IV U54284 ( .A(n41323), .Z(n41324) );
  NOR U54285 ( .A(n41325), .B(n41324), .Z(n44660) );
  IV U54286 ( .A(n41326), .Z(n41330) );
  NOR U54287 ( .A(n41327), .B(n41332), .Z(n41328) );
  IV U54288 ( .A(n41328), .Z(n41329) );
  NOR U54289 ( .A(n41330), .B(n41329), .Z(n47380) );
  IV U54290 ( .A(n41331), .Z(n41333) );
  NOR U54291 ( .A(n41333), .B(n41332), .Z(n48049) );
  IV U54292 ( .A(n41334), .Z(n41335) );
  NOR U54293 ( .A(n41336), .B(n41335), .Z(n48040) );
  NOR U54294 ( .A(n48049), .B(n48040), .Z(n47379) );
  IV U54295 ( .A(n41337), .Z(n44013) );
  IV U54296 ( .A(n41338), .Z(n41339) );
  NOR U54297 ( .A(n44013), .B(n41339), .Z(n47365) );
  IV U54298 ( .A(n41340), .Z(n41341) );
  NOR U54299 ( .A(n41341), .B(n44000), .Z(n44670) );
  NOR U54300 ( .A(n41342), .B(n44677), .Z(n41346) );
  IV U54301 ( .A(n41343), .Z(n41345) );
  NOR U54302 ( .A(n41345), .B(n41344), .Z(n44673) );
  NOR U54303 ( .A(n41346), .B(n44673), .Z(n41347) );
  IV U54304 ( .A(n41347), .Z(n43998) );
  IV U54305 ( .A(n41348), .Z(n41353) );
  IV U54306 ( .A(n41349), .Z(n41350) );
  NOR U54307 ( .A(n41353), .B(n41350), .Z(n47350) );
  IV U54308 ( .A(n41351), .Z(n41352) );
  NOR U54309 ( .A(n41353), .B(n41352), .Z(n47347) );
  XOR U54310 ( .A(n41355), .B(n41354), .Z(n41356) );
  NOR U54311 ( .A(n43989), .B(n41356), .Z(n41357) );
  IV U54312 ( .A(n41357), .Z(n41358) );
  NOR U54313 ( .A(n41359), .B(n41358), .Z(n43992) );
  IV U54314 ( .A(n43992), .Z(n43986) );
  IV U54315 ( .A(n41360), .Z(n41362) );
  IV U54316 ( .A(n41361), .Z(n41366) );
  NOR U54317 ( .A(n41362), .B(n41366), .Z(n47342) );
  IV U54318 ( .A(n41363), .Z(n41364) );
  NOR U54319 ( .A(n41364), .B(n41372), .Z(n48080) );
  IV U54320 ( .A(n41365), .Z(n41367) );
  NOR U54321 ( .A(n41367), .B(n41366), .Z(n48074) );
  NOR U54322 ( .A(n48080), .B(n48074), .Z(n47341) );
  IV U54323 ( .A(n41368), .Z(n41370) );
  NOR U54324 ( .A(n41370), .B(n41369), .Z(n47332) );
  IV U54325 ( .A(n41371), .Z(n41373) );
  NOR U54326 ( .A(n41373), .B(n41372), .Z(n47337) );
  NOR U54327 ( .A(n47332), .B(n47337), .Z(n43983) );
  IV U54328 ( .A(n41374), .Z(n41376) );
  NOR U54329 ( .A(n41376), .B(n41375), .Z(n41377) );
  IV U54330 ( .A(n41377), .Z(n44697) );
  IV U54331 ( .A(n41378), .Z(n41379) );
  NOR U54332 ( .A(n43963), .B(n41379), .Z(n41380) );
  IV U54333 ( .A(n41380), .Z(n43964) );
  IV U54334 ( .A(n41381), .Z(n41383) );
  IV U54335 ( .A(n41382), .Z(n43959) );
  NOR U54336 ( .A(n41383), .B(n43959), .Z(n44704) );
  IV U54337 ( .A(n41384), .Z(n41385) );
  NOR U54338 ( .A(n41386), .B(n41385), .Z(n44701) );
  IV U54339 ( .A(n41387), .Z(n41389) );
  IV U54340 ( .A(n41388), .Z(n41393) );
  NOR U54341 ( .A(n41389), .B(n41393), .Z(n44710) );
  IV U54342 ( .A(n41390), .Z(n41391) );
  NOR U54343 ( .A(n41391), .B(n41393), .Z(n44707) );
  IV U54344 ( .A(n41392), .Z(n41394) );
  NOR U54345 ( .A(n41394), .B(n41393), .Z(n47323) );
  IV U54346 ( .A(n41395), .Z(n41396) );
  NOR U54347 ( .A(n41399), .B(n41396), .Z(n47320) );
  IV U54348 ( .A(n41397), .Z(n41398) );
  NOR U54349 ( .A(n41399), .B(n41398), .Z(n44713) );
  IV U54350 ( .A(n41400), .Z(n41405) );
  IV U54351 ( .A(n41401), .Z(n41402) );
  NOR U54352 ( .A(n41403), .B(n41402), .Z(n41404) );
  IV U54353 ( .A(n41404), .Z(n43956) );
  NOR U54354 ( .A(n41405), .B(n43956), .Z(n44716) );
  IV U54355 ( .A(n41406), .Z(n41408) );
  NOR U54356 ( .A(n41408), .B(n41407), .Z(n47294) );
  IV U54357 ( .A(n41409), .Z(n41419) );
  IV U54358 ( .A(n41410), .Z(n41411) );
  NOR U54359 ( .A(n41419), .B(n41411), .Z(n47297) );
  XOR U54360 ( .A(n41412), .B(n41419), .Z(n41415) );
  IV U54361 ( .A(n41413), .Z(n41414) );
  NOR U54362 ( .A(n41415), .B(n41414), .Z(n47298) );
  XOR U54363 ( .A(n47297), .B(n47298), .Z(n41416) );
  NOR U54364 ( .A(n47294), .B(n41416), .Z(n43944) );
  IV U54365 ( .A(n41417), .Z(n41421) );
  NOR U54366 ( .A(n41419), .B(n41418), .Z(n41420) );
  IV U54367 ( .A(n41420), .Z(n41423) );
  NOR U54368 ( .A(n41421), .B(n41423), .Z(n47289) );
  IV U54369 ( .A(n41422), .Z(n41424) );
  NOR U54370 ( .A(n41424), .B(n41423), .Z(n47285) );
  IV U54371 ( .A(n41425), .Z(n41427) );
  NOR U54372 ( .A(n41427), .B(n41426), .Z(n47282) );
  IV U54373 ( .A(n41428), .Z(n41429) );
  NOR U54374 ( .A(n43940), .B(n41429), .Z(n44724) );
  NOR U54375 ( .A(n41431), .B(n41430), .Z(n50681) );
  IV U54376 ( .A(n41432), .Z(n41434) );
  IV U54377 ( .A(n41433), .Z(n43942) );
  NOR U54378 ( .A(n41434), .B(n43942), .Z(n50689) );
  NOR U54379 ( .A(n50681), .B(n50689), .Z(n44727) );
  IV U54380 ( .A(n41435), .Z(n44734) );
  IV U54381 ( .A(n41436), .Z(n41437) );
  NOR U54382 ( .A(n44734), .B(n41437), .Z(n47274) );
  NOR U54383 ( .A(n41438), .B(n44734), .Z(n43937) );
  NOR U54384 ( .A(n41439), .B(n43935), .Z(n41440) );
  IV U54385 ( .A(n41440), .Z(n41441) );
  NOR U54386 ( .A(n41442), .B(n41441), .Z(n47267) );
  IV U54387 ( .A(n41443), .Z(n43929) );
  IV U54388 ( .A(n41444), .Z(n41445) );
  NOR U54389 ( .A(n43929), .B(n41445), .Z(n41446) );
  IV U54390 ( .A(n41446), .Z(n47259) );
  IV U54391 ( .A(n41447), .Z(n41448) );
  NOR U54392 ( .A(n41448), .B(n41452), .Z(n44742) );
  IV U54393 ( .A(n41449), .Z(n47242) );
  NOR U54394 ( .A(n47242), .B(n41450), .Z(n47232) );
  IV U54395 ( .A(n41451), .Z(n41453) );
  NOR U54396 ( .A(n41453), .B(n41452), .Z(n47238) );
  NOR U54397 ( .A(n47232), .B(n47238), .Z(n41454) );
  IV U54398 ( .A(n41454), .Z(n43926) );
  IV U54399 ( .A(n41455), .Z(n41456) );
  NOR U54400 ( .A(n41456), .B(n41462), .Z(n44746) );
  IV U54401 ( .A(n41457), .Z(n41458) );
  NOR U54402 ( .A(n41459), .B(n41458), .Z(n44750) );
  IV U54403 ( .A(n41460), .Z(n41461) );
  NOR U54404 ( .A(n41462), .B(n41461), .Z(n44748) );
  NOR U54405 ( .A(n44750), .B(n44748), .Z(n43924) );
  IV U54406 ( .A(n41463), .Z(n41466) );
  IV U54407 ( .A(n41464), .Z(n41465) );
  NOR U54408 ( .A(n41466), .B(n41465), .Z(n44754) );
  NOR U54409 ( .A(n41467), .B(n41474), .Z(n41468) );
  IV U54410 ( .A(n41468), .Z(n41471) );
  NOR U54411 ( .A(n41469), .B(n41471), .Z(n47226) );
  NOR U54412 ( .A(n44754), .B(n47226), .Z(n43923) );
  IV U54413 ( .A(n41470), .Z(n41472) );
  NOR U54414 ( .A(n41472), .B(n41471), .Z(n43919) );
  IV U54415 ( .A(n41473), .Z(n41475) );
  NOR U54416 ( .A(n41475), .B(n41474), .Z(n47219) );
  NOR U54417 ( .A(n41477), .B(n41476), .Z(n44756) );
  NOR U54418 ( .A(n47219), .B(n44756), .Z(n43917) );
  IV U54419 ( .A(n41478), .Z(n41479) );
  NOR U54420 ( .A(n41480), .B(n41479), .Z(n47222) );
  IV U54421 ( .A(n41481), .Z(n41485) );
  IV U54422 ( .A(n41482), .Z(n41483) );
  NOR U54423 ( .A(n41485), .B(n41483), .Z(n47216) );
  NOR U54424 ( .A(n47222), .B(n47216), .Z(n43916) );
  IV U54425 ( .A(n41484), .Z(n41486) );
  NOR U54426 ( .A(n41486), .B(n41485), .Z(n47212) );
  NOR U54427 ( .A(n47200), .B(n47212), .Z(n43915) );
  IV U54428 ( .A(n41487), .Z(n41491) );
  NOR U54429 ( .A(n43911), .B(n41488), .Z(n41489) );
  IV U54430 ( .A(n41489), .Z(n41490) );
  NOR U54431 ( .A(n41491), .B(n41490), .Z(n41492) );
  IV U54432 ( .A(n41492), .Z(n44765) );
  IV U54433 ( .A(n41493), .Z(n41494) );
  NOR U54434 ( .A(n41494), .B(n41496), .Z(n44761) );
  IV U54435 ( .A(n41495), .Z(n41499) );
  NOR U54436 ( .A(n41497), .B(n41496), .Z(n41498) );
  IV U54437 ( .A(n41498), .Z(n41504) );
  NOR U54438 ( .A(n41499), .B(n41504), .Z(n44767) );
  IV U54439 ( .A(n41500), .Z(n41502) );
  IV U54440 ( .A(n41501), .Z(n41508) );
  NOR U54441 ( .A(n41502), .B(n41508), .Z(n48188) );
  IV U54442 ( .A(n41503), .Z(n41505) );
  NOR U54443 ( .A(n41505), .B(n41504), .Z(n48184) );
  NOR U54444 ( .A(n48188), .B(n48184), .Z(n44766) );
  IV U54445 ( .A(n44766), .Z(n43906) );
  IV U54446 ( .A(n41506), .Z(n41507) );
  NOR U54447 ( .A(n41508), .B(n41507), .Z(n44771) );
  IV U54448 ( .A(n41509), .Z(n41510) );
  NOR U54449 ( .A(n43901), .B(n41510), .Z(n44777) );
  IV U54450 ( .A(n41511), .Z(n41512) );
  NOR U54451 ( .A(n41513), .B(n41512), .Z(n44785) );
  IV U54452 ( .A(n41514), .Z(n41515) );
  NOR U54453 ( .A(n41518), .B(n41515), .Z(n44788) );
  IV U54454 ( .A(n41516), .Z(n41520) );
  NOR U54455 ( .A(n41518), .B(n41517), .Z(n41519) );
  IV U54456 ( .A(n41519), .Z(n43893) );
  NOR U54457 ( .A(n41520), .B(n43893), .Z(n47190) );
  IV U54458 ( .A(n41521), .Z(n41522) );
  NOR U54459 ( .A(n41523), .B(n41522), .Z(n47182) );
  IV U54460 ( .A(n41524), .Z(n41525) );
  NOR U54461 ( .A(n43890), .B(n41525), .Z(n44791) );
  NOR U54462 ( .A(n47182), .B(n44791), .Z(n43887) );
  IV U54463 ( .A(n41526), .Z(n41529) );
  IV U54464 ( .A(n41527), .Z(n41528) );
  NOR U54465 ( .A(n41529), .B(n41528), .Z(n44797) );
  IV U54466 ( .A(n41530), .Z(n41533) );
  NOR U54467 ( .A(n41531), .B(n43881), .Z(n41532) );
  IV U54468 ( .A(n41532), .Z(n43884) );
  NOR U54469 ( .A(n41533), .B(n43884), .Z(n44794) );
  IV U54470 ( .A(n41534), .Z(n41535) );
  IV U54471 ( .A(n43836), .Z(n43834) );
  NOR U54472 ( .A(n41535), .B(n43834), .Z(n47148) );
  IV U54473 ( .A(n41536), .Z(n41537) );
  NOR U54474 ( .A(n41537), .B(n43844), .Z(n47152) );
  NOR U54475 ( .A(n47148), .B(n47152), .Z(n43841) );
  IV U54476 ( .A(n41538), .Z(n41539) );
  NOR U54477 ( .A(n43832), .B(n41539), .Z(n44826) );
  IV U54478 ( .A(n41540), .Z(n41545) );
  IV U54479 ( .A(n41541), .Z(n41542) );
  NOR U54480 ( .A(n41543), .B(n41542), .Z(n41544) );
  IV U54481 ( .A(n41544), .Z(n43824) );
  NOR U54482 ( .A(n41545), .B(n43824), .Z(n48233) );
  NOR U54483 ( .A(n48239), .B(n48233), .Z(n47140) );
  IV U54484 ( .A(n41546), .Z(n41547) );
  NOR U54485 ( .A(n41550), .B(n41547), .Z(n47133) );
  IV U54486 ( .A(n41548), .Z(n41552) );
  NOR U54487 ( .A(n41550), .B(n41549), .Z(n41551) );
  IV U54488 ( .A(n41551), .Z(n41554) );
  NOR U54489 ( .A(n41552), .B(n41554), .Z(n47130) );
  IV U54490 ( .A(n41553), .Z(n41555) );
  NOR U54491 ( .A(n41555), .B(n41554), .Z(n44838) );
  IV U54492 ( .A(n41556), .Z(n41559) );
  NOR U54493 ( .A(n41557), .B(n43820), .Z(n41558) );
  IV U54494 ( .A(n41558), .Z(n41561) );
  NOR U54495 ( .A(n41559), .B(n41561), .Z(n44844) );
  IV U54496 ( .A(n41560), .Z(n41562) );
  NOR U54497 ( .A(n41562), .B(n41561), .Z(n44841) );
  IV U54498 ( .A(n41563), .Z(n41564) );
  NOR U54499 ( .A(n43816), .B(n41564), .Z(n41565) );
  IV U54500 ( .A(n41565), .Z(n44851) );
  IV U54501 ( .A(n41566), .Z(n41567) );
  NOR U54502 ( .A(n43816), .B(n41567), .Z(n44847) );
  IV U54503 ( .A(n41568), .Z(n41572) );
  IV U54504 ( .A(n41569), .Z(n41576) );
  NOR U54505 ( .A(n41570), .B(n41576), .Z(n41571) );
  IV U54506 ( .A(n41571), .Z(n43797) );
  NOR U54507 ( .A(n41572), .B(n43797), .Z(n47108) );
  IV U54508 ( .A(n41573), .Z(n41574) );
  NOR U54509 ( .A(n41581), .B(n41574), .Z(n44871) );
  IV U54510 ( .A(n41575), .Z(n41577) );
  NOR U54511 ( .A(n41577), .B(n41576), .Z(n47111) );
  NOR U54512 ( .A(n44871), .B(n47111), .Z(n41578) );
  IV U54513 ( .A(n41578), .Z(n43794) );
  IV U54514 ( .A(n41579), .Z(n41580) );
  NOR U54515 ( .A(n41581), .B(n41580), .Z(n47105) );
  IV U54516 ( .A(n41582), .Z(n41584) );
  IV U54517 ( .A(n41583), .Z(n41586) );
  NOR U54518 ( .A(n41584), .B(n41586), .Z(n47102) );
  IV U54519 ( .A(n41585), .Z(n41587) );
  NOR U54520 ( .A(n41587), .B(n41586), .Z(n48271) );
  IV U54521 ( .A(n41588), .Z(n41591) );
  NOR U54522 ( .A(n41597), .B(n41589), .Z(n41590) );
  IV U54523 ( .A(n41590), .Z(n41593) );
  NOR U54524 ( .A(n41591), .B(n41593), .Z(n50496) );
  NOR U54525 ( .A(n48271), .B(n50496), .Z(n47099) );
  IV U54526 ( .A(n41592), .Z(n41594) );
  NOR U54527 ( .A(n41594), .B(n41593), .Z(n47095) );
  IV U54528 ( .A(n41595), .Z(n41596) );
  NOR U54529 ( .A(n41597), .B(n41596), .Z(n44874) );
  NOR U54530 ( .A(n47095), .B(n44874), .Z(n43793) );
  IV U54531 ( .A(n41598), .Z(n41600) );
  IV U54532 ( .A(n41599), .Z(n41604) );
  NOR U54533 ( .A(n41600), .B(n41604), .Z(n47084) );
  IV U54534 ( .A(n41601), .Z(n41602) );
  NOR U54535 ( .A(n41608), .B(n41602), .Z(n47079) );
  IV U54536 ( .A(n41603), .Z(n41605) );
  NOR U54537 ( .A(n41605), .B(n41604), .Z(n47077) );
  NOR U54538 ( .A(n47079), .B(n47077), .Z(n43792) );
  IV U54539 ( .A(n41606), .Z(n41607) );
  NOR U54540 ( .A(n41608), .B(n41607), .Z(n44876) );
  IV U54541 ( .A(n41609), .Z(n41613) );
  IV U54542 ( .A(n41610), .Z(n43785) );
  NOR U54543 ( .A(n41611), .B(n43785), .Z(n41612) );
  IV U54544 ( .A(n41612), .Z(n43789) );
  NOR U54545 ( .A(n41613), .B(n43789), .Z(n47065) );
  NOR U54546 ( .A(n44876), .B(n47065), .Z(n43791) );
  IV U54547 ( .A(n41614), .Z(n41615) );
  NOR U54548 ( .A(n41615), .B(n41617), .Z(n50453) );
  IV U54549 ( .A(n41616), .Z(n41618) );
  NOR U54550 ( .A(n41618), .B(n41617), .Z(n48286) );
  NOR U54551 ( .A(n50453), .B(n48286), .Z(n47050) );
  IV U54552 ( .A(n41619), .Z(n41621) );
  NOR U54553 ( .A(n41621), .B(n41620), .Z(n47047) );
  IV U54554 ( .A(n41622), .Z(n41623) );
  NOR U54555 ( .A(n41623), .B(n41625), .Z(n47043) );
  IV U54556 ( .A(n41624), .Z(n41626) );
  NOR U54557 ( .A(n41626), .B(n41625), .Z(n47040) );
  IV U54558 ( .A(n41627), .Z(n41630) );
  NOR U54559 ( .A(n41634), .B(n41628), .Z(n41629) );
  IV U54560 ( .A(n41629), .Z(n43769) );
  NOR U54561 ( .A(n41630), .B(n43769), .Z(n41631) );
  IV U54562 ( .A(n41631), .Z(n47034) );
  IV U54563 ( .A(n41632), .Z(n41633) );
  NOR U54564 ( .A(n41634), .B(n41633), .Z(n47030) );
  IV U54565 ( .A(n41635), .Z(n41637) );
  IV U54566 ( .A(n41636), .Z(n41639) );
  NOR U54567 ( .A(n41637), .B(n41639), .Z(n44887) );
  IV U54568 ( .A(n41638), .Z(n41640) );
  NOR U54569 ( .A(n41640), .B(n41639), .Z(n44881) );
  XOR U54570 ( .A(n44887), .B(n44881), .Z(n41641) );
  NOR U54571 ( .A(n47030), .B(n41641), .Z(n41642) );
  IV U54572 ( .A(n41642), .Z(n43767) );
  IV U54573 ( .A(n41643), .Z(n41644) );
  NOR U54574 ( .A(n41647), .B(n41644), .Z(n44884) );
  IV U54575 ( .A(n41645), .Z(n41646) );
  NOR U54576 ( .A(n41647), .B(n41646), .Z(n44890) );
  IV U54577 ( .A(n41651), .Z(n41659) );
  IV U54578 ( .A(n41650), .Z(n41648) );
  NOR U54579 ( .A(n41659), .B(n41648), .Z(n41656) );
  IV U54580 ( .A(n41649), .Z(n41654) );
  NOR U54581 ( .A(n41657), .B(n41650), .Z(n41652) );
  XOR U54582 ( .A(n41652), .B(n41651), .Z(n41653) );
  NOR U54583 ( .A(n41654), .B(n41653), .Z(n41655) );
  NOR U54584 ( .A(n41656), .B(n41655), .Z(n44894) );
  IV U54585 ( .A(n41657), .Z(n41658) );
  NOR U54586 ( .A(n41659), .B(n41658), .Z(n47025) );
  IV U54587 ( .A(n41660), .Z(n41661) );
  NOR U54588 ( .A(n41661), .B(n41663), .Z(n47022) );
  IV U54589 ( .A(n41662), .Z(n41664) );
  NOR U54590 ( .A(n41664), .B(n41663), .Z(n44895) );
  NOR U54591 ( .A(n41666), .B(n41665), .Z(n44902) );
  IV U54592 ( .A(n41667), .Z(n41668) );
  NOR U54593 ( .A(n41669), .B(n41668), .Z(n44911) );
  NOR U54594 ( .A(n41671), .B(n41670), .Z(n44906) );
  NOR U54595 ( .A(n44911), .B(n44906), .Z(n41672) );
  IV U54596 ( .A(n41672), .Z(n43765) );
  IV U54597 ( .A(n41673), .Z(n41675) );
  IV U54598 ( .A(n41674), .Z(n41677) );
  NOR U54599 ( .A(n41675), .B(n41677), .Z(n44908) );
  IV U54600 ( .A(n41676), .Z(n41678) );
  NOR U54601 ( .A(n41678), .B(n41677), .Z(n47016) );
  IV U54602 ( .A(n41679), .Z(n41680) );
  NOR U54603 ( .A(n41683), .B(n41680), .Z(n47013) );
  IV U54604 ( .A(n41681), .Z(n41682) );
  NOR U54605 ( .A(n41683), .B(n41682), .Z(n44917) );
  IV U54606 ( .A(n41684), .Z(n41685) );
  NOR U54607 ( .A(n41686), .B(n41685), .Z(n47003) );
  IV U54608 ( .A(n41687), .Z(n41688) );
  NOR U54609 ( .A(n41688), .B(n43756), .Z(n44920) );
  NOR U54610 ( .A(n47003), .B(n44920), .Z(n43754) );
  IV U54611 ( .A(n41689), .Z(n41692) );
  IV U54612 ( .A(n41690), .Z(n41691) );
  NOR U54613 ( .A(n41692), .B(n41691), .Z(n47000) );
  IV U54614 ( .A(n41693), .Z(n41694) );
  NOR U54615 ( .A(n41694), .B(n43738), .Z(n46996) );
  IV U54616 ( .A(n41695), .Z(n41696) );
  NOR U54617 ( .A(n43721), .B(n41696), .Z(n46984) );
  IV U54618 ( .A(n41697), .Z(n41698) );
  NOR U54619 ( .A(n41699), .B(n41698), .Z(n44944) );
  IV U54620 ( .A(n41700), .Z(n41702) );
  NOR U54621 ( .A(n41702), .B(n41701), .Z(n44938) );
  NOR U54622 ( .A(n44944), .B(n44938), .Z(n41703) );
  IV U54623 ( .A(n41703), .Z(n43718) );
  IV U54624 ( .A(n41704), .Z(n41708) );
  NOR U54625 ( .A(n41706), .B(n41705), .Z(n41707) );
  IV U54626 ( .A(n41707), .Z(n41710) );
  NOR U54627 ( .A(n41708), .B(n41710), .Z(n44941) );
  IV U54628 ( .A(n41709), .Z(n41711) );
  NOR U54629 ( .A(n41711), .B(n41710), .Z(n46979) );
  IV U54630 ( .A(n41712), .Z(n41714) );
  IV U54631 ( .A(n41713), .Z(n41716) );
  NOR U54632 ( .A(n41714), .B(n41716), .Z(n46976) );
  IV U54633 ( .A(n41715), .Z(n41717) );
  NOR U54634 ( .A(n41717), .B(n41716), .Z(n46972) );
  IV U54635 ( .A(n41718), .Z(n41719) );
  NOR U54636 ( .A(n41722), .B(n41719), .Z(n46969) );
  IV U54637 ( .A(n41720), .Z(n41721) );
  NOR U54638 ( .A(n41722), .B(n41721), .Z(n46965) );
  IV U54639 ( .A(n41723), .Z(n41725) );
  NOR U54640 ( .A(n41725), .B(n41724), .Z(n43707) );
  IV U54641 ( .A(n43707), .Z(n43702) );
  IV U54642 ( .A(n41726), .Z(n41728) );
  IV U54643 ( .A(n41727), .Z(n43690) );
  NOR U54644 ( .A(n41728), .B(n43690), .Z(n44947) );
  NOR U54645 ( .A(n41730), .B(n41729), .Z(n46918) );
  IV U54646 ( .A(n41731), .Z(n41734) );
  IV U54647 ( .A(n41732), .Z(n41733) );
  NOR U54648 ( .A(n41734), .B(n41733), .Z(n44951) );
  NOR U54649 ( .A(n46918), .B(n44951), .Z(n41735) );
  IV U54650 ( .A(n41735), .Z(n43688) );
  IV U54651 ( .A(n41736), .Z(n41737) );
  NOR U54652 ( .A(n41738), .B(n41737), .Z(n46896) );
  IV U54653 ( .A(n41739), .Z(n41740) );
  NOR U54654 ( .A(n41740), .B(n43676), .Z(n44955) );
  NOR U54655 ( .A(n46896), .B(n44955), .Z(n43674) );
  IV U54656 ( .A(n41741), .Z(n43667) );
  NOR U54657 ( .A(n41742), .B(n43667), .Z(n43665) );
  IV U54658 ( .A(n41743), .Z(n41746) );
  IV U54659 ( .A(n41744), .Z(n41745) );
  NOR U54660 ( .A(n41746), .B(n41745), .Z(n41747) );
  IV U54661 ( .A(n41747), .Z(n44958) );
  IV U54662 ( .A(n41748), .Z(n41750) );
  NOR U54663 ( .A(n41750), .B(n41749), .Z(n52135) );
  NOR U54664 ( .A(n41751), .B(n54159), .Z(n41752) );
  NOR U54665 ( .A(n52135), .B(n41752), .Z(n44971) );
  IV U54666 ( .A(n41753), .Z(n41754) );
  NOR U54667 ( .A(n41755), .B(n41754), .Z(n48426) );
  IV U54668 ( .A(n41756), .Z(n41757) );
  NOR U54669 ( .A(n41758), .B(n41757), .Z(n48421) );
  NOR U54670 ( .A(n48426), .B(n48421), .Z(n44969) );
  IV U54671 ( .A(n41759), .Z(n41761) );
  NOR U54672 ( .A(n41761), .B(n41760), .Z(n46859) );
  NOR U54673 ( .A(n41762), .B(n44974), .Z(n41763) );
  NOR U54674 ( .A(n46859), .B(n41763), .Z(n43633) );
  IV U54675 ( .A(n41764), .Z(n41765) );
  NOR U54676 ( .A(n43629), .B(n41765), .Z(n46856) );
  IV U54677 ( .A(n41766), .Z(n41767) );
  NOR U54678 ( .A(n41773), .B(n41767), .Z(n48450) );
  IV U54679 ( .A(n41768), .Z(n41770) );
  IV U54680 ( .A(n41769), .Z(n43631) );
  NOR U54681 ( .A(n41770), .B(n43631), .Z(n48444) );
  NOR U54682 ( .A(n48450), .B(n48444), .Z(n46850) );
  IV U54683 ( .A(n41771), .Z(n41772) );
  NOR U54684 ( .A(n41773), .B(n41772), .Z(n44977) );
  IV U54685 ( .A(n41774), .Z(n41776) );
  IV U54686 ( .A(n41775), .Z(n41779) );
  NOR U54687 ( .A(n41776), .B(n41779), .Z(n41777) );
  IV U54688 ( .A(n41777), .Z(n44991) );
  IV U54689 ( .A(n41778), .Z(n41780) );
  NOR U54690 ( .A(n41780), .B(n41779), .Z(n44993) );
  IV U54691 ( .A(n41781), .Z(n41782) );
  NOR U54692 ( .A(n41788), .B(n41782), .Z(n44996) );
  NOR U54693 ( .A(n44993), .B(n44996), .Z(n41783) );
  IV U54694 ( .A(n41783), .Z(n43617) );
  IV U54695 ( .A(n41784), .Z(n41785) );
  NOR U54696 ( .A(n41788), .B(n41785), .Z(n46838) );
  IV U54697 ( .A(n41786), .Z(n41787) );
  NOR U54698 ( .A(n41788), .B(n41787), .Z(n46825) );
  IV U54699 ( .A(n41789), .Z(n41791) );
  IV U54700 ( .A(n41790), .Z(n41795) );
  NOR U54701 ( .A(n41791), .B(n41795), .Z(n46822) );
  IV U54702 ( .A(n41792), .Z(n41793) );
  NOR U54703 ( .A(n41793), .B(n41798), .Z(n52204) );
  IV U54704 ( .A(n41794), .Z(n41796) );
  NOR U54705 ( .A(n41796), .B(n41795), .Z(n52192) );
  NOR U54706 ( .A(n52204), .B(n52192), .Z(n44998) );
  IV U54707 ( .A(n41797), .Z(n41799) );
  NOR U54708 ( .A(n41799), .B(n41798), .Z(n41800) );
  IV U54709 ( .A(n41800), .Z(n45006) );
  IV U54710 ( .A(n41801), .Z(n41802) );
  NOR U54711 ( .A(n41803), .B(n41802), .Z(n41804) );
  IV U54712 ( .A(n41804), .Z(n43612) );
  IV U54713 ( .A(n41805), .Z(n41806) );
  NOR U54714 ( .A(n41806), .B(n43603), .Z(n45007) );
  IV U54715 ( .A(n41807), .Z(n41808) );
  NOR U54716 ( .A(n41809), .B(n41808), .Z(n41810) );
  IV U54717 ( .A(n41810), .Z(n45022) );
  IV U54718 ( .A(n41811), .Z(n43582) );
  IV U54719 ( .A(n41812), .Z(n41813) );
  NOR U54720 ( .A(n43582), .B(n41813), .Z(n46812) );
  IV U54721 ( .A(n41814), .Z(n41815) );
  NOR U54722 ( .A(n41820), .B(n41815), .Z(n46809) );
  IV U54723 ( .A(n41816), .Z(n41817) );
  NOR U54724 ( .A(n41818), .B(n41817), .Z(n45037) );
  IV U54725 ( .A(n41819), .Z(n41821) );
  NOR U54726 ( .A(n41821), .B(n41820), .Z(n45031) );
  NOR U54727 ( .A(n45037), .B(n45031), .Z(n41822) );
  IV U54728 ( .A(n41822), .Z(n43580) );
  IV U54729 ( .A(n41823), .Z(n41826) );
  IV U54730 ( .A(n41824), .Z(n41825) );
  NOR U54731 ( .A(n41826), .B(n41825), .Z(n45035) );
  IV U54732 ( .A(n41827), .Z(n41831) );
  NOR U54733 ( .A(n41828), .B(n41836), .Z(n41829) );
  IV U54734 ( .A(n41829), .Z(n41830) );
  NOR U54735 ( .A(n41831), .B(n41830), .Z(n46803) );
  IV U54736 ( .A(n41832), .Z(n41834) );
  NOR U54737 ( .A(n41834), .B(n41833), .Z(n48507) );
  IV U54738 ( .A(n41835), .Z(n41840) );
  NOR U54739 ( .A(n41837), .B(n41836), .Z(n41838) );
  IV U54740 ( .A(n41838), .Z(n41839) );
  NOR U54741 ( .A(n41840), .B(n41839), .Z(n48497) );
  NOR U54742 ( .A(n48507), .B(n48497), .Z(n46802) );
  IV U54743 ( .A(n41841), .Z(n41842) );
  NOR U54744 ( .A(n41843), .B(n41842), .Z(n45044) );
  IV U54745 ( .A(n41844), .Z(n41846) );
  NOR U54746 ( .A(n41846), .B(n41845), .Z(n46797) );
  NOR U54747 ( .A(n45044), .B(n46797), .Z(n43579) );
  IV U54748 ( .A(n41847), .Z(n41849) );
  NOR U54749 ( .A(n41849), .B(n41848), .Z(n46793) );
  IV U54750 ( .A(n41850), .Z(n41851) );
  NOR U54751 ( .A(n41852), .B(n41851), .Z(n46790) );
  IV U54752 ( .A(n41853), .Z(n43547) );
  IV U54753 ( .A(n41854), .Z(n41855) );
  NOR U54754 ( .A(n43547), .B(n41855), .Z(n48543) );
  IV U54755 ( .A(n41856), .Z(n41858) );
  NOR U54756 ( .A(n41858), .B(n41857), .Z(n48536) );
  NOR U54757 ( .A(n48543), .B(n48536), .Z(n45058) );
  IV U54758 ( .A(n41859), .Z(n41860) );
  NOR U54759 ( .A(n41861), .B(n41860), .Z(n48546) );
  IV U54760 ( .A(n41862), .Z(n41864) );
  NOR U54761 ( .A(n41864), .B(n41863), .Z(n50213) );
  NOR U54762 ( .A(n48546), .B(n50213), .Z(n45066) );
  IV U54763 ( .A(n41865), .Z(n41867) );
  NOR U54764 ( .A(n41867), .B(n41866), .Z(n41868) );
  IV U54765 ( .A(n41868), .Z(n46759) );
  IV U54766 ( .A(n41869), .Z(n41870) );
  NOR U54767 ( .A(n41871), .B(n41870), .Z(n45070) );
  IV U54768 ( .A(n41872), .Z(n41873) );
  NOR U54769 ( .A(n41874), .B(n41873), .Z(n45067) );
  NOR U54770 ( .A(n45070), .B(n45067), .Z(n41875) );
  IV U54771 ( .A(n41875), .Z(n43532) );
  IV U54772 ( .A(n41876), .Z(n41879) );
  NOR U54773 ( .A(n43520), .B(n41877), .Z(n41878) );
  IV U54774 ( .A(n41878), .Z(n43516) );
  NOR U54775 ( .A(n41879), .B(n43516), .Z(n45073) );
  IV U54776 ( .A(n41880), .Z(n41881) );
  NOR U54777 ( .A(n41881), .B(n43507), .Z(n46727) );
  IV U54778 ( .A(n41882), .Z(n45078) );
  NOR U54779 ( .A(n45078), .B(n41883), .Z(n41885) );
  IV U54780 ( .A(n43508), .Z(n41884) );
  NOR U54781 ( .A(n43507), .B(n41884), .Z(n46724) );
  NOR U54782 ( .A(n41885), .B(n46724), .Z(n41886) );
  IV U54783 ( .A(n41886), .Z(n43505) );
  IV U54784 ( .A(n41887), .Z(n41890) );
  IV U54785 ( .A(n41888), .Z(n41889) );
  NOR U54786 ( .A(n41890), .B(n41889), .Z(n41891) );
  IV U54787 ( .A(n41891), .Z(n46718) );
  IV U54788 ( .A(n41892), .Z(n41893) );
  NOR U54789 ( .A(n41893), .B(n41898), .Z(n52363) );
  IV U54790 ( .A(n41894), .Z(n41896) );
  NOR U54791 ( .A(n41896), .B(n41895), .Z(n52355) );
  NOR U54792 ( .A(n52363), .B(n52355), .Z(n45094) );
  IV U54793 ( .A(n45094), .Z(n43495) );
  IV U54794 ( .A(n41897), .Z(n41899) );
  NOR U54795 ( .A(n41899), .B(n41898), .Z(n45096) );
  NOR U54796 ( .A(n41900), .B(n43490), .Z(n41901) );
  IV U54797 ( .A(n41901), .Z(n41904) );
  IV U54798 ( .A(n41902), .Z(n43489) );
  XOR U54799 ( .A(n41906), .B(n43489), .Z(n41903) );
  NOR U54800 ( .A(n41904), .B(n41903), .Z(n41905) );
  IV U54801 ( .A(n41905), .Z(n45106) );
  IV U54802 ( .A(n41906), .Z(n41907) );
  NOR U54803 ( .A(n41907), .B(n43489), .Z(n45108) );
  NOR U54804 ( .A(n45113), .B(n45108), .Z(n41908) );
  IV U54805 ( .A(n41908), .Z(n43484) );
  IV U54806 ( .A(n41909), .Z(n41910) );
  NOR U54807 ( .A(n41910), .B(n43475), .Z(n45120) );
  IV U54808 ( .A(n41911), .Z(n41913) );
  NOR U54809 ( .A(n41913), .B(n41912), .Z(n45117) );
  NOR U54810 ( .A(n45120), .B(n45117), .Z(n43477) );
  IV U54811 ( .A(n41914), .Z(n41915) );
  NOR U54812 ( .A(n41916), .B(n41915), .Z(n41917) );
  IV U54813 ( .A(n41917), .Z(n41918) );
  NOR U54814 ( .A(n41919), .B(n41918), .Z(n46694) );
  NOR U54815 ( .A(n41920), .B(n43469), .Z(n45127) );
  IV U54816 ( .A(n41921), .Z(n41922) );
  NOR U54817 ( .A(n41922), .B(n41924), .Z(n45124) );
  IV U54818 ( .A(n41923), .Z(n41925) );
  NOR U54819 ( .A(n41925), .B(n41924), .Z(n46689) );
  IV U54820 ( .A(n41926), .Z(n41927) );
  NOR U54821 ( .A(n41927), .B(n45142), .Z(n45137) );
  IV U54822 ( .A(n41928), .Z(n41929) );
  NOR U54823 ( .A(n41935), .B(n41929), .Z(n41930) );
  IV U54824 ( .A(n41930), .Z(n45148) );
  IV U54825 ( .A(n41931), .Z(n41932) );
  NOR U54826 ( .A(n41932), .B(n45142), .Z(n43457) );
  IV U54827 ( .A(n41933), .Z(n41934) );
  NOR U54828 ( .A(n41935), .B(n41934), .Z(n50128) );
  IV U54829 ( .A(n41936), .Z(n41939) );
  IV U54830 ( .A(n41937), .Z(n41938) );
  NOR U54831 ( .A(n41939), .B(n41938), .Z(n48637) );
  NOR U54832 ( .A(n50128), .B(n48637), .Z(n45153) );
  IV U54833 ( .A(n41940), .Z(n41943) );
  IV U54834 ( .A(n41941), .Z(n41942) );
  NOR U54835 ( .A(n41943), .B(n41942), .Z(n46679) );
  IV U54836 ( .A(n41944), .Z(n41945) );
  NOR U54837 ( .A(n41945), .B(n41947), .Z(n46676) );
  IV U54838 ( .A(n41946), .Z(n41948) );
  NOR U54839 ( .A(n41948), .B(n41947), .Z(n46665) );
  IV U54840 ( .A(n41949), .Z(n41954) );
  IV U54841 ( .A(n41950), .Z(n41951) );
  NOR U54842 ( .A(n41951), .B(n41956), .Z(n41952) );
  IV U54843 ( .A(n41952), .Z(n41953) );
  NOR U54844 ( .A(n41954), .B(n41953), .Z(n46661) );
  IV U54845 ( .A(n41955), .Z(n41960) );
  NOR U54846 ( .A(n41957), .B(n41956), .Z(n41958) );
  IV U54847 ( .A(n41958), .Z(n41959) );
  NOR U54848 ( .A(n41960), .B(n41959), .Z(n46668) );
  IV U54849 ( .A(n41961), .Z(n41966) );
  IV U54850 ( .A(n41962), .Z(n41963) );
  NOR U54851 ( .A(n41964), .B(n41963), .Z(n41965) );
  IV U54852 ( .A(n41965), .Z(n43453) );
  NOR U54853 ( .A(n41966), .B(n43453), .Z(n46657) );
  IV U54854 ( .A(n41967), .Z(n41974) );
  IV U54855 ( .A(n41968), .Z(n41969) );
  NOR U54856 ( .A(n41974), .B(n41969), .Z(n46642) );
  IV U54857 ( .A(n41970), .Z(n41971) );
  NOR U54858 ( .A(n41971), .B(n43438), .Z(n46627) );
  IV U54859 ( .A(n41972), .Z(n41973) );
  NOR U54860 ( .A(n41974), .B(n41973), .Z(n45166) );
  NOR U54861 ( .A(n46627), .B(n45166), .Z(n43440) );
  IV U54862 ( .A(n41975), .Z(n41978) );
  NOR U54863 ( .A(n41976), .B(n43428), .Z(n41977) );
  IV U54864 ( .A(n41977), .Z(n43431) );
  NOR U54865 ( .A(n41978), .B(n43431), .Z(n46624) );
  IV U54866 ( .A(n41979), .Z(n41984) );
  IV U54867 ( .A(n41980), .Z(n41981) );
  NOR U54868 ( .A(n41984), .B(n41981), .Z(n46621) );
  NOR U54869 ( .A(n46624), .B(n46621), .Z(n43426) );
  IV U54870 ( .A(n41982), .Z(n41983) );
  NOR U54871 ( .A(n41984), .B(n41983), .Z(n46618) );
  IV U54872 ( .A(n41985), .Z(n41987) );
  NOR U54873 ( .A(n41987), .B(n41986), .Z(n45176) );
  IV U54874 ( .A(n41988), .Z(n41991) );
  IV U54875 ( .A(n41989), .Z(n42001) );
  XOR U54876 ( .A(n41995), .B(n42001), .Z(n41990) );
  NOR U54877 ( .A(n41991), .B(n41990), .Z(n45180) );
  IV U54878 ( .A(n41992), .Z(n41993) );
  NOR U54879 ( .A(n42001), .B(n41993), .Z(n45183) );
  IV U54880 ( .A(n41994), .Z(n41999) );
  IV U54881 ( .A(n41995), .Z(n41996) );
  NOR U54882 ( .A(n42001), .B(n41996), .Z(n41997) );
  IV U54883 ( .A(n41997), .Z(n41998) );
  NOR U54884 ( .A(n41999), .B(n41998), .Z(n45186) );
  IV U54885 ( .A(n42000), .Z(n42005) );
  NOR U54886 ( .A(n42002), .B(n42001), .Z(n42003) );
  IV U54887 ( .A(n42003), .Z(n42004) );
  NOR U54888 ( .A(n42005), .B(n42004), .Z(n45192) );
  IV U54889 ( .A(n42006), .Z(n42007) );
  NOR U54890 ( .A(n42007), .B(n43415), .Z(n46613) );
  IV U54891 ( .A(n42008), .Z(n42009) );
  NOR U54892 ( .A(n42010), .B(n42009), .Z(n46610) );
  IV U54893 ( .A(n42011), .Z(n42012) );
  NOR U54894 ( .A(n42013), .B(n42012), .Z(n42014) );
  IV U54895 ( .A(n42014), .Z(n43421) );
  IV U54896 ( .A(n42015), .Z(n43419) );
  IV U54897 ( .A(n42016), .Z(n42017) );
  NOR U54898 ( .A(n43419), .B(n42017), .Z(n45205) );
  IV U54899 ( .A(n42018), .Z(n42019) );
  NOR U54900 ( .A(n42020), .B(n42019), .Z(n43395) );
  IV U54901 ( .A(n43395), .Z(n43390) );
  IV U54902 ( .A(n42021), .Z(n42022) );
  NOR U54903 ( .A(n42022), .B(n42024), .Z(n50044) );
  IV U54904 ( .A(n42023), .Z(n42027) );
  NOR U54905 ( .A(n42025), .B(n42024), .Z(n42026) );
  IV U54906 ( .A(n42026), .Z(n43392) );
  NOR U54907 ( .A(n42027), .B(n43392), .Z(n50049) );
  NOR U54908 ( .A(n50044), .B(n50049), .Z(n45215) );
  IV U54909 ( .A(n42028), .Z(n42030) );
  IV U54910 ( .A(n42029), .Z(n42033) );
  NOR U54911 ( .A(n42030), .B(n42033), .Z(n46597) );
  NOR U54912 ( .A(n42031), .B(n48713), .Z(n45216) );
  NOR U54913 ( .A(n46597), .B(n45216), .Z(n43389) );
  IV U54914 ( .A(n42032), .Z(n42034) );
  NOR U54915 ( .A(n42034), .B(n42033), .Z(n46590) );
  IV U54916 ( .A(n42035), .Z(n42036) );
  NOR U54917 ( .A(n42037), .B(n42036), .Z(n52494) );
  IV U54918 ( .A(n42038), .Z(n42039) );
  NOR U54919 ( .A(n42039), .B(n43377), .Z(n53920) );
  NOR U54920 ( .A(n52494), .B(n53920), .Z(n49992) );
  IV U54921 ( .A(n42040), .Z(n42043) );
  IV U54922 ( .A(n42041), .Z(n42042) );
  NOR U54923 ( .A(n42043), .B(n42042), .Z(n46569) );
  IV U54924 ( .A(n42044), .Z(n42046) );
  IV U54925 ( .A(n42045), .Z(n42051) );
  NOR U54926 ( .A(n42046), .B(n42051), .Z(n42047) );
  IV U54927 ( .A(n42047), .Z(n45226) );
  IV U54928 ( .A(n42048), .Z(n42049) );
  NOR U54929 ( .A(n42049), .B(n42055), .Z(n46547) );
  IV U54930 ( .A(n42050), .Z(n42052) );
  NOR U54931 ( .A(n42052), .B(n42051), .Z(n45228) );
  NOR U54932 ( .A(n46547), .B(n45228), .Z(n42053) );
  IV U54933 ( .A(n42053), .Z(n43368) );
  IV U54934 ( .A(n42054), .Z(n42056) );
  NOR U54935 ( .A(n42056), .B(n42055), .Z(n45230) );
  NOR U54936 ( .A(n42058), .B(n42057), .Z(n48749) );
  IV U54937 ( .A(n42059), .Z(n43363) );
  IV U54938 ( .A(n42060), .Z(n42061) );
  NOR U54939 ( .A(n43363), .B(n42061), .Z(n48754) );
  NOR U54940 ( .A(n48749), .B(n48754), .Z(n45237) );
  IV U54941 ( .A(n42062), .Z(n42064) );
  IV U54942 ( .A(n42063), .Z(n42067) );
  NOR U54943 ( .A(n42064), .B(n42067), .Z(n45240) );
  IV U54944 ( .A(n42065), .Z(n42066) );
  NOR U54945 ( .A(n42067), .B(n42066), .Z(n45246) );
  IV U54946 ( .A(n42068), .Z(n42071) );
  IV U54947 ( .A(n42069), .Z(n42070) );
  NOR U54948 ( .A(n42071), .B(n42070), .Z(n46538) );
  NOR U54949 ( .A(n42073), .B(n42072), .Z(n49972) );
  NOR U54950 ( .A(n49972), .B(n48770), .Z(n46537) );
  IV U54951 ( .A(n46537), .Z(n43355) );
  IV U54952 ( .A(n42074), .Z(n42078) );
  IV U54953 ( .A(n42075), .Z(n42084) );
  NOR U54954 ( .A(n42084), .B(n42076), .Z(n42077) );
  IV U54955 ( .A(n42077), .Z(n42080) );
  NOR U54956 ( .A(n42078), .B(n42080), .Z(n45252) );
  IV U54957 ( .A(n42079), .Z(n42081) );
  NOR U54958 ( .A(n42081), .B(n42080), .Z(n45249) );
  IV U54959 ( .A(n42082), .Z(n42083) );
  NOR U54960 ( .A(n42084), .B(n42083), .Z(n45255) );
  IV U54961 ( .A(n42085), .Z(n42088) );
  NOR U54962 ( .A(n42086), .B(n43345), .Z(n42087) );
  IV U54963 ( .A(n42087), .Z(n43352) );
  NOR U54964 ( .A(n42088), .B(n43352), .Z(n42089) );
  IV U54965 ( .A(n42089), .Z(n42090) );
  NOR U54966 ( .A(n42091), .B(n42090), .Z(n43348) );
  IV U54967 ( .A(n42092), .Z(n42093) );
  NOR U54968 ( .A(n43338), .B(n42093), .Z(n42094) );
  IV U54969 ( .A(n42094), .Z(n42095) );
  NOR U54970 ( .A(n42096), .B(n42095), .Z(n42097) );
  IV U54971 ( .A(n42097), .Z(n46523) );
  IV U54972 ( .A(n42098), .Z(n42099) );
  NOR U54973 ( .A(n42100), .B(n42099), .Z(n46516) );
  IV U54974 ( .A(n42101), .Z(n42111) );
  NOR U54975 ( .A(n42111), .B(n42102), .Z(n42103) );
  IV U54976 ( .A(n42103), .Z(n42107) );
  NOR U54977 ( .A(n43333), .B(n42104), .Z(n42105) );
  IV U54978 ( .A(n42105), .Z(n42106) );
  NOR U54979 ( .A(n42107), .B(n42106), .Z(n45263) );
  NOR U54980 ( .A(n42109), .B(n42108), .Z(n46511) );
  IV U54981 ( .A(n42110), .Z(n42112) );
  NOR U54982 ( .A(n42112), .B(n42111), .Z(n45266) );
  NOR U54983 ( .A(n46511), .B(n45266), .Z(n42113) );
  IV U54984 ( .A(n42113), .Z(n43331) );
  IV U54985 ( .A(n42114), .Z(n42116) );
  NOR U54986 ( .A(n42116), .B(n42115), .Z(n45271) );
  IV U54987 ( .A(n42117), .Z(n42118) );
  NOR U54988 ( .A(n42118), .B(n42120), .Z(n45268) );
  IV U54989 ( .A(n42119), .Z(n42121) );
  NOR U54990 ( .A(n42121), .B(n42120), .Z(n45274) );
  NOR U54991 ( .A(n42122), .B(n48815), .Z(n42126) );
  IV U54992 ( .A(n42123), .Z(n42125) );
  IV U54993 ( .A(n42124), .Z(n43309) );
  NOR U54994 ( .A(n42125), .B(n43309), .Z(n48797) );
  NOR U54995 ( .A(n42126), .B(n48797), .Z(n45287) );
  IV U54996 ( .A(n45287), .Z(n43306) );
  IV U54997 ( .A(n42127), .Z(n42132) );
  IV U54998 ( .A(n42128), .Z(n42129) );
  NOR U54999 ( .A(n43295), .B(n42129), .Z(n42130) );
  IV U55000 ( .A(n42130), .Z(n42131) );
  NOR U55001 ( .A(n42132), .B(n42131), .Z(n45284) );
  IV U55002 ( .A(n42133), .Z(n42134) );
  NOR U55003 ( .A(n42134), .B(n42140), .Z(n46476) );
  IV U55004 ( .A(n42135), .Z(n42137) );
  NOR U55005 ( .A(n42137), .B(n42136), .Z(n45297) );
  IV U55006 ( .A(n42138), .Z(n42139) );
  NOR U55007 ( .A(n42140), .B(n42139), .Z(n46479) );
  NOR U55008 ( .A(n45297), .B(n46479), .Z(n43280) );
  IV U55009 ( .A(n42141), .Z(n42143) );
  IV U55010 ( .A(n42142), .Z(n43277) );
  NOR U55011 ( .A(n42143), .B(n43277), .Z(n46469) );
  IV U55012 ( .A(n42144), .Z(n42145) );
  NOR U55013 ( .A(n42148), .B(n42145), .Z(n45302) );
  IV U55014 ( .A(n42146), .Z(n42147) );
  NOR U55015 ( .A(n42148), .B(n42147), .Z(n45305) );
  IV U55016 ( .A(n42149), .Z(n42153) );
  IV U55017 ( .A(n42150), .Z(n42159) );
  NOR U55018 ( .A(n42151), .B(n42159), .Z(n42152) );
  IV U55019 ( .A(n42152), .Z(n42156) );
  NOR U55020 ( .A(n42153), .B(n42156), .Z(n45300) );
  NOR U55021 ( .A(n45305), .B(n45300), .Z(n42154) );
  IV U55022 ( .A(n42154), .Z(n43272) );
  IV U55023 ( .A(n42155), .Z(n42157) );
  NOR U55024 ( .A(n42157), .B(n42156), .Z(n45311) );
  IV U55025 ( .A(n42158), .Z(n42162) );
  NOR U55026 ( .A(n42160), .B(n42159), .Z(n42161) );
  IV U55027 ( .A(n42161), .Z(n42164) );
  NOR U55028 ( .A(n42162), .B(n42164), .Z(n45308) );
  IV U55029 ( .A(n42163), .Z(n42165) );
  NOR U55030 ( .A(n42165), .B(n42164), .Z(n46462) );
  IV U55031 ( .A(n42166), .Z(n42167) );
  NOR U55032 ( .A(n42167), .B(n42169), .Z(n46459) );
  IV U55033 ( .A(n42168), .Z(n42170) );
  NOR U55034 ( .A(n42170), .B(n42169), .Z(n45314) );
  IV U55035 ( .A(n42171), .Z(n48857) );
  IV U55036 ( .A(n42172), .Z(n42173) );
  NOR U55037 ( .A(n48857), .B(n42173), .Z(n42174) );
  IV U55038 ( .A(n42174), .Z(n45326) );
  NOR U55039 ( .A(n42175), .B(n48857), .Z(n45323) );
  IV U55040 ( .A(n42176), .Z(n42178) );
  IV U55041 ( .A(n42177), .Z(n42184) );
  NOR U55042 ( .A(n42178), .B(n42184), .Z(n46451) );
  NOR U55043 ( .A(n42180), .B(n42179), .Z(n46455) );
  NOR U55044 ( .A(n46451), .B(n46455), .Z(n42181) );
  IV U55045 ( .A(n42181), .Z(n43264) );
  IV U55046 ( .A(n42182), .Z(n42183) );
  NOR U55047 ( .A(n42184), .B(n42183), .Z(n46449) );
  IV U55048 ( .A(n42185), .Z(n42186) );
  NOR U55049 ( .A(n42187), .B(n42186), .Z(n42188) );
  IV U55050 ( .A(n42188), .Z(n45329) );
  IV U55051 ( .A(n42189), .Z(n42190) );
  NOR U55052 ( .A(n43251), .B(n42190), .Z(n45344) );
  IV U55053 ( .A(n42191), .Z(n42193) );
  IV U55054 ( .A(n42192), .Z(n42195) );
  NOR U55055 ( .A(n42193), .B(n42195), .Z(n46438) );
  NOR U55056 ( .A(n45344), .B(n46438), .Z(n43247) );
  IV U55057 ( .A(n42194), .Z(n42196) );
  NOR U55058 ( .A(n42196), .B(n42195), .Z(n46435) );
  IV U55059 ( .A(n42197), .Z(n42198) );
  NOR U55060 ( .A(n42198), .B(n43244), .Z(n45346) );
  IV U55061 ( .A(n42199), .Z(n42204) );
  IV U55062 ( .A(n42200), .Z(n42201) );
  NOR U55063 ( .A(n42201), .B(n43223), .Z(n42202) );
  IV U55064 ( .A(n42202), .Z(n42203) );
  NOR U55065 ( .A(n42204), .B(n42203), .Z(n46418) );
  IV U55066 ( .A(n42205), .Z(n42206) );
  NOR U55067 ( .A(n42206), .B(n42211), .Z(n42207) );
  IV U55068 ( .A(n42207), .Z(n42208) );
  NOR U55069 ( .A(n42215), .B(n42208), .Z(n42209) );
  IV U55070 ( .A(n42209), .Z(n45362) );
  IV U55071 ( .A(n42210), .Z(n42212) );
  NOR U55072 ( .A(n42212), .B(n42211), .Z(n42213) );
  IV U55073 ( .A(n42213), .Z(n42214) );
  NOR U55074 ( .A(n42215), .B(n42214), .Z(n45366) );
  IV U55075 ( .A(n42216), .Z(n42217) );
  NOR U55076 ( .A(n42217), .B(n43215), .Z(n45369) );
  IV U55077 ( .A(n42218), .Z(n42219) );
  NOR U55078 ( .A(n42220), .B(n42219), .Z(n45377) );
  NOR U55079 ( .A(n42221), .B(n46401), .Z(n42224) );
  IV U55080 ( .A(n42222), .Z(n45381) );
  NOR U55081 ( .A(n45383), .B(n45381), .Z(n42223) );
  NOR U55082 ( .A(n42224), .B(n42223), .Z(n42225) );
  IV U55083 ( .A(n42225), .Z(n43212) );
  IV U55084 ( .A(n42226), .Z(n42230) );
  NOR U55085 ( .A(n42228), .B(n42227), .Z(n42229) );
  IV U55086 ( .A(n42229), .Z(n42232) );
  NOR U55087 ( .A(n42230), .B(n42232), .Z(n46396) );
  IV U55088 ( .A(n42231), .Z(n42233) );
  NOR U55089 ( .A(n42233), .B(n42232), .Z(n45384) );
  IV U55090 ( .A(n42234), .Z(n43207) );
  IV U55091 ( .A(n42235), .Z(n42236) );
  NOR U55092 ( .A(n42236), .B(n42241), .Z(n46381) );
  IV U55093 ( .A(n42237), .Z(n42238) );
  NOR U55094 ( .A(n42239), .B(n42238), .Z(n45392) );
  IV U55095 ( .A(n42240), .Z(n42242) );
  NOR U55096 ( .A(n42242), .B(n42241), .Z(n46384) );
  NOR U55097 ( .A(n45392), .B(n46384), .Z(n43199) );
  IV U55098 ( .A(n42243), .Z(n42244) );
  NOR U55099 ( .A(n42245), .B(n42244), .Z(n45397) );
  IV U55100 ( .A(n42246), .Z(n42247) );
  NOR U55101 ( .A(n42248), .B(n42247), .Z(n45394) );
  NOR U55102 ( .A(n45397), .B(n45394), .Z(n43198) );
  IV U55103 ( .A(n42249), .Z(n42252) );
  IV U55104 ( .A(n42250), .Z(n42251) );
  NOR U55105 ( .A(n42252), .B(n42251), .Z(n42253) );
  IV U55106 ( .A(n42253), .Z(n46376) );
  IV U55107 ( .A(n42254), .Z(n42255) );
  NOR U55108 ( .A(n45413), .B(n42255), .Z(n46359) );
  NOR U55109 ( .A(n42256), .B(n42257), .Z(n42262) );
  IV U55110 ( .A(n42257), .Z(n42258) );
  NOR U55111 ( .A(n42259), .B(n42258), .Z(n45418) );
  NOR U55112 ( .A(n42260), .B(n45418), .Z(n42261) );
  NOR U55113 ( .A(n42262), .B(n42261), .Z(n45408) );
  IV U55114 ( .A(n42263), .Z(n42266) );
  IV U55115 ( .A(n42264), .Z(n42265) );
  NOR U55116 ( .A(n42266), .B(n42265), .Z(n45415) );
  NOR U55117 ( .A(n42268), .B(n42267), .Z(n46351) );
  IV U55118 ( .A(n42269), .Z(n42272) );
  IV U55119 ( .A(n42270), .Z(n42271) );
  NOR U55120 ( .A(n42272), .B(n42271), .Z(n45420) );
  IV U55121 ( .A(n42273), .Z(n42274) );
  XOR U55122 ( .A(n42277), .B(n42278), .Z(n45425) );
  NOR U55123 ( .A(n42274), .B(n45425), .Z(n43169) );
  IV U55124 ( .A(n42275), .Z(n42276) );
  NOR U55125 ( .A(n42276), .B(n42278), .Z(n46344) );
  IV U55126 ( .A(n42277), .Z(n42279) );
  NOR U55127 ( .A(n42279), .B(n42278), .Z(n46341) );
  IV U55128 ( .A(n42280), .Z(n43164) );
  IV U55129 ( .A(n42281), .Z(n42282) );
  NOR U55130 ( .A(n43164), .B(n42282), .Z(n46337) );
  IV U55131 ( .A(n42283), .Z(n42285) );
  NOR U55132 ( .A(n42285), .B(n42284), .Z(n43158) );
  IV U55133 ( .A(n43158), .Z(n43152) );
  IV U55134 ( .A(n42286), .Z(n42289) );
  IV U55135 ( .A(n42287), .Z(n42288) );
  NOR U55136 ( .A(n42289), .B(n42288), .Z(n45436) );
  IV U55137 ( .A(n42290), .Z(n42291) );
  NOR U55138 ( .A(n42292), .B(n42291), .Z(n42293) );
  IV U55139 ( .A(n42293), .Z(n46320) );
  IV U55140 ( .A(n42294), .Z(n42305) );
  IV U55141 ( .A(n42295), .Z(n42296) );
  NOR U55142 ( .A(n42305), .B(n42296), .Z(n46316) );
  IV U55143 ( .A(n42297), .Z(n42298) );
  NOR U55144 ( .A(n42300), .B(n42298), .Z(n49704) );
  IV U55145 ( .A(n42299), .Z(n42301) );
  NOR U55146 ( .A(n42301), .B(n42300), .Z(n49711) );
  NOR U55147 ( .A(n49704), .B(n49711), .Z(n42302) );
  IV U55148 ( .A(n42302), .Z(n46309) );
  IV U55149 ( .A(n42303), .Z(n42304) );
  NOR U55150 ( .A(n42305), .B(n42304), .Z(n46313) );
  NOR U55151 ( .A(n46309), .B(n46313), .Z(n42306) );
  IV U55152 ( .A(n42306), .Z(n43140) );
  IV U55153 ( .A(n42307), .Z(n42308) );
  NOR U55154 ( .A(n42309), .B(n42308), .Z(n46306) );
  IV U55155 ( .A(n42310), .Z(n45445) );
  NOR U55156 ( .A(n42311), .B(n45445), .Z(n42314) );
  IV U55157 ( .A(n42312), .Z(n42313) );
  NOR U55158 ( .A(n42325), .B(n42313), .Z(n46299) );
  NOR U55159 ( .A(n42314), .B(n46299), .Z(n43139) );
  IV U55160 ( .A(n42324), .Z(n42319) );
  NOR U55161 ( .A(n42316), .B(n42315), .Z(n42317) );
  IV U55162 ( .A(n42317), .Z(n42318) );
  NOR U55163 ( .A(n42319), .B(n42318), .Z(n46282) );
  IV U55164 ( .A(n46282), .Z(n42320) );
  NOR U55165 ( .A(n42325), .B(n42320), .Z(n46287) );
  XOR U55166 ( .A(n42322), .B(n42321), .Z(n42323) );
  NOR U55167 ( .A(n42324), .B(n42323), .Z(n42326) );
  NOR U55168 ( .A(n42326), .B(n42325), .Z(n42327) );
  IV U55169 ( .A(n42327), .Z(n42333) );
  IV U55170 ( .A(n42328), .Z(n42330) );
  NOR U55171 ( .A(n42330), .B(n42329), .Z(n42331) );
  IV U55172 ( .A(n42331), .Z(n42332) );
  NOR U55173 ( .A(n42333), .B(n42332), .Z(n46280) );
  NOR U55174 ( .A(n46287), .B(n46280), .Z(n42334) );
  IV U55175 ( .A(n42334), .Z(n43138) );
  IV U55176 ( .A(n42335), .Z(n43130) );
  IV U55177 ( .A(n42336), .Z(n43125) );
  IV U55178 ( .A(n42337), .Z(n42338) );
  NOR U55179 ( .A(n42338), .B(n45455), .Z(n45448) );
  IV U55180 ( .A(n42340), .Z(n45465) );
  IV U55181 ( .A(n42342), .Z(n42344) );
  NOR U55182 ( .A(n42344), .B(n42343), .Z(n45477) );
  NOR U55183 ( .A(n42346), .B(n42345), .Z(n45473) );
  NOR U55184 ( .A(n45477), .B(n45473), .Z(n43124) );
  NOR U55185 ( .A(n42347), .B(n45483), .Z(n43117) );
  IV U55186 ( .A(n42348), .Z(n43101) );
  IV U55187 ( .A(n42349), .Z(n42350) );
  NOR U55188 ( .A(n43101), .B(n42350), .Z(n45498) );
  IV U55189 ( .A(n42351), .Z(n42353) );
  NOR U55190 ( .A(n42353), .B(n42352), .Z(n45507) );
  IV U55191 ( .A(n42354), .Z(n42355) );
  NOR U55192 ( .A(n42355), .B(n43097), .Z(n45504) );
  NOR U55193 ( .A(n45507), .B(n45504), .Z(n43095) );
  IV U55194 ( .A(n42356), .Z(n42358) );
  NOR U55195 ( .A(n42358), .B(n42357), .Z(n49019) );
  NOR U55196 ( .A(n49023), .B(n49019), .Z(n45506) );
  IV U55197 ( .A(n42359), .Z(n42360) );
  NOR U55198 ( .A(n42360), .B(n42363), .Z(n42361) );
  IV U55199 ( .A(n42361), .Z(n45513) );
  IV U55200 ( .A(n42362), .Z(n42364) );
  NOR U55201 ( .A(n42364), .B(n42363), .Z(n43091) );
  IV U55202 ( .A(n42365), .Z(n42368) );
  IV U55203 ( .A(n42366), .Z(n42367) );
  NOR U55204 ( .A(n42368), .B(n42367), .Z(n45523) );
  IV U55205 ( .A(n42369), .Z(n42374) );
  XOR U55206 ( .A(n42370), .B(n43073), .Z(n42371) );
  NOR U55207 ( .A(n42372), .B(n42371), .Z(n42373) );
  IV U55208 ( .A(n42373), .Z(n43081) );
  NOR U55209 ( .A(n42374), .B(n43081), .Z(n45520) );
  IV U55210 ( .A(n42375), .Z(n42381) );
  NOR U55211 ( .A(n42376), .B(n43052), .Z(n42377) );
  IV U55212 ( .A(n42377), .Z(n42378) );
  NOR U55213 ( .A(n42379), .B(n42378), .Z(n42380) );
  IV U55214 ( .A(n42380), .Z(n43049) );
  NOR U55215 ( .A(n42381), .B(n43049), .Z(n46244) );
  IV U55216 ( .A(n42382), .Z(n42384) );
  NOR U55217 ( .A(n42384), .B(n42383), .Z(n45547) );
  IV U55218 ( .A(n42385), .Z(n42387) );
  NOR U55219 ( .A(n42387), .B(n42386), .Z(n45543) );
  NOR U55220 ( .A(n45547), .B(n45543), .Z(n43047) );
  IV U55221 ( .A(n42388), .Z(n42389) );
  NOR U55222 ( .A(n42389), .B(n43035), .Z(n43033) );
  IV U55223 ( .A(n42390), .Z(n42392) );
  NOR U55224 ( .A(n42392), .B(n42391), .Z(n42393) );
  IV U55225 ( .A(n42393), .Z(n46240) );
  IV U55226 ( .A(n42394), .Z(n42396) );
  XOR U55227 ( .A(n42397), .B(n42400), .Z(n42395) );
  NOR U55228 ( .A(n42396), .B(n42395), .Z(n46208) );
  IV U55229 ( .A(n42397), .Z(n42398) );
  NOR U55230 ( .A(n42400), .B(n42398), .Z(n46200) );
  IV U55231 ( .A(n42399), .Z(n42401) );
  NOR U55232 ( .A(n42401), .B(n42400), .Z(n46198) );
  IV U55233 ( .A(n42402), .Z(n45562) );
  NOR U55234 ( .A(n45562), .B(n42403), .Z(n42404) );
  NOR U55235 ( .A(n46198), .B(n42404), .Z(n42405) );
  IV U55236 ( .A(n42405), .Z(n42406) );
  NOR U55237 ( .A(n46200), .B(n42406), .Z(n42407) );
  IV U55238 ( .A(n42407), .Z(n43017) );
  IV U55239 ( .A(n42408), .Z(n42411) );
  NOR U55240 ( .A(n42409), .B(n42416), .Z(n42410) );
  IV U55241 ( .A(n42410), .Z(n42413) );
  NOR U55242 ( .A(n42411), .B(n42413), .Z(n45568) );
  IV U55243 ( .A(n42412), .Z(n42414) );
  NOR U55244 ( .A(n42414), .B(n42413), .Z(n45565) );
  IV U55245 ( .A(n42415), .Z(n42417) );
  NOR U55246 ( .A(n42417), .B(n42416), .Z(n43012) );
  IV U55247 ( .A(n42418), .Z(n42423) );
  IV U55248 ( .A(n42419), .Z(n42995) );
  XOR U55249 ( .A(n42988), .B(n42995), .Z(n42420) );
  NOR U55250 ( .A(n42421), .B(n42420), .Z(n42422) );
  IV U55251 ( .A(n42422), .Z(n43002) );
  NOR U55252 ( .A(n42423), .B(n43002), .Z(n46186) );
  IV U55253 ( .A(n42424), .Z(n42430) );
  IV U55254 ( .A(n42425), .Z(n42426) );
  NOR U55255 ( .A(n42427), .B(n42426), .Z(n42428) );
  IV U55256 ( .A(n42428), .Z(n42429) );
  NOR U55257 ( .A(n42430), .B(n42429), .Z(n45587) );
  IV U55258 ( .A(n42431), .Z(n42432) );
  NOR U55259 ( .A(n42433), .B(n42432), .Z(n45595) );
  NOR U55260 ( .A(n45595), .B(n45590), .Z(n42434) );
  IV U55261 ( .A(n42434), .Z(n42986) );
  IV U55262 ( .A(n42435), .Z(n42436) );
  NOR U55263 ( .A(n42437), .B(n42436), .Z(n45592) );
  IV U55264 ( .A(n42438), .Z(n46172) );
  IV U55265 ( .A(n42439), .Z(n42443) );
  NOR U55266 ( .A(n42441), .B(n42440), .Z(n42442) );
  IV U55267 ( .A(n42442), .Z(n42447) );
  NOR U55268 ( .A(n42443), .B(n42447), .Z(n46155) );
  XOR U55269 ( .A(n46154), .B(n46155), .Z(n42444) );
  NOR U55270 ( .A(n46168), .B(n42444), .Z(n42445) );
  IV U55271 ( .A(n42445), .Z(n42979) );
  IV U55272 ( .A(n42446), .Z(n42448) );
  NOR U55273 ( .A(n42448), .B(n42447), .Z(n45598) );
  IV U55274 ( .A(n42449), .Z(n42451) );
  IV U55275 ( .A(n42450), .Z(n42976) );
  NOR U55276 ( .A(n42451), .B(n42976), .Z(n45602) );
  IV U55277 ( .A(n42452), .Z(n42453) );
  NOR U55278 ( .A(n42953), .B(n42453), .Z(n45622) );
  IV U55279 ( .A(n45622), .Z(n45620) );
  IV U55280 ( .A(n42454), .Z(n42455) );
  NOR U55281 ( .A(n42456), .B(n42455), .Z(n46135) );
  IV U55282 ( .A(n42457), .Z(n42458) );
  NOR U55283 ( .A(n42459), .B(n42458), .Z(n42460) );
  IV U55284 ( .A(n42460), .Z(n42461) );
  NOR U55285 ( .A(n42461), .B(n42946), .Z(n46138) );
  NOR U55286 ( .A(n46135), .B(n46138), .Z(n42944) );
  IV U55287 ( .A(n42462), .Z(n42935) );
  IV U55288 ( .A(n42463), .Z(n42464) );
  NOR U55289 ( .A(n42935), .B(n42464), .Z(n46132) );
  IV U55290 ( .A(n42465), .Z(n42467) );
  IV U55291 ( .A(n42466), .Z(n42931) );
  NOR U55292 ( .A(n42467), .B(n42931), .Z(n42468) );
  IV U55293 ( .A(n42468), .Z(n46117) );
  IV U55294 ( .A(n42469), .Z(n42470) );
  NOR U55295 ( .A(n42470), .B(n42931), .Z(n46107) );
  IV U55296 ( .A(n42471), .Z(n42474) );
  NOR U55297 ( .A(n42476), .B(n42472), .Z(n42473) );
  IV U55298 ( .A(n42473), .Z(n42928) );
  NOR U55299 ( .A(n42474), .B(n42928), .Z(n46099) );
  IV U55300 ( .A(n42475), .Z(n49136) );
  NOR U55301 ( .A(n42476), .B(n49136), .Z(n46096) );
  IV U55302 ( .A(n42477), .Z(n42478) );
  NOR U55303 ( .A(n42909), .B(n42478), .Z(n46077) );
  IV U55304 ( .A(n42479), .Z(n42480) );
  NOR U55305 ( .A(n42481), .B(n42480), .Z(n45652) );
  IV U55306 ( .A(n42482), .Z(n42484) );
  NOR U55307 ( .A(n42484), .B(n42483), .Z(n45648) );
  NOR U55308 ( .A(n45652), .B(n45648), .Z(n42896) );
  NOR U55309 ( .A(n42485), .B(n42492), .Z(n46069) );
  IV U55310 ( .A(n42486), .Z(n42487) );
  NOR U55311 ( .A(n42487), .B(n42492), .Z(n46066) );
  IV U55312 ( .A(n42488), .Z(n42490) );
  NOR U55313 ( .A(n42490), .B(n42489), .Z(n45659) );
  IV U55314 ( .A(n42491), .Z(n42493) );
  NOR U55315 ( .A(n42493), .B(n42492), .Z(n45656) );
  NOR U55316 ( .A(n45659), .B(n45656), .Z(n42895) );
  IV U55317 ( .A(n42494), .Z(n42495) );
  NOR U55318 ( .A(n42496), .B(n42495), .Z(n46061) );
  IV U55319 ( .A(n42497), .Z(n42499) );
  NOR U55320 ( .A(n42499), .B(n42498), .Z(n45662) );
  NOR U55321 ( .A(n46061), .B(n45662), .Z(n42894) );
  IV U55322 ( .A(n42500), .Z(n42502) );
  NOR U55323 ( .A(n42502), .B(n42501), .Z(n46058) );
  IV U55324 ( .A(n42503), .Z(n42504) );
  NOR U55325 ( .A(n42504), .B(n42891), .Z(n45668) );
  IV U55326 ( .A(n42505), .Z(n46048) );
  IV U55327 ( .A(n42506), .Z(n42510) );
  IV U55328 ( .A(n42507), .Z(n42518) );
  NOR U55329 ( .A(n42508), .B(n42518), .Z(n42509) );
  IV U55330 ( .A(n42509), .Z(n42879) );
  NOR U55331 ( .A(n42510), .B(n42879), .Z(n45671) );
  IV U55332 ( .A(n42511), .Z(n42512) );
  NOR U55333 ( .A(n42512), .B(n42514), .Z(n45675) );
  IV U55334 ( .A(n42513), .Z(n42515) );
  NOR U55335 ( .A(n42515), .B(n42514), .Z(n45677) );
  NOR U55336 ( .A(n45675), .B(n45677), .Z(n42516) );
  IV U55337 ( .A(n42516), .Z(n42520) );
  IV U55338 ( .A(n42517), .Z(n42519) );
  NOR U55339 ( .A(n42519), .B(n42518), .Z(n46026) );
  NOR U55340 ( .A(n42520), .B(n46026), .Z(n42521) );
  IV U55341 ( .A(n42521), .Z(n42876) );
  IV U55342 ( .A(n42522), .Z(n42524) );
  IV U55343 ( .A(n42523), .Z(n42530) );
  NOR U55344 ( .A(n42524), .B(n42530), .Z(n45682) );
  IV U55345 ( .A(n42525), .Z(n42527) );
  NOR U55346 ( .A(n42527), .B(n42526), .Z(n45680) );
  NOR U55347 ( .A(n45682), .B(n45680), .Z(n42875) );
  IV U55348 ( .A(n42531), .Z(n42528) );
  NOR U55349 ( .A(n42528), .B(n42530), .Z(n46012) );
  IV U55350 ( .A(n42529), .Z(n42533) );
  XOR U55351 ( .A(n42531), .B(n42530), .Z(n42532) );
  NOR U55352 ( .A(n42533), .B(n42532), .Z(n46022) );
  NOR U55353 ( .A(n46012), .B(n46022), .Z(n42874) );
  IV U55354 ( .A(n42534), .Z(n42535) );
  NOR U55355 ( .A(n42535), .B(n42540), .Z(n45685) );
  IV U55356 ( .A(n42536), .Z(n42538) );
  NOR U55357 ( .A(n42538), .B(n42537), .Z(n45689) );
  IV U55358 ( .A(n42539), .Z(n42541) );
  NOR U55359 ( .A(n42541), .B(n42540), .Z(n46014) );
  NOR U55360 ( .A(n45689), .B(n46014), .Z(n42872) );
  IV U55361 ( .A(n42542), .Z(n42550) );
  IV U55362 ( .A(n42543), .Z(n42544) );
  NOR U55363 ( .A(n42550), .B(n42544), .Z(n46005) );
  IV U55364 ( .A(n42545), .Z(n42547) );
  NOR U55365 ( .A(n42547), .B(n42546), .Z(n46009) );
  NOR U55366 ( .A(n46005), .B(n46009), .Z(n42871) );
  IV U55367 ( .A(n42548), .Z(n42549) );
  NOR U55368 ( .A(n42550), .B(n42549), .Z(n46002) );
  IV U55369 ( .A(n42551), .Z(n42553) );
  NOR U55370 ( .A(n42553), .B(n42552), .Z(n45691) );
  NOR U55371 ( .A(n46002), .B(n45691), .Z(n42870) );
  IV U55372 ( .A(n42554), .Z(n42556) );
  NOR U55373 ( .A(n42556), .B(n42555), .Z(n45694) );
  IV U55374 ( .A(n42557), .Z(n42561) );
  XOR U55375 ( .A(n42855), .B(n42863), .Z(n42558) );
  NOR U55376 ( .A(n42559), .B(n42558), .Z(n42560) );
  IV U55377 ( .A(n42560), .Z(n42859) );
  NOR U55378 ( .A(n42561), .B(n42859), .Z(n45701) );
  NOR U55379 ( .A(n45694), .B(n45701), .Z(n42869) );
  IV U55380 ( .A(n42562), .Z(n42563) );
  NOR U55381 ( .A(n42564), .B(n42563), .Z(n42565) );
  IV U55382 ( .A(n42565), .Z(n42865) );
  IV U55383 ( .A(n42566), .Z(n42571) );
  IV U55384 ( .A(n42567), .Z(n42568) );
  NOR U55385 ( .A(n42571), .B(n42568), .Z(n45710) );
  IV U55386 ( .A(n42569), .Z(n42570) );
  NOR U55387 ( .A(n42571), .B(n42570), .Z(n45716) );
  IV U55388 ( .A(n42572), .Z(n42574) );
  IV U55389 ( .A(n42573), .Z(n42576) );
  NOR U55390 ( .A(n42574), .B(n42576), .Z(n45976) );
  IV U55391 ( .A(n42575), .Z(n42577) );
  NOR U55392 ( .A(n42577), .B(n42576), .Z(n45973) );
  NOR U55393 ( .A(n42578), .B(n45966), .Z(n42579) );
  NOR U55394 ( .A(n42580), .B(n42579), .Z(n42581) );
  IV U55395 ( .A(n42581), .Z(n42835) );
  NOR U55396 ( .A(n42583), .B(n42582), .Z(n45726) );
  IV U55397 ( .A(n42584), .Z(n42588) );
  IV U55398 ( .A(n42585), .Z(n42586) );
  NOR U55399 ( .A(n42588), .B(n42586), .Z(n45732) );
  IV U55400 ( .A(n42587), .Z(n42589) );
  NOR U55401 ( .A(n42589), .B(n42588), .Z(n45959) );
  IV U55402 ( .A(n42590), .Z(n42592) );
  IV U55403 ( .A(n42591), .Z(n42817) );
  NOR U55404 ( .A(n42592), .B(n42817), .Z(n42814) );
  IV U55405 ( .A(n42814), .Z(n42809) );
  IV U55406 ( .A(n42593), .Z(n42594) );
  NOR U55407 ( .A(n42597), .B(n42594), .Z(n49279) );
  IV U55408 ( .A(n42595), .Z(n42599) );
  NOR U55409 ( .A(n42597), .B(n42596), .Z(n42598) );
  IV U55410 ( .A(n42598), .Z(n42811) );
  NOR U55411 ( .A(n42599), .B(n42811), .Z(n49432) );
  NOR U55412 ( .A(n49279), .B(n49432), .Z(n45933) );
  IV U55413 ( .A(n42610), .Z(n42601) );
  IV U55414 ( .A(n42600), .Z(n42609) );
  NOR U55415 ( .A(n42601), .B(n42609), .Z(n45747) );
  XOR U55416 ( .A(n42603), .B(n42602), .Z(n42604) );
  NOR U55417 ( .A(n42605), .B(n42604), .Z(n42606) );
  IV U55418 ( .A(n42606), .Z(n42615) );
  XOR U55419 ( .A(n42608), .B(n42607), .Z(n42612) );
  XOR U55420 ( .A(n42610), .B(n42609), .Z(n42611) );
  NOR U55421 ( .A(n42612), .B(n42611), .Z(n42613) );
  IV U55422 ( .A(n42613), .Z(n42614) );
  NOR U55423 ( .A(n42615), .B(n42614), .Z(n45929) );
  NOR U55424 ( .A(n45747), .B(n45929), .Z(n42808) );
  IV U55425 ( .A(n42616), .Z(n42617) );
  NOR U55426 ( .A(n42617), .B(n42787), .Z(n42790) );
  IV U55427 ( .A(n42618), .Z(n42619) );
  NOR U55428 ( .A(n42619), .B(n42787), .Z(n42794) );
  NOR U55429 ( .A(n42790), .B(n42794), .Z(n42620) );
  IV U55430 ( .A(n42620), .Z(n42789) );
  IV U55431 ( .A(n42621), .Z(n42624) );
  IV U55432 ( .A(n42622), .Z(n42623) );
  NOR U55433 ( .A(n42624), .B(n42623), .Z(n45910) );
  IV U55434 ( .A(n42625), .Z(n42627) );
  NOR U55435 ( .A(n42627), .B(n42626), .Z(n45753) );
  IV U55436 ( .A(n42628), .Z(n42630) );
  NOR U55437 ( .A(n42630), .B(n42629), .Z(n45900) );
  NOR U55438 ( .A(n45753), .B(n45900), .Z(n42631) );
  IV U55439 ( .A(n42631), .Z(n42778) );
  IV U55440 ( .A(n42632), .Z(n42633) );
  NOR U55441 ( .A(n42636), .B(n42633), .Z(n45758) );
  IV U55442 ( .A(n42634), .Z(n42635) );
  NOR U55443 ( .A(n42636), .B(n42635), .Z(n45755) );
  IV U55444 ( .A(n42637), .Z(n42639) );
  IV U55445 ( .A(n42638), .Z(n42776) );
  NOR U55446 ( .A(n42639), .B(n42776), .Z(n45887) );
  IV U55447 ( .A(n42640), .Z(n42642) );
  NOR U55448 ( .A(n42642), .B(n42641), .Z(n42643) );
  IV U55449 ( .A(n42643), .Z(n42770) );
  IV U55450 ( .A(n42644), .Z(n42648) );
  IV U55451 ( .A(n42645), .Z(n45770) );
  NOR U55452 ( .A(n45770), .B(n42646), .Z(n42647) );
  IV U55453 ( .A(n42647), .Z(n42650) );
  NOR U55454 ( .A(n42648), .B(n42650), .Z(n45881) );
  IV U55455 ( .A(n42649), .Z(n42651) );
  NOR U55456 ( .A(n42651), .B(n42650), .Z(n45766) );
  NOR U55457 ( .A(n42652), .B(n45770), .Z(n42764) );
  IV U55458 ( .A(n42653), .Z(n42655) );
  NOR U55459 ( .A(n42655), .B(n42654), .Z(n45874) );
  IV U55460 ( .A(n42656), .Z(n42658) );
  NOR U55461 ( .A(n42658), .B(n42657), .Z(n42745) );
  IV U55462 ( .A(n42745), .Z(n42739) );
  IV U55463 ( .A(n42659), .Z(n42663) );
  NOR U55464 ( .A(n42661), .B(n42660), .Z(n42662) );
  IV U55465 ( .A(n42662), .Z(n42665) );
  NOR U55466 ( .A(n42663), .B(n42665), .Z(n45857) );
  IV U55467 ( .A(n42664), .Z(n42666) );
  NOR U55468 ( .A(n42666), .B(n42665), .Z(n45781) );
  IV U55469 ( .A(n42667), .Z(n42668) );
  NOR U55470 ( .A(n42670), .B(n42668), .Z(n45850) );
  NOR U55471 ( .A(n42670), .B(n42669), .Z(n42671) );
  IV U55472 ( .A(n42671), .Z(n42676) );
  NOR U55473 ( .A(n42673), .B(n42672), .Z(n42674) );
  IV U55474 ( .A(n42674), .Z(n42675) );
  NOR U55475 ( .A(n42676), .B(n42675), .Z(n45785) );
  IV U55476 ( .A(n42677), .Z(n42679) );
  IV U55477 ( .A(n42678), .Z(n42682) );
  NOR U55478 ( .A(n42679), .B(n42682), .Z(n45839) );
  NOR U55479 ( .A(n45785), .B(n45839), .Z(n42738) );
  NOR U55480 ( .A(n42680), .B(n45788), .Z(n42684) );
  IV U55481 ( .A(n42681), .Z(n42683) );
  NOR U55482 ( .A(n42683), .B(n42682), .Z(n45842) );
  NOR U55483 ( .A(n42684), .B(n45842), .Z(n42737) );
  IV U55484 ( .A(n42685), .Z(n42736) );
  IV U55485 ( .A(n42686), .Z(n42687) );
  NOR U55486 ( .A(n42736), .B(n42687), .Z(n45795) );
  IV U55487 ( .A(n42688), .Z(n42691) );
  NOR U55488 ( .A(n42689), .B(n42697), .Z(n42690) );
  IV U55489 ( .A(n42690), .Z(n42725) );
  NOR U55490 ( .A(n42691), .B(n42725), .Z(n45811) );
  IV U55491 ( .A(n42692), .Z(n42701) );
  IV U55492 ( .A(n42693), .Z(n42694) );
  NOR U55493 ( .A(n42701), .B(n42694), .Z(n45814) );
  IV U55494 ( .A(n42695), .Z(n42696) );
  NOR U55495 ( .A(n42697), .B(n42696), .Z(n45809) );
  NOR U55496 ( .A(n45814), .B(n45809), .Z(n42698) );
  IV U55497 ( .A(n42698), .Z(n42723) );
  IV U55498 ( .A(n42699), .Z(n42700) );
  NOR U55499 ( .A(n42701), .B(n42700), .Z(n45825) );
  IV U55500 ( .A(n42702), .Z(n42703) );
  NOR U55501 ( .A(n42703), .B(n42708), .Z(n45820) );
  IV U55502 ( .A(n42704), .Z(n42705) );
  NOR U55503 ( .A(n42706), .B(n42705), .Z(n42711) );
  IV U55504 ( .A(n42707), .Z(n42709) );
  NOR U55505 ( .A(n42709), .B(n42708), .Z(n42710) );
  NOR U55506 ( .A(n42711), .B(n42710), .Z(n45818) );
  XOR U55507 ( .A(n45818), .B(n45817), .Z(n45819) );
  XOR U55508 ( .A(n45820), .B(n45819), .Z(n42719) );
  IV U55509 ( .A(n42715), .Z(n42716) );
  NOR U55510 ( .A(n42716), .B(n42721), .Z(n42717) );
  NOR U55511 ( .A(n42718), .B(n42717), .Z(n45821) );
  XOR U55512 ( .A(n42719), .B(n45821), .Z(n45824) );
  IV U55513 ( .A(n42720), .Z(n42722) );
  NOR U55514 ( .A(n42722), .B(n42721), .Z(n45822) );
  XOR U55515 ( .A(n45824), .B(n45822), .Z(n45826) );
  XOR U55516 ( .A(n45825), .B(n45826), .Z(n45815) );
  XOR U55517 ( .A(n42723), .B(n45815), .Z(n45812) );
  XOR U55518 ( .A(n45811), .B(n45812), .Z(n45803) );
  IV U55519 ( .A(n42724), .Z(n42726) );
  NOR U55520 ( .A(n42726), .B(n42725), .Z(n42727) );
  IV U55521 ( .A(n42727), .Z(n45802) );
  XOR U55522 ( .A(n45803), .B(n45802), .Z(n45799) );
  IV U55523 ( .A(n42728), .Z(n42729) );
  NOR U55524 ( .A(n42736), .B(n42729), .Z(n45800) );
  IV U55525 ( .A(n42730), .Z(n42731) );
  NOR U55526 ( .A(n42732), .B(n42731), .Z(n45804) );
  NOR U55527 ( .A(n45800), .B(n45804), .Z(n42733) );
  XOR U55528 ( .A(n45799), .B(n42733), .Z(n45794) );
  IV U55529 ( .A(n42734), .Z(n42735) );
  NOR U55530 ( .A(n42736), .B(n42735), .Z(n45792) );
  XOR U55531 ( .A(n45794), .B(n45792), .Z(n45797) );
  XOR U55532 ( .A(n45795), .B(n45797), .Z(n45844) );
  XOR U55533 ( .A(n42737), .B(n45844), .Z(n45784) );
  XOR U55534 ( .A(n42738), .B(n45784), .Z(n45852) );
  XOR U55535 ( .A(n45850), .B(n45852), .Z(n45783) );
  XOR U55536 ( .A(n45781), .B(n45783), .Z(n45859) );
  XOR U55537 ( .A(n45857), .B(n45859), .Z(n45860) );
  NOR U55538 ( .A(n42739), .B(n45860), .Z(n49343) );
  IV U55539 ( .A(n42740), .Z(n42742) );
  NOR U55540 ( .A(n42742), .B(n42741), .Z(n42743) );
  IV U55541 ( .A(n42743), .Z(n45861) );
  XOR U55542 ( .A(n45861), .B(n45860), .Z(n42744) );
  NOR U55543 ( .A(n42745), .B(n42744), .Z(n45869) );
  IV U55544 ( .A(n42746), .Z(n42748) );
  NOR U55545 ( .A(n42748), .B(n42747), .Z(n45867) );
  XOR U55546 ( .A(n45869), .B(n45867), .Z(n42749) );
  NOR U55547 ( .A(n49343), .B(n42749), .Z(n42750) );
  IV U55548 ( .A(n42750), .Z(n45865) );
  IV U55549 ( .A(n42751), .Z(n42752) );
  NOR U55550 ( .A(n42752), .B(n42754), .Z(n45863) );
  XOR U55551 ( .A(n45865), .B(n45863), .Z(n45777) );
  IV U55552 ( .A(n42753), .Z(n42755) );
  NOR U55553 ( .A(n42755), .B(n42754), .Z(n42756) );
  IV U55554 ( .A(n42756), .Z(n45776) );
  XOR U55555 ( .A(n45777), .B(n45776), .Z(n45773) );
  IV U55556 ( .A(n42757), .Z(n42758) );
  NOR U55557 ( .A(n42761), .B(n42758), .Z(n45778) );
  IV U55558 ( .A(n42759), .Z(n42760) );
  NOR U55559 ( .A(n42761), .B(n42760), .Z(n45774) );
  NOR U55560 ( .A(n45778), .B(n45774), .Z(n42762) );
  XOR U55561 ( .A(n45773), .B(n42762), .Z(n45875) );
  XOR U55562 ( .A(n45874), .B(n45875), .Z(n42763) );
  XOR U55563 ( .A(n42764), .B(n42763), .Z(n45767) );
  XOR U55564 ( .A(n45766), .B(n45767), .Z(n45883) );
  XOR U55565 ( .A(n45881), .B(n45883), .Z(n45884) );
  NOR U55566 ( .A(n42770), .B(n45884), .Z(n45765) );
  NOR U55567 ( .A(n42765), .B(n49411), .Z(n45890) );
  IV U55568 ( .A(n42766), .Z(n42767) );
  NOR U55569 ( .A(n42768), .B(n42767), .Z(n42769) );
  IV U55570 ( .A(n42769), .Z(n45885) );
  XOR U55571 ( .A(n45885), .B(n45884), .Z(n45891) );
  XOR U55572 ( .A(n45890), .B(n45891), .Z(n42772) );
  NOR U55573 ( .A(n45891), .B(n42770), .Z(n42771) );
  NOR U55574 ( .A(n42772), .B(n42771), .Z(n42773) );
  NOR U55575 ( .A(n45765), .B(n42773), .Z(n45761) );
  IV U55576 ( .A(n42774), .Z(n42775) );
  NOR U55577 ( .A(n42776), .B(n42775), .Z(n42777) );
  IV U55578 ( .A(n42777), .Z(n45762) );
  XOR U55579 ( .A(n45761), .B(n45762), .Z(n45889) );
  XOR U55580 ( .A(n45887), .B(n45889), .Z(n45757) );
  XOR U55581 ( .A(n45755), .B(n45757), .Z(n45760) );
  XOR U55582 ( .A(n45758), .B(n45760), .Z(n45901) );
  XOR U55583 ( .A(n42778), .B(n45901), .Z(n45905) );
  XOR U55584 ( .A(n45903), .B(n45905), .Z(n45907) );
  XOR U55585 ( .A(n45906), .B(n45907), .Z(n45911) );
  XOR U55586 ( .A(n45910), .B(n45911), .Z(n45915) );
  IV U55587 ( .A(n42779), .Z(n42782) );
  IV U55588 ( .A(n42780), .Z(n42781) );
  NOR U55589 ( .A(n42782), .B(n42781), .Z(n45913) );
  XOR U55590 ( .A(n45915), .B(n45913), .Z(n49287) );
  IV U55591 ( .A(n42783), .Z(n42784) );
  NOR U55592 ( .A(n42785), .B(n42784), .Z(n49286) );
  IV U55593 ( .A(n42786), .Z(n42788) );
  NOR U55594 ( .A(n42788), .B(n42787), .Z(n49423) );
  NOR U55595 ( .A(n49286), .B(n49423), .Z(n45917) );
  XOR U55596 ( .A(n49287), .B(n45917), .Z(n42791) );
  NOR U55597 ( .A(n42789), .B(n42791), .Z(n42798) );
  IV U55598 ( .A(n42790), .Z(n42793) );
  IV U55599 ( .A(n42791), .Z(n42792) );
  NOR U55600 ( .A(n42793), .B(n42792), .Z(n49421) );
  IV U55601 ( .A(n42794), .Z(n42795) );
  NOR U55602 ( .A(n42795), .B(n49287), .Z(n45924) );
  NOR U55603 ( .A(n49421), .B(n45924), .Z(n42796) );
  IV U55604 ( .A(n42796), .Z(n42797) );
  NOR U55605 ( .A(n42798), .B(n42797), .Z(n45750) );
  XOR U55606 ( .A(n42800), .B(n42799), .Z(n42803) );
  IV U55607 ( .A(n42801), .Z(n42802) );
  NOR U55608 ( .A(n42803), .B(n42802), .Z(n42804) );
  IV U55609 ( .A(n42804), .Z(n42805) );
  NOR U55610 ( .A(n42806), .B(n42805), .Z(n42807) );
  IV U55611 ( .A(n42807), .Z(n45751) );
  XOR U55612 ( .A(n45750), .B(n45751), .Z(n45931) );
  XOR U55613 ( .A(n42808), .B(n45931), .Z(n45932) );
  XOR U55614 ( .A(n45933), .B(n45932), .Z(n45934) );
  NOR U55615 ( .A(n42809), .B(n45934), .Z(n49271) );
  IV U55616 ( .A(n42810), .Z(n42812) );
  NOR U55617 ( .A(n42812), .B(n42811), .Z(n42813) );
  IV U55618 ( .A(n42813), .Z(n45935) );
  XOR U55619 ( .A(n45935), .B(n45934), .Z(n45941) );
  NOR U55620 ( .A(n42814), .B(n45941), .Z(n42815) );
  NOR U55621 ( .A(n49271), .B(n42815), .Z(n45949) );
  IV U55622 ( .A(n42816), .Z(n42818) );
  NOR U55623 ( .A(n42818), .B(n42817), .Z(n45940) );
  IV U55624 ( .A(n42819), .Z(n42821) );
  NOR U55625 ( .A(n42821), .B(n42820), .Z(n45948) );
  NOR U55626 ( .A(n45940), .B(n45948), .Z(n42822) );
  XOR U55627 ( .A(n45949), .B(n42822), .Z(n45746) );
  IV U55628 ( .A(n42823), .Z(n42824) );
  NOR U55629 ( .A(n42825), .B(n42824), .Z(n45744) );
  IV U55630 ( .A(n42826), .Z(n42828) );
  NOR U55631 ( .A(n42828), .B(n42827), .Z(n45741) );
  NOR U55632 ( .A(n45744), .B(n45741), .Z(n42829) );
  XOR U55633 ( .A(n45746), .B(n42829), .Z(n45739) );
  IV U55634 ( .A(n42830), .Z(n42831) );
  NOR U55635 ( .A(n42831), .B(n42833), .Z(n49259) );
  IV U55636 ( .A(n42832), .Z(n42834) );
  NOR U55637 ( .A(n42834), .B(n42833), .Z(n49255) );
  NOR U55638 ( .A(n49259), .B(n49255), .Z(n45740) );
  XOR U55639 ( .A(n45739), .B(n45740), .Z(n45737) );
  XOR U55640 ( .A(n45736), .B(n45737), .Z(n45957) );
  XOR U55641 ( .A(n45956), .B(n45957), .Z(n45960) );
  XOR U55642 ( .A(n45959), .B(n45960), .Z(n45733) );
  XOR U55643 ( .A(n45732), .B(n45733), .Z(n45727) );
  XOR U55644 ( .A(n45726), .B(n45727), .Z(n45965) );
  XOR U55645 ( .A(n42835), .B(n45965), .Z(n45975) );
  XOR U55646 ( .A(n45973), .B(n45975), .Z(n45977) );
  XOR U55647 ( .A(n45976), .B(n45977), .Z(n45720) );
  IV U55648 ( .A(n42836), .Z(n42838) );
  NOR U55649 ( .A(n42838), .B(n42837), .Z(n45722) );
  IV U55650 ( .A(n42839), .Z(n42841) );
  NOR U55651 ( .A(n42841), .B(n42840), .Z(n45719) );
  NOR U55652 ( .A(n45722), .B(n45719), .Z(n42842) );
  XOR U55653 ( .A(n45720), .B(n42842), .Z(n45981) );
  IV U55654 ( .A(n42843), .Z(n42844) );
  NOR U55655 ( .A(n42844), .B(n42846), .Z(n45982) );
  IV U55656 ( .A(n42845), .Z(n42847) );
  NOR U55657 ( .A(n42847), .B(n42846), .Z(n45989) );
  NOR U55658 ( .A(n45982), .B(n45989), .Z(n42848) );
  XOR U55659 ( .A(n45981), .B(n42848), .Z(n45988) );
  IV U55660 ( .A(n42849), .Z(n42850) );
  NOR U55661 ( .A(n42851), .B(n42850), .Z(n45986) );
  XOR U55662 ( .A(n45988), .B(n45986), .Z(n45717) );
  XOR U55663 ( .A(n45716), .B(n45717), .Z(n45711) );
  XOR U55664 ( .A(n45710), .B(n45711), .Z(n45714) );
  IV U55665 ( .A(n42852), .Z(n42854) );
  NOR U55666 ( .A(n42854), .B(n42853), .Z(n45713) );
  IV U55667 ( .A(n42855), .Z(n42856) );
  NOR U55668 ( .A(n42863), .B(n42856), .Z(n45705) );
  NOR U55669 ( .A(n45713), .B(n45705), .Z(n42857) );
  XOR U55670 ( .A(n45714), .B(n42857), .Z(n42864) );
  IV U55671 ( .A(n42864), .Z(n45708) );
  NOR U55672 ( .A(n42865), .B(n45708), .Z(n49231) );
  IV U55673 ( .A(n42858), .Z(n42860) );
  NOR U55674 ( .A(n42860), .B(n42859), .Z(n45697) );
  IV U55675 ( .A(n42861), .Z(n42862) );
  NOR U55676 ( .A(n42863), .B(n42862), .Z(n45707) );
  XOR U55677 ( .A(n45707), .B(n42864), .Z(n45698) );
  XOR U55678 ( .A(n45697), .B(n45698), .Z(n42867) );
  NOR U55679 ( .A(n45698), .B(n42865), .Z(n42866) );
  NOR U55680 ( .A(n42867), .B(n42866), .Z(n42868) );
  NOR U55681 ( .A(n49231), .B(n42868), .Z(n45695) );
  XOR U55682 ( .A(n42869), .B(n45695), .Z(n46004) );
  XOR U55683 ( .A(n42870), .B(n46004), .Z(n46006) );
  XOR U55684 ( .A(n42871), .B(n46006), .Z(n46016) );
  XOR U55685 ( .A(n42872), .B(n46016), .Z(n42873) );
  IV U55686 ( .A(n42873), .Z(n45686) );
  XOR U55687 ( .A(n45685), .B(n45686), .Z(n46023) );
  XOR U55688 ( .A(n42874), .B(n46023), .Z(n45679) );
  XOR U55689 ( .A(n42875), .B(n45679), .Z(n46027) );
  XOR U55690 ( .A(n42876), .B(n46027), .Z(n45673) );
  XOR U55691 ( .A(n45671), .B(n45673), .Z(n46038) );
  IV U55692 ( .A(n49185), .Z(n42877) );
  NOR U55693 ( .A(n49184), .B(n42877), .Z(n46037) );
  IV U55694 ( .A(n42878), .Z(n42880) );
  NOR U55695 ( .A(n42880), .B(n42879), .Z(n46029) );
  NOR U55696 ( .A(n46037), .B(n46029), .Z(n42881) );
  XOR U55697 ( .A(n46038), .B(n42881), .Z(n46040) );
  IV U55698 ( .A(n42882), .Z(n49187) );
  NOR U55699 ( .A(n49184), .B(n49187), .Z(n42885) );
  NOR U55700 ( .A(n42884), .B(n42883), .Z(n49188) );
  NOR U55701 ( .A(n42885), .B(n49188), .Z(n46041) );
  XOR U55702 ( .A(n46040), .B(n46041), .Z(n46047) );
  XOR U55703 ( .A(n46048), .B(n46047), .Z(n45666) );
  IV U55704 ( .A(n42886), .Z(n42889) );
  IV U55705 ( .A(n42887), .Z(n42888) );
  NOR U55706 ( .A(n42889), .B(n42888), .Z(n46044) );
  IV U55707 ( .A(n42890), .Z(n42892) );
  NOR U55708 ( .A(n42892), .B(n42891), .Z(n45665) );
  NOR U55709 ( .A(n46044), .B(n45665), .Z(n42893) );
  XOR U55710 ( .A(n45666), .B(n42893), .Z(n45669) );
  XOR U55711 ( .A(n45668), .B(n45669), .Z(n46060) );
  XOR U55712 ( .A(n46058), .B(n46060), .Z(n46062) );
  XOR U55713 ( .A(n42894), .B(n46062), .Z(n45655) );
  XOR U55714 ( .A(n42895), .B(n45655), .Z(n46068) );
  XOR U55715 ( .A(n46066), .B(n46068), .Z(n46070) );
  XOR U55716 ( .A(n46069), .B(n46070), .Z(n45653) );
  XOR U55717 ( .A(n42896), .B(n45653), .Z(n42897) );
  IV U55718 ( .A(n42897), .Z(n46074) );
  IV U55719 ( .A(n42898), .Z(n42899) );
  NOR U55720 ( .A(n42900), .B(n42899), .Z(n45650) );
  IV U55721 ( .A(n42901), .Z(n42902) );
  NOR U55722 ( .A(n42903), .B(n42902), .Z(n46073) );
  NOR U55723 ( .A(n45650), .B(n46073), .Z(n42904) );
  XOR U55724 ( .A(n46074), .B(n42904), .Z(n45646) );
  IV U55725 ( .A(n42905), .Z(n42906) );
  NOR U55726 ( .A(n42907), .B(n42906), .Z(n49509) );
  IV U55727 ( .A(n42908), .Z(n42910) );
  NOR U55728 ( .A(n42910), .B(n42909), .Z(n49154) );
  NOR U55729 ( .A(n49509), .B(n49154), .Z(n45647) );
  XOR U55730 ( .A(n45646), .B(n45647), .Z(n46078) );
  XOR U55731 ( .A(n46077), .B(n46078), .Z(n46081) );
  NOR U55732 ( .A(n42913), .B(n42911), .Z(n46080) );
  IV U55733 ( .A(n42912), .Z(n42916) );
  NOR U55734 ( .A(n42914), .B(n42913), .Z(n42915) );
  IV U55735 ( .A(n42915), .Z(n42922) );
  NOR U55736 ( .A(n42916), .B(n42922), .Z(n45641) );
  NOR U55737 ( .A(n46080), .B(n45641), .Z(n42917) );
  XOR U55738 ( .A(n46081), .B(n42917), .Z(n45643) );
  IV U55739 ( .A(n42918), .Z(n42920) );
  IV U55740 ( .A(n42919), .Z(n42925) );
  NOR U55741 ( .A(n42920), .B(n42925), .Z(n46093) );
  IV U55742 ( .A(n42921), .Z(n42923) );
  NOR U55743 ( .A(n42923), .B(n42922), .Z(n45644) );
  NOR U55744 ( .A(n46093), .B(n45644), .Z(n42924) );
  XOR U55745 ( .A(n45643), .B(n42924), .Z(n49142) );
  IV U55746 ( .A(n49139), .Z(n42926) );
  NOR U55747 ( .A(n42926), .B(n42925), .Z(n45638) );
  XOR U55748 ( .A(n49142), .B(n45638), .Z(n46097) );
  XOR U55749 ( .A(n46096), .B(n46097), .Z(n46100) );
  XOR U55750 ( .A(n46099), .B(n46100), .Z(n46106) );
  IV U55751 ( .A(n42927), .Z(n42929) );
  NOR U55752 ( .A(n42929), .B(n42928), .Z(n46104) );
  XOR U55753 ( .A(n46106), .B(n46104), .Z(n46108) );
  XOR U55754 ( .A(n46107), .B(n46108), .Z(n45637) );
  IV U55755 ( .A(n42930), .Z(n42932) );
  NOR U55756 ( .A(n42932), .B(n42931), .Z(n45635) );
  XOR U55757 ( .A(n45637), .B(n45635), .Z(n46116) );
  XOR U55758 ( .A(n46117), .B(n46116), .Z(n45630) );
  NOR U55759 ( .A(n46121), .B(n42933), .Z(n42939) );
  IV U55760 ( .A(n42934), .Z(n42938) );
  NOR U55761 ( .A(n42936), .B(n42935), .Z(n42937) );
  IV U55762 ( .A(n42937), .Z(n42942) );
  NOR U55763 ( .A(n42938), .B(n42942), .Z(n46125) );
  NOR U55764 ( .A(n42939), .B(n46125), .Z(n42940) );
  XOR U55765 ( .A(n45630), .B(n42940), .Z(n45628) );
  IV U55766 ( .A(n42941), .Z(n42943) );
  NOR U55767 ( .A(n42943), .B(n42942), .Z(n45626) );
  XOR U55768 ( .A(n45628), .B(n45626), .Z(n46133) );
  XOR U55769 ( .A(n46132), .B(n46133), .Z(n46140) );
  XOR U55770 ( .A(n42944), .B(n46140), .Z(n46141) );
  IV U55771 ( .A(n42945), .Z(n42950) );
  NOR U55772 ( .A(n42947), .B(n42946), .Z(n42948) );
  IV U55773 ( .A(n42948), .Z(n42949) );
  NOR U55774 ( .A(n42950), .B(n42949), .Z(n46142) );
  XOR U55775 ( .A(n46141), .B(n46142), .Z(n45621) );
  XOR U55776 ( .A(n45620), .B(n45621), .Z(n46147) );
  IV U55777 ( .A(n42951), .Z(n42952) );
  NOR U55778 ( .A(n42953), .B(n42952), .Z(n45623) );
  IV U55779 ( .A(n42954), .Z(n42965) );
  IV U55780 ( .A(n42955), .Z(n42956) );
  NOR U55781 ( .A(n42965), .B(n42956), .Z(n46146) );
  NOR U55782 ( .A(n45623), .B(n46146), .Z(n42957) );
  XOR U55783 ( .A(n46147), .B(n42957), .Z(n42967) );
  IV U55784 ( .A(n42967), .Z(n45618) );
  IV U55785 ( .A(n42958), .Z(n42960) );
  NOR U55786 ( .A(n42960), .B(n42959), .Z(n42961) );
  IV U55787 ( .A(n42961), .Z(n42968) );
  NOR U55788 ( .A(n45618), .B(n42968), .Z(n49539) );
  IV U55789 ( .A(n42962), .Z(n42963) );
  NOR U55790 ( .A(n42973), .B(n42963), .Z(n45609) );
  IV U55791 ( .A(n42964), .Z(n42966) );
  NOR U55792 ( .A(n42966), .B(n42965), .Z(n45616) );
  XOR U55793 ( .A(n45616), .B(n42967), .Z(n45610) );
  XOR U55794 ( .A(n45609), .B(n45610), .Z(n42970) );
  NOR U55795 ( .A(n45610), .B(n42968), .Z(n42969) );
  NOR U55796 ( .A(n42970), .B(n42969), .Z(n42971) );
  NOR U55797 ( .A(n49539), .B(n42971), .Z(n45606) );
  IV U55798 ( .A(n42972), .Z(n42974) );
  NOR U55799 ( .A(n42974), .B(n42973), .Z(n45613) );
  IV U55800 ( .A(n42975), .Z(n42977) );
  NOR U55801 ( .A(n42977), .B(n42976), .Z(n45605) );
  NOR U55802 ( .A(n45613), .B(n45605), .Z(n42978) );
  XOR U55803 ( .A(n45606), .B(n42978), .Z(n45604) );
  XOR U55804 ( .A(n45602), .B(n45604), .Z(n45600) );
  XOR U55805 ( .A(n45598), .B(n45600), .Z(n46169) );
  XOR U55806 ( .A(n42979), .B(n46169), .Z(n46171) );
  XOR U55807 ( .A(n46172), .B(n46171), .Z(n46175) );
  IV U55808 ( .A(n42980), .Z(n42981) );
  NOR U55809 ( .A(n42985), .B(n42981), .Z(n46180) );
  NOR U55810 ( .A(n46174), .B(n46180), .Z(n42982) );
  XOR U55811 ( .A(n46175), .B(n42982), .Z(n46179) );
  IV U55812 ( .A(n42983), .Z(n42984) );
  NOR U55813 ( .A(n42985), .B(n42984), .Z(n46177) );
  XOR U55814 ( .A(n46179), .B(n46177), .Z(n45594) );
  XOR U55815 ( .A(n45592), .B(n45594), .Z(n45596) );
  XOR U55816 ( .A(n42986), .B(n45596), .Z(n45589) );
  XOR U55817 ( .A(n45587), .B(n45589), .Z(n45582) );
  IV U55818 ( .A(n42987), .Z(n42992) );
  IV U55819 ( .A(n42988), .Z(n42989) );
  NOR U55820 ( .A(n42989), .B(n42995), .Z(n42990) );
  IV U55821 ( .A(n42990), .Z(n42991) );
  NOR U55822 ( .A(n42992), .B(n42991), .Z(n42993) );
  IV U55823 ( .A(n42993), .Z(n45581) );
  XOR U55824 ( .A(n45582), .B(n45581), .Z(n45579) );
  IV U55825 ( .A(n42994), .Z(n42996) );
  NOR U55826 ( .A(n42996), .B(n42995), .Z(n45583) );
  IV U55827 ( .A(n42997), .Z(n42999) );
  NOR U55828 ( .A(n42999), .B(n42998), .Z(n45578) );
  NOR U55829 ( .A(n45583), .B(n45578), .Z(n43000) );
  XOR U55830 ( .A(n45579), .B(n43000), .Z(n45576) );
  IV U55831 ( .A(n43001), .Z(n43003) );
  NOR U55832 ( .A(n43003), .B(n43002), .Z(n45574) );
  XOR U55833 ( .A(n45576), .B(n45574), .Z(n46188) );
  XOR U55834 ( .A(n46186), .B(n46188), .Z(n46191) );
  IV U55835 ( .A(n43004), .Z(n43006) );
  NOR U55836 ( .A(n43006), .B(n43005), .Z(n45572) );
  IV U55837 ( .A(n43007), .Z(n43009) );
  NOR U55838 ( .A(n43009), .B(n43008), .Z(n46189) );
  NOR U55839 ( .A(n45572), .B(n46189), .Z(n43010) );
  XOR U55840 ( .A(n46191), .B(n43010), .Z(n43011) );
  NOR U55841 ( .A(n43012), .B(n43011), .Z(n43015) );
  IV U55842 ( .A(n43012), .Z(n43014) );
  XOR U55843 ( .A(n46189), .B(n46191), .Z(n43013) );
  NOR U55844 ( .A(n43014), .B(n43013), .Z(n49597) );
  NOR U55845 ( .A(n43015), .B(n49597), .Z(n43016) );
  IV U55846 ( .A(n43016), .Z(n45566) );
  XOR U55847 ( .A(n45565), .B(n45566), .Z(n45570) );
  XOR U55848 ( .A(n45568), .B(n45570), .Z(n46201) );
  XOR U55849 ( .A(n43017), .B(n46201), .Z(n46210) );
  XOR U55850 ( .A(n46208), .B(n46210), .Z(n46206) );
  IV U55851 ( .A(n43018), .Z(n43020) );
  IV U55852 ( .A(n43019), .Z(n43026) );
  NOR U55853 ( .A(n43020), .B(n43026), .Z(n46204) );
  XOR U55854 ( .A(n46206), .B(n46204), .Z(n46220) );
  IV U55855 ( .A(n43021), .Z(n43022) );
  NOR U55856 ( .A(n43023), .B(n43022), .Z(n46219) );
  IV U55857 ( .A(n43024), .Z(n43025) );
  NOR U55858 ( .A(n43026), .B(n43025), .Z(n45559) );
  NOR U55859 ( .A(n46219), .B(n45559), .Z(n43027) );
  XOR U55860 ( .A(n46220), .B(n43027), .Z(n45552) );
  IV U55861 ( .A(n43028), .Z(n43029) );
  NOR U55862 ( .A(n43029), .B(n46235), .Z(n46233) );
  NOR U55863 ( .A(n43031), .B(n43030), .Z(n45553) );
  NOR U55864 ( .A(n46233), .B(n45553), .Z(n43032) );
  XOR U55865 ( .A(n45552), .B(n43032), .Z(n46239) );
  XOR U55866 ( .A(n46240), .B(n46239), .Z(n45548) );
  NOR U55867 ( .A(n43033), .B(n45548), .Z(n43046) );
  IV U55868 ( .A(n43034), .Z(n43040) );
  NOR U55869 ( .A(n43035), .B(n46239), .Z(n43036) );
  IV U55870 ( .A(n43036), .Z(n43037) );
  NOR U55871 ( .A(n43038), .B(n43037), .Z(n43039) );
  IV U55872 ( .A(n43039), .Z(n43042) );
  NOR U55873 ( .A(n43040), .B(n43042), .Z(n53545) );
  IV U55874 ( .A(n43041), .Z(n43043) );
  NOR U55875 ( .A(n43043), .B(n43042), .Z(n49046) );
  NOR U55876 ( .A(n53545), .B(n49046), .Z(n43044) );
  IV U55877 ( .A(n43044), .Z(n43045) );
  NOR U55878 ( .A(n43046), .B(n43045), .Z(n45544) );
  XOR U55879 ( .A(n43047), .B(n45544), .Z(n46246) );
  XOR U55880 ( .A(n46244), .B(n46246), .Z(n45541) );
  IV U55881 ( .A(n43048), .Z(n43050) );
  NOR U55882 ( .A(n43050), .B(n43049), .Z(n45539) );
  XOR U55883 ( .A(n45541), .B(n45539), .Z(n46243) );
  IV U55884 ( .A(n43051), .Z(n43053) );
  NOR U55885 ( .A(n43053), .B(n43052), .Z(n46241) );
  XOR U55886 ( .A(n46243), .B(n46241), .Z(n46256) );
  IV U55887 ( .A(n43054), .Z(n43063) );
  IV U55888 ( .A(n43055), .Z(n43056) );
  NOR U55889 ( .A(n43063), .B(n43056), .Z(n46255) );
  IV U55890 ( .A(n43057), .Z(n43059) );
  NOR U55891 ( .A(n43059), .B(n43058), .Z(n45537) );
  NOR U55892 ( .A(n46255), .B(n45537), .Z(n43060) );
  XOR U55893 ( .A(n46256), .B(n43060), .Z(n45534) );
  IV U55894 ( .A(n43061), .Z(n43062) );
  NOR U55895 ( .A(n43063), .B(n43062), .Z(n46252) );
  IV U55896 ( .A(n43064), .Z(n43070) );
  NOR U55897 ( .A(n43065), .B(n43073), .Z(n43066) );
  IV U55898 ( .A(n43066), .Z(n43067) );
  NOR U55899 ( .A(n43068), .B(n43067), .Z(n43069) );
  IV U55900 ( .A(n43069), .Z(n43076) );
  NOR U55901 ( .A(n43070), .B(n43076), .Z(n45535) );
  NOR U55902 ( .A(n46252), .B(n45535), .Z(n43071) );
  XOR U55903 ( .A(n45534), .B(n43071), .Z(n45532) );
  IV U55904 ( .A(n43072), .Z(n43074) );
  NOR U55905 ( .A(n43074), .B(n43073), .Z(n45529) );
  IV U55906 ( .A(n43075), .Z(n43077) );
  NOR U55907 ( .A(n43077), .B(n43076), .Z(n45531) );
  NOR U55908 ( .A(n45529), .B(n45531), .Z(n43078) );
  XOR U55909 ( .A(n45532), .B(n43078), .Z(n43079) );
  IV U55910 ( .A(n43079), .Z(n45528) );
  IV U55911 ( .A(n43080), .Z(n43082) );
  NOR U55912 ( .A(n43082), .B(n43081), .Z(n45526) );
  XOR U55913 ( .A(n45528), .B(n45526), .Z(n45522) );
  XOR U55914 ( .A(n45520), .B(n45522), .Z(n45524) );
  XOR U55915 ( .A(n45523), .B(n45524), .Z(n45518) );
  IV U55916 ( .A(n43083), .Z(n43084) );
  NOR U55917 ( .A(n43085), .B(n43084), .Z(n45517) );
  IV U55918 ( .A(n43086), .Z(n43087) );
  NOR U55919 ( .A(n43088), .B(n43087), .Z(n45515) );
  NOR U55920 ( .A(n45517), .B(n45515), .Z(n43089) );
  XOR U55921 ( .A(n45518), .B(n43089), .Z(n43090) );
  NOR U55922 ( .A(n43091), .B(n43090), .Z(n43094) );
  IV U55923 ( .A(n43091), .Z(n43093) );
  XOR U55924 ( .A(n45517), .B(n45518), .Z(n43092) );
  NOR U55925 ( .A(n43093), .B(n43092), .Z(n49031) );
  NOR U55926 ( .A(n43094), .B(n49031), .Z(n45511) );
  XOR U55927 ( .A(n45513), .B(n45511), .Z(n49020) );
  XOR U55928 ( .A(n45506), .B(n49020), .Z(n45503) );
  XOR U55929 ( .A(n43095), .B(n45503), .Z(n46267) );
  IV U55930 ( .A(n46267), .Z(n43105) );
  IV U55931 ( .A(n43096), .Z(n43098) );
  NOR U55932 ( .A(n43098), .B(n43097), .Z(n46265) );
  IV U55933 ( .A(n43099), .Z(n43103) );
  NOR U55934 ( .A(n43101), .B(n43100), .Z(n43102) );
  IV U55935 ( .A(n43102), .Z(n43107) );
  NOR U55936 ( .A(n43103), .B(n43107), .Z(n45501) );
  NOR U55937 ( .A(n46265), .B(n45501), .Z(n43104) );
  XOR U55938 ( .A(n43105), .B(n43104), .Z(n45497) );
  IV U55939 ( .A(n43106), .Z(n43108) );
  NOR U55940 ( .A(n43108), .B(n43107), .Z(n45495) );
  XOR U55941 ( .A(n45497), .B(n45495), .Z(n45499) );
  XOR U55942 ( .A(n45498), .B(n45499), .Z(n45491) );
  IV U55943 ( .A(n43113), .Z(n43111) );
  IV U55944 ( .A(n43109), .Z(n43110) );
  NOR U55945 ( .A(n43111), .B(n43110), .Z(n45489) );
  XOR U55946 ( .A(n45491), .B(n45489), .Z(n45494) );
  IV U55947 ( .A(n43112), .Z(n43116) );
  XOR U55948 ( .A(n43114), .B(n43113), .Z(n43115) );
  NOR U55949 ( .A(n43116), .B(n43115), .Z(n45492) );
  XOR U55950 ( .A(n45494), .B(n45492), .Z(n45482) );
  XOR U55951 ( .A(n43117), .B(n45482), .Z(n49007) );
  IV U55952 ( .A(n43118), .Z(n43120) );
  NOR U55953 ( .A(n43120), .B(n43119), .Z(n49006) );
  IV U55954 ( .A(n43121), .Z(n43122) );
  NOR U55955 ( .A(n43123), .B(n43122), .Z(n49685) );
  NOR U55956 ( .A(n49006), .B(n49685), .Z(n45476) );
  XOR U55957 ( .A(n49007), .B(n45476), .Z(n45474) );
  XOR U55958 ( .A(n43124), .B(n45474), .Z(n45466) );
  XOR U55959 ( .A(n45448), .B(n45450), .Z(n45452) );
  XOR U55960 ( .A(n45451), .B(n45452), .Z(n43128) );
  NOR U55961 ( .A(n43125), .B(n43128), .Z(n43126) );
  IV U55962 ( .A(n43126), .Z(n43127) );
  NOR U55963 ( .A(n43130), .B(n43127), .Z(n48990) );
  IV U55964 ( .A(n43128), .Z(n43132) );
  IV U55965 ( .A(n43129), .Z(n43135) );
  NOR U55966 ( .A(n43130), .B(n43135), .Z(n43131) );
  NOR U55967 ( .A(n43132), .B(n43131), .Z(n43133) );
  NOR U55968 ( .A(n48990), .B(n43133), .Z(n46276) );
  IV U55969 ( .A(n43134), .Z(n43136) );
  NOR U55970 ( .A(n43136), .B(n43135), .Z(n43137) );
  IV U55971 ( .A(n43137), .Z(n46277) );
  XOR U55972 ( .A(n46276), .B(n46277), .Z(n46289) );
  XOR U55973 ( .A(n43138), .B(n46289), .Z(n46301) );
  XOR U55974 ( .A(n43139), .B(n46301), .Z(n46305) );
  IV U55975 ( .A(n46305), .Z(n46307) );
  XOR U55976 ( .A(n46306), .B(n46307), .Z(n49706) );
  XOR U55977 ( .A(n43140), .B(n49706), .Z(n46318) );
  XOR U55978 ( .A(n46316), .B(n46318), .Z(n46319) );
  XOR U55979 ( .A(n46320), .B(n46319), .Z(n45438) );
  NOR U55980 ( .A(n43141), .B(n43143), .Z(n45442) );
  IV U55981 ( .A(n43142), .Z(n43146) );
  NOR U55982 ( .A(n43144), .B(n43143), .Z(n43145) );
  IV U55983 ( .A(n43145), .Z(n43149) );
  NOR U55984 ( .A(n43146), .B(n43149), .Z(n45439) );
  NOR U55985 ( .A(n45442), .B(n45439), .Z(n43147) );
  XOR U55986 ( .A(n45438), .B(n43147), .Z(n45435) );
  IV U55987 ( .A(n43148), .Z(n43150) );
  NOR U55988 ( .A(n43150), .B(n43149), .Z(n45433) );
  XOR U55989 ( .A(n45435), .B(n45433), .Z(n46323) );
  XOR U55990 ( .A(n45436), .B(n46323), .Z(n43151) );
  NOR U55991 ( .A(n43152), .B(n43151), .Z(n48963) );
  IV U55992 ( .A(n43153), .Z(n43154) );
  NOR U55993 ( .A(n43155), .B(n43154), .Z(n46322) );
  NOR U55994 ( .A(n46322), .B(n45436), .Z(n43156) );
  XOR U55995 ( .A(n46323), .B(n43156), .Z(n43157) );
  NOR U55996 ( .A(n43158), .B(n43157), .Z(n43159) );
  NOR U55997 ( .A(n48963), .B(n43159), .Z(n46326) );
  IV U55998 ( .A(n43160), .Z(n43161) );
  NOR U55999 ( .A(n43167), .B(n43161), .Z(n46327) );
  XOR U56000 ( .A(n46326), .B(n46327), .Z(n46330) );
  IV U56001 ( .A(n43162), .Z(n43163) );
  NOR U56002 ( .A(n43164), .B(n43163), .Z(n46334) );
  IV U56003 ( .A(n43165), .Z(n43166) );
  NOR U56004 ( .A(n43167), .B(n43166), .Z(n46331) );
  NOR U56005 ( .A(n46334), .B(n46331), .Z(n43168) );
  XOR U56006 ( .A(n46330), .B(n43168), .Z(n46339) );
  XOR U56007 ( .A(n46337), .B(n46339), .Z(n46342) );
  XOR U56008 ( .A(n46341), .B(n46342), .Z(n46345) );
  XOR U56009 ( .A(n46344), .B(n46345), .Z(n45424) );
  XOR U56010 ( .A(n43169), .B(n45424), .Z(n45421) );
  XOR U56011 ( .A(n45420), .B(n45421), .Z(n46352) );
  XOR U56012 ( .A(n46351), .B(n46352), .Z(n46355) );
  XOR U56013 ( .A(n46354), .B(n46355), .Z(n45416) );
  XOR U56014 ( .A(n45415), .B(n45416), .Z(n45410) );
  XOR U56015 ( .A(n45408), .B(n45410), .Z(n46361) );
  XOR U56016 ( .A(n46359), .B(n46361), .Z(n46362) );
  IV U56017 ( .A(n43170), .Z(n43171) );
  NOR U56018 ( .A(n43171), .B(n43173), .Z(n43172) );
  IV U56019 ( .A(n43172), .Z(n43179) );
  NOR U56020 ( .A(n46362), .B(n43179), .Z(n45402) );
  NOR U56021 ( .A(n43174), .B(n43173), .Z(n45403) );
  IV U56022 ( .A(n43175), .Z(n43176) );
  NOR U56023 ( .A(n43177), .B(n43176), .Z(n43178) );
  IV U56024 ( .A(n43178), .Z(n46363) );
  XOR U56025 ( .A(n46363), .B(n46362), .Z(n45404) );
  XOR U56026 ( .A(n45403), .B(n45404), .Z(n43181) );
  NOR U56027 ( .A(n45404), .B(n43179), .Z(n43180) );
  NOR U56028 ( .A(n43181), .B(n43180), .Z(n43182) );
  NOR U56029 ( .A(n45402), .B(n43182), .Z(n46374) );
  XOR U56030 ( .A(n46376), .B(n46374), .Z(n46378) );
  IV U56031 ( .A(n43183), .Z(n43184) );
  NOR U56032 ( .A(n43185), .B(n43184), .Z(n46377) );
  NOR U56033 ( .A(n43187), .B(n43186), .Z(n43188) );
  IV U56034 ( .A(n43188), .Z(n43193) );
  NOR U56035 ( .A(n43190), .B(n43189), .Z(n43191) );
  IV U56036 ( .A(n43191), .Z(n43192) );
  NOR U56037 ( .A(n43193), .B(n43192), .Z(n43194) );
  IV U56038 ( .A(n43194), .Z(n43195) );
  NOR U56039 ( .A(n43196), .B(n43195), .Z(n45400) );
  NOR U56040 ( .A(n46377), .B(n45400), .Z(n43197) );
  XOR U56041 ( .A(n46378), .B(n43197), .Z(n45395) );
  XOR U56042 ( .A(n43198), .B(n45395), .Z(n46386) );
  XOR U56043 ( .A(n43199), .B(n46386), .Z(n43200) );
  IV U56044 ( .A(n43200), .Z(n46382) );
  XOR U56045 ( .A(n46381), .B(n46382), .Z(n45390) );
  NOR U56046 ( .A(n43207), .B(n45390), .Z(n49775) );
  IV U56047 ( .A(n43201), .Z(n43203) );
  NOR U56048 ( .A(n43203), .B(n43202), .Z(n45389) );
  NOR U56049 ( .A(n43205), .B(n43204), .Z(n45387) );
  NOR U56050 ( .A(n45389), .B(n45387), .Z(n43206) );
  XOR U56051 ( .A(n43206), .B(n45390), .Z(n46389) );
  XOR U56052 ( .A(n46388), .B(n46389), .Z(n43209) );
  NOR U56053 ( .A(n46389), .B(n43207), .Z(n43208) );
  NOR U56054 ( .A(n43209), .B(n43208), .Z(n43210) );
  NOR U56055 ( .A(n49775), .B(n43210), .Z(n43211) );
  IV U56056 ( .A(n43211), .Z(n46400) );
  XOR U56057 ( .A(n45384), .B(n46400), .Z(n46397) );
  XOR U56058 ( .A(n46396), .B(n46397), .Z(n45380) );
  XOR U56059 ( .A(n43212), .B(n45380), .Z(n45379) );
  XOR U56060 ( .A(n45377), .B(n45379), .Z(n45374) );
  IV U56061 ( .A(n43213), .Z(n43214) );
  NOR U56062 ( .A(n43215), .B(n43214), .Z(n45372) );
  XOR U56063 ( .A(n45374), .B(n45372), .Z(n45370) );
  XOR U56064 ( .A(n45369), .B(n45370), .Z(n45367) );
  XOR U56065 ( .A(n45366), .B(n45367), .Z(n45361) );
  XOR U56066 ( .A(n45362), .B(n45361), .Z(n45359) );
  IV U56067 ( .A(n43216), .Z(n43217) );
  NOR U56068 ( .A(n43218), .B(n43217), .Z(n45363) );
  IV U56069 ( .A(n43219), .Z(n43220) );
  NOR U56070 ( .A(n43221), .B(n43220), .Z(n45358) );
  NOR U56071 ( .A(n45363), .B(n45358), .Z(n43222) );
  XOR U56072 ( .A(n45359), .B(n43222), .Z(n45357) );
  NOR U56073 ( .A(n43224), .B(n43223), .Z(n43225) );
  IV U56074 ( .A(n43225), .Z(n43233) );
  IV U56075 ( .A(n43226), .Z(n43230) );
  XOR U56076 ( .A(n43228), .B(n43227), .Z(n43229) );
  NOR U56077 ( .A(n43230), .B(n43229), .Z(n43231) );
  IV U56078 ( .A(n43231), .Z(n43232) );
  NOR U56079 ( .A(n43233), .B(n43232), .Z(n45355) );
  XOR U56080 ( .A(n45357), .B(n45355), .Z(n46419) );
  XOR U56081 ( .A(n46418), .B(n46419), .Z(n46431) );
  NOR U56082 ( .A(n43234), .B(n46411), .Z(n43238) );
  IV U56083 ( .A(n43235), .Z(n43237) );
  IV U56084 ( .A(n43236), .Z(n43241) );
  NOR U56085 ( .A(n43237), .B(n43241), .Z(n46430) );
  NOR U56086 ( .A(n43238), .B(n46430), .Z(n43239) );
  XOR U56087 ( .A(n46431), .B(n43239), .Z(n45349) );
  IV U56088 ( .A(n43240), .Z(n43242) );
  NOR U56089 ( .A(n43242), .B(n43241), .Z(n45352) );
  IV U56090 ( .A(n43243), .Z(n43245) );
  NOR U56091 ( .A(n43245), .B(n43244), .Z(n45350) );
  NOR U56092 ( .A(n45352), .B(n45350), .Z(n43246) );
  XOR U56093 ( .A(n45349), .B(n43246), .Z(n45347) );
  XOR U56094 ( .A(n45346), .B(n45347), .Z(n46437) );
  XOR U56095 ( .A(n46435), .B(n46437), .Z(n46440) );
  XOR U56096 ( .A(n43247), .B(n46440), .Z(n43248) );
  IV U56097 ( .A(n43248), .Z(n45339) );
  IV U56098 ( .A(n43249), .Z(n43250) );
  NOR U56099 ( .A(n43251), .B(n43250), .Z(n45337) );
  XOR U56100 ( .A(n45339), .B(n45337), .Z(n45342) );
  IV U56101 ( .A(n43252), .Z(n43254) );
  IV U56102 ( .A(n43253), .Z(n43256) );
  NOR U56103 ( .A(n43254), .B(n43256), .Z(n45340) );
  XOR U56104 ( .A(n45342), .B(n45340), .Z(n45335) );
  IV U56105 ( .A(n43255), .Z(n43257) );
  NOR U56106 ( .A(n43257), .B(n43256), .Z(n45333) );
  XOR U56107 ( .A(n45335), .B(n45333), .Z(n45331) );
  XOR U56108 ( .A(n45329), .B(n45331), .Z(n46446) );
  IV U56109 ( .A(n43258), .Z(n43259) );
  NOR U56110 ( .A(n43260), .B(n43259), .Z(n45330) );
  NOR U56111 ( .A(n43262), .B(n43261), .Z(n46445) );
  NOR U56112 ( .A(n45330), .B(n46445), .Z(n43263) );
  XOR U56113 ( .A(n46446), .B(n43263), .Z(n46457) );
  XOR U56114 ( .A(n46449), .B(n46457), .Z(n46452) );
  XOR U56115 ( .A(n43264), .B(n46452), .Z(n48854) );
  XOR U56116 ( .A(n45323), .B(n48854), .Z(n45325) );
  XOR U56117 ( .A(n45326), .B(n45325), .Z(n45318) );
  IV U56118 ( .A(n43265), .Z(n43266) );
  NOR U56119 ( .A(n43267), .B(n43266), .Z(n45321) );
  IV U56120 ( .A(n43268), .Z(n43270) );
  NOR U56121 ( .A(n43270), .B(n43269), .Z(n45317) );
  NOR U56122 ( .A(n45321), .B(n45317), .Z(n43271) );
  XOR U56123 ( .A(n45318), .B(n43271), .Z(n45316) );
  XOR U56124 ( .A(n45314), .B(n45316), .Z(n46460) );
  XOR U56125 ( .A(n46459), .B(n46460), .Z(n46464) );
  XOR U56126 ( .A(n46462), .B(n46464), .Z(n45310) );
  XOR U56127 ( .A(n45308), .B(n45310), .Z(n45313) );
  XOR U56128 ( .A(n45311), .B(n45313), .Z(n45307) );
  XOR U56129 ( .A(n43272), .B(n45307), .Z(n45303) );
  XOR U56130 ( .A(n45302), .B(n45303), .Z(n46470) );
  XOR U56131 ( .A(n46469), .B(n46470), .Z(n46474) );
  IV U56132 ( .A(n43273), .Z(n43274) );
  NOR U56133 ( .A(n43275), .B(n43274), .Z(n45295) );
  IV U56134 ( .A(n43276), .Z(n43278) );
  NOR U56135 ( .A(n43278), .B(n43277), .Z(n46472) );
  NOR U56136 ( .A(n45295), .B(n46472), .Z(n43279) );
  XOR U56137 ( .A(n46474), .B(n43279), .Z(n45298) );
  XOR U56138 ( .A(n43280), .B(n45298), .Z(n46478) );
  XOR U56139 ( .A(n46476), .B(n46478), .Z(n46485) );
  IV U56140 ( .A(n46485), .Z(n43289) );
  IV U56141 ( .A(n43281), .Z(n43282) );
  NOR U56142 ( .A(n43283), .B(n43282), .Z(n46484) );
  NOR U56143 ( .A(n43285), .B(n43284), .Z(n45293) );
  NOR U56144 ( .A(n46484), .B(n45293), .Z(n43286) );
  IV U56145 ( .A(n43286), .Z(n43287) );
  NOR U56146 ( .A(n45291), .B(n43287), .Z(n43288) );
  XOR U56147 ( .A(n43289), .B(n43288), .Z(n45290) );
  IV U56148 ( .A(n43290), .Z(n43292) );
  IV U56149 ( .A(n43291), .Z(n43304) );
  NOR U56150 ( .A(n43292), .B(n43304), .Z(n43293) );
  IV U56151 ( .A(n43293), .Z(n45289) );
  XOR U56152 ( .A(n45290), .B(n45289), .Z(n48808) );
  NOR U56153 ( .A(n43295), .B(n43294), .Z(n43296) );
  IV U56154 ( .A(n43296), .Z(n43302) );
  IV U56155 ( .A(n43297), .Z(n43299) );
  NOR U56156 ( .A(n43299), .B(n43298), .Z(n43300) );
  IV U56157 ( .A(n43300), .Z(n43301) );
  NOR U56158 ( .A(n43302), .B(n43301), .Z(n49914) );
  IV U56159 ( .A(n43303), .Z(n43305) );
  NOR U56160 ( .A(n43305), .B(n43304), .Z(n48824) );
  NOR U56161 ( .A(n49914), .B(n48824), .Z(n48806) );
  XOR U56162 ( .A(n48808), .B(n48806), .Z(n45286) );
  XOR U56163 ( .A(n45284), .B(n45286), .Z(n48799) );
  XOR U56164 ( .A(n43306), .B(n48799), .Z(n46491) );
  IV U56165 ( .A(n43307), .Z(n43308) );
  NOR U56166 ( .A(n43309), .B(n43308), .Z(n46489) );
  XOR U56167 ( .A(n46491), .B(n46489), .Z(n46493) );
  IV U56168 ( .A(n43310), .Z(n43311) );
  NOR U56169 ( .A(n43312), .B(n43311), .Z(n45282) );
  IV U56170 ( .A(n43313), .Z(n43315) );
  NOR U56171 ( .A(n43315), .B(n43314), .Z(n46492) );
  NOR U56172 ( .A(n45282), .B(n46492), .Z(n43316) );
  XOR U56173 ( .A(n46493), .B(n43316), .Z(n45278) );
  NOR U56174 ( .A(n43318), .B(n43317), .Z(n45279) );
  IV U56175 ( .A(n43319), .Z(n43321) );
  IV U56176 ( .A(n43320), .Z(n43325) );
  NOR U56177 ( .A(n43321), .B(n43325), .Z(n46501) );
  NOR U56178 ( .A(n45279), .B(n46501), .Z(n43322) );
  XOR U56179 ( .A(n45278), .B(n43322), .Z(n46507) );
  IV U56180 ( .A(n43323), .Z(n43324) );
  NOR U56181 ( .A(n43325), .B(n43324), .Z(n46504) );
  IV U56182 ( .A(n43326), .Z(n43327) );
  NOR U56183 ( .A(n43328), .B(n43327), .Z(n46506) );
  NOR U56184 ( .A(n46504), .B(n46506), .Z(n43329) );
  XOR U56185 ( .A(n46507), .B(n43329), .Z(n43330) );
  IV U56186 ( .A(n43330), .Z(n45276) );
  XOR U56187 ( .A(n45274), .B(n45276), .Z(n45270) );
  XOR U56188 ( .A(n45268), .B(n45270), .Z(n45272) );
  XOR U56189 ( .A(n45271), .B(n45272), .Z(n46512) );
  XOR U56190 ( .A(n43331), .B(n46512), .Z(n45265) );
  XOR U56191 ( .A(n45263), .B(n45265), .Z(n46517) );
  XOR U56192 ( .A(n46516), .B(n46517), .Z(n45262) );
  IV U56193 ( .A(n43332), .Z(n43336) );
  NOR U56194 ( .A(n43333), .B(n43338), .Z(n43334) );
  IV U56195 ( .A(n43334), .Z(n43335) );
  NOR U56196 ( .A(n43336), .B(n43335), .Z(n45260) );
  XOR U56197 ( .A(n45262), .B(n45260), .Z(n46522) );
  XOR U56198 ( .A(n46523), .B(n46522), .Z(n46525) );
  IV U56199 ( .A(n43337), .Z(n43339) );
  NOR U56200 ( .A(n43339), .B(n43338), .Z(n46524) );
  NOR U56201 ( .A(n43341), .B(n43340), .Z(n46531) );
  NOR U56202 ( .A(n46524), .B(n46531), .Z(n43342) );
  XOR U56203 ( .A(n46525), .B(n43342), .Z(n46530) );
  IV U56204 ( .A(n43343), .Z(n43344) );
  NOR U56205 ( .A(n43345), .B(n43344), .Z(n45258) );
  NOR U56206 ( .A(n46528), .B(n45258), .Z(n43346) );
  XOR U56207 ( .A(n46530), .B(n43346), .Z(n43347) );
  NOR U56208 ( .A(n43348), .B(n43347), .Z(n43351) );
  IV U56209 ( .A(n43348), .Z(n43350) );
  XOR U56210 ( .A(n46528), .B(n46530), .Z(n43349) );
  NOR U56211 ( .A(n43350), .B(n43349), .Z(n49952) );
  NOR U56212 ( .A(n43351), .B(n49952), .Z(n46534) );
  NOR U56213 ( .A(n43353), .B(n43352), .Z(n43354) );
  IV U56214 ( .A(n43354), .Z(n46535) );
  XOR U56215 ( .A(n46534), .B(n46535), .Z(n45257) );
  XOR U56216 ( .A(n45255), .B(n45257), .Z(n45250) );
  XOR U56217 ( .A(n45249), .B(n45250), .Z(n45253) );
  XOR U56218 ( .A(n45252), .B(n45253), .Z(n48772) );
  XOR U56219 ( .A(n43355), .B(n48772), .Z(n46539) );
  XOR U56220 ( .A(n46538), .B(n46539), .Z(n45247) );
  XOR U56221 ( .A(n45246), .B(n45247), .Z(n45241) );
  XOR U56222 ( .A(n45240), .B(n45241), .Z(n45245) );
  IV U56223 ( .A(n43356), .Z(n43357) );
  NOR U56224 ( .A(n43357), .B(n43359), .Z(n45243) );
  XOR U56225 ( .A(n45245), .B(n45243), .Z(n48758) );
  IV U56226 ( .A(n43358), .Z(n43360) );
  NOR U56227 ( .A(n43360), .B(n43359), .Z(n48762) );
  IV U56228 ( .A(n43361), .Z(n43362) );
  NOR U56229 ( .A(n43363), .B(n43362), .Z(n48757) );
  NOR U56230 ( .A(n48762), .B(n48757), .Z(n45235) );
  XOR U56231 ( .A(n48758), .B(n45235), .Z(n45236) );
  XOR U56232 ( .A(n45237), .B(n45236), .Z(n48746) );
  IV U56233 ( .A(n43364), .Z(n43366) );
  NOR U56234 ( .A(n43366), .B(n43365), .Z(n53894) );
  NOR U56235 ( .A(n52508), .B(n53894), .Z(n48748) );
  XOR U56236 ( .A(n48746), .B(n48748), .Z(n43367) );
  IV U56237 ( .A(n43367), .Z(n45231) );
  XOR U56238 ( .A(n45230), .B(n45231), .Z(n46548) );
  XOR U56239 ( .A(n43368), .B(n46548), .Z(n45227) );
  XOR U56240 ( .A(n45226), .B(n45227), .Z(n46554) );
  IV U56241 ( .A(n43369), .Z(n43370) );
  NOR U56242 ( .A(n43371), .B(n43370), .Z(n46561) );
  NOR U56243 ( .A(n43372), .B(n46555), .Z(n43373) );
  NOR U56244 ( .A(n46561), .B(n43373), .Z(n43374) );
  XOR U56245 ( .A(n46554), .B(n43374), .Z(n45225) );
  XOR U56246 ( .A(n45223), .B(n45225), .Z(n46570) );
  XOR U56247 ( .A(n46569), .B(n46570), .Z(n49990) );
  XOR U56248 ( .A(n49992), .B(n49990), .Z(n43375) );
  IV U56249 ( .A(n43375), .Z(n45222) );
  IV U56250 ( .A(n43376), .Z(n43378) );
  NOR U56251 ( .A(n43378), .B(n43377), .Z(n45220) );
  XOR U56252 ( .A(n45222), .B(n45220), .Z(n46580) );
  IV U56253 ( .A(n43379), .Z(n43381) );
  NOR U56254 ( .A(n43381), .B(n43380), .Z(n43382) );
  IV U56255 ( .A(n43382), .Z(n46579) );
  XOR U56256 ( .A(n46580), .B(n46579), .Z(n46575) );
  IV U56257 ( .A(n43383), .Z(n43384) );
  NOR U56258 ( .A(n43385), .B(n43384), .Z(n46574) );
  NOR U56259 ( .A(n43386), .B(n46587), .Z(n43387) );
  NOR U56260 ( .A(n46574), .B(n43387), .Z(n43388) );
  XOR U56261 ( .A(n46575), .B(n43388), .Z(n46592) );
  XOR U56262 ( .A(n46590), .B(n46592), .Z(n48714) );
  XOR U56263 ( .A(n43389), .B(n48714), .Z(n45214) );
  XOR U56264 ( .A(n45215), .B(n45214), .Z(n45213) );
  NOR U56265 ( .A(n43390), .B(n45213), .Z(n50056) );
  NOR U56266 ( .A(n43397), .B(n50056), .Z(n45209) );
  IV U56267 ( .A(n45209), .Z(n43396) );
  IV U56268 ( .A(n43391), .Z(n43393) );
  NOR U56269 ( .A(n43393), .B(n43392), .Z(n43394) );
  IV U56270 ( .A(n43394), .Z(n45212) );
  XOR U56271 ( .A(n45213), .B(n45212), .Z(n43398) );
  NOR U56272 ( .A(n43395), .B(n43398), .Z(n45210) );
  NOR U56273 ( .A(n43396), .B(n45210), .Z(n43401) );
  IV U56274 ( .A(n43397), .Z(n43399) );
  NOR U56275 ( .A(n43399), .B(n43398), .Z(n43400) );
  NOR U56276 ( .A(n43401), .B(n43400), .Z(n46601) );
  NOR U56277 ( .A(n43403), .B(n43402), .Z(n43404) );
  IV U56278 ( .A(n43404), .Z(n46600) );
  XOR U56279 ( .A(n46601), .B(n46600), .Z(n46603) );
  IV U56280 ( .A(n43405), .Z(n43406) );
  NOR U56281 ( .A(n43407), .B(n43406), .Z(n46602) );
  IV U56282 ( .A(n43408), .Z(n43409) );
  NOR U56283 ( .A(n43409), .B(n43413), .Z(n46606) );
  NOR U56284 ( .A(n46602), .B(n46606), .Z(n43410) );
  XOR U56285 ( .A(n46603), .B(n43410), .Z(n45204) );
  IV U56286 ( .A(n43411), .Z(n43412) );
  NOR U56287 ( .A(n43413), .B(n43412), .Z(n45202) );
  XOR U56288 ( .A(n45204), .B(n45202), .Z(n45207) );
  XOR U56289 ( .A(n45205), .B(n45207), .Z(n45201) );
  NOR U56290 ( .A(n43421), .B(n45201), .Z(n50068) );
  IV U56291 ( .A(n43414), .Z(n43416) );
  NOR U56292 ( .A(n43416), .B(n43415), .Z(n45195) );
  IV U56293 ( .A(n43417), .Z(n43418) );
  NOR U56294 ( .A(n43419), .B(n43418), .Z(n43420) );
  IV U56295 ( .A(n43420), .Z(n45200) );
  XOR U56296 ( .A(n45201), .B(n45200), .Z(n45196) );
  XOR U56297 ( .A(n45195), .B(n45196), .Z(n43423) );
  NOR U56298 ( .A(n45196), .B(n43421), .Z(n43422) );
  NOR U56299 ( .A(n43423), .B(n43422), .Z(n43424) );
  NOR U56300 ( .A(n50068), .B(n43424), .Z(n43425) );
  IV U56301 ( .A(n43425), .Z(n46611) );
  XOR U56302 ( .A(n46610), .B(n46611), .Z(n46615) );
  XOR U56303 ( .A(n46613), .B(n46615), .Z(n45194) );
  XOR U56304 ( .A(n45192), .B(n45194), .Z(n45187) );
  XOR U56305 ( .A(n45186), .B(n45187), .Z(n45184) );
  XOR U56306 ( .A(n45183), .B(n45184), .Z(n45181) );
  XOR U56307 ( .A(n45180), .B(n45181), .Z(n45178) );
  XOR U56308 ( .A(n45176), .B(n45178), .Z(n46620) );
  XOR U56309 ( .A(n46618), .B(n46620), .Z(n46626) );
  XOR U56310 ( .A(n43426), .B(n46626), .Z(n45170) );
  IV U56311 ( .A(n43427), .Z(n43429) );
  NOR U56312 ( .A(n43429), .B(n43428), .Z(n45171) );
  IV U56313 ( .A(n43430), .Z(n43432) );
  NOR U56314 ( .A(n43432), .B(n43431), .Z(n45173) );
  NOR U56315 ( .A(n45171), .B(n45173), .Z(n43433) );
  XOR U56316 ( .A(n45170), .B(n43433), .Z(n48665) );
  IV U56317 ( .A(n43434), .Z(n48668) );
  NOR U56318 ( .A(n48668), .B(n43435), .Z(n46633) );
  IV U56319 ( .A(n43436), .Z(n43437) );
  NOR U56320 ( .A(n43438), .B(n43437), .Z(n46631) );
  NOR U56321 ( .A(n46633), .B(n46631), .Z(n43439) );
  XOR U56322 ( .A(n48665), .B(n43439), .Z(n45167) );
  XOR U56323 ( .A(n43440), .B(n45167), .Z(n46644) );
  XOR U56324 ( .A(n46642), .B(n46644), .Z(n45164) );
  NOR U56325 ( .A(n43441), .B(n45160), .Z(n43444) );
  IV U56326 ( .A(n43442), .Z(n43443) );
  NOR U56327 ( .A(n43443), .B(n43447), .Z(n45163) );
  NOR U56328 ( .A(n43444), .B(n45163), .Z(n43445) );
  XOR U56329 ( .A(n45164), .B(n43445), .Z(n45156) );
  IV U56330 ( .A(n43446), .Z(n43448) );
  NOR U56331 ( .A(n43448), .B(n43447), .Z(n45157) );
  NOR U56332 ( .A(n43450), .B(n43449), .Z(n46651) );
  NOR U56333 ( .A(n45157), .B(n46651), .Z(n43451) );
  XOR U56334 ( .A(n45156), .B(n43451), .Z(n46656) );
  IV U56335 ( .A(n43452), .Z(n43454) );
  NOR U56336 ( .A(n43454), .B(n43453), .Z(n46654) );
  NOR U56337 ( .A(n45154), .B(n46654), .Z(n43455) );
  XOR U56338 ( .A(n46656), .B(n43455), .Z(n43456) );
  IV U56339 ( .A(n43456), .Z(n46658) );
  XOR U56340 ( .A(n46657), .B(n46658), .Z(n46669) );
  XOR U56341 ( .A(n46668), .B(n46669), .Z(n46663) );
  XOR U56342 ( .A(n46661), .B(n46663), .Z(n46667) );
  XOR U56343 ( .A(n46665), .B(n46667), .Z(n46677) );
  XOR U56344 ( .A(n46676), .B(n46677), .Z(n46681) );
  XOR U56345 ( .A(n46679), .B(n46681), .Z(n48638) );
  XOR U56346 ( .A(n45153), .B(n48638), .Z(n45141) );
  XOR U56347 ( .A(n43457), .B(n45141), .Z(n43458) );
  XOR U56348 ( .A(n45148), .B(n43458), .Z(n45138) );
  XOR U56349 ( .A(n45137), .B(n45138), .Z(n45133) );
  IV U56350 ( .A(n43459), .Z(n43461) );
  NOR U56351 ( .A(n43461), .B(n43460), .Z(n45131) );
  XOR U56352 ( .A(n45133), .B(n45131), .Z(n45136) );
  IV U56353 ( .A(n43462), .Z(n43467) );
  IV U56354 ( .A(n43463), .Z(n43464) );
  NOR U56355 ( .A(n43467), .B(n43464), .Z(n45134) );
  XOR U56356 ( .A(n45136), .B(n45134), .Z(n46688) );
  IV U56357 ( .A(n43465), .Z(n43466) );
  NOR U56358 ( .A(n43467), .B(n43466), .Z(n46686) );
  XOR U56359 ( .A(n46688), .B(n46686), .Z(n46690) );
  XOR U56360 ( .A(n46689), .B(n46690), .Z(n45125) );
  XOR U56361 ( .A(n45124), .B(n45125), .Z(n45128) );
  XOR U56362 ( .A(n45127), .B(n45128), .Z(n46701) );
  IV U56363 ( .A(n43468), .Z(n43470) );
  NOR U56364 ( .A(n43470), .B(n43469), .Z(n46699) );
  XOR U56365 ( .A(n46701), .B(n46699), .Z(n46695) );
  XOR U56366 ( .A(n46694), .B(n46695), .Z(n48622) );
  IV U56367 ( .A(n43471), .Z(n43472) );
  NOR U56368 ( .A(n43473), .B(n43472), .Z(n50158) );
  IV U56369 ( .A(n43474), .Z(n43476) );
  NOR U56370 ( .A(n43476), .B(n43475), .Z(n48619) );
  NOR U56371 ( .A(n50158), .B(n48619), .Z(n45123) );
  XOR U56372 ( .A(n48622), .B(n45123), .Z(n45118) );
  XOR U56373 ( .A(n43477), .B(n45118), .Z(n48609) );
  IV U56374 ( .A(n43478), .Z(n43479) );
  NOR U56375 ( .A(n43479), .B(n43481), .Z(n50163) );
  IV U56376 ( .A(n43480), .Z(n43482) );
  NOR U56377 ( .A(n43482), .B(n43481), .Z(n48608) );
  NOR U56378 ( .A(n50163), .B(n48608), .Z(n45116) );
  XOR U56379 ( .A(n48609), .B(n45116), .Z(n43483) );
  IV U56380 ( .A(n43483), .Z(n45111) );
  XOR U56381 ( .A(n45110), .B(n45111), .Z(n45114) );
  XOR U56382 ( .A(n43484), .B(n45114), .Z(n45107) );
  XOR U56383 ( .A(n45106), .B(n45107), .Z(n45100) );
  IV U56384 ( .A(n43485), .Z(n43486) );
  NOR U56385 ( .A(n43487), .B(n43486), .Z(n45099) );
  IV U56386 ( .A(n43488), .Z(n43493) );
  NOR U56387 ( .A(n43490), .B(n43489), .Z(n43491) );
  IV U56388 ( .A(n43491), .Z(n43492) );
  NOR U56389 ( .A(n43493), .B(n43492), .Z(n45103) );
  NOR U56390 ( .A(n45099), .B(n45103), .Z(n43494) );
  XOR U56391 ( .A(n45100), .B(n43494), .Z(n45098) );
  XOR U56392 ( .A(n45096), .B(n45098), .Z(n52360) );
  XOR U56393 ( .A(n43495), .B(n52360), .Z(n46715) );
  XOR U56394 ( .A(n46714), .B(n46715), .Z(n46717) );
  XOR U56395 ( .A(n46718), .B(n46717), .Z(n45091) );
  IV U56396 ( .A(n43496), .Z(n43498) );
  NOR U56397 ( .A(n43498), .B(n43497), .Z(n46720) );
  IV U56398 ( .A(n43499), .Z(n43500) );
  NOR U56399 ( .A(n43500), .B(n43503), .Z(n45092) );
  NOR U56400 ( .A(n46720), .B(n45092), .Z(n43501) );
  XOR U56401 ( .A(n45091), .B(n43501), .Z(n45086) );
  IV U56402 ( .A(n43502), .Z(n43504) );
  NOR U56403 ( .A(n43504), .B(n43503), .Z(n45084) );
  XOR U56404 ( .A(n45086), .B(n45084), .Z(n46725) );
  XOR U56405 ( .A(n43505), .B(n46725), .Z(n46729) );
  XOR U56406 ( .A(n46727), .B(n46729), .Z(n46732) );
  IV U56407 ( .A(n43506), .Z(n43510) );
  XOR U56408 ( .A(n43508), .B(n43507), .Z(n43509) );
  NOR U56409 ( .A(n43510), .B(n43509), .Z(n46730) );
  XOR U56410 ( .A(n46732), .B(n46730), .Z(n46736) );
  IV U56411 ( .A(n43511), .Z(n43514) );
  IV U56412 ( .A(n43512), .Z(n43513) );
  NOR U56413 ( .A(n43514), .B(n43513), .Z(n46734) );
  XOR U56414 ( .A(n46736), .B(n46734), .Z(n46739) );
  IV U56415 ( .A(n43515), .Z(n43517) );
  NOR U56416 ( .A(n43517), .B(n43516), .Z(n46737) );
  XOR U56417 ( .A(n46739), .B(n46737), .Z(n45074) );
  XOR U56418 ( .A(n45073), .B(n45074), .Z(n46742) );
  IV U56419 ( .A(n43518), .Z(n43519) );
  NOR U56420 ( .A(n43520), .B(n43519), .Z(n43521) );
  IV U56421 ( .A(n43521), .Z(n46741) );
  XOR U56422 ( .A(n46742), .B(n46741), .Z(n46743) );
  IV U56423 ( .A(n43522), .Z(n43524) );
  IV U56424 ( .A(n43523), .Z(n43530) );
  NOR U56425 ( .A(n43524), .B(n43530), .Z(n46747) );
  IV U56426 ( .A(n43525), .Z(n43526) );
  NOR U56427 ( .A(n43527), .B(n43526), .Z(n46744) );
  NOR U56428 ( .A(n46747), .B(n46744), .Z(n43528) );
  XOR U56429 ( .A(n46743), .B(n43528), .Z(n46754) );
  IV U56430 ( .A(n43529), .Z(n43531) );
  NOR U56431 ( .A(n43531), .B(n43530), .Z(n46752) );
  XOR U56432 ( .A(n46754), .B(n46752), .Z(n45071) );
  XOR U56433 ( .A(n43532), .B(n45071), .Z(n46758) );
  XOR U56434 ( .A(n46759), .B(n46758), .Z(n46761) );
  NOR U56435 ( .A(n43534), .B(n43533), .Z(n46760) );
  IV U56436 ( .A(n43535), .Z(n43541) );
  IV U56437 ( .A(n43536), .Z(n43537) );
  NOR U56438 ( .A(n43541), .B(n43537), .Z(n46767) );
  NOR U56439 ( .A(n46760), .B(n46767), .Z(n43538) );
  XOR U56440 ( .A(n46761), .B(n43538), .Z(n46766) );
  IV U56441 ( .A(n43539), .Z(n43540) );
  NOR U56442 ( .A(n43541), .B(n43540), .Z(n46764) );
  XOR U56443 ( .A(n46766), .B(n46764), .Z(n48547) );
  XOR U56444 ( .A(n45066), .B(n48547), .Z(n43542) );
  IV U56445 ( .A(n43542), .Z(n46774) );
  IV U56446 ( .A(n43543), .Z(n43544) );
  NOR U56447 ( .A(n43544), .B(n43549), .Z(n46772) );
  XOR U56448 ( .A(n46774), .B(n46772), .Z(n46777) );
  IV U56449 ( .A(n43545), .Z(n43546) );
  NOR U56450 ( .A(n43547), .B(n43546), .Z(n45064) );
  IV U56451 ( .A(n43548), .Z(n43550) );
  NOR U56452 ( .A(n43550), .B(n43549), .Z(n46775) );
  NOR U56453 ( .A(n45064), .B(n46775), .Z(n43551) );
  XOR U56454 ( .A(n46777), .B(n43551), .Z(n45057) );
  XOR U56455 ( .A(n45058), .B(n45057), .Z(n45061) );
  IV U56456 ( .A(n43552), .Z(n43553) );
  NOR U56457 ( .A(n43553), .B(n43555), .Z(n45059) );
  XOR U56458 ( .A(n45061), .B(n45059), .Z(n45055) );
  IV U56459 ( .A(n43554), .Z(n43558) );
  NOR U56460 ( .A(n43556), .B(n43555), .Z(n43557) );
  IV U56461 ( .A(n43557), .Z(n43560) );
  NOR U56462 ( .A(n43558), .B(n43560), .Z(n45053) );
  XOR U56463 ( .A(n45055), .B(n45053), .Z(n46783) );
  IV U56464 ( .A(n43559), .Z(n43561) );
  NOR U56465 ( .A(n43561), .B(n43560), .Z(n46781) );
  XOR U56466 ( .A(n46783), .B(n46781), .Z(n46785) );
  IV U56467 ( .A(n43562), .Z(n43565) );
  NOR U56468 ( .A(n43572), .B(n43563), .Z(n43564) );
  IV U56469 ( .A(n43564), .Z(n43568) );
  NOR U56470 ( .A(n43565), .B(n43568), .Z(n43566) );
  IV U56471 ( .A(n43566), .Z(n46784) );
  XOR U56472 ( .A(n46785), .B(n46784), .Z(n45050) );
  IV U56473 ( .A(n43567), .Z(n43569) );
  NOR U56474 ( .A(n43569), .B(n43568), .Z(n46787) );
  IV U56475 ( .A(n43570), .Z(n43574) );
  NOR U56476 ( .A(n43572), .B(n43571), .Z(n43573) );
  IV U56477 ( .A(n43573), .Z(n43577) );
  NOR U56478 ( .A(n43574), .B(n43577), .Z(n45051) );
  NOR U56479 ( .A(n46787), .B(n45051), .Z(n43575) );
  XOR U56480 ( .A(n45050), .B(n43575), .Z(n45049) );
  IV U56481 ( .A(n43576), .Z(n43578) );
  NOR U56482 ( .A(n43578), .B(n43577), .Z(n45047) );
  XOR U56483 ( .A(n45049), .B(n45047), .Z(n46792) );
  XOR U56484 ( .A(n46790), .B(n46792), .Z(n46794) );
  XOR U56485 ( .A(n46793), .B(n46794), .Z(n46798) );
  XOR U56486 ( .A(n43579), .B(n46798), .Z(n46801) );
  XOR U56487 ( .A(n46802), .B(n46801), .Z(n46804) );
  XOR U56488 ( .A(n46803), .B(n46804), .Z(n45042) );
  XOR U56489 ( .A(n45041), .B(n45042), .Z(n45038) );
  XOR U56490 ( .A(n45035), .B(n45038), .Z(n45032) );
  XOR U56491 ( .A(n43580), .B(n45032), .Z(n46811) );
  XOR U56492 ( .A(n46809), .B(n46811), .Z(n46813) );
  XOR U56493 ( .A(n46812), .B(n46813), .Z(n46817) );
  IV U56494 ( .A(n43581), .Z(n43583) );
  NOR U56495 ( .A(n43583), .B(n43582), .Z(n46816) );
  IV U56496 ( .A(n43584), .Z(n43586) );
  NOR U56497 ( .A(n43586), .B(n43585), .Z(n45029) );
  NOR U56498 ( .A(n46816), .B(n45029), .Z(n43587) );
  XOR U56499 ( .A(n46817), .B(n43587), .Z(n45023) );
  IV U56500 ( .A(n43588), .Z(n43589) );
  NOR U56501 ( .A(n43590), .B(n43589), .Z(n45026) );
  IV U56502 ( .A(n43591), .Z(n43592) );
  NOR U56503 ( .A(n43593), .B(n43592), .Z(n45024) );
  NOR U56504 ( .A(n45026), .B(n45024), .Z(n43594) );
  XOR U56505 ( .A(n45023), .B(n43594), .Z(n45021) );
  XOR U56506 ( .A(n45022), .B(n45021), .Z(n45016) );
  IV U56507 ( .A(n43595), .Z(n43596) );
  NOR U56508 ( .A(n43597), .B(n43596), .Z(n45019) );
  IV U56509 ( .A(n43598), .Z(n43599) );
  NOR U56510 ( .A(n43600), .B(n43599), .Z(n45015) );
  NOR U56511 ( .A(n45019), .B(n45015), .Z(n43601) );
  XOR U56512 ( .A(n45016), .B(n43601), .Z(n45014) );
  IV U56513 ( .A(n43602), .Z(n43604) );
  NOR U56514 ( .A(n43604), .B(n43603), .Z(n45012) );
  XOR U56515 ( .A(n45014), .B(n45012), .Z(n45009) );
  XOR U56516 ( .A(n45007), .B(n45009), .Z(n45010) );
  NOR U56517 ( .A(n43612), .B(n45010), .Z(n50253) );
  IV U56518 ( .A(n43605), .Z(n43607) );
  NOR U56519 ( .A(n43607), .B(n43606), .Z(n45000) );
  IV U56520 ( .A(n43608), .Z(n43609) );
  NOR U56521 ( .A(n43610), .B(n43609), .Z(n43611) );
  IV U56522 ( .A(n43611), .Z(n45011) );
  XOR U56523 ( .A(n45011), .B(n45010), .Z(n45001) );
  XOR U56524 ( .A(n45000), .B(n45001), .Z(n43614) );
  NOR U56525 ( .A(n45001), .B(n43612), .Z(n43613) );
  NOR U56526 ( .A(n43614), .B(n43613), .Z(n43615) );
  NOR U56527 ( .A(n50253), .B(n43615), .Z(n45004) );
  XOR U56528 ( .A(n45006), .B(n45004), .Z(n52196) );
  XOR U56529 ( .A(n44998), .B(n52196), .Z(n43616) );
  IV U56530 ( .A(n43616), .Z(n46824) );
  XOR U56531 ( .A(n46822), .B(n46824), .Z(n46826) );
  XOR U56532 ( .A(n46825), .B(n46826), .Z(n46840) );
  XOR U56533 ( .A(n46838), .B(n46840), .Z(n44995) );
  XOR U56534 ( .A(n43617), .B(n44995), .Z(n44992) );
  XOR U56535 ( .A(n44991), .B(n44992), .Z(n44980) );
  NOR U56536 ( .A(n43618), .B(n44985), .Z(n43622) );
  IV U56537 ( .A(n43619), .Z(n43621) );
  IV U56538 ( .A(n43620), .Z(n43626) );
  NOR U56539 ( .A(n43621), .B(n43626), .Z(n44981) );
  NOR U56540 ( .A(n43622), .B(n44981), .Z(n43623) );
  XOR U56541 ( .A(n44980), .B(n43623), .Z(n46846) );
  IV U56542 ( .A(n43624), .Z(n43625) );
  NOR U56543 ( .A(n43626), .B(n43625), .Z(n46844) );
  XOR U56544 ( .A(n46846), .B(n46844), .Z(n44978) );
  XOR U56545 ( .A(n44977), .B(n44978), .Z(n48447) );
  XOR U56546 ( .A(n46850), .B(n48447), .Z(n46851) );
  IV U56547 ( .A(n43627), .Z(n43628) );
  NOR U56548 ( .A(n43629), .B(n43628), .Z(n48435) );
  IV U56549 ( .A(n43630), .Z(n43632) );
  NOR U56550 ( .A(n43632), .B(n43631), .Z(n48441) );
  NOR U56551 ( .A(n48435), .B(n48441), .Z(n46852) );
  XOR U56552 ( .A(n46851), .B(n46852), .Z(n46857) );
  XOR U56553 ( .A(n46856), .B(n46857), .Z(n46860) );
  XOR U56554 ( .A(n43633), .B(n46860), .Z(n44968) );
  XOR U56555 ( .A(n44969), .B(n44968), .Z(n44970) );
  XOR U56556 ( .A(n44971), .B(n44970), .Z(n43634) );
  IV U56557 ( .A(n43634), .Z(n46875) );
  IV U56558 ( .A(n43635), .Z(n43638) );
  IV U56559 ( .A(n43636), .Z(n43637) );
  NOR U56560 ( .A(n43638), .B(n43637), .Z(n46873) );
  XOR U56561 ( .A(n46875), .B(n46873), .Z(n46878) );
  IV U56562 ( .A(n43639), .Z(n43640) );
  NOR U56563 ( .A(n43640), .B(n54159), .Z(n46876) );
  XOR U56564 ( .A(n46878), .B(n46876), .Z(n44966) );
  IV U56565 ( .A(n43641), .Z(n43642) );
  NOR U56566 ( .A(n43643), .B(n43642), .Z(n44965) );
  IV U56567 ( .A(n43644), .Z(n43646) );
  NOR U56568 ( .A(n43646), .B(n43645), .Z(n44963) );
  NOR U56569 ( .A(n44965), .B(n44963), .Z(n43647) );
  XOR U56570 ( .A(n44966), .B(n43647), .Z(n46883) );
  NOR U56571 ( .A(n43649), .B(n43648), .Z(n50301) );
  NOR U56572 ( .A(n43651), .B(n43650), .Z(n43656) );
  IV U56573 ( .A(n43652), .Z(n43654) );
  NOR U56574 ( .A(n43654), .B(n43653), .Z(n43655) );
  IV U56575 ( .A(n43655), .Z(n48411) );
  NOR U56576 ( .A(n43656), .B(n48411), .Z(n43657) );
  NOR U56577 ( .A(n50301), .B(n43657), .Z(n46884) );
  XOR U56578 ( .A(n46883), .B(n46884), .Z(n44961) );
  IV U56579 ( .A(n43658), .Z(n43663) );
  NOR U56580 ( .A(n43660), .B(n43659), .Z(n43661) );
  IV U56581 ( .A(n43661), .Z(n43662) );
  NOR U56582 ( .A(n43663), .B(n43662), .Z(n44959) );
  XOR U56583 ( .A(n44961), .B(n44959), .Z(n46881) );
  XOR U56584 ( .A(n46880), .B(n46881), .Z(n44957) );
  XOR U56585 ( .A(n44958), .B(n44957), .Z(n43664) );
  NOR U56586 ( .A(n43665), .B(n43664), .Z(n43673) );
  IV U56587 ( .A(n43666), .Z(n54207) );
  NOR U56588 ( .A(n43667), .B(n46881), .Z(n43668) );
  IV U56589 ( .A(n43668), .Z(n43670) );
  NOR U56590 ( .A(n54207), .B(n43670), .Z(n46899) );
  IV U56591 ( .A(n43669), .Z(n43671) );
  NOR U56592 ( .A(n43671), .B(n43670), .Z(n54196) );
  NOR U56593 ( .A(n46899), .B(n54196), .Z(n48400) );
  IV U56594 ( .A(n48400), .Z(n43672) );
  NOR U56595 ( .A(n43673), .B(n43672), .Z(n44954) );
  XOR U56596 ( .A(n43674), .B(n44954), .Z(n46907) );
  IV U56597 ( .A(n43675), .Z(n43679) );
  NOR U56598 ( .A(n43677), .B(n43676), .Z(n43678) );
  IV U56599 ( .A(n43678), .Z(n43685) );
  NOR U56600 ( .A(n43679), .B(n43685), .Z(n43680) );
  IV U56601 ( .A(n43680), .Z(n46906) );
  XOR U56602 ( .A(n46907), .B(n46906), .Z(n46901) );
  IV U56603 ( .A(n43681), .Z(n43683) );
  NOR U56604 ( .A(n43683), .B(n43682), .Z(n46913) );
  IV U56605 ( .A(n43684), .Z(n43686) );
  NOR U56606 ( .A(n43686), .B(n43685), .Z(n46902) );
  NOR U56607 ( .A(n46913), .B(n46902), .Z(n43687) );
  XOR U56608 ( .A(n46901), .B(n43687), .Z(n46920) );
  XOR U56609 ( .A(n46916), .B(n46920), .Z(n44952) );
  XOR U56610 ( .A(n43688), .B(n44952), .Z(n44949) );
  XOR U56611 ( .A(n44947), .B(n44949), .Z(n46930) );
  IV U56612 ( .A(n43689), .Z(n43691) );
  NOR U56613 ( .A(n43691), .B(n43690), .Z(n43692) );
  IV U56614 ( .A(n43692), .Z(n46929) );
  XOR U56615 ( .A(n46930), .B(n46929), .Z(n46924) );
  NOR U56616 ( .A(n46925), .B(n43693), .Z(n48383) );
  IV U56617 ( .A(n43694), .Z(n43696) );
  IV U56618 ( .A(n43695), .Z(n43699) );
  NOR U56619 ( .A(n43696), .B(n43699), .Z(n46939) );
  NOR U56620 ( .A(n48383), .B(n46939), .Z(n43697) );
  XOR U56621 ( .A(n46924), .B(n43697), .Z(n46950) );
  IV U56622 ( .A(n43698), .Z(n43700) );
  NOR U56623 ( .A(n43700), .B(n43699), .Z(n46948) );
  XOR U56624 ( .A(n46950), .B(n46948), .Z(n43701) );
  NOR U56625 ( .A(n43702), .B(n43701), .Z(n48373) );
  IV U56626 ( .A(n43703), .Z(n43704) );
  NOR U56627 ( .A(n43705), .B(n43704), .Z(n46946) );
  NOR U56628 ( .A(n46946), .B(n46948), .Z(n43706) );
  XOR U56629 ( .A(n46950), .B(n43706), .Z(n46955) );
  NOR U56630 ( .A(n43707), .B(n46955), .Z(n43708) );
  NOR U56631 ( .A(n48373), .B(n43708), .Z(n46958) );
  IV U56632 ( .A(n43709), .Z(n43710) );
  NOR U56633 ( .A(n43710), .B(n43716), .Z(n46954) );
  IV U56634 ( .A(n43711), .Z(n43712) );
  NOR U56635 ( .A(n43713), .B(n43712), .Z(n46959) );
  NOR U56636 ( .A(n46954), .B(n46959), .Z(n43714) );
  XOR U56637 ( .A(n46958), .B(n43714), .Z(n46964) );
  IV U56638 ( .A(n43715), .Z(n43717) );
  NOR U56639 ( .A(n43717), .B(n43716), .Z(n46962) );
  XOR U56640 ( .A(n46964), .B(n46962), .Z(n46966) );
  XOR U56641 ( .A(n46965), .B(n46966), .Z(n46970) );
  XOR U56642 ( .A(n46969), .B(n46970), .Z(n46973) );
  XOR U56643 ( .A(n46972), .B(n46973), .Z(n46978) );
  XOR U56644 ( .A(n46976), .B(n46978), .Z(n46980) );
  XOR U56645 ( .A(n46979), .B(n46980), .Z(n44943) );
  XOR U56646 ( .A(n44941), .B(n44943), .Z(n44945) );
  XOR U56647 ( .A(n43718), .B(n44945), .Z(n46985) );
  XOR U56648 ( .A(n46984), .B(n46985), .Z(n46988) );
  IV U56649 ( .A(n43719), .Z(n43720) );
  NOR U56650 ( .A(n43721), .B(n43720), .Z(n46987) );
  IV U56651 ( .A(n43722), .Z(n43724) );
  IV U56652 ( .A(n43723), .Z(n43727) );
  NOR U56653 ( .A(n43724), .B(n43727), .Z(n44936) );
  NOR U56654 ( .A(n46987), .B(n44936), .Z(n43725) );
  XOR U56655 ( .A(n46988), .B(n43725), .Z(n44929) );
  IV U56656 ( .A(n43726), .Z(n43728) );
  NOR U56657 ( .A(n43728), .B(n43727), .Z(n48336) );
  IV U56658 ( .A(n43729), .Z(n43730) );
  NOR U56659 ( .A(n43735), .B(n43730), .Z(n48332) );
  NOR U56660 ( .A(n48336), .B(n48332), .Z(n44930) );
  XOR U56661 ( .A(n44929), .B(n44930), .Z(n44932) );
  IV U56662 ( .A(n43731), .Z(n44926) );
  NOR U56663 ( .A(n43732), .B(n44926), .Z(n43736) );
  IV U56664 ( .A(n43733), .Z(n43734) );
  NOR U56665 ( .A(n43735), .B(n43734), .Z(n44931) );
  NOR U56666 ( .A(n43736), .B(n44931), .Z(n43737) );
  XOR U56667 ( .A(n44932), .B(n43737), .Z(n43747) );
  IV U56668 ( .A(n43747), .Z(n43741) );
  NOR U56669 ( .A(n43739), .B(n43738), .Z(n43751) );
  IV U56670 ( .A(n43751), .Z(n43740) );
  NOR U56671 ( .A(n43741), .B(n43740), .Z(n50374) );
  IV U56672 ( .A(n43742), .Z(n43744) );
  NOR U56673 ( .A(n43744), .B(n43743), .Z(n43748) );
  IV U56674 ( .A(n43748), .Z(n43746) );
  XOR U56675 ( .A(n44931), .B(n44932), .Z(n43745) );
  NOR U56676 ( .A(n43746), .B(n43745), .Z(n50358) );
  NOR U56677 ( .A(n43748), .B(n43747), .Z(n43749) );
  NOR U56678 ( .A(n50358), .B(n43749), .Z(n43750) );
  NOR U56679 ( .A(n43751), .B(n43750), .Z(n43752) );
  NOR U56680 ( .A(n50374), .B(n43752), .Z(n43753) );
  IV U56681 ( .A(n43753), .Z(n46997) );
  XOR U56682 ( .A(n46996), .B(n46997), .Z(n47002) );
  XOR U56683 ( .A(n47000), .B(n47002), .Z(n47004) );
  XOR U56684 ( .A(n43754), .B(n47004), .Z(n44923) );
  IV U56685 ( .A(n43755), .Z(n43757) );
  NOR U56686 ( .A(n43757), .B(n43756), .Z(n47008) );
  IV U56687 ( .A(n43758), .Z(n43760) );
  IV U56688 ( .A(n43759), .Z(n43763) );
  NOR U56689 ( .A(n43760), .B(n43763), .Z(n44922) );
  NOR U56690 ( .A(n47008), .B(n44922), .Z(n43761) );
  XOR U56691 ( .A(n44923), .B(n43761), .Z(n44916) );
  IV U56692 ( .A(n43762), .Z(n43764) );
  NOR U56693 ( .A(n43764), .B(n43763), .Z(n44914) );
  XOR U56694 ( .A(n44916), .B(n44914), .Z(n44919) );
  XOR U56695 ( .A(n44917), .B(n44919), .Z(n47014) );
  XOR U56696 ( .A(n47013), .B(n47014), .Z(n47018) );
  XOR U56697 ( .A(n47016), .B(n47018), .Z(n44910) );
  XOR U56698 ( .A(n44908), .B(n44910), .Z(n44912) );
  XOR U56699 ( .A(n43765), .B(n44912), .Z(n44901) );
  XOR U56700 ( .A(n44899), .B(n44901), .Z(n44903) );
  XOR U56701 ( .A(n44902), .B(n44903), .Z(n44896) );
  XOR U56702 ( .A(n44895), .B(n44896), .Z(n47023) );
  XOR U56703 ( .A(n47022), .B(n47023), .Z(n47026) );
  XOR U56704 ( .A(n47025), .B(n47026), .Z(n44893) );
  XOR U56705 ( .A(n44894), .B(n44893), .Z(n43766) );
  IV U56706 ( .A(n43766), .Z(n44892) );
  XOR U56707 ( .A(n44890), .B(n44892), .Z(n44886) );
  XOR U56708 ( .A(n44884), .B(n44886), .Z(n47031) );
  XOR U56709 ( .A(n43767), .B(n47031), .Z(n47033) );
  XOR U56710 ( .A(n47034), .B(n47033), .Z(n44879) );
  IV U56711 ( .A(n43768), .Z(n43770) );
  NOR U56712 ( .A(n43770), .B(n43769), .Z(n44878) );
  XOR U56713 ( .A(n44879), .B(n44878), .Z(n47037) );
  IV U56714 ( .A(n43771), .Z(n43773) );
  NOR U56715 ( .A(n43773), .B(n43772), .Z(n47036) );
  NOR U56716 ( .A(n44880), .B(n47036), .Z(n43774) );
  XOR U56717 ( .A(n47037), .B(n43774), .Z(n47042) );
  XOR U56718 ( .A(n47040), .B(n47042), .Z(n47044) );
  XOR U56719 ( .A(n47043), .B(n47044), .Z(n47048) );
  XOR U56720 ( .A(n47047), .B(n47048), .Z(n48288) );
  XOR U56721 ( .A(n47050), .B(n48288), .Z(n47054) );
  NOR U56722 ( .A(n47056), .B(n47053), .Z(n43775) );
  XOR U56723 ( .A(n47054), .B(n43775), .Z(n48283) );
  IV U56724 ( .A(n43776), .Z(n43777) );
  NOR U56725 ( .A(n43778), .B(n43777), .Z(n48282) );
  IV U56726 ( .A(n43779), .Z(n43780) );
  NOR U56727 ( .A(n43780), .B(n43782), .Z(n50465) );
  NOR U56728 ( .A(n48282), .B(n50465), .Z(n47059) );
  XOR U56729 ( .A(n48283), .B(n47059), .Z(n47061) );
  IV U56730 ( .A(n43781), .Z(n43783) );
  NOR U56731 ( .A(n43783), .B(n43782), .Z(n47060) );
  IV U56732 ( .A(n43784), .Z(n43786) );
  NOR U56733 ( .A(n43786), .B(n43785), .Z(n47071) );
  NOR U56734 ( .A(n47060), .B(n47071), .Z(n43787) );
  XOR U56735 ( .A(n47061), .B(n43787), .Z(n47070) );
  IV U56736 ( .A(n43788), .Z(n43790) );
  NOR U56737 ( .A(n43790), .B(n43789), .Z(n47068) );
  XOR U56738 ( .A(n47070), .B(n47068), .Z(n47067) );
  XOR U56739 ( .A(n43791), .B(n47067), .Z(n47076) );
  XOR U56740 ( .A(n43792), .B(n47076), .Z(n47085) );
  XOR U56741 ( .A(n47084), .B(n47085), .Z(n47096) );
  XOR U56742 ( .A(n43793), .B(n47096), .Z(n47098) );
  XOR U56743 ( .A(n47099), .B(n47098), .Z(n47104) );
  XOR U56744 ( .A(n47102), .B(n47104), .Z(n47107) );
  XOR U56745 ( .A(n47105), .B(n47107), .Z(n47113) );
  XOR U56746 ( .A(n43794), .B(n47113), .Z(n47110) );
  XOR U56747 ( .A(n47108), .B(n47110), .Z(n44867) );
  NOR U56748 ( .A(n43795), .B(n44862), .Z(n43799) );
  IV U56749 ( .A(n43796), .Z(n43798) );
  NOR U56750 ( .A(n43798), .B(n43797), .Z(n44865) );
  NOR U56751 ( .A(n43799), .B(n44865), .Z(n43800) );
  XOR U56752 ( .A(n44867), .B(n43800), .Z(n44855) );
  IV U56753 ( .A(n43801), .Z(n43805) );
  IV U56754 ( .A(n43802), .Z(n43807) );
  NOR U56755 ( .A(n43803), .B(n43807), .Z(n43804) );
  IV U56756 ( .A(n43804), .Z(n43811) );
  NOR U56757 ( .A(n43805), .B(n43811), .Z(n44856) );
  IV U56758 ( .A(n43806), .Z(n43808) );
  NOR U56759 ( .A(n43808), .B(n43807), .Z(n44858) );
  NOR U56760 ( .A(n44856), .B(n44858), .Z(n43809) );
  XOR U56761 ( .A(n44855), .B(n43809), .Z(n44854) );
  IV U56762 ( .A(n43810), .Z(n43812) );
  NOR U56763 ( .A(n43812), .B(n43811), .Z(n44852) );
  XOR U56764 ( .A(n44854), .B(n44852), .Z(n44848) );
  XOR U56765 ( .A(n44847), .B(n44848), .Z(n44850) );
  XOR U56766 ( .A(n44851), .B(n44850), .Z(n47118) );
  IV U56767 ( .A(n43813), .Z(n47125) );
  NOR U56768 ( .A(n47125), .B(n47127), .Z(n43817) );
  IV U56769 ( .A(n43814), .Z(n43815) );
  NOR U56770 ( .A(n43816), .B(n43815), .Z(n47119) );
  NOR U56771 ( .A(n43817), .B(n47119), .Z(n43818) );
  XOR U56772 ( .A(n47118), .B(n43818), .Z(n47123) );
  IV U56773 ( .A(n43819), .Z(n43821) );
  NOR U56774 ( .A(n43821), .B(n43820), .Z(n47121) );
  XOR U56775 ( .A(n47123), .B(n47121), .Z(n44843) );
  XOR U56776 ( .A(n44841), .B(n44843), .Z(n44845) );
  XOR U56777 ( .A(n44844), .B(n44845), .Z(n44840) );
  XOR U56778 ( .A(n44838), .B(n44840), .Z(n47132) );
  XOR U56779 ( .A(n47130), .B(n47132), .Z(n47134) );
  XOR U56780 ( .A(n47133), .B(n47134), .Z(n47138) );
  XOR U56781 ( .A(n47137), .B(n47138), .Z(n48235) );
  XOR U56782 ( .A(n47140), .B(n48235), .Z(n43822) );
  IV U56783 ( .A(n43822), .Z(n44834) );
  IV U56784 ( .A(n43823), .Z(n43825) );
  NOR U56785 ( .A(n43825), .B(n43824), .Z(n44832) );
  XOR U56786 ( .A(n44834), .B(n44832), .Z(n44837) );
  IV U56787 ( .A(n43826), .Z(n43829) );
  IV U56788 ( .A(n43827), .Z(n43828) );
  NOR U56789 ( .A(n43829), .B(n43828), .Z(n44835) );
  XOR U56790 ( .A(n44837), .B(n44835), .Z(n44827) );
  XOR U56791 ( .A(n44826), .B(n44827), .Z(n44831) );
  IV U56792 ( .A(n43830), .Z(n43831) );
  NOR U56793 ( .A(n43832), .B(n43831), .Z(n44829) );
  XOR U56794 ( .A(n44831), .B(n44829), .Z(n47146) );
  IV U56795 ( .A(n43833), .Z(n43837) );
  NOR U56796 ( .A(n43834), .B(n43837), .Z(n44824) );
  IV U56797 ( .A(n43835), .Z(n43839) );
  XOR U56798 ( .A(n43837), .B(n43836), .Z(n43838) );
  NOR U56799 ( .A(n43839), .B(n43838), .Z(n47145) );
  NOR U56800 ( .A(n44824), .B(n47145), .Z(n43840) );
  XOR U56801 ( .A(n47146), .B(n43840), .Z(n47149) );
  XOR U56802 ( .A(n43841), .B(n47149), .Z(n47159) );
  IV U56803 ( .A(n43842), .Z(n43843) );
  NOR U56804 ( .A(n43844), .B(n43843), .Z(n47155) );
  XOR U56805 ( .A(n47159), .B(n47155), .Z(n47162) );
  IV U56806 ( .A(n43845), .Z(n43846) );
  NOR U56807 ( .A(n43847), .B(n43846), .Z(n47158) );
  IV U56808 ( .A(n43848), .Z(n43849) );
  NOR U56809 ( .A(n43849), .B(n43852), .Z(n47161) );
  NOR U56810 ( .A(n47158), .B(n47161), .Z(n43850) );
  XOR U56811 ( .A(n47162), .B(n43850), .Z(n47164) );
  IV U56812 ( .A(n43851), .Z(n43853) );
  NOR U56813 ( .A(n43853), .B(n43852), .Z(n47165) );
  IV U56814 ( .A(n43854), .Z(n43856) );
  NOR U56815 ( .A(n43856), .B(n43855), .Z(n47171) );
  NOR U56816 ( .A(n47165), .B(n47171), .Z(n43857) );
  XOR U56817 ( .A(n47164), .B(n43857), .Z(n47169) );
  IV U56818 ( .A(n43858), .Z(n43859) );
  NOR U56819 ( .A(n43860), .B(n43859), .Z(n47168) );
  IV U56820 ( .A(n43861), .Z(n43862) );
  NOR U56821 ( .A(n43863), .B(n43862), .Z(n44822) );
  NOR U56822 ( .A(n47168), .B(n44822), .Z(n43864) );
  XOR U56823 ( .A(n47169), .B(n43864), .Z(n44816) );
  IV U56824 ( .A(n43865), .Z(n43866) );
  NOR U56825 ( .A(n43867), .B(n43866), .Z(n44819) );
  IV U56826 ( .A(n43868), .Z(n43869) );
  NOR U56827 ( .A(n43869), .B(n43872), .Z(n44817) );
  NOR U56828 ( .A(n44819), .B(n44817), .Z(n43870) );
  XOR U56829 ( .A(n44816), .B(n43870), .Z(n44811) );
  IV U56830 ( .A(n43871), .Z(n43873) );
  NOR U56831 ( .A(n43873), .B(n43872), .Z(n44809) );
  XOR U56832 ( .A(n44811), .B(n44809), .Z(n44814) );
  IV U56833 ( .A(n43874), .Z(n43879) );
  IV U56834 ( .A(n43875), .Z(n43876) );
  NOR U56835 ( .A(n43879), .B(n43876), .Z(n44812) );
  XOR U56836 ( .A(n44814), .B(n44812), .Z(n44802) );
  IV U56837 ( .A(n43877), .Z(n43878) );
  NOR U56838 ( .A(n43879), .B(n43878), .Z(n43880) );
  IV U56839 ( .A(n43880), .Z(n44801) );
  XOR U56840 ( .A(n44802), .B(n44801), .Z(n44804) );
  NOR U56841 ( .A(n43882), .B(n43881), .Z(n44803) );
  IV U56842 ( .A(n43883), .Z(n43885) );
  NOR U56843 ( .A(n43885), .B(n43884), .Z(n44806) );
  NOR U56844 ( .A(n44803), .B(n44806), .Z(n43886) );
  XOR U56845 ( .A(n44804), .B(n43886), .Z(n44796) );
  XOR U56846 ( .A(n44794), .B(n44796), .Z(n44799) );
  XOR U56847 ( .A(n44797), .B(n44799), .Z(n47183) );
  XOR U56848 ( .A(n43887), .B(n47183), .Z(n43888) );
  IV U56849 ( .A(n43888), .Z(n47181) );
  IV U56850 ( .A(n43889), .Z(n43891) );
  NOR U56851 ( .A(n43891), .B(n43890), .Z(n47179) );
  XOR U56852 ( .A(n47181), .B(n47179), .Z(n47191) );
  XOR U56853 ( .A(n47190), .B(n47191), .Z(n47195) );
  IV U56854 ( .A(n43892), .Z(n43894) );
  NOR U56855 ( .A(n43894), .B(n43893), .Z(n47193) );
  XOR U56856 ( .A(n47195), .B(n47193), .Z(n44789) );
  XOR U56857 ( .A(n44788), .B(n44789), .Z(n44786) );
  XOR U56858 ( .A(n44785), .B(n44786), .Z(n44781) );
  IV U56859 ( .A(n43895), .Z(n43897) );
  IV U56860 ( .A(n43896), .Z(n43903) );
  NOR U56861 ( .A(n43897), .B(n43903), .Z(n43898) );
  IV U56862 ( .A(n43898), .Z(n44780) );
  XOR U56863 ( .A(n44781), .B(n44780), .Z(n44775) );
  IV U56864 ( .A(n43899), .Z(n43900) );
  NOR U56865 ( .A(n43901), .B(n43900), .Z(n44774) );
  IV U56866 ( .A(n43902), .Z(n43904) );
  NOR U56867 ( .A(n43904), .B(n43903), .Z(n44782) );
  NOR U56868 ( .A(n44774), .B(n44782), .Z(n43905) );
  XOR U56869 ( .A(n44775), .B(n43905), .Z(n44779) );
  XOR U56870 ( .A(n44777), .B(n44779), .Z(n44772) );
  XOR U56871 ( .A(n44771), .B(n44772), .Z(n48185) );
  XOR U56872 ( .A(n43906), .B(n48185), .Z(n44768) );
  XOR U56873 ( .A(n44767), .B(n44768), .Z(n44762) );
  XOR U56874 ( .A(n44761), .B(n44762), .Z(n44764) );
  XOR U56875 ( .A(n44765), .B(n44764), .Z(n44759) );
  IV U56876 ( .A(n43907), .Z(n43908) );
  NOR U56877 ( .A(n43911), .B(n43908), .Z(n48175) );
  IV U56878 ( .A(n43909), .Z(n43914) );
  NOR U56879 ( .A(n43911), .B(n43910), .Z(n43912) );
  IV U56880 ( .A(n43912), .Z(n43913) );
  NOR U56881 ( .A(n43914), .B(n43913), .Z(n50640) );
  NOR U56882 ( .A(n48175), .B(n50640), .Z(n44760) );
  XOR U56883 ( .A(n44759), .B(n44760), .Z(n47205) );
  XOR U56884 ( .A(n47204), .B(n47205), .Z(n47214) );
  XOR U56885 ( .A(n43915), .B(n47214), .Z(n47215) );
  XOR U56886 ( .A(n43916), .B(n47215), .Z(n47220) );
  XOR U56887 ( .A(n43917), .B(n47220), .Z(n43918) );
  NOR U56888 ( .A(n43919), .B(n43918), .Z(n43922) );
  IV U56889 ( .A(n43919), .Z(n43921) );
  XOR U56890 ( .A(n47219), .B(n47220), .Z(n43920) );
  NOR U56891 ( .A(n43921), .B(n43920), .Z(n50658) );
  NOR U56892 ( .A(n43922), .B(n50658), .Z(n44753) );
  XOR U56893 ( .A(n43923), .B(n44753), .Z(n44752) );
  XOR U56894 ( .A(n43924), .B(n44752), .Z(n43925) );
  IV U56895 ( .A(n43925), .Z(n47241) );
  XOR U56896 ( .A(n44746), .B(n47241), .Z(n47239) );
  XOR U56897 ( .A(n43926), .B(n47239), .Z(n44744) );
  XOR U56898 ( .A(n44742), .B(n44744), .Z(n47258) );
  XOR U56899 ( .A(n47259), .B(n47258), .Z(n44740) );
  IV U56900 ( .A(n43927), .Z(n43928) );
  NOR U56901 ( .A(n43929), .B(n43928), .Z(n47260) );
  IV U56902 ( .A(n43930), .Z(n43931) );
  NOR U56903 ( .A(n43932), .B(n43931), .Z(n44739) );
  NOR U56904 ( .A(n47260), .B(n44739), .Z(n43933) );
  XOR U56905 ( .A(n44740), .B(n43933), .Z(n47266) );
  IV U56906 ( .A(n43934), .Z(n43936) );
  NOR U56907 ( .A(n43936), .B(n43935), .Z(n47264) );
  XOR U56908 ( .A(n47266), .B(n47264), .Z(n47268) );
  XOR U56909 ( .A(n47267), .B(n47268), .Z(n44733) );
  XOR U56910 ( .A(n43937), .B(n44733), .Z(n47276) );
  XOR U56911 ( .A(n47274), .B(n47276), .Z(n50685) );
  XOR U56912 ( .A(n44727), .B(n50685), .Z(n44728) );
  IV U56913 ( .A(n43938), .Z(n43939) );
  NOR U56914 ( .A(n43940), .B(n43939), .Z(n48122) );
  IV U56915 ( .A(n43941), .Z(n43943) );
  NOR U56916 ( .A(n43943), .B(n43942), .Z(n48128) );
  NOR U56917 ( .A(n48122), .B(n48128), .Z(n44729) );
  XOR U56918 ( .A(n44728), .B(n44729), .Z(n44726) );
  XOR U56919 ( .A(n44724), .B(n44726), .Z(n47283) );
  XOR U56920 ( .A(n47282), .B(n47283), .Z(n47286) );
  XOR U56921 ( .A(n47285), .B(n47286), .Z(n47290) );
  XOR U56922 ( .A(n47289), .B(n47290), .Z(n47296) );
  XOR U56923 ( .A(n43944), .B(n47296), .Z(n44719) );
  IV U56924 ( .A(n43945), .Z(n43946) );
  NOR U56925 ( .A(n43946), .B(n43950), .Z(n44720) );
  IV U56926 ( .A(n43947), .Z(n43948) );
  NOR U56927 ( .A(n43949), .B(n43948), .Z(n47303) );
  NOR U56928 ( .A(n43951), .B(n43950), .Z(n44722) );
  NOR U56929 ( .A(n47303), .B(n44722), .Z(n43952) );
  IV U56930 ( .A(n43952), .Z(n43953) );
  NOR U56931 ( .A(n44720), .B(n43953), .Z(n43954) );
  XOR U56932 ( .A(n44719), .B(n43954), .Z(n47310) );
  IV U56933 ( .A(n43955), .Z(n43957) );
  NOR U56934 ( .A(n43957), .B(n43956), .Z(n47308) );
  XOR U56935 ( .A(n47310), .B(n47308), .Z(n44717) );
  XOR U56936 ( .A(n44716), .B(n44717), .Z(n44715) );
  XOR U56937 ( .A(n44713), .B(n44715), .Z(n47322) );
  XOR U56938 ( .A(n47320), .B(n47322), .Z(n47325) );
  XOR U56939 ( .A(n47323), .B(n47325), .Z(n44709) );
  XOR U56940 ( .A(n44707), .B(n44709), .Z(n44712) );
  XOR U56941 ( .A(n44710), .B(n44712), .Z(n44702) );
  XOR U56942 ( .A(n44701), .B(n44702), .Z(n44706) );
  XOR U56943 ( .A(n44704), .B(n44706), .Z(n44699) );
  NOR U56944 ( .A(n43964), .B(n44699), .Z(n50734) );
  IV U56945 ( .A(n43958), .Z(n43960) );
  NOR U56946 ( .A(n43960), .B(n43959), .Z(n44698) );
  XOR U56947 ( .A(n44698), .B(n44699), .Z(n44694) );
  IV U56948 ( .A(n43961), .Z(n43962) );
  NOR U56949 ( .A(n43963), .B(n43962), .Z(n43965) );
  IV U56950 ( .A(n43965), .Z(n44693) );
  XOR U56951 ( .A(n44694), .B(n44693), .Z(n43967) );
  NOR U56952 ( .A(n43965), .B(n43964), .Z(n43966) );
  NOR U56953 ( .A(n43967), .B(n43966), .Z(n43968) );
  NOR U56954 ( .A(n50734), .B(n43968), .Z(n44695) );
  XOR U56955 ( .A(n44697), .B(n44695), .Z(n48093) );
  IV U56956 ( .A(n43969), .Z(n43976) );
  IV U56957 ( .A(n43970), .Z(n43971) );
  NOR U56958 ( .A(n43976), .B(n43971), .Z(n44691) );
  XOR U56959 ( .A(n48093), .B(n44691), .Z(n44686) );
  IV U56960 ( .A(n43972), .Z(n43973) );
  NOR U56961 ( .A(n43976), .B(n43973), .Z(n44685) );
  XOR U56962 ( .A(n44686), .B(n44685), .Z(n44689) );
  IV U56963 ( .A(n43974), .Z(n43975) );
  NOR U56964 ( .A(n43976), .B(n43975), .Z(n44687) );
  XOR U56965 ( .A(n44689), .B(n44687), .Z(n50747) );
  IV U56966 ( .A(n43977), .Z(n43978) );
  NOR U56967 ( .A(n43979), .B(n43978), .Z(n50746) );
  IV U56968 ( .A(n43980), .Z(n43982) );
  NOR U56969 ( .A(n43982), .B(n43981), .Z(n50751) );
  NOR U56970 ( .A(n50746), .B(n50751), .Z(n47331) );
  XOR U56971 ( .A(n50747), .B(n47331), .Z(n47333) );
  XOR U56972 ( .A(n43983), .B(n47333), .Z(n48075) );
  XOR U56973 ( .A(n47341), .B(n48075), .Z(n43984) );
  IV U56974 ( .A(n43984), .Z(n47343) );
  XOR U56975 ( .A(n47342), .B(n47343), .Z(n43985) );
  NOR U56976 ( .A(n43986), .B(n43985), .Z(n51732) );
  IV U56977 ( .A(n43987), .Z(n43988) );
  NOR U56978 ( .A(n43989), .B(n43988), .Z(n44683) );
  NOR U56979 ( .A(n44683), .B(n47342), .Z(n43990) );
  XOR U56980 ( .A(n47343), .B(n43990), .Z(n43991) );
  NOR U56981 ( .A(n43992), .B(n43991), .Z(n43993) );
  NOR U56982 ( .A(n51732), .B(n43993), .Z(n44680) );
  IV U56983 ( .A(n43994), .Z(n43996) );
  NOR U56984 ( .A(n43996), .B(n43995), .Z(n43997) );
  IV U56985 ( .A(n43997), .Z(n44681) );
  XOR U56986 ( .A(n44680), .B(n44681), .Z(n47348) );
  XOR U56987 ( .A(n47347), .B(n47348), .Z(n47351) );
  XOR U56988 ( .A(n47350), .B(n47351), .Z(n44674) );
  XOR U56989 ( .A(n43998), .B(n44674), .Z(n44672) );
  XOR U56990 ( .A(n44670), .B(n44672), .Z(n47361) );
  IV U56991 ( .A(n43999), .Z(n44003) );
  NOR U56992 ( .A(n44001), .B(n44000), .Z(n44002) );
  IV U56993 ( .A(n44002), .Z(n44005) );
  NOR U56994 ( .A(n44003), .B(n44005), .Z(n47359) );
  XOR U56995 ( .A(n47361), .B(n47359), .Z(n44669) );
  IV U56996 ( .A(n44004), .Z(n44006) );
  NOR U56997 ( .A(n44006), .B(n44005), .Z(n44667) );
  XOR U56998 ( .A(n44669), .B(n44667), .Z(n47366) );
  XOR U56999 ( .A(n47365), .B(n47366), .Z(n47370) );
  IV U57000 ( .A(n44007), .Z(n44011) );
  NOR U57001 ( .A(n44013), .B(n44008), .Z(n44009) );
  IV U57002 ( .A(n44009), .Z(n44010) );
  NOR U57003 ( .A(n44011), .B(n44010), .Z(n47368) );
  XOR U57004 ( .A(n47370), .B(n47368), .Z(n50783) );
  NOR U57005 ( .A(n44013), .B(n44012), .Z(n44014) );
  IV U57006 ( .A(n44014), .Z(n44021) );
  XOR U57007 ( .A(n44016), .B(n44015), .Z(n44017) );
  NOR U57008 ( .A(n44018), .B(n44017), .Z(n44019) );
  IV U57009 ( .A(n44019), .Z(n44020) );
  NOR U57010 ( .A(n44021), .B(n44020), .Z(n44022) );
  IV U57011 ( .A(n44022), .Z(n50778) );
  NOR U57012 ( .A(n44023), .B(n50778), .Z(n47372) );
  XOR U57013 ( .A(n50783), .B(n47372), .Z(n48046) );
  IV U57014 ( .A(n44024), .Z(n44026) );
  NOR U57015 ( .A(n44026), .B(n44025), .Z(n48053) );
  IV U57016 ( .A(n44027), .Z(n44029) );
  NOR U57017 ( .A(n44029), .B(n44028), .Z(n48045) );
  NOR U57018 ( .A(n48053), .B(n48045), .Z(n47374) );
  XOR U57019 ( .A(n48046), .B(n47374), .Z(n47378) );
  XOR U57020 ( .A(n47379), .B(n47378), .Z(n47381) );
  XOR U57021 ( .A(n47380), .B(n47381), .Z(n44661) );
  XOR U57022 ( .A(n44660), .B(n44661), .Z(n44664) );
  IV U57023 ( .A(n44030), .Z(n44032) );
  NOR U57024 ( .A(n44032), .B(n44031), .Z(n44663) );
  IV U57025 ( .A(n44033), .Z(n44034) );
  NOR U57026 ( .A(n44035), .B(n44034), .Z(n44657) );
  NOR U57027 ( .A(n44663), .B(n44657), .Z(n44036) );
  XOR U57028 ( .A(n44664), .B(n44036), .Z(n44046) );
  IV U57029 ( .A(n44046), .Z(n44656) );
  IV U57030 ( .A(n44037), .Z(n44038) );
  NOR U57031 ( .A(n44039), .B(n44038), .Z(n44040) );
  IV U57032 ( .A(n44040), .Z(n44047) );
  NOR U57033 ( .A(n44656), .B(n44047), .Z(n54611) );
  NOR U57034 ( .A(n44042), .B(n44041), .Z(n44648) );
  IV U57035 ( .A(n44043), .Z(n44045) );
  NOR U57036 ( .A(n44045), .B(n44044), .Z(n44654) );
  XOR U57037 ( .A(n44654), .B(n44046), .Z(n44649) );
  XOR U57038 ( .A(n44648), .B(n44649), .Z(n44049) );
  NOR U57039 ( .A(n44649), .B(n44047), .Z(n44048) );
  NOR U57040 ( .A(n44049), .B(n44048), .Z(n44050) );
  NOR U57041 ( .A(n54611), .B(n44050), .Z(n44051) );
  IV U57042 ( .A(n44051), .Z(n50810) );
  NOR U57043 ( .A(n44052), .B(n50810), .Z(n50825) );
  IV U57044 ( .A(n44053), .Z(n44054) );
  NOR U57045 ( .A(n44054), .B(n51650), .Z(n50808) );
  NOR U57046 ( .A(n44055), .B(n50808), .Z(n44056) );
  XOR U57047 ( .A(n44056), .B(n50810), .Z(n51645) );
  NOR U57048 ( .A(n47388), .B(n51645), .Z(n44057) );
  NOR U57049 ( .A(n50825), .B(n44057), .Z(n47391) );
  XOR U57050 ( .A(n47393), .B(n47391), .Z(n47396) );
  IV U57051 ( .A(n44058), .Z(n44061) );
  IV U57052 ( .A(n44059), .Z(n44060) );
  NOR U57053 ( .A(n44061), .B(n44060), .Z(n47394) );
  XOR U57054 ( .A(n47396), .B(n47394), .Z(n44643) );
  IV U57055 ( .A(n44062), .Z(n44065) );
  IV U57056 ( .A(n44063), .Z(n44064) );
  NOR U57057 ( .A(n44065), .B(n44064), .Z(n44641) );
  XOR U57058 ( .A(n44643), .B(n44641), .Z(n44644) );
  XOR U57059 ( .A(n44645), .B(n44644), .Z(n50837) );
  XOR U57060 ( .A(n47398), .B(n50837), .Z(n50830) );
  XOR U57061 ( .A(n47399), .B(n50830), .Z(n44639) );
  XOR U57062 ( .A(n44640), .B(n44639), .Z(n47404) );
  XOR U57063 ( .A(n47405), .B(n47404), .Z(n47407) );
  IV U57064 ( .A(n44066), .Z(n44068) );
  NOR U57065 ( .A(n44068), .B(n44067), .Z(n47406) );
  IV U57066 ( .A(n44069), .Z(n44071) );
  NOR U57067 ( .A(n44071), .B(n44070), .Z(n47410) );
  NOR U57068 ( .A(n47406), .B(n47410), .Z(n44072) );
  XOR U57069 ( .A(n47407), .B(n44072), .Z(n47415) );
  XOR U57070 ( .A(n47413), .B(n47415), .Z(n44634) );
  XOR U57071 ( .A(n44633), .B(n44634), .Z(n44637) );
  XOR U57072 ( .A(n44636), .B(n44637), .Z(n47418) );
  XOR U57073 ( .A(n47417), .B(n47418), .Z(n47422) );
  XOR U57074 ( .A(n47420), .B(n47422), .Z(n48001) );
  XOR U57075 ( .A(n47427), .B(n48001), .Z(n44073) );
  IV U57076 ( .A(n44073), .Z(n44631) );
  IV U57077 ( .A(n44074), .Z(n44075) );
  NOR U57078 ( .A(n44076), .B(n44075), .Z(n44629) );
  XOR U57079 ( .A(n44631), .B(n44629), .Z(n47425) );
  XOR U57080 ( .A(n47424), .B(n47425), .Z(n44627) );
  XOR U57081 ( .A(n44626), .B(n44627), .Z(n47435) );
  XOR U57082 ( .A(n47434), .B(n47435), .Z(n47437) );
  XOR U57083 ( .A(n47438), .B(n47437), .Z(n44624) );
  IV U57084 ( .A(n44077), .Z(n44078) );
  NOR U57085 ( .A(n44079), .B(n44078), .Z(n47440) );
  IV U57086 ( .A(n44084), .Z(n44080) );
  NOR U57087 ( .A(n44080), .B(n44083), .Z(n44623) );
  NOR U57088 ( .A(n47440), .B(n44623), .Z(n44081) );
  XOR U57089 ( .A(n44624), .B(n44081), .Z(n44618) );
  IV U57090 ( .A(n44082), .Z(n44086) );
  XOR U57091 ( .A(n44084), .B(n44083), .Z(n44085) );
  NOR U57092 ( .A(n44086), .B(n44085), .Z(n44616) );
  XOR U57093 ( .A(n44618), .B(n44616), .Z(n44620) );
  XOR U57094 ( .A(n44087), .B(n44620), .Z(n47445) );
  XOR U57095 ( .A(n47444), .B(n47445), .Z(n47447) );
  IV U57096 ( .A(n44088), .Z(n44089) );
  NOR U57097 ( .A(n44090), .B(n44089), .Z(n47446) );
  IV U57098 ( .A(n44091), .Z(n44093) );
  IV U57099 ( .A(n44092), .Z(n44096) );
  NOR U57100 ( .A(n44093), .B(n44096), .Z(n47453) );
  NOR U57101 ( .A(n47446), .B(n47453), .Z(n44094) );
  XOR U57102 ( .A(n47447), .B(n44094), .Z(n47452) );
  IV U57103 ( .A(n44095), .Z(n44097) );
  NOR U57104 ( .A(n44097), .B(n44096), .Z(n47450) );
  XOR U57105 ( .A(n47452), .B(n47450), .Z(n47458) );
  XOR U57106 ( .A(n47457), .B(n47458), .Z(n47980) );
  XOR U57107 ( .A(n44098), .B(n47980), .Z(n47464) );
  XOR U57108 ( .A(n47463), .B(n47464), .Z(n47467) );
  XOR U57109 ( .A(n47466), .B(n47467), .Z(n47471) );
  XOR U57110 ( .A(n47470), .B(n47471), .Z(n47474) );
  IV U57111 ( .A(n44099), .Z(n44102) );
  IV U57112 ( .A(n44100), .Z(n44101) );
  NOR U57113 ( .A(n44102), .B(n44101), .Z(n44103) );
  IV U57114 ( .A(n44103), .Z(n47473) );
  XOR U57115 ( .A(n47474), .B(n47473), .Z(n44611) );
  IV U57116 ( .A(n44104), .Z(n44106) );
  IV U57117 ( .A(n44105), .Z(n44116) );
  NOR U57118 ( .A(n44106), .B(n44116), .Z(n47479) );
  IV U57119 ( .A(n44107), .Z(n44108) );
  NOR U57120 ( .A(n44111), .B(n44108), .Z(n47476) );
  IV U57121 ( .A(n44109), .Z(n44110) );
  NOR U57122 ( .A(n44111), .B(n44110), .Z(n44610) );
  NOR U57123 ( .A(n47476), .B(n44610), .Z(n44112) );
  IV U57124 ( .A(n44112), .Z(n44113) );
  NOR U57125 ( .A(n47479), .B(n44113), .Z(n44114) );
  XOR U57126 ( .A(n44611), .B(n44114), .Z(n44609) );
  IV U57127 ( .A(n44115), .Z(n44117) );
  NOR U57128 ( .A(n44117), .B(n44116), .Z(n44607) );
  XOR U57129 ( .A(n44609), .B(n44607), .Z(n47486) );
  XOR U57130 ( .A(n47485), .B(n47486), .Z(n47488) );
  NOR U57131 ( .A(n44125), .B(n47488), .Z(n50942) );
  IV U57132 ( .A(n44118), .Z(n44120) );
  NOR U57133 ( .A(n44120), .B(n44119), .Z(n44603) );
  IV U57134 ( .A(n44121), .Z(n44122) );
  NOR U57135 ( .A(n44123), .B(n44122), .Z(n44124) );
  IV U57136 ( .A(n44124), .Z(n47489) );
  XOR U57137 ( .A(n47489), .B(n47488), .Z(n44604) );
  XOR U57138 ( .A(n44603), .B(n44604), .Z(n44127) );
  NOR U57139 ( .A(n44604), .B(n44125), .Z(n44126) );
  NOR U57140 ( .A(n44127), .B(n44126), .Z(n44128) );
  NOR U57141 ( .A(n50942), .B(n44128), .Z(n44596) );
  IV U57142 ( .A(n44129), .Z(n44131) );
  NOR U57143 ( .A(n44131), .B(n44130), .Z(n44601) );
  XOR U57144 ( .A(n44596), .B(n44601), .Z(n44132) );
  XOR U57145 ( .A(n44133), .B(n44132), .Z(n44134) );
  IV U57146 ( .A(n44134), .Z(n47500) );
  IV U57147 ( .A(n44135), .Z(n47494) );
  IV U57148 ( .A(n44136), .Z(n44137) );
  NOR U57149 ( .A(n47494), .B(n44137), .Z(n47498) );
  XOR U57150 ( .A(n47500), .B(n47498), .Z(n47502) );
  XOR U57151 ( .A(n47501), .B(n47502), .Z(n47508) );
  IV U57152 ( .A(n44138), .Z(n44140) );
  NOR U57153 ( .A(n44140), .B(n44139), .Z(n47506) );
  XOR U57154 ( .A(n47508), .B(n47506), .Z(n44593) );
  XOR U57155 ( .A(n44592), .B(n44593), .Z(n47519) );
  IV U57156 ( .A(n44141), .Z(n44148) );
  IV U57157 ( .A(n44142), .Z(n44143) );
  NOR U57158 ( .A(n44148), .B(n44143), .Z(n44144) );
  IV U57159 ( .A(n44144), .Z(n47505) );
  XOR U57160 ( .A(n47519), .B(n47505), .Z(n47514) );
  NOR U57161 ( .A(n44145), .B(n47520), .Z(n44149) );
  IV U57162 ( .A(n44146), .Z(n44147) );
  NOR U57163 ( .A(n44148), .B(n44147), .Z(n47515) );
  NOR U57164 ( .A(n44149), .B(n47515), .Z(n44150) );
  XOR U57165 ( .A(n47514), .B(n44150), .Z(n47535) );
  XOR U57166 ( .A(n47524), .B(n47535), .Z(n44156) );
  IV U57167 ( .A(n44151), .Z(n44154) );
  NOR U57168 ( .A(n44152), .B(n44159), .Z(n44153) );
  IV U57169 ( .A(n44153), .Z(n44165) );
  NOR U57170 ( .A(n44154), .B(n44165), .Z(n44162) );
  IV U57171 ( .A(n44162), .Z(n44155) );
  NOR U57172 ( .A(n44156), .B(n44155), .Z(n47944) );
  IV U57173 ( .A(n44157), .Z(n44158) );
  NOR U57174 ( .A(n44159), .B(n44158), .Z(n47533) );
  NOR U57175 ( .A(n47524), .B(n47533), .Z(n44160) );
  XOR U57176 ( .A(n47535), .B(n44160), .Z(n44161) );
  NOR U57177 ( .A(n44162), .B(n44161), .Z(n44163) );
  NOR U57178 ( .A(n47944), .B(n44163), .Z(n47538) );
  IV U57179 ( .A(n44164), .Z(n44166) );
  NOR U57180 ( .A(n44166), .B(n44165), .Z(n44167) );
  IV U57181 ( .A(n44167), .Z(n47539) );
  XOR U57182 ( .A(n47538), .B(n47539), .Z(n47542) );
  XOR U57183 ( .A(n47541), .B(n47542), .Z(n47548) );
  XOR U57184 ( .A(n47547), .B(n47548), .Z(n50996) );
  XOR U57185 ( .A(n50997), .B(n50996), .Z(n44168) );
  IV U57186 ( .A(n44168), .Z(n47558) );
  IV U57187 ( .A(n44169), .Z(n44171) );
  NOR U57188 ( .A(n44171), .B(n44170), .Z(n47556) );
  XOR U57189 ( .A(n47558), .B(n47556), .Z(n47938) );
  XOR U57190 ( .A(n47559), .B(n47938), .Z(n44172) );
  IV U57191 ( .A(n44172), .Z(n47570) );
  XOR U57192 ( .A(n47569), .B(n47570), .Z(n47563) );
  XOR U57193 ( .A(n47562), .B(n47563), .Z(n47568) );
  XOR U57194 ( .A(n47566), .B(n47568), .Z(n44590) );
  XOR U57195 ( .A(n44173), .B(n44590), .Z(n44581) );
  IV U57196 ( .A(n44174), .Z(n44175) );
  NOR U57197 ( .A(n44176), .B(n44175), .Z(n44180) );
  NOR U57198 ( .A(n44178), .B(n44177), .Z(n44179) );
  NOR U57199 ( .A(n44180), .B(n44179), .Z(n44584) );
  IV U57200 ( .A(n44584), .Z(n44188) );
  IV U57201 ( .A(n44181), .Z(n44183) );
  IV U57202 ( .A(n44182), .Z(n44192) );
  NOR U57203 ( .A(n44183), .B(n44192), .Z(n47582) );
  IV U57204 ( .A(n44184), .Z(n44185) );
  NOR U57205 ( .A(n44192), .B(n44185), .Z(n44582) );
  NOR U57206 ( .A(n47582), .B(n44582), .Z(n44186) );
  IV U57207 ( .A(n44186), .Z(n44187) );
  NOR U57208 ( .A(n44188), .B(n44187), .Z(n44189) );
  XOR U57209 ( .A(n44581), .B(n44189), .Z(n47591) );
  IV U57210 ( .A(n44190), .Z(n44191) );
  NOR U57211 ( .A(n44192), .B(n44191), .Z(n47585) );
  IV U57212 ( .A(n44193), .Z(n44194) );
  NOR U57213 ( .A(n44197), .B(n44194), .Z(n47589) );
  IV U57214 ( .A(n44195), .Z(n44196) );
  NOR U57215 ( .A(n44197), .B(n44196), .Z(n44579) );
  NOR U57216 ( .A(n47589), .B(n44579), .Z(n44198) );
  IV U57217 ( .A(n44198), .Z(n44199) );
  NOR U57218 ( .A(n47585), .B(n44199), .Z(n44200) );
  XOR U57219 ( .A(n47591), .B(n44200), .Z(n44568) );
  IV U57220 ( .A(n44201), .Z(n44204) );
  IV U57221 ( .A(n44202), .Z(n44203) );
  NOR U57222 ( .A(n44204), .B(n44203), .Z(n44571) );
  NOR U57223 ( .A(n44576), .B(n44571), .Z(n44205) );
  XOR U57224 ( .A(n44568), .B(n44205), .Z(n44575) );
  XOR U57225 ( .A(n44573), .B(n44575), .Z(n47598) );
  XOR U57226 ( .A(n44206), .B(n47598), .Z(n47601) );
  IV U57227 ( .A(n44207), .Z(n44209) );
  NOR U57228 ( .A(n44209), .B(n44208), .Z(n47599) );
  NOR U57229 ( .A(n44211), .B(n44210), .Z(n44215) );
  IV U57230 ( .A(n44211), .Z(n47604) );
  NOR U57231 ( .A(n47602), .B(n47604), .Z(n44212) );
  NOR U57232 ( .A(n44213), .B(n44212), .Z(n44214) );
  NOR U57233 ( .A(n44215), .B(n44214), .Z(n44216) );
  XOR U57234 ( .A(n47599), .B(n44216), .Z(n44217) );
  XOR U57235 ( .A(n47601), .B(n44217), .Z(n47617) );
  XOR U57236 ( .A(n47616), .B(n47617), .Z(n44565) );
  IV U57237 ( .A(n44218), .Z(n44220) );
  NOR U57238 ( .A(n44220), .B(n44219), .Z(n44563) );
  XOR U57239 ( .A(n44565), .B(n44563), .Z(n47614) );
  XOR U57240 ( .A(n47613), .B(n47614), .Z(n47625) );
  XOR U57241 ( .A(n47624), .B(n47625), .Z(n47630) );
  IV U57242 ( .A(n47630), .Z(n44228) );
  IV U57243 ( .A(n44221), .Z(n44223) );
  NOR U57244 ( .A(n44223), .B(n44222), .Z(n47629) );
  IV U57245 ( .A(n44224), .Z(n44226) );
  NOR U57246 ( .A(n44226), .B(n44225), .Z(n47627) );
  NOR U57247 ( .A(n47629), .B(n47627), .Z(n44227) );
  XOR U57248 ( .A(n44228), .B(n44227), .Z(n44560) );
  XOR U57249 ( .A(n44558), .B(n44560), .Z(n44561) );
  NOR U57250 ( .A(n44236), .B(n44561), .Z(n51052) );
  IV U57251 ( .A(n44229), .Z(n44230) );
  NOR U57252 ( .A(n44231), .B(n44230), .Z(n44554) );
  IV U57253 ( .A(n44232), .Z(n44233) );
  NOR U57254 ( .A(n44234), .B(n44233), .Z(n44235) );
  IV U57255 ( .A(n44235), .Z(n44562) );
  XOR U57256 ( .A(n44562), .B(n44561), .Z(n44555) );
  XOR U57257 ( .A(n44554), .B(n44555), .Z(n44238) );
  NOR U57258 ( .A(n44555), .B(n44236), .Z(n44237) );
  NOR U57259 ( .A(n44238), .B(n44237), .Z(n44239) );
  NOR U57260 ( .A(n51052), .B(n44239), .Z(n44548) );
  XOR U57261 ( .A(n44549), .B(n44548), .Z(n44551) );
  IV U57262 ( .A(n44240), .Z(n44241) );
  NOR U57263 ( .A(n44242), .B(n44241), .Z(n44550) );
  IV U57264 ( .A(n44243), .Z(n44245) );
  NOR U57265 ( .A(n44245), .B(n44244), .Z(n44546) );
  NOR U57266 ( .A(n44550), .B(n44546), .Z(n44246) );
  XOR U57267 ( .A(n44551), .B(n44246), .Z(n44540) );
  XOR U57268 ( .A(n44247), .B(n44540), .Z(n47642) );
  XOR U57269 ( .A(n47641), .B(n47642), .Z(n44538) );
  XOR U57270 ( .A(n44536), .B(n44538), .Z(n47639) );
  XOR U57271 ( .A(n44248), .B(n47639), .Z(n44249) );
  IV U57272 ( .A(n44249), .Z(n44529) );
  IV U57273 ( .A(n44250), .Z(n44251) );
  NOR U57274 ( .A(n44251), .B(n44253), .Z(n44527) );
  XOR U57275 ( .A(n44529), .B(n44527), .Z(n44532) );
  IV U57276 ( .A(n44252), .Z(n44254) );
  NOR U57277 ( .A(n44254), .B(n44253), .Z(n44530) );
  XOR U57278 ( .A(n44532), .B(n44530), .Z(n44525) );
  IV U57279 ( .A(n44255), .Z(n44256) );
  NOR U57280 ( .A(n44257), .B(n44256), .Z(n44522) );
  NOR U57281 ( .A(n44522), .B(n44524), .Z(n44258) );
  XOR U57282 ( .A(n44525), .B(n44258), .Z(n47652) );
  XOR U57283 ( .A(n44259), .B(n47652), .Z(n47662) );
  XOR U57284 ( .A(n44260), .B(n47662), .Z(n44261) );
  IV U57285 ( .A(n44261), .Z(n47664) );
  IV U57286 ( .A(n44262), .Z(n44264) );
  NOR U57287 ( .A(n44264), .B(n44263), .Z(n47663) );
  IV U57288 ( .A(n44265), .Z(n44266) );
  NOR U57289 ( .A(n44267), .B(n44266), .Z(n44519) );
  NOR U57290 ( .A(n47663), .B(n44519), .Z(n44268) );
  XOR U57291 ( .A(n47664), .B(n44268), .Z(n44269) );
  NOR U57292 ( .A(n44270), .B(n44269), .Z(n44273) );
  IV U57293 ( .A(n44270), .Z(n44272) );
  XOR U57294 ( .A(n47663), .B(n47664), .Z(n44271) );
  NOR U57295 ( .A(n44272), .B(n44271), .Z(n51465) );
  NOR U57296 ( .A(n44273), .B(n51465), .Z(n44511) );
  XOR U57297 ( .A(n44274), .B(n44511), .Z(n44515) );
  XOR U57298 ( .A(n44514), .B(n44515), .Z(n44510) );
  IV U57299 ( .A(n44275), .Z(n44276) );
  NOR U57300 ( .A(n44277), .B(n44276), .Z(n44508) );
  XOR U57301 ( .A(n44510), .B(n44508), .Z(n47670) );
  XOR U57302 ( .A(n47671), .B(n47670), .Z(n44500) );
  NOR U57303 ( .A(n44278), .B(n44505), .Z(n44284) );
  IV U57304 ( .A(n44279), .Z(n44283) );
  NOR U57305 ( .A(n44281), .B(n44280), .Z(n44282) );
  IV U57306 ( .A(n44282), .Z(n44287) );
  NOR U57307 ( .A(n44283), .B(n44287), .Z(n44501) );
  NOR U57308 ( .A(n44284), .B(n44501), .Z(n44285) );
  XOR U57309 ( .A(n44500), .B(n44285), .Z(n47678) );
  IV U57310 ( .A(n44286), .Z(n44288) );
  NOR U57311 ( .A(n44288), .B(n44287), .Z(n47676) );
  XOR U57312 ( .A(n47678), .B(n47676), .Z(n47680) );
  XOR U57313 ( .A(n47679), .B(n47680), .Z(n44498) );
  XOR U57314 ( .A(n44497), .B(n44498), .Z(n44492) );
  XOR U57315 ( .A(n44491), .B(n44492), .Z(n44496) );
  XOR U57316 ( .A(n44494), .B(n44496), .Z(n44487) );
  XOR U57317 ( .A(n44485), .B(n44487), .Z(n44489) );
  XOR U57318 ( .A(n44289), .B(n44489), .Z(n44477) );
  IV U57319 ( .A(n44290), .Z(n44292) );
  NOR U57320 ( .A(n44292), .B(n44291), .Z(n44480) );
  NOR U57321 ( .A(n44294), .B(n44293), .Z(n44478) );
  NOR U57322 ( .A(n44480), .B(n44478), .Z(n44295) );
  XOR U57323 ( .A(n44477), .B(n44295), .Z(n47815) );
  XOR U57324 ( .A(n44296), .B(n47815), .Z(n44473) );
  IV U57325 ( .A(n44297), .Z(n44299) );
  NOR U57326 ( .A(n44299), .B(n44298), .Z(n44471) );
  XOR U57327 ( .A(n44473), .B(n44471), .Z(n47688) );
  IV U57328 ( .A(n44300), .Z(n44301) );
  NOR U57329 ( .A(n44302), .B(n44301), .Z(n44474) );
  NOR U57330 ( .A(n44474), .B(n47687), .Z(n44303) );
  XOR U57331 ( .A(n47688), .B(n44303), .Z(n44465) );
  IV U57332 ( .A(n44304), .Z(n44307) );
  IV U57333 ( .A(n44305), .Z(n44306) );
  NOR U57334 ( .A(n44307), .B(n44306), .Z(n44468) );
  IV U57335 ( .A(n44308), .Z(n44312) );
  NOR U57336 ( .A(n44310), .B(n44309), .Z(n44311) );
  IV U57337 ( .A(n44311), .Z(n44318) );
  NOR U57338 ( .A(n44312), .B(n44318), .Z(n44466) );
  NOR U57339 ( .A(n44468), .B(n44466), .Z(n44313) );
  XOR U57340 ( .A(n44465), .B(n44313), .Z(n47694) );
  IV U57341 ( .A(n44314), .Z(n44315) );
  NOR U57342 ( .A(n44316), .B(n44315), .Z(n47693) );
  IV U57343 ( .A(n44317), .Z(n44319) );
  NOR U57344 ( .A(n44319), .B(n44318), .Z(n44462) );
  NOR U57345 ( .A(n47693), .B(n44462), .Z(n44320) );
  XOR U57346 ( .A(n47694), .B(n44320), .Z(n44321) );
  IV U57347 ( .A(n44321), .Z(n47692) );
  XOR U57348 ( .A(n47690), .B(n47692), .Z(n44460) );
  XOR U57349 ( .A(n44322), .B(n44460), .Z(n44451) );
  XOR U57350 ( .A(n44323), .B(n44451), .Z(n47707) );
  XOR U57351 ( .A(n44324), .B(n47707), .Z(n44325) );
  IV U57352 ( .A(n44325), .Z(n47710) );
  XOR U57353 ( .A(n47708), .B(n47710), .Z(n44447) );
  XOR U57354 ( .A(n44446), .B(n44447), .Z(n44444) );
  XOR U57355 ( .A(n44442), .B(n44444), .Z(n51173) );
  XOR U57356 ( .A(n44326), .B(n51173), .Z(n44437) );
  XOR U57357 ( .A(n44438), .B(n44437), .Z(n44435) );
  IV U57358 ( .A(n44327), .Z(n44329) );
  NOR U57359 ( .A(n44329), .B(n44328), .Z(n44439) );
  NOR U57360 ( .A(n44331), .B(n44330), .Z(n44434) );
  NOR U57361 ( .A(n44439), .B(n44434), .Z(n44332) );
  XOR U57362 ( .A(n44435), .B(n44332), .Z(n44432) );
  XOR U57363 ( .A(n44431), .B(n44432), .Z(n47723) );
  XOR U57364 ( .A(n47722), .B(n47723), .Z(n44429) );
  IV U57365 ( .A(n44333), .Z(n44334) );
  NOR U57366 ( .A(n44335), .B(n44334), .Z(n44428) );
  NOR U57367 ( .A(n44337), .B(n44336), .Z(n44364) );
  IV U57368 ( .A(n44364), .Z(n44338) );
  NOR U57369 ( .A(n44338), .B(n44365), .Z(n44426) );
  NOR U57370 ( .A(n44428), .B(n44426), .Z(n44339) );
  XOR U57371 ( .A(n44429), .B(n44339), .Z(n44423) );
  XOR U57372 ( .A(n44424), .B(n44423), .Z(n44418) );
  XOR U57373 ( .A(n44417), .B(n44418), .Z(n44422) );
  XOR U57374 ( .A(n44340), .B(n44342), .Z(n44344) );
  NOR U57375 ( .A(n44342), .B(n44341), .Z(n44343) );
  NOR U57376 ( .A(n44344), .B(n44343), .Z(n44345) );
  NOR U57377 ( .A(n44363), .B(n44345), .Z(n44396) );
  IV U57378 ( .A(n44396), .Z(n44362) );
  XOR U57379 ( .A(n44375), .B(n44346), .Z(n44360) );
  XOR U57380 ( .A(n44348), .B(n44347), .Z(n44380) );
  IV U57381 ( .A(n44349), .Z(n44351) );
  NOR U57382 ( .A(n44351), .B(n44350), .Z(n44378) );
  IV U57383 ( .A(n44378), .Z(n44352) );
  NOR U57384 ( .A(n44380), .B(n44352), .Z(n44391) );
  IV U57385 ( .A(n44391), .Z(n44358) );
  NOR U57386 ( .A(n44354), .B(n44353), .Z(n44355) );
  NOR U57387 ( .A(n44356), .B(n44355), .Z(n44385) );
  IV U57388 ( .A(n44385), .Z(n44357) );
  NOR U57389 ( .A(n44358), .B(n44357), .Z(n44393) );
  IV U57390 ( .A(n44393), .Z(n44359) );
  NOR U57391 ( .A(n44360), .B(n44359), .Z(n44395) );
  IV U57392 ( .A(n44395), .Z(n44361) );
  NOR U57393 ( .A(n44362), .B(n44361), .Z(n44405) );
  IV U57394 ( .A(n44405), .Z(n44368) );
  NOR U57395 ( .A(n44364), .B(n44363), .Z(n44366) );
  XOR U57396 ( .A(n44366), .B(n44365), .Z(n44369) );
  IV U57397 ( .A(n44369), .Z(n44367) );
  NOR U57398 ( .A(n44368), .B(n44367), .Z(n44420) );
  XOR U57399 ( .A(n44422), .B(n44420), .Z(n44415) );
  NOR U57400 ( .A(n44370), .B(n44369), .Z(n44371) );
  NOR U57401 ( .A(n44417), .B(n44371), .Z(n44407) );
  IV U57402 ( .A(n44407), .Z(n44402) );
  IV U57403 ( .A(n44372), .Z(n44374) );
  NOR U57404 ( .A(n44374), .B(n44373), .Z(n47732) );
  IV U57405 ( .A(n47732), .Z(n44400) );
  NOR U57406 ( .A(n44375), .B(n44393), .Z(n44376) );
  XOR U57407 ( .A(n44377), .B(n44376), .Z(n47759) );
  NOR U57408 ( .A(n44379), .B(n44378), .Z(n44381) );
  XOR U57409 ( .A(n44381), .B(n44380), .Z(n47735) );
  IV U57410 ( .A(n47735), .Z(n47748) );
  NOR U57411 ( .A(n44383), .B(n44382), .Z(n44387) );
  IV U57412 ( .A(n44387), .Z(n44384) );
  NOR U57413 ( .A(n44385), .B(n44384), .Z(n44389) );
  NOR U57414 ( .A(n44387), .B(n44386), .Z(n44388) );
  NOR U57415 ( .A(n44389), .B(n44388), .Z(n44390) );
  NOR U57416 ( .A(n44391), .B(n44390), .Z(n44392) );
  NOR U57417 ( .A(n44393), .B(n44392), .Z(n47750) );
  IV U57418 ( .A(n47750), .Z(n47741) );
  NOR U57419 ( .A(n47748), .B(n47741), .Z(n44394) );
  IV U57420 ( .A(n44394), .Z(n47733) );
  XOR U57421 ( .A(n44396), .B(n44395), .Z(n47746) );
  IV U57422 ( .A(n47746), .Z(n47765) );
  NOR U57423 ( .A(n47733), .B(n47765), .Z(n44397) );
  IV U57424 ( .A(n44397), .Z(n44398) );
  NOR U57425 ( .A(n47759), .B(n44398), .Z(n44399) );
  IV U57426 ( .A(n44399), .Z(n44411) );
  NOR U57427 ( .A(n44400), .B(n44411), .Z(n44404) );
  IV U57428 ( .A(n44404), .Z(n44401) );
  NOR U57429 ( .A(n44402), .B(n44401), .Z(n44414) );
  IV U57430 ( .A(n44414), .Z(n44403) );
  NOR U57431 ( .A(n44415), .B(n44403), .Z(n47775) );
  NOR U57432 ( .A(n44405), .B(n44404), .Z(n44406) );
  XOR U57433 ( .A(n44407), .B(n44406), .Z(n51210) );
  IV U57434 ( .A(n44408), .Z(n44410) );
  NOR U57435 ( .A(n44410), .B(n44409), .Z(n47731) );
  IV U57436 ( .A(n47731), .Z(n44412) );
  NOR U57437 ( .A(n44412), .B(n44411), .Z(n51207) );
  IV U57438 ( .A(n51207), .Z(n44413) );
  NOR U57439 ( .A(n51210), .B(n44413), .Z(n47768) );
  IV U57440 ( .A(n47768), .Z(n44416) );
  XOR U57441 ( .A(n44415), .B(n44414), .Z(n47767) );
  NOR U57442 ( .A(n44416), .B(n47767), .Z(n51201) );
  NOR U57443 ( .A(n47775), .B(n51201), .Z(n47730) );
  IV U57444 ( .A(n44417), .Z(n44419) );
  NOR U57445 ( .A(n44419), .B(n44418), .Z(n47780) );
  IV U57446 ( .A(n44420), .Z(n44421) );
  NOR U57447 ( .A(n44422), .B(n44421), .Z(n47778) );
  NOR U57448 ( .A(n47780), .B(n47778), .Z(n47729) );
  IV U57449 ( .A(n44423), .Z(n44425) );
  NOR U57450 ( .A(n44425), .B(n44424), .Z(n51195) );
  IV U57451 ( .A(n44426), .Z(n44427) );
  NOR U57452 ( .A(n44427), .B(n44429), .Z(n51190) );
  NOR U57453 ( .A(n51195), .B(n51190), .Z(n47728) );
  IV U57454 ( .A(n44428), .Z(n44430) );
  NOR U57455 ( .A(n44430), .B(n44429), .Z(n47726) );
  IV U57456 ( .A(n47726), .Z(n47721) );
  IV U57457 ( .A(n44431), .Z(n44433) );
  NOR U57458 ( .A(n44433), .B(n44432), .Z(n51185) );
  IV U57459 ( .A(n44434), .Z(n44436) );
  IV U57460 ( .A(n44435), .Z(n44440) );
  NOR U57461 ( .A(n44436), .B(n44440), .Z(n51176) );
  NOR U57462 ( .A(n44438), .B(n44437), .Z(n47783) );
  IV U57463 ( .A(n44439), .Z(n44441) );
  NOR U57464 ( .A(n44441), .B(n44440), .Z(n51179) );
  NOR U57465 ( .A(n47783), .B(n51179), .Z(n47718) );
  IV U57466 ( .A(n44442), .Z(n44443) );
  NOR U57467 ( .A(n44444), .B(n44443), .Z(n47785) );
  NOR U57468 ( .A(n44445), .B(n51173), .Z(n47788) );
  NOR U57469 ( .A(n47785), .B(n47788), .Z(n47717) );
  IV U57470 ( .A(n44446), .Z(n44448) );
  NOR U57471 ( .A(n44448), .B(n44447), .Z(n47713) );
  IV U57472 ( .A(n44449), .Z(n44453) );
  NOR U57473 ( .A(n44451), .B(n44450), .Z(n44452) );
  IV U57474 ( .A(n44452), .Z(n44455) );
  NOR U57475 ( .A(n44453), .B(n44455), .Z(n47700) );
  IV U57476 ( .A(n47700), .Z(n47697) );
  IV U57477 ( .A(n44454), .Z(n44456) );
  NOR U57478 ( .A(n44456), .B(n44455), .Z(n51149) );
  IV U57479 ( .A(n44457), .Z(n44458) );
  NOR U57480 ( .A(n44458), .B(n44460), .Z(n51146) );
  IV U57481 ( .A(n44459), .Z(n44461) );
  NOR U57482 ( .A(n44461), .B(n44460), .Z(n47796) );
  IV U57483 ( .A(n44462), .Z(n44463) );
  NOR U57484 ( .A(n44463), .B(n47694), .Z(n44464) );
  IV U57485 ( .A(n44464), .Z(n47806) );
  IV U57486 ( .A(n44465), .Z(n44470) );
  IV U57487 ( .A(n44466), .Z(n44467) );
  NOR U57488 ( .A(n44470), .B(n44467), .Z(n47802) );
  IV U57489 ( .A(n44468), .Z(n44469) );
  NOR U57490 ( .A(n44470), .B(n44469), .Z(n47810) );
  IV U57491 ( .A(n44471), .Z(n44472) );
  NOR U57492 ( .A(n44473), .B(n44472), .Z(n51414) );
  IV U57493 ( .A(n44474), .Z(n44475) );
  NOR U57494 ( .A(n44475), .B(n47688), .Z(n51409) );
  NOR U57495 ( .A(n51414), .B(n51409), .Z(n47813) );
  NOR U57496 ( .A(n44476), .B(n47815), .Z(n47685) );
  IV U57497 ( .A(n44477), .Z(n44482) );
  IV U57498 ( .A(n44478), .Z(n44479) );
  NOR U57499 ( .A(n44482), .B(n44479), .Z(n51136) );
  IV U57500 ( .A(n44480), .Z(n44481) );
  NOR U57501 ( .A(n44482), .B(n44481), .Z(n47826) );
  IV U57502 ( .A(n44483), .Z(n44484) );
  NOR U57503 ( .A(n44484), .B(n44489), .Z(n47829) );
  IV U57504 ( .A(n44485), .Z(n44486) );
  NOR U57505 ( .A(n44487), .B(n44486), .Z(n51123) );
  IV U57506 ( .A(n44488), .Z(n44490) );
  NOR U57507 ( .A(n44490), .B(n44489), .Z(n51125) );
  NOR U57508 ( .A(n51123), .B(n51125), .Z(n47684) );
  IV U57509 ( .A(n44491), .Z(n44493) );
  NOR U57510 ( .A(n44493), .B(n44492), .Z(n51110) );
  IV U57511 ( .A(n44494), .Z(n44495) );
  NOR U57512 ( .A(n44496), .B(n44495), .Z(n51107) );
  NOR U57513 ( .A(n51110), .B(n51107), .Z(n47683) );
  IV U57514 ( .A(n44497), .Z(n44499) );
  NOR U57515 ( .A(n44499), .B(n44498), .Z(n51103) );
  IV U57516 ( .A(n44500), .Z(n44503) );
  IV U57517 ( .A(n44501), .Z(n44502) );
  NOR U57518 ( .A(n44503), .B(n44502), .Z(n51447) );
  IV U57519 ( .A(n44504), .Z(n44507) );
  NOR U57520 ( .A(n44505), .B(n44510), .Z(n44506) );
  IV U57521 ( .A(n44506), .Z(n47673) );
  NOR U57522 ( .A(n44507), .B(n47673), .Z(n51452) );
  NOR U57523 ( .A(n51447), .B(n51452), .Z(n51096) );
  IV U57524 ( .A(n44508), .Z(n44509) );
  NOR U57525 ( .A(n44510), .B(n44509), .Z(n47835) );
  IV U57526 ( .A(n44511), .Z(n47668) );
  IV U57527 ( .A(n44512), .Z(n44513) );
  NOR U57528 ( .A(n47668), .B(n44513), .Z(n44518) );
  IV U57529 ( .A(n44514), .Z(n44516) );
  NOR U57530 ( .A(n44516), .B(n44515), .Z(n44517) );
  NOR U57531 ( .A(n44518), .B(n44517), .Z(n54827) );
  IV U57532 ( .A(n54827), .Z(n47838) );
  IV U57533 ( .A(n44519), .Z(n44520) );
  NOR U57534 ( .A(n44520), .B(n47664), .Z(n44521) );
  IV U57535 ( .A(n44521), .Z(n47846) );
  IV U57536 ( .A(n44522), .Z(n44523) );
  NOR U57537 ( .A(n44523), .B(n44525), .Z(n47853) );
  IV U57538 ( .A(n44524), .Z(n44526) );
  NOR U57539 ( .A(n44526), .B(n44525), .Z(n47859) );
  IV U57540 ( .A(n44527), .Z(n44528) );
  NOR U57541 ( .A(n44529), .B(n44528), .Z(n47865) );
  IV U57542 ( .A(n44530), .Z(n44531) );
  NOR U57543 ( .A(n44532), .B(n44531), .Z(n47862) );
  NOR U57544 ( .A(n47865), .B(n47862), .Z(n44533) );
  IV U57545 ( .A(n44533), .Z(n47650) );
  IV U57546 ( .A(n44534), .Z(n44535) );
  NOR U57547 ( .A(n44535), .B(n47639), .Z(n47867) );
  IV U57548 ( .A(n44536), .Z(n44537) );
  NOR U57549 ( .A(n44538), .B(n44537), .Z(n44539) );
  IV U57550 ( .A(n44539), .Z(n47645) );
  IV U57551 ( .A(n44540), .Z(n44545) );
  IV U57552 ( .A(n44541), .Z(n44542) );
  NOR U57553 ( .A(n44545), .B(n44542), .Z(n51066) );
  IV U57554 ( .A(n44543), .Z(n44544) );
  NOR U57555 ( .A(n44545), .B(n44544), .Z(n54808) );
  IV U57556 ( .A(n44546), .Z(n44547) );
  NOR U57557 ( .A(n44551), .B(n44547), .Z(n54802) );
  NOR U57558 ( .A(n54808), .B(n54802), .Z(n47878) );
  IV U57559 ( .A(n44548), .Z(n47880) );
  NOR U57560 ( .A(n44549), .B(n47880), .Z(n44553) );
  IV U57561 ( .A(n44550), .Z(n44552) );
  NOR U57562 ( .A(n44552), .B(n44551), .Z(n47874) );
  NOR U57563 ( .A(n44553), .B(n47874), .Z(n47637) );
  IV U57564 ( .A(n44554), .Z(n44557) );
  IV U57565 ( .A(n44555), .Z(n44556) );
  NOR U57566 ( .A(n44557), .B(n44556), .Z(n51055) );
  IV U57567 ( .A(n44558), .Z(n44559) );
  NOR U57568 ( .A(n44560), .B(n44559), .Z(n47886) );
  NOR U57569 ( .A(n44562), .B(n44561), .Z(n47891) );
  NOR U57570 ( .A(n47886), .B(n47891), .Z(n47635) );
  IV U57571 ( .A(n44563), .Z(n44564) );
  NOR U57572 ( .A(n44565), .B(n44564), .Z(n44566) );
  IV U57573 ( .A(n44566), .Z(n47620) );
  IV U57574 ( .A(n44567), .Z(n44570) );
  IV U57575 ( .A(n44568), .Z(n44577) );
  XOR U57576 ( .A(n44576), .B(n44577), .Z(n44569) );
  NOR U57577 ( .A(n44570), .B(n44569), .Z(n51030) );
  IV U57578 ( .A(n44571), .Z(n44572) );
  NOR U57579 ( .A(n44577), .B(n44572), .Z(n51026) );
  IV U57580 ( .A(n44573), .Z(n44574) );
  NOR U57581 ( .A(n44575), .B(n44574), .Z(n47910) );
  NOR U57582 ( .A(n51026), .B(n47910), .Z(n47595) );
  IV U57583 ( .A(n44576), .Z(n44578) );
  NOR U57584 ( .A(n44578), .B(n44577), .Z(n47593) );
  IV U57585 ( .A(n47593), .Z(n47588) );
  IV U57586 ( .A(n44579), .Z(n44580) );
  NOR U57587 ( .A(n47591), .B(n44580), .Z(n47915) );
  IV U57588 ( .A(n44581), .Z(n47584) );
  IV U57589 ( .A(n44582), .Z(n44583) );
  NOR U57590 ( .A(n47584), .B(n44583), .Z(n47921) );
  NOR U57591 ( .A(n44584), .B(n47584), .Z(n44585) );
  IV U57592 ( .A(n44585), .Z(n47931) );
  IV U57593 ( .A(n44586), .Z(n44587) );
  NOR U57594 ( .A(n44587), .B(n44590), .Z(n47932) );
  IV U57595 ( .A(n44588), .Z(n44589) );
  NOR U57596 ( .A(n44590), .B(n44589), .Z(n44591) );
  IV U57597 ( .A(n44591), .Z(n51020) );
  IV U57598 ( .A(n44592), .Z(n44594) );
  NOR U57599 ( .A(n44594), .B(n44593), .Z(n44595) );
  IV U57600 ( .A(n44595), .Z(n47510) );
  IV U57601 ( .A(n44596), .Z(n47493) );
  NOR U57602 ( .A(n47493), .B(n44597), .Z(n44598) );
  IV U57603 ( .A(n44598), .Z(n44599) );
  NOR U57604 ( .A(n44600), .B(n44599), .Z(n47960) );
  IV U57605 ( .A(n44601), .Z(n44602) );
  NOR U57606 ( .A(n47493), .B(n44602), .Z(n50951) );
  IV U57607 ( .A(n44603), .Z(n44606) );
  IV U57608 ( .A(n44604), .Z(n44605) );
  NOR U57609 ( .A(n44606), .B(n44605), .Z(n50945) );
  IV U57610 ( .A(n44607), .Z(n44608) );
  NOR U57611 ( .A(n44609), .B(n44608), .Z(n47483) );
  IV U57612 ( .A(n47483), .Z(n47478) );
  IV U57613 ( .A(n44610), .Z(n44612) );
  IV U57614 ( .A(n44611), .Z(n47481) );
  NOR U57615 ( .A(n44612), .B(n47481), .Z(n47974) );
  IV U57616 ( .A(n44613), .Z(n44614) );
  NOR U57617 ( .A(n44620), .B(n44614), .Z(n44615) );
  IV U57618 ( .A(n44615), .Z(n50899) );
  IV U57619 ( .A(n44616), .Z(n44617) );
  NOR U57620 ( .A(n44618), .B(n44617), .Z(n50896) );
  IV U57621 ( .A(n44619), .Z(n44621) );
  NOR U57622 ( .A(n44621), .B(n44620), .Z(n50901) );
  NOR U57623 ( .A(n50896), .B(n50901), .Z(n44622) );
  IV U57624 ( .A(n44622), .Z(n47443) );
  IV U57625 ( .A(n44623), .Z(n44625) );
  IV U57626 ( .A(n44624), .Z(n47441) );
  NOR U57627 ( .A(n44625), .B(n47441), .Z(n50893) );
  IV U57628 ( .A(n44626), .Z(n44628) );
  NOR U57629 ( .A(n44628), .B(n44627), .Z(n50879) );
  IV U57630 ( .A(n44629), .Z(n44630) );
  NOR U57631 ( .A(n44631), .B(n44630), .Z(n44632) );
  IV U57632 ( .A(n44632), .Z(n47429) );
  IV U57633 ( .A(n44633), .Z(n44635) );
  NOR U57634 ( .A(n44635), .B(n44634), .Z(n48009) );
  IV U57635 ( .A(n44636), .Z(n44638) );
  NOR U57636 ( .A(n44638), .B(n44637), .Z(n48007) );
  NOR U57637 ( .A(n48009), .B(n48007), .Z(n51623) );
  IV U57638 ( .A(n44639), .Z(n48023) );
  NOR U57639 ( .A(n44640), .B(n48023), .Z(n47403) );
  IV U57640 ( .A(n44641), .Z(n44642) );
  NOR U57641 ( .A(n44643), .B(n44642), .Z(n44647) );
  NOR U57642 ( .A(n44645), .B(n44644), .Z(n44646) );
  NOR U57643 ( .A(n44647), .B(n44646), .Z(n54624) );
  IV U57644 ( .A(n54624), .Z(n50821) );
  IV U57645 ( .A(n44648), .Z(n44651) );
  IV U57646 ( .A(n44649), .Z(n44650) );
  NOR U57647 ( .A(n44651), .B(n44650), .Z(n48027) );
  IV U57648 ( .A(n44652), .Z(n44653) );
  NOR U57649 ( .A(n44653), .B(n50810), .Z(n50805) );
  NOR U57650 ( .A(n48027), .B(n50805), .Z(n51671) );
  IV U57651 ( .A(n44654), .Z(n44655) );
  NOR U57652 ( .A(n44656), .B(n44655), .Z(n54594) );
  NOR U57653 ( .A(n54594), .B(n54611), .Z(n48028) );
  IV U57654 ( .A(n44657), .Z(n44658) );
  NOR U57655 ( .A(n44658), .B(n44664), .Z(n44659) );
  IV U57656 ( .A(n44659), .Z(n50795) );
  IV U57657 ( .A(n44660), .Z(n44662) );
  NOR U57658 ( .A(n44662), .B(n44661), .Z(n48033) );
  IV U57659 ( .A(n44663), .Z(n44665) );
  NOR U57660 ( .A(n44665), .B(n44664), .Z(n50797) );
  NOR U57661 ( .A(n48033), .B(n50797), .Z(n44666) );
  IV U57662 ( .A(n44666), .Z(n47384) );
  IV U57663 ( .A(n44667), .Z(n44668) );
  NOR U57664 ( .A(n44669), .B(n44668), .Z(n47363) );
  IV U57665 ( .A(n47363), .Z(n47358) );
  IV U57666 ( .A(n44670), .Z(n44671) );
  NOR U57667 ( .A(n44672), .B(n44671), .Z(n48059) );
  IV U57668 ( .A(n44673), .Z(n44675) );
  NOR U57669 ( .A(n44675), .B(n44674), .Z(n48056) );
  IV U57670 ( .A(n44676), .Z(n44679) );
  NOR U57671 ( .A(n44677), .B(n47348), .Z(n44678) );
  IV U57672 ( .A(n44678), .Z(n47355) );
  NOR U57673 ( .A(n44679), .B(n47355), .Z(n48068) );
  IV U57674 ( .A(n44680), .Z(n44682) );
  NOR U57675 ( .A(n44682), .B(n44681), .Z(n51727) );
  NOR U57676 ( .A(n51732), .B(n51727), .Z(n50764) );
  IV U57677 ( .A(n44683), .Z(n44684) );
  NOR U57678 ( .A(n44684), .B(n47343), .Z(n50756) );
  IV U57679 ( .A(n44685), .Z(n48090) );
  NOR U57680 ( .A(n44686), .B(n48090), .Z(n44690) );
  IV U57681 ( .A(n44687), .Z(n44688) );
  NOR U57682 ( .A(n44689), .B(n44688), .Z(n48087) );
  NOR U57683 ( .A(n44690), .B(n48087), .Z(n47330) );
  IV U57684 ( .A(n44691), .Z(n44692) );
  NOR U57685 ( .A(n48093), .B(n44692), .Z(n50741) );
  NOR U57686 ( .A(n44694), .B(n44693), .Z(n50732) );
  IV U57687 ( .A(n44695), .Z(n44696) );
  NOR U57688 ( .A(n44697), .B(n44696), .Z(n50738) );
  NOR U57689 ( .A(n50732), .B(n50738), .Z(n47329) );
  IV U57690 ( .A(n44698), .Z(n44700) );
  NOR U57691 ( .A(n44700), .B(n44699), .Z(n50727) );
  NOR U57692 ( .A(n50727), .B(n50734), .Z(n47328) );
  IV U57693 ( .A(n44701), .Z(n44703) );
  NOR U57694 ( .A(n44703), .B(n44702), .Z(n51758) );
  IV U57695 ( .A(n44704), .Z(n44705) );
  NOR U57696 ( .A(n44706), .B(n44705), .Z(n51754) );
  NOR U57697 ( .A(n51758), .B(n51754), .Z(n50726) );
  IV U57698 ( .A(n44707), .Z(n44708) );
  NOR U57699 ( .A(n44709), .B(n44708), .Z(n50722) );
  IV U57700 ( .A(n44710), .Z(n44711) );
  NOR U57701 ( .A(n44712), .B(n44711), .Z(n48094) );
  NOR U57702 ( .A(n50722), .B(n48094), .Z(n47327) );
  IV U57703 ( .A(n44713), .Z(n44714) );
  NOR U57704 ( .A(n44715), .B(n44714), .Z(n47315) );
  IV U57705 ( .A(n44716), .Z(n44718) );
  NOR U57706 ( .A(n44718), .B(n44717), .Z(n47312) );
  IV U57707 ( .A(n47312), .Z(n47307) );
  IV U57708 ( .A(n44719), .Z(n47304) );
  IV U57709 ( .A(n44720), .Z(n44721) );
  NOR U57710 ( .A(n47304), .B(n44721), .Z(n48109) );
  IV U57711 ( .A(n44722), .Z(n44723) );
  NOR U57712 ( .A(n44723), .B(n47304), .Z(n48106) );
  IV U57713 ( .A(n44724), .Z(n44725) );
  NOR U57714 ( .A(n44726), .B(n44725), .Z(n48117) );
  NOR U57715 ( .A(n44727), .B(n50685), .Z(n44731) );
  IV U57716 ( .A(n44728), .Z(n48125) );
  NOR U57717 ( .A(n44729), .B(n48125), .Z(n44730) );
  NOR U57718 ( .A(n44731), .B(n44730), .Z(n47281) );
  IV U57719 ( .A(n44732), .Z(n44738) );
  NOR U57720 ( .A(n44734), .B(n44733), .Z(n44735) );
  IV U57721 ( .A(n44735), .Z(n47278) );
  NOR U57722 ( .A(n44736), .B(n47278), .Z(n44737) );
  IV U57723 ( .A(n44737), .Z(n47272) );
  NOR U57724 ( .A(n44738), .B(n47272), .Z(n48135) );
  IV U57725 ( .A(n44739), .Z(n44741) );
  IV U57726 ( .A(n44740), .Z(n47261) );
  NOR U57727 ( .A(n44741), .B(n47261), .Z(n50669) );
  IV U57728 ( .A(n44742), .Z(n44743) );
  NOR U57729 ( .A(n44744), .B(n44743), .Z(n44745) );
  IV U57730 ( .A(n44745), .Z(n48139) );
  IV U57731 ( .A(n44746), .Z(n44747) );
  NOR U57732 ( .A(n47241), .B(n44747), .Z(n48150) );
  IV U57733 ( .A(n44748), .Z(n44749) );
  NOR U57734 ( .A(n44752), .B(n44749), .Z(n48152) );
  NOR U57735 ( .A(n48150), .B(n48152), .Z(n47231) );
  IV U57736 ( .A(n44750), .Z(n44751) );
  NOR U57737 ( .A(n44752), .B(n44751), .Z(n50659) );
  IV U57738 ( .A(n44753), .Z(n47228) );
  IV U57739 ( .A(n44754), .Z(n44755) );
  NOR U57740 ( .A(n47228), .B(n44755), .Z(n50654) );
  NOR U57741 ( .A(n50659), .B(n50654), .Z(n47230) );
  IV U57742 ( .A(n44756), .Z(n44757) );
  NOR U57743 ( .A(n44757), .B(n47220), .Z(n44758) );
  IV U57744 ( .A(n44758), .Z(n48159) );
  IV U57745 ( .A(n44759), .Z(n48177) );
  NOR U57746 ( .A(n44760), .B(n48177), .Z(n47207) );
  IV U57747 ( .A(n44761), .Z(n44763) );
  NOR U57748 ( .A(n44763), .B(n44762), .Z(n51875) );
  NOR U57749 ( .A(n44765), .B(n44764), .Z(n54464) );
  NOR U57750 ( .A(n51875), .B(n54464), .Z(n48174) );
  NOR U57751 ( .A(n44766), .B(n48185), .Z(n44770) );
  IV U57752 ( .A(n44767), .Z(n44769) );
  NOR U57753 ( .A(n44769), .B(n44768), .Z(n48181) );
  NOR U57754 ( .A(n44770), .B(n48181), .Z(n47199) );
  IV U57755 ( .A(n44771), .Z(n44773) );
  NOR U57756 ( .A(n44773), .B(n44772), .Z(n50632) );
  IV U57757 ( .A(n44774), .Z(n44776) );
  IV U57758 ( .A(n44775), .Z(n44784) );
  NOR U57759 ( .A(n44776), .B(n44784), .Z(n48192) );
  IV U57760 ( .A(n44777), .Z(n44778) );
  NOR U57761 ( .A(n44779), .B(n44778), .Z(n50635) );
  NOR U57762 ( .A(n48192), .B(n50635), .Z(n47198) );
  NOR U57763 ( .A(n44781), .B(n44780), .Z(n50626) );
  IV U57764 ( .A(n44782), .Z(n44783) );
  NOR U57765 ( .A(n44784), .B(n44783), .Z(n50629) );
  NOR U57766 ( .A(n50626), .B(n50629), .Z(n47197) );
  IV U57767 ( .A(n44785), .Z(n44787) );
  NOR U57768 ( .A(n44787), .B(n44786), .Z(n48198) );
  IV U57769 ( .A(n44788), .Z(n44790) );
  NOR U57770 ( .A(n44790), .B(n44789), .Z(n48195) );
  IV U57771 ( .A(n44791), .Z(n44792) );
  NOR U57772 ( .A(n47183), .B(n44792), .Z(n44793) );
  IV U57773 ( .A(n44793), .Z(n47186) );
  IV U57774 ( .A(n44794), .Z(n44795) );
  NOR U57775 ( .A(n44796), .B(n44795), .Z(n50615) );
  IV U57776 ( .A(n44797), .Z(n44798) );
  NOR U57777 ( .A(n44799), .B(n44798), .Z(n50619) );
  NOR U57778 ( .A(n50615), .B(n50619), .Z(n44800) );
  IV U57779 ( .A(n44800), .Z(n47178) );
  NOR U57780 ( .A(n44802), .B(n44801), .Z(n50602) );
  IV U57781 ( .A(n44803), .Z(n44805) );
  IV U57782 ( .A(n44804), .Z(n44807) );
  NOR U57783 ( .A(n44805), .B(n44807), .Z(n51897) );
  NOR U57784 ( .A(n50602), .B(n51897), .Z(n47177) );
  IV U57785 ( .A(n44806), .Z(n44808) );
  NOR U57786 ( .A(n44808), .B(n44807), .Z(n50612) );
  IV U57787 ( .A(n50612), .Z(n51893) );
  IV U57788 ( .A(n44809), .Z(n44810) );
  NOR U57789 ( .A(n44811), .B(n44810), .Z(n50604) );
  IV U57790 ( .A(n44812), .Z(n44813) );
  NOR U57791 ( .A(n44814), .B(n44813), .Z(n50606) );
  NOR U57792 ( .A(n50604), .B(n50606), .Z(n44815) );
  IV U57793 ( .A(n44815), .Z(n47175) );
  IV U57794 ( .A(n44816), .Z(n44821) );
  IV U57795 ( .A(n44817), .Z(n44818) );
  NOR U57796 ( .A(n44821), .B(n44818), .Z(n50598) );
  IV U57797 ( .A(n44819), .Z(n44820) );
  NOR U57798 ( .A(n44821), .B(n44820), .Z(n50595) );
  IV U57799 ( .A(n44822), .Z(n44823) );
  NOR U57800 ( .A(n44823), .B(n47169), .Z(n48216) );
  IV U57801 ( .A(n44824), .Z(n44825) );
  NOR U57802 ( .A(n44825), .B(n47146), .Z(n48224) );
  IV U57803 ( .A(n44826), .Z(n44828) );
  NOR U57804 ( .A(n44828), .B(n44827), .Z(n50560) );
  IV U57805 ( .A(n44829), .Z(n44830) );
  NOR U57806 ( .A(n44831), .B(n44830), .Z(n48229) );
  NOR U57807 ( .A(n50560), .B(n48229), .Z(n47144) );
  IV U57808 ( .A(n44832), .Z(n44833) );
  NOR U57809 ( .A(n44834), .B(n44833), .Z(n50562) );
  IV U57810 ( .A(n44835), .Z(n44836) );
  NOR U57811 ( .A(n44837), .B(n44836), .Z(n50557) );
  NOR U57812 ( .A(n50562), .B(n50557), .Z(n47143) );
  IV U57813 ( .A(n44838), .Z(n44839) );
  NOR U57814 ( .A(n44840), .B(n44839), .Z(n50544) );
  IV U57815 ( .A(n44841), .Z(n44842) );
  NOR U57816 ( .A(n44843), .B(n44842), .Z(n54369) );
  IV U57817 ( .A(n44844), .Z(n44846) );
  NOR U57818 ( .A(n44846), .B(n44845), .Z(n51947) );
  NOR U57819 ( .A(n54369), .B(n51947), .Z(n48251) );
  IV U57820 ( .A(n44847), .Z(n44849) );
  NOR U57821 ( .A(n44849), .B(n44848), .Z(n54353) );
  NOR U57822 ( .A(n44851), .B(n44850), .Z(n54358) );
  NOR U57823 ( .A(n54353), .B(n54358), .Z(n48259) );
  IV U57824 ( .A(n44852), .Z(n44853) );
  NOR U57825 ( .A(n44854), .B(n44853), .Z(n50529) );
  IV U57826 ( .A(n44855), .Z(n44860) );
  IV U57827 ( .A(n44856), .Z(n44857) );
  NOR U57828 ( .A(n44860), .B(n44857), .Z(n50526) );
  IV U57829 ( .A(n44858), .Z(n44859) );
  NOR U57830 ( .A(n44860), .B(n44859), .Z(n48265) );
  IV U57831 ( .A(n44861), .Z(n44864) );
  NOR U57832 ( .A(n44862), .B(n47110), .Z(n44863) );
  IV U57833 ( .A(n44863), .Z(n44869) );
  NOR U57834 ( .A(n44864), .B(n44869), .Z(n48260) );
  NOR U57835 ( .A(n48265), .B(n48260), .Z(n47115) );
  IV U57836 ( .A(n44865), .Z(n44866) );
  NOR U57837 ( .A(n44867), .B(n44866), .Z(n50519) );
  IV U57838 ( .A(n44868), .Z(n44870) );
  NOR U57839 ( .A(n44870), .B(n44869), .Z(n48263) );
  NOR U57840 ( .A(n50519), .B(n48263), .Z(n47114) );
  IV U57841 ( .A(n44871), .Z(n44872) );
  NOR U57842 ( .A(n47113), .B(n44872), .Z(n44873) );
  IV U57843 ( .A(n44873), .Z(n48270) );
  IV U57844 ( .A(n44874), .Z(n44875) );
  NOR U57845 ( .A(n47096), .B(n44875), .Z(n47093) );
  IV U57846 ( .A(n47093), .Z(n47083) );
  IV U57847 ( .A(n44876), .Z(n44877) );
  NOR U57848 ( .A(n44877), .B(n47067), .Z(n50484) );
  XOR U57849 ( .A(n44887), .B(n47031), .Z(n44883) );
  IV U57850 ( .A(n44881), .Z(n44882) );
  NOR U57851 ( .A(n44883), .B(n44882), .Z(n50413) );
  IV U57852 ( .A(n44884), .Z(n44885) );
  NOR U57853 ( .A(n44886), .B(n44885), .Z(n48297) );
  IV U57854 ( .A(n44887), .Z(n44888) );
  NOR U57855 ( .A(n47031), .B(n44888), .Z(n50407) );
  NOR U57856 ( .A(n48297), .B(n50407), .Z(n44889) );
  IV U57857 ( .A(n44889), .Z(n47029) );
  IV U57858 ( .A(n44890), .Z(n44891) );
  NOR U57859 ( .A(n44892), .B(n44891), .Z(n48295) );
  NOR U57860 ( .A(n44894), .B(n44893), .Z(n48300) );
  IV U57861 ( .A(n44895), .Z(n44897) );
  NOR U57862 ( .A(n44897), .B(n44896), .Z(n44898) );
  IV U57863 ( .A(n44898), .Z(n48306) );
  IV U57864 ( .A(n44899), .Z(n44900) );
  NOR U57865 ( .A(n44901), .B(n44900), .Z(n50403) );
  IV U57866 ( .A(n44902), .Z(n44904) );
  NOR U57867 ( .A(n44904), .B(n44903), .Z(n48312) );
  NOR U57868 ( .A(n50403), .B(n48312), .Z(n44905) );
  IV U57869 ( .A(n44905), .Z(n47021) );
  IV U57870 ( .A(n44906), .Z(n44907) );
  NOR U57871 ( .A(n44907), .B(n44912), .Z(n50398) );
  IV U57872 ( .A(n44908), .Z(n44909) );
  NOR U57873 ( .A(n44910), .B(n44909), .Z(n48315) );
  IV U57874 ( .A(n44911), .Z(n44913) );
  NOR U57875 ( .A(n44913), .B(n44912), .Z(n50395) );
  NOR U57876 ( .A(n48315), .B(n50395), .Z(n47020) );
  IV U57877 ( .A(n44914), .Z(n44915) );
  NOR U57878 ( .A(n44916), .B(n44915), .Z(n52047) );
  IV U57879 ( .A(n44917), .Z(n44918) );
  NOR U57880 ( .A(n44919), .B(n44918), .Z(n52042) );
  NOR U57881 ( .A(n52047), .B(n52042), .Z(n48320) );
  IV U57882 ( .A(n44920), .Z(n44921) );
  NOR U57883 ( .A(n44921), .B(n47004), .Z(n50387) );
  IV U57884 ( .A(n44922), .Z(n44924) );
  IV U57885 ( .A(n44923), .Z(n47009) );
  NOR U57886 ( .A(n44924), .B(n47009), .Z(n48325) );
  NOR U57887 ( .A(n50387), .B(n48325), .Z(n47012) );
  IV U57888 ( .A(n44925), .Z(n44928) );
  NOR U57889 ( .A(n44926), .B(n44932), .Z(n44927) );
  IV U57890 ( .A(n44927), .Z(n46993) );
  NOR U57891 ( .A(n44928), .B(n46993), .Z(n50362) );
  IV U57892 ( .A(n44929), .Z(n48333) );
  NOR U57893 ( .A(n48333), .B(n44930), .Z(n44934) );
  IV U57894 ( .A(n44931), .Z(n44933) );
  NOR U57895 ( .A(n44933), .B(n44932), .Z(n48329) );
  NOR U57896 ( .A(n44934), .B(n48329), .Z(n44935) );
  IV U57897 ( .A(n44935), .Z(n46991) );
  IV U57898 ( .A(n44936), .Z(n44937) );
  NOR U57899 ( .A(n46988), .B(n44937), .Z(n50354) );
  IV U57900 ( .A(n44938), .Z(n44939) );
  NOR U57901 ( .A(n44939), .B(n44945), .Z(n44940) );
  IV U57902 ( .A(n44940), .Z(n48340) );
  IV U57903 ( .A(n44941), .Z(n44942) );
  NOR U57904 ( .A(n44943), .B(n44942), .Z(n50347) );
  IV U57905 ( .A(n44944), .Z(n44946) );
  NOR U57906 ( .A(n44946), .B(n44945), .Z(n48346) );
  NOR U57907 ( .A(n50347), .B(n48346), .Z(n46983) );
  IV U57908 ( .A(n44947), .Z(n44948) );
  NOR U57909 ( .A(n44949), .B(n44948), .Z(n44950) );
  IV U57910 ( .A(n44950), .Z(n50328) );
  IV U57911 ( .A(n44951), .Z(n44953) );
  NOR U57912 ( .A(n44953), .B(n44952), .Z(n50330) );
  IV U57913 ( .A(n44954), .Z(n46897) );
  IV U57914 ( .A(n44955), .Z(n44956) );
  NOR U57915 ( .A(n46897), .B(n44956), .Z(n50317) );
  NOR U57916 ( .A(n44958), .B(n44957), .Z(n48406) );
  NOR U57917 ( .A(n48406), .B(n54196), .Z(n46895) );
  IV U57918 ( .A(n44959), .Z(n44960) );
  NOR U57919 ( .A(n44961), .B(n44960), .Z(n44962) );
  IV U57920 ( .A(n44962), .Z(n46890) );
  IV U57921 ( .A(n44963), .Z(n44964) );
  NOR U57922 ( .A(n44964), .B(n44966), .Z(n50295) );
  IV U57923 ( .A(n44965), .Z(n44967) );
  NOR U57924 ( .A(n44967), .B(n44966), .Z(n50293) );
  IV U57925 ( .A(n44968), .Z(n48423) );
  NOR U57926 ( .A(n44969), .B(n48423), .Z(n44972) );
  NOR U57927 ( .A(n44971), .B(n44970), .Z(n48418) );
  NOR U57928 ( .A(n44972), .B(n48418), .Z(n46872) );
  IV U57929 ( .A(n44973), .Z(n44976) );
  NOR U57930 ( .A(n44974), .B(n46860), .Z(n44975) );
  IV U57931 ( .A(n44975), .Z(n46869) );
  NOR U57932 ( .A(n44976), .B(n46869), .Z(n46864) );
  IV U57933 ( .A(n44977), .Z(n44979) );
  NOR U57934 ( .A(n44979), .B(n44978), .Z(n46848) );
  IV U57935 ( .A(n46848), .Z(n46843) );
  IV U57936 ( .A(n44980), .Z(n44983) );
  IV U57937 ( .A(n44981), .Z(n44982) );
  NOR U57938 ( .A(n44983), .B(n44982), .Z(n50279) );
  IV U57939 ( .A(n44984), .Z(n44987) );
  NOR U57940 ( .A(n44985), .B(n44992), .Z(n44986) );
  IV U57941 ( .A(n44986), .Z(n44989) );
  NOR U57942 ( .A(n44987), .B(n44989), .Z(n50276) );
  IV U57943 ( .A(n44988), .Z(n44990) );
  NOR U57944 ( .A(n44990), .B(n44989), .Z(n48453) );
  NOR U57945 ( .A(n44992), .B(n44991), .Z(n50267) );
  IV U57946 ( .A(n44993), .Z(n44994) );
  NOR U57947 ( .A(n44995), .B(n44994), .Z(n50264) );
  IV U57948 ( .A(n44996), .Z(n44997) );
  NOR U57949 ( .A(n46826), .B(n44997), .Z(n48459) );
  NOR U57950 ( .A(n44998), .B(n52196), .Z(n44999) );
  IV U57951 ( .A(n44999), .Z(n48462) );
  IV U57952 ( .A(n45000), .Z(n45003) );
  IV U57953 ( .A(n45001), .Z(n45002) );
  NOR U57954 ( .A(n45003), .B(n45002), .Z(n54110) );
  IV U57955 ( .A(n45004), .Z(n45005) );
  NOR U57956 ( .A(n45006), .B(n45005), .Z(n52199) );
  NOR U57957 ( .A(n54110), .B(n52199), .Z(n48465) );
  IV U57958 ( .A(n48465), .Z(n46821) );
  IV U57959 ( .A(n45007), .Z(n45008) );
  NOR U57960 ( .A(n45009), .B(n45008), .Z(n48467) );
  NOR U57961 ( .A(n45011), .B(n45010), .Z(n50256) );
  NOR U57962 ( .A(n48467), .B(n50256), .Z(n46820) );
  IV U57963 ( .A(n45012), .Z(n45013) );
  NOR U57964 ( .A(n45014), .B(n45013), .Z(n48469) );
  IV U57965 ( .A(n45015), .Z(n45018) );
  IV U57966 ( .A(n45016), .Z(n45017) );
  NOR U57967 ( .A(n45018), .B(n45017), .Z(n50250) );
  NOR U57968 ( .A(n48469), .B(n50250), .Z(n46819) );
  IV U57969 ( .A(n45019), .Z(n45020) );
  NOR U57970 ( .A(n45020), .B(n45021), .Z(n48472) );
  NOR U57971 ( .A(n45022), .B(n45021), .Z(n48478) );
  IV U57972 ( .A(n45023), .Z(n45028) );
  IV U57973 ( .A(n45024), .Z(n45025) );
  NOR U57974 ( .A(n45028), .B(n45025), .Z(n48475) );
  IV U57975 ( .A(n45026), .Z(n45027) );
  NOR U57976 ( .A(n45028), .B(n45027), .Z(n50245) );
  IV U57977 ( .A(n45029), .Z(n45030) );
  NOR U57978 ( .A(n45030), .B(n46817), .Z(n50242) );
  IV U57979 ( .A(n45031), .Z(n45033) );
  NOR U57980 ( .A(n45033), .B(n45032), .Z(n45034) );
  IV U57981 ( .A(n45034), .Z(n48492) );
  IV U57982 ( .A(n45035), .Z(n45036) );
  NOR U57983 ( .A(n45036), .B(n45038), .Z(n50237) );
  IV U57984 ( .A(n45037), .Z(n45039) );
  NOR U57985 ( .A(n45039), .B(n45038), .Z(n48494) );
  NOR U57986 ( .A(n50237), .B(n48494), .Z(n45040) );
  IV U57987 ( .A(n45040), .Z(n46808) );
  IV U57988 ( .A(n45041), .Z(n45043) );
  NOR U57989 ( .A(n45043), .B(n45042), .Z(n50235) );
  IV U57990 ( .A(n45044), .Z(n45045) );
  NOR U57991 ( .A(n45045), .B(n46794), .Z(n45046) );
  IV U57992 ( .A(n45046), .Z(n48502) );
  IV U57993 ( .A(n45047), .Z(n45048) );
  NOR U57994 ( .A(n45049), .B(n45048), .Z(n48516) );
  IV U57995 ( .A(n45050), .Z(n46789) );
  IV U57996 ( .A(n45051), .Z(n45052) );
  NOR U57997 ( .A(n46789), .B(n45052), .Z(n48519) );
  IV U57998 ( .A(n45053), .Z(n45054) );
  NOR U57999 ( .A(n45055), .B(n45054), .Z(n45056) );
  IV U58000 ( .A(n45056), .Z(n48534) );
  IV U58001 ( .A(n45057), .Z(n48537) );
  NOR U58002 ( .A(n45058), .B(n48537), .Z(n45062) );
  IV U58003 ( .A(n45059), .Z(n45060) );
  NOR U58004 ( .A(n45061), .B(n45060), .Z(n48540) );
  NOR U58005 ( .A(n45062), .B(n48540), .Z(n45063) );
  IV U58006 ( .A(n45063), .Z(n46780) );
  IV U58007 ( .A(n45064), .Z(n45065) );
  NOR U58008 ( .A(n45065), .B(n46777), .Z(n50220) );
  NOR U58009 ( .A(n45066), .B(n48547), .Z(n46771) );
  IV U58010 ( .A(n45067), .Z(n45068) );
  NOR U58011 ( .A(n45068), .B(n45071), .Z(n45069) );
  IV U58012 ( .A(n45069), .Z(n48570) );
  IV U58013 ( .A(n45070), .Z(n45072) );
  NOR U58014 ( .A(n45072), .B(n45071), .Z(n46756) );
  IV U58015 ( .A(n46756), .Z(n46751) );
  IV U58016 ( .A(n45073), .Z(n45075) );
  NOR U58017 ( .A(n45075), .B(n45074), .Z(n45076) );
  IV U58018 ( .A(n45076), .Z(n50203) );
  IV U58019 ( .A(n45077), .Z(n45083) );
  NOR U58020 ( .A(n45078), .B(n45086), .Z(n45079) );
  IV U58021 ( .A(n45079), .Z(n45080) );
  NOR U58022 ( .A(n45081), .B(n45080), .Z(n45082) );
  IV U58023 ( .A(n45082), .Z(n45088) );
  NOR U58024 ( .A(n45083), .B(n45088), .Z(n50193) );
  IV U58025 ( .A(n45084), .Z(n45085) );
  NOR U58026 ( .A(n45086), .B(n45085), .Z(n50187) );
  IV U58027 ( .A(n45087), .Z(n45089) );
  NOR U58028 ( .A(n45089), .B(n45088), .Z(n50189) );
  NOR U58029 ( .A(n50187), .B(n50189), .Z(n45090) );
  IV U58030 ( .A(n45090), .Z(n46723) );
  IV U58031 ( .A(n45091), .Z(n46721) );
  IV U58032 ( .A(n45092), .Z(n45093) );
  NOR U58033 ( .A(n46721), .B(n45093), .Z(n48594) );
  NOR U58034 ( .A(n45094), .B(n52360), .Z(n45095) );
  IV U58035 ( .A(n45095), .Z(n50179) );
  IV U58036 ( .A(n45096), .Z(n45097) );
  NOR U58037 ( .A(n45098), .B(n45097), .Z(n50173) );
  IV U58038 ( .A(n45099), .Z(n45101) );
  IV U58039 ( .A(n45100), .Z(n45105) );
  NOR U58040 ( .A(n45101), .B(n45105), .Z(n48601) );
  NOR U58041 ( .A(n50173), .B(n48601), .Z(n45102) );
  IV U58042 ( .A(n45102), .Z(n46713) );
  IV U58043 ( .A(n45103), .Z(n45104) );
  NOR U58044 ( .A(n45105), .B(n45104), .Z(n48598) );
  NOR U58045 ( .A(n45107), .B(n45106), .Z(n50170) );
  IV U58046 ( .A(n45108), .Z(n45109) );
  NOR U58047 ( .A(n45109), .B(n45114), .Z(n48603) );
  NOR U58048 ( .A(n50170), .B(n48603), .Z(n46712) );
  IV U58049 ( .A(n45110), .Z(n45112) );
  NOR U58050 ( .A(n45112), .B(n45111), .Z(n50166) );
  IV U58051 ( .A(n45113), .Z(n45115) );
  NOR U58052 ( .A(n45115), .B(n45114), .Z(n48605) );
  NOR U58053 ( .A(n50166), .B(n48605), .Z(n46711) );
  NOR U58054 ( .A(n45116), .B(n48609), .Z(n46710) );
  IV U58055 ( .A(n45117), .Z(n45119) );
  IV U58056 ( .A(n45118), .Z(n45121) );
  NOR U58057 ( .A(n45119), .B(n45121), .Z(n48615) );
  IV U58058 ( .A(n45120), .Z(n45122) );
  NOR U58059 ( .A(n45122), .B(n45121), .Z(n48612) );
  NOR U58060 ( .A(n45123), .B(n48622), .Z(n46706) );
  IV U58061 ( .A(n45124), .Z(n45126) );
  NOR U58062 ( .A(n45126), .B(n45125), .Z(n50151) );
  IV U58063 ( .A(n45127), .Z(n45129) );
  NOR U58064 ( .A(n45129), .B(n45128), .Z(n48627) );
  NOR U58065 ( .A(n50151), .B(n48627), .Z(n45130) );
  IV U58066 ( .A(n45130), .Z(n46693) );
  IV U58067 ( .A(n45131), .Z(n45132) );
  NOR U58068 ( .A(n45133), .B(n45132), .Z(n48629) );
  IV U58069 ( .A(n45134), .Z(n45135) );
  NOR U58070 ( .A(n45136), .B(n45135), .Z(n50137) );
  NOR U58071 ( .A(n48629), .B(n50137), .Z(n46685) );
  IV U58072 ( .A(n45137), .Z(n45139) );
  NOR U58073 ( .A(n45139), .B(n45138), .Z(n48632) );
  IV U58074 ( .A(n45140), .Z(n45147) );
  IV U58075 ( .A(n45141), .Z(n45149) );
  NOR U58076 ( .A(n45142), .B(n45149), .Z(n45143) );
  IV U58077 ( .A(n45143), .Z(n45144) );
  NOR U58078 ( .A(n45145), .B(n45144), .Z(n45146) );
  IV U58079 ( .A(n45146), .Z(n45151) );
  NOR U58080 ( .A(n45147), .B(n45151), .Z(n48634) );
  NOR U58081 ( .A(n48632), .B(n48634), .Z(n46684) );
  NOR U58082 ( .A(n45149), .B(n45148), .Z(n50131) );
  IV U58083 ( .A(n45150), .Z(n45152) );
  NOR U58084 ( .A(n45152), .B(n45151), .Z(n50134) );
  NOR U58085 ( .A(n50131), .B(n50134), .Z(n46683) );
  NOR U58086 ( .A(n45153), .B(n48638), .Z(n46682) );
  IV U58087 ( .A(n45154), .Z(n45155) );
  NOR U58088 ( .A(n45155), .B(n46656), .Z(n50114) );
  IV U58089 ( .A(n45156), .Z(n46653) );
  IV U58090 ( .A(n45157), .Z(n45158) );
  NOR U58091 ( .A(n46653), .B(n45158), .Z(n50104) );
  IV U58092 ( .A(n45159), .Z(n45162) );
  NOR U58093 ( .A(n46644), .B(n45160), .Z(n45161) );
  IV U58094 ( .A(n45161), .Z(n46646) );
  NOR U58095 ( .A(n45162), .B(n46646), .Z(n48652) );
  IV U58096 ( .A(n45163), .Z(n45165) );
  NOR U58097 ( .A(n45165), .B(n45164), .Z(n50107) );
  NOR U58098 ( .A(n48652), .B(n50107), .Z(n46650) );
  IV U58099 ( .A(n45166), .Z(n45168) );
  IV U58100 ( .A(n45167), .Z(n46628) );
  NOR U58101 ( .A(n45168), .B(n46628), .Z(n45169) );
  IV U58102 ( .A(n45169), .Z(n48657) );
  IV U58103 ( .A(n45170), .Z(n45175) );
  IV U58104 ( .A(n45171), .Z(n45172) );
  NOR U58105 ( .A(n45175), .B(n45172), .Z(n50090) );
  IV U58106 ( .A(n45173), .Z(n45174) );
  NOR U58107 ( .A(n45175), .B(n45174), .Z(n48674) );
  IV U58108 ( .A(n45176), .Z(n45177) );
  NOR U58109 ( .A(n45178), .B(n45177), .Z(n45179) );
  IV U58110 ( .A(n45179), .Z(n50082) );
  IV U58111 ( .A(n45180), .Z(n45182) );
  NOR U58112 ( .A(n45182), .B(n45181), .Z(n50084) );
  IV U58113 ( .A(n45183), .Z(n45185) );
  NOR U58114 ( .A(n45185), .B(n45184), .Z(n50080) );
  IV U58115 ( .A(n45186), .Z(n45188) );
  NOR U58116 ( .A(n45188), .B(n45187), .Z(n50076) );
  NOR U58117 ( .A(n50080), .B(n50076), .Z(n45189) );
  IV U58118 ( .A(n45189), .Z(n45190) );
  NOR U58119 ( .A(n50084), .B(n45190), .Z(n45191) );
  IV U58120 ( .A(n45191), .Z(n46617) );
  IV U58121 ( .A(n45192), .Z(n45193) );
  NOR U58122 ( .A(n45194), .B(n45193), .Z(n50074) );
  IV U58123 ( .A(n45195), .Z(n45198) );
  IV U58124 ( .A(n45196), .Z(n45197) );
  NOR U58125 ( .A(n45198), .B(n45197), .Z(n45199) );
  IV U58126 ( .A(n45199), .Z(n48691) );
  NOR U58127 ( .A(n45201), .B(n45200), .Z(n50065) );
  IV U58128 ( .A(n45202), .Z(n45203) );
  NOR U58129 ( .A(n45204), .B(n45203), .Z(n50062) );
  IV U58130 ( .A(n45205), .Z(n45206) );
  NOR U58131 ( .A(n45207), .B(n45206), .Z(n48695) );
  NOR U58132 ( .A(n50062), .B(n48695), .Z(n45208) );
  IV U58133 ( .A(n45208), .Z(n46609) );
  NOR U58134 ( .A(n45210), .B(n45209), .Z(n45211) );
  IV U58135 ( .A(n45211), .Z(n48706) );
  NOR U58136 ( .A(n45213), .B(n45212), .Z(n50053) );
  IV U58137 ( .A(n45214), .Z(n50046) );
  NOR U58138 ( .A(n50046), .B(n45215), .Z(n45218) );
  IV U58139 ( .A(n45216), .Z(n45217) );
  NOR U58140 ( .A(n45217), .B(n48714), .Z(n50036) );
  NOR U58141 ( .A(n45218), .B(n50036), .Z(n45219) );
  IV U58142 ( .A(n45219), .Z(n46599) );
  IV U58143 ( .A(n45220), .Z(n45221) );
  NOR U58144 ( .A(n45222), .B(n45221), .Z(n49994) );
  IV U58145 ( .A(n45223), .Z(n45224) );
  NOR U58146 ( .A(n45225), .B(n45224), .Z(n48721) );
  NOR U58147 ( .A(n45227), .B(n45226), .Z(n48734) );
  IV U58148 ( .A(n45228), .Z(n45229) );
  NOR U58149 ( .A(n46548), .B(n45229), .Z(n48738) );
  NOR U58150 ( .A(n48734), .B(n48738), .Z(n46552) );
  NOR U58151 ( .A(n48748), .B(n48746), .Z(n45233) );
  IV U58152 ( .A(n45230), .Z(n45232) );
  NOR U58153 ( .A(n45232), .B(n45231), .Z(n48736) );
  NOR U58154 ( .A(n45233), .B(n48736), .Z(n45234) );
  IV U58155 ( .A(n45234), .Z(n46546) );
  NOR U58156 ( .A(n45235), .B(n48758), .Z(n45239) );
  IV U58157 ( .A(n45236), .Z(n48751) );
  NOR U58158 ( .A(n45237), .B(n48751), .Z(n45238) );
  NOR U58159 ( .A(n45239), .B(n45238), .Z(n46545) );
  IV U58160 ( .A(n45240), .Z(n45242) );
  NOR U58161 ( .A(n45242), .B(n45241), .Z(n49975) );
  IV U58162 ( .A(n45243), .Z(n45244) );
  NOR U58163 ( .A(n45245), .B(n45244), .Z(n49980) );
  NOR U58164 ( .A(n49975), .B(n49980), .Z(n46544) );
  IV U58165 ( .A(n45246), .Z(n45248) );
  NOR U58166 ( .A(n45248), .B(n45247), .Z(n48765) );
  IV U58167 ( .A(n45249), .Z(n45251) );
  NOR U58168 ( .A(n45251), .B(n45250), .Z(n52534) );
  IV U58169 ( .A(n45252), .Z(n45254) );
  NOR U58170 ( .A(n45254), .B(n45253), .Z(n53877) );
  NOR U58171 ( .A(n52534), .B(n53877), .Z(n48775) );
  IV U58172 ( .A(n45255), .Z(n45256) );
  NOR U58173 ( .A(n45257), .B(n45256), .Z(n49960) );
  IV U58174 ( .A(n45258), .Z(n45259) );
  NOR U58175 ( .A(n46530), .B(n45259), .Z(n49954) );
  IV U58176 ( .A(n45260), .Z(n45261) );
  NOR U58177 ( .A(n45262), .B(n45261), .Z(n46520) );
  IV U58178 ( .A(n46520), .Z(n46515) );
  IV U58179 ( .A(n45263), .Z(n45264) );
  NOR U58180 ( .A(n45265), .B(n45264), .Z(n49934) );
  IV U58181 ( .A(n45266), .Z(n45267) );
  NOR U58182 ( .A(n46512), .B(n45267), .Z(n49930) );
  IV U58183 ( .A(n45268), .Z(n45269) );
  NOR U58184 ( .A(n45270), .B(n45269), .Z(n48780) );
  IV U58185 ( .A(n45271), .Z(n45273) );
  NOR U58186 ( .A(n45273), .B(n45272), .Z(n48778) );
  NOR U58187 ( .A(n48780), .B(n48778), .Z(n46510) );
  IV U58188 ( .A(n45274), .Z(n45275) );
  NOR U58189 ( .A(n45276), .B(n45275), .Z(n45277) );
  IV U58190 ( .A(n45277), .Z(n48783) );
  IV U58191 ( .A(n45278), .Z(n46503) );
  IV U58192 ( .A(n45279), .Z(n45280) );
  NOR U58193 ( .A(n46503), .B(n45280), .Z(n45281) );
  IV U58194 ( .A(n45281), .Z(n48791) );
  IV U58195 ( .A(n45282), .Z(n45283) );
  NOR U58196 ( .A(n45283), .B(n46491), .Z(n46497) );
  IV U58197 ( .A(n45284), .Z(n45285) );
  NOR U58198 ( .A(n45286), .B(n45285), .Z(n48821) );
  NOR U58199 ( .A(n45287), .B(n48799), .Z(n45288) );
  NOR U58200 ( .A(n48821), .B(n45288), .Z(n46488) );
  NOR U58201 ( .A(n45290), .B(n45289), .Z(n49901) );
  IV U58202 ( .A(n48808), .Z(n48825) );
  NOR U58203 ( .A(n48806), .B(n48825), .Z(n48809) );
  NOR U58204 ( .A(n49901), .B(n48809), .Z(n46487) );
  IV U58205 ( .A(n45291), .Z(n45292) );
  NOR U58206 ( .A(n45292), .B(n46485), .Z(n49898) );
  IV U58207 ( .A(n45293), .Z(n45294) );
  NOR U58208 ( .A(n45294), .B(n46485), .Z(n49887) );
  IV U58209 ( .A(n45295), .Z(n45296) );
  NOR U58210 ( .A(n45296), .B(n46474), .Z(n52605) );
  IV U58211 ( .A(n45297), .Z(n45299) );
  IV U58212 ( .A(n45298), .Z(n46480) );
  NOR U58213 ( .A(n45299), .B(n46480), .Z(n53790) );
  NOR U58214 ( .A(n52605), .B(n53790), .Z(n49878) );
  IV U58215 ( .A(n45300), .Z(n45301) );
  NOR U58216 ( .A(n45307), .B(n45301), .Z(n53776) );
  IV U58217 ( .A(n45302), .Z(n45304) );
  NOR U58218 ( .A(n45304), .B(n45303), .Z(n48828) );
  NOR U58219 ( .A(n53776), .B(n48828), .Z(n46468) );
  IV U58220 ( .A(n45305), .Z(n45306) );
  NOR U58221 ( .A(n45307), .B(n45306), .Z(n48830) );
  IV U58222 ( .A(n48830), .Z(n53784) );
  IV U58223 ( .A(n45308), .Z(n45309) );
  NOR U58224 ( .A(n45310), .B(n45309), .Z(n53773) );
  IV U58225 ( .A(n45311), .Z(n45312) );
  NOR U58226 ( .A(n45313), .B(n45312), .Z(n52618) );
  NOR U58227 ( .A(n53773), .B(n52618), .Z(n48835) );
  IV U58228 ( .A(n45314), .Z(n45315) );
  NOR U58229 ( .A(n45316), .B(n45315), .Z(n48841) );
  IV U58230 ( .A(n45317), .Z(n45320) );
  IV U58231 ( .A(n45318), .Z(n45319) );
  NOR U58232 ( .A(n45320), .B(n45319), .Z(n48838) );
  IV U58233 ( .A(n45321), .Z(n45322) );
  NOR U58234 ( .A(n45322), .B(n45325), .Z(n48844) );
  IV U58235 ( .A(n45323), .Z(n45324) );
  NOR U58236 ( .A(n48854), .B(n45324), .Z(n45327) );
  NOR U58237 ( .A(n45326), .B(n45325), .Z(n48847) );
  NOR U58238 ( .A(n45327), .B(n48847), .Z(n45328) );
  IV U58239 ( .A(n45328), .Z(n46458) );
  NOR U58240 ( .A(n45329), .B(n45331), .Z(n49853) );
  IV U58241 ( .A(n45330), .Z(n45332) );
  NOR U58242 ( .A(n45332), .B(n45331), .Z(n48871) );
  NOR U58243 ( .A(n49853), .B(n48871), .Z(n46444) );
  IV U58244 ( .A(n45333), .Z(n45334) );
  NOR U58245 ( .A(n45335), .B(n45334), .Z(n45336) );
  IV U58246 ( .A(n45336), .Z(n49852) );
  IV U58247 ( .A(n45337), .Z(n45338) );
  NOR U58248 ( .A(n45339), .B(n45338), .Z(n48874) );
  IV U58249 ( .A(n45340), .Z(n45341) );
  NOR U58250 ( .A(n45342), .B(n45341), .Z(n48869) );
  NOR U58251 ( .A(n48874), .B(n48869), .Z(n45343) );
  IV U58252 ( .A(n45343), .Z(n46442) );
  IV U58253 ( .A(n45344), .Z(n45345) );
  NOR U58254 ( .A(n45345), .B(n46440), .Z(n49846) );
  IV U58255 ( .A(n45346), .Z(n45348) );
  NOR U58256 ( .A(n45348), .B(n45347), .Z(n48883) );
  IV U58257 ( .A(n45349), .Z(n45354) );
  IV U58258 ( .A(n45350), .Z(n45351) );
  NOR U58259 ( .A(n45354), .B(n45351), .Z(n49839) );
  NOR U58260 ( .A(n48883), .B(n49839), .Z(n46434) );
  IV U58261 ( .A(n45352), .Z(n45353) );
  NOR U58262 ( .A(n45354), .B(n45353), .Z(n49836) );
  IV U58263 ( .A(n45355), .Z(n45356) );
  NOR U58264 ( .A(n45357), .B(n45356), .Z(n48889) );
  IV U58265 ( .A(n45358), .Z(n45360) );
  IV U58266 ( .A(n45359), .Z(n45364) );
  NOR U58267 ( .A(n45360), .B(n45364), .Z(n48892) );
  NOR U58268 ( .A(n45362), .B(n45361), .Z(n49819) );
  IV U58269 ( .A(n45363), .Z(n45365) );
  NOR U58270 ( .A(n45365), .B(n45364), .Z(n49821) );
  NOR U58271 ( .A(n49819), .B(n49821), .Z(n46409) );
  IV U58272 ( .A(n45366), .Z(n45368) );
  NOR U58273 ( .A(n45368), .B(n45367), .Z(n49814) );
  IV U58274 ( .A(n45369), .Z(n45371) );
  NOR U58275 ( .A(n45371), .B(n45370), .Z(n49809) );
  IV U58276 ( .A(n45372), .Z(n45373) );
  NOR U58277 ( .A(n45374), .B(n45373), .Z(n49804) );
  NOR U58278 ( .A(n49809), .B(n49804), .Z(n45375) );
  IV U58279 ( .A(n45375), .Z(n45376) );
  NOR U58280 ( .A(n49814), .B(n45376), .Z(n46408) );
  IV U58281 ( .A(n45377), .Z(n45378) );
  NOR U58282 ( .A(n45379), .B(n45378), .Z(n49806) );
  NOR U58283 ( .A(n45381), .B(n45380), .Z(n45382) );
  IV U58284 ( .A(n45382), .Z(n48897) );
  NOR U58285 ( .A(n45383), .B(n48897), .Z(n49798) );
  IV U58286 ( .A(n45384), .Z(n45385) );
  NOR U58287 ( .A(n46400), .B(n45385), .Z(n45386) );
  IV U58288 ( .A(n45386), .Z(n46392) );
  IV U58289 ( .A(n45387), .Z(n45388) );
  NOR U58290 ( .A(n45388), .B(n45390), .Z(n49771) );
  IV U58291 ( .A(n45389), .Z(n45391) );
  NOR U58292 ( .A(n45391), .B(n45390), .Z(n49768) );
  IV U58293 ( .A(n45392), .Z(n45393) );
  NOR U58294 ( .A(n46386), .B(n45393), .Z(n48915) );
  IV U58295 ( .A(n45394), .Z(n45396) );
  IV U58296 ( .A(n45395), .Z(n45398) );
  NOR U58297 ( .A(n45396), .B(n45398), .Z(n48921) );
  NOR U58298 ( .A(n48915), .B(n48921), .Z(n46380) );
  IV U58299 ( .A(n45397), .Z(n45399) );
  NOR U58300 ( .A(n45399), .B(n45398), .Z(n48927) );
  IV U58301 ( .A(n45400), .Z(n45401) );
  NOR U58302 ( .A(n45401), .B(n46378), .Z(n48924) );
  IV U58303 ( .A(n45402), .Z(n48936) );
  IV U58304 ( .A(n45403), .Z(n45406) );
  IV U58305 ( .A(n45404), .Z(n45405) );
  NOR U58306 ( .A(n45406), .B(n45405), .Z(n45407) );
  IV U58307 ( .A(n45407), .Z(n48934) );
  IV U58308 ( .A(n45408), .Z(n45409) );
  NOR U58309 ( .A(n45410), .B(n45409), .Z(n45411) );
  IV U58310 ( .A(n45411), .Z(n45412) );
  NOR U58311 ( .A(n45413), .B(n45412), .Z(n45414) );
  IV U58312 ( .A(n45414), .Z(n48937) );
  IV U58313 ( .A(n45415), .Z(n45417) );
  NOR U58314 ( .A(n45417), .B(n45416), .Z(n48945) );
  IV U58315 ( .A(n45418), .Z(n45419) );
  NOR U58316 ( .A(n45419), .B(n46355), .Z(n48940) );
  NOR U58317 ( .A(n48945), .B(n48940), .Z(n46358) );
  IV U58318 ( .A(n45420), .Z(n45422) );
  NOR U58319 ( .A(n45422), .B(n45421), .Z(n49755) );
  IV U58320 ( .A(n45423), .Z(n45430) );
  NOR U58321 ( .A(n45425), .B(n45424), .Z(n45426) );
  IV U58322 ( .A(n45426), .Z(n45427) );
  NOR U58323 ( .A(n45428), .B(n45427), .Z(n45429) );
  IV U58324 ( .A(n45429), .Z(n48953) );
  NOR U58325 ( .A(n45430), .B(n48953), .Z(n48950) );
  NOR U58326 ( .A(n49755), .B(n48950), .Z(n46350) );
  IV U58327 ( .A(n45431), .Z(n45432) );
  NOR U58328 ( .A(n45432), .B(n48953), .Z(n46349) );
  IV U58329 ( .A(n45433), .Z(n45434) );
  NOR U58330 ( .A(n45435), .B(n45434), .Z(n48973) );
  IV U58331 ( .A(n45436), .Z(n45437) );
  NOR U58332 ( .A(n46323), .B(n45437), .Z(n49728) );
  NOR U58333 ( .A(n48973), .B(n49728), .Z(n46321) );
  IV U58334 ( .A(n45438), .Z(n45441) );
  IV U58335 ( .A(n45439), .Z(n45440) );
  NOR U58336 ( .A(n45441), .B(n45440), .Z(n48975) );
  IV U58337 ( .A(n45442), .Z(n45443) );
  NOR U58338 ( .A(n45443), .B(n46319), .Z(n49718) );
  IV U58339 ( .A(n45444), .Z(n45447) );
  NOR U58340 ( .A(n46301), .B(n45445), .Z(n45446) );
  IV U58341 ( .A(n45446), .Z(n46303) );
  NOR U58342 ( .A(n45447), .B(n46303), .Z(n48982) );
  IV U58343 ( .A(n45448), .Z(n45449) );
  NOR U58344 ( .A(n45450), .B(n45449), .Z(n48996) );
  IV U58345 ( .A(n45451), .Z(n45453) );
  NOR U58346 ( .A(n45453), .B(n45452), .Z(n48993) );
  NOR U58347 ( .A(n48996), .B(n48993), .Z(n46275) );
  IV U58348 ( .A(n45454), .Z(n45460) );
  NOR U58349 ( .A(n45466), .B(n45455), .Z(n45456) );
  IV U58350 ( .A(n45456), .Z(n45457) );
  NOR U58351 ( .A(n45458), .B(n45457), .Z(n45459) );
  IV U58352 ( .A(n45459), .Z(n45462) );
  NOR U58353 ( .A(n45460), .B(n45462), .Z(n49691) );
  IV U58354 ( .A(n45461), .Z(n45463) );
  NOR U58355 ( .A(n45463), .B(n45462), .Z(n49693) );
  IV U58356 ( .A(n45464), .Z(n45468) );
  NOR U58357 ( .A(n45466), .B(n45465), .Z(n45467) );
  IV U58358 ( .A(n45467), .Z(n45471) );
  NOR U58359 ( .A(n45468), .B(n45471), .Z(n49695) );
  XOR U58360 ( .A(n49693), .B(n49695), .Z(n45469) );
  NOR U58361 ( .A(n49691), .B(n45469), .Z(n46274) );
  IV U58362 ( .A(n45470), .Z(n45472) );
  NOR U58363 ( .A(n45472), .B(n45471), .Z(n49001) );
  IV U58364 ( .A(n45473), .Z(n45475) );
  IV U58365 ( .A(n45474), .Z(n45478) );
  NOR U58366 ( .A(n45475), .B(n45478), .Z(n49003) );
  NOR U58367 ( .A(n49001), .B(n49003), .Z(n46273) );
  NOR U58368 ( .A(n45476), .B(n49007), .Z(n45480) );
  IV U58369 ( .A(n45477), .Z(n45479) );
  NOR U58370 ( .A(n45479), .B(n45478), .Z(n49688) );
  NOR U58371 ( .A(n45480), .B(n49688), .Z(n46272) );
  IV U58372 ( .A(n45481), .Z(n45485) );
  NOR U58373 ( .A(n45483), .B(n45482), .Z(n45484) );
  IV U58374 ( .A(n45484), .Z(n45487) );
  NOR U58375 ( .A(n45485), .B(n45487), .Z(n49675) );
  IV U58376 ( .A(n45486), .Z(n45488) );
  NOR U58377 ( .A(n45488), .B(n45487), .Z(n49672) );
  IV U58378 ( .A(n45489), .Z(n45490) );
  NOR U58379 ( .A(n45491), .B(n45490), .Z(n49013) );
  IV U58380 ( .A(n45492), .Z(n45493) );
  NOR U58381 ( .A(n45494), .B(n45493), .Z(n49011) );
  NOR U58382 ( .A(n49013), .B(n49011), .Z(n46271) );
  IV U58383 ( .A(n45495), .Z(n45496) );
  NOR U58384 ( .A(n45497), .B(n45496), .Z(n49669) );
  IV U58385 ( .A(n45498), .Z(n45500) );
  NOR U58386 ( .A(n45500), .B(n45499), .Z(n49016) );
  NOR U58387 ( .A(n49669), .B(n49016), .Z(n46270) );
  IV U58388 ( .A(n45501), .Z(n45502) );
  NOR U58389 ( .A(n46267), .B(n45502), .Z(n49661) );
  IV U58390 ( .A(n45503), .Z(n45508) );
  IV U58391 ( .A(n45504), .Z(n45505) );
  NOR U58392 ( .A(n45508), .B(n45505), .Z(n46264) );
  IV U58393 ( .A(n46264), .Z(n46262) );
  NOR U58394 ( .A(n45506), .B(n49020), .Z(n45510) );
  IV U58395 ( .A(n45507), .Z(n45509) );
  NOR U58396 ( .A(n45509), .B(n45508), .Z(n49657) );
  NOR U58397 ( .A(n45510), .B(n49657), .Z(n46260) );
  IV U58398 ( .A(n45511), .Z(n45512) );
  NOR U58399 ( .A(n45513), .B(n45512), .Z(n49026) );
  NOR U58400 ( .A(n49031), .B(n49026), .Z(n45514) );
  IV U58401 ( .A(n45514), .Z(n46259) );
  IV U58402 ( .A(n45515), .Z(n45516) );
  NOR U58403 ( .A(n45516), .B(n45518), .Z(n49028) );
  IV U58404 ( .A(n45517), .Z(n45519) );
  NOR U58405 ( .A(n45519), .B(n45518), .Z(n49034) );
  IV U58406 ( .A(n45520), .Z(n45521) );
  NOR U58407 ( .A(n45522), .B(n45521), .Z(n52813) );
  IV U58408 ( .A(n45523), .Z(n45525) );
  NOR U58409 ( .A(n45525), .B(n45524), .Z(n52809) );
  NOR U58410 ( .A(n52813), .B(n52809), .Z(n49650) );
  IV U58411 ( .A(n45526), .Z(n45527) );
  NOR U58412 ( .A(n45528), .B(n45527), .Z(n49645) );
  IV U58413 ( .A(n45529), .Z(n45530) );
  NOR U58414 ( .A(n45530), .B(n45532), .Z(n49642) );
  NOR U58415 ( .A(n49645), .B(n49642), .Z(n46258) );
  IV U58416 ( .A(n45531), .Z(n45533) );
  NOR U58417 ( .A(n45533), .B(n45532), .Z(n49639) );
  IV U58418 ( .A(n45534), .Z(n46254) );
  IV U58419 ( .A(n45535), .Z(n45536) );
  NOR U58420 ( .A(n46254), .B(n45536), .Z(n49037) );
  IV U58421 ( .A(n45537), .Z(n45538) );
  NOR U58422 ( .A(n46256), .B(n45538), .Z(n49626) );
  IV U58423 ( .A(n45539), .Z(n45540) );
  NOR U58424 ( .A(n45541), .B(n45540), .Z(n45542) );
  IV U58425 ( .A(n45542), .Z(n46248) );
  IV U58426 ( .A(n45543), .Z(n45546) );
  IV U58427 ( .A(n45544), .Z(n45545) );
  NOR U58428 ( .A(n45546), .B(n45545), .Z(n49040) );
  IV U58429 ( .A(n45547), .Z(n45550) );
  IV U58430 ( .A(n45548), .Z(n45549) );
  NOR U58431 ( .A(n45550), .B(n45549), .Z(n49049) );
  IV U58432 ( .A(n45551), .Z(n45557) );
  IV U58433 ( .A(n45552), .Z(n46232) );
  IV U58434 ( .A(n45553), .Z(n45554) );
  NOR U58435 ( .A(n46232), .B(n45554), .Z(n45555) );
  IV U58436 ( .A(n45555), .Z(n45556) );
  NOR U58437 ( .A(n45557), .B(n45556), .Z(n45558) );
  IV U58438 ( .A(n45558), .Z(n49060) );
  IV U58439 ( .A(n45559), .Z(n45560) );
  NOR U58440 ( .A(n46220), .B(n45560), .Z(n46215) );
  IV U58441 ( .A(n45561), .Z(n45564) );
  NOR U58442 ( .A(n45562), .B(n46201), .Z(n45563) );
  IV U58443 ( .A(n45563), .Z(n46195) );
  NOR U58444 ( .A(n45564), .B(n46195), .Z(n49066) );
  IV U58445 ( .A(n45565), .Z(n45567) );
  NOR U58446 ( .A(n45567), .B(n45566), .Z(n49600) );
  IV U58447 ( .A(n45568), .Z(n45569) );
  NOR U58448 ( .A(n45570), .B(n45569), .Z(n49069) );
  NOR U58449 ( .A(n49600), .B(n49069), .Z(n45571) );
  IV U58450 ( .A(n45571), .Z(n46193) );
  IV U58451 ( .A(n45572), .Z(n45573) );
  NOR U58452 ( .A(n45573), .B(n46191), .Z(n49594) );
  IV U58453 ( .A(n45574), .Z(n45575) );
  NOR U58454 ( .A(n45576), .B(n45575), .Z(n45577) );
  IV U58455 ( .A(n45577), .Z(n49083) );
  IV U58456 ( .A(n45578), .Z(n45580) );
  IV U58457 ( .A(n45579), .Z(n45584) );
  NOR U58458 ( .A(n45580), .B(n45584), .Z(n49079) );
  NOR U58459 ( .A(n45582), .B(n45581), .Z(n49088) );
  IV U58460 ( .A(n45583), .Z(n45585) );
  NOR U58461 ( .A(n45585), .B(n45584), .Z(n49085) );
  NOR U58462 ( .A(n49088), .B(n49085), .Z(n45586) );
  IV U58463 ( .A(n45586), .Z(n46185) );
  IV U58464 ( .A(n45587), .Z(n45588) );
  NOR U58465 ( .A(n45589), .B(n45588), .Z(n49093) );
  IV U58466 ( .A(n45590), .Z(n45591) );
  NOR U58467 ( .A(n45591), .B(n45596), .Z(n49090) );
  IV U58468 ( .A(n45592), .Z(n45593) );
  NOR U58469 ( .A(n45594), .B(n45593), .Z(n49581) );
  IV U58470 ( .A(n45595), .Z(n45597) );
  NOR U58471 ( .A(n45597), .B(n45596), .Z(n49097) );
  NOR U58472 ( .A(n49581), .B(n49097), .Z(n46184) );
  IV U58473 ( .A(n45598), .Z(n45599) );
  NOR U58474 ( .A(n45600), .B(n45599), .Z(n45601) );
  IV U58475 ( .A(n45601), .Z(n49560) );
  IV U58476 ( .A(n45602), .Z(n45603) );
  NOR U58477 ( .A(n45604), .B(n45603), .Z(n49099) );
  IV U58478 ( .A(n45605), .Z(n45607) );
  IV U58479 ( .A(n45606), .Z(n45614) );
  NOR U58480 ( .A(n45607), .B(n45614), .Z(n49551) );
  NOR U58481 ( .A(n49099), .B(n49551), .Z(n45608) );
  IV U58482 ( .A(n45608), .Z(n46152) );
  IV U58483 ( .A(n45609), .Z(n45612) );
  IV U58484 ( .A(n45610), .Z(n45611) );
  NOR U58485 ( .A(n45612), .B(n45611), .Z(n49550) );
  IV U58486 ( .A(n45613), .Z(n45615) );
  NOR U58487 ( .A(n45615), .B(n45614), .Z(n49543) );
  NOR U58488 ( .A(n49550), .B(n49543), .Z(n46151) );
  IV U58489 ( .A(n45616), .Z(n45617) );
  NOR U58490 ( .A(n45618), .B(n45617), .Z(n49102) );
  NOR U58491 ( .A(n49102), .B(n49539), .Z(n46150) );
  IV U58492 ( .A(n45621), .Z(n45619) );
  NOR U58493 ( .A(n45620), .B(n45619), .Z(n53450) );
  NOR U58494 ( .A(n45622), .B(n45621), .Z(n45625) );
  IV U58495 ( .A(n45623), .Z(n45624) );
  NOR U58496 ( .A(n45625), .B(n45624), .Z(n53462) );
  NOR U58497 ( .A(n53450), .B(n53462), .Z(n49105) );
  IV U58498 ( .A(n45626), .Z(n45627) );
  NOR U58499 ( .A(n45628), .B(n45627), .Z(n46130) );
  IV U58500 ( .A(n46130), .Z(n46119) );
  IV U58501 ( .A(n45629), .Z(n45634) );
  IV U58502 ( .A(n45630), .Z(n46127) );
  NOR U58503 ( .A(n45631), .B(n46127), .Z(n45632) );
  IV U58504 ( .A(n45632), .Z(n45633) );
  NOR U58505 ( .A(n45634), .B(n45633), .Z(n49118) );
  IV U58506 ( .A(n45635), .Z(n45636) );
  NOR U58507 ( .A(n45637), .B(n45636), .Z(n46112) );
  IV U58508 ( .A(n45638), .Z(n45639) );
  NOR U58509 ( .A(n49142), .B(n45639), .Z(n45640) );
  IV U58510 ( .A(n45640), .Z(n49147) );
  IV U58511 ( .A(n45641), .Z(n45642) );
  NOR U58512 ( .A(n46081), .B(n45642), .Z(n52957) );
  IV U58513 ( .A(n45643), .Z(n46095) );
  IV U58514 ( .A(n45644), .Z(n45645) );
  NOR U58515 ( .A(n46095), .B(n45645), .Z(n52953) );
  NOR U58516 ( .A(n52957), .B(n52953), .Z(n49149) );
  IV U58517 ( .A(n45646), .Z(n49510) );
  NOR U58518 ( .A(n49510), .B(n45647), .Z(n46076) );
  IV U58519 ( .A(n45648), .Z(n45649) );
  NOR U58520 ( .A(n45649), .B(n45653), .Z(n53389) );
  IV U58521 ( .A(n45650), .Z(n45651) );
  NOR U58522 ( .A(n45651), .B(n46074), .Z(n53399) );
  NOR U58523 ( .A(n53389), .B(n53399), .Z(n49502) );
  IV U58524 ( .A(n45652), .Z(n45654) );
  NOR U58525 ( .A(n45654), .B(n45653), .Z(n49499) );
  IV U58526 ( .A(n45655), .Z(n45661) );
  IV U58527 ( .A(n45656), .Z(n45657) );
  NOR U58528 ( .A(n45661), .B(n45657), .Z(n45658) );
  IV U58529 ( .A(n45658), .Z(n49159) );
  IV U58530 ( .A(n45659), .Z(n45660) );
  NOR U58531 ( .A(n45661), .B(n45660), .Z(n49168) );
  IV U58532 ( .A(n45662), .Z(n45663) );
  NOR U58533 ( .A(n45663), .B(n46062), .Z(n49494) );
  NOR U58534 ( .A(n49168), .B(n49494), .Z(n45664) );
  IV U58535 ( .A(n45664), .Z(n46065) );
  IV U58536 ( .A(n45665), .Z(n45667) );
  IV U58537 ( .A(n45666), .Z(n46045) );
  NOR U58538 ( .A(n45667), .B(n46045), .Z(n53374) );
  IV U58539 ( .A(n45668), .Z(n45670) );
  NOR U58540 ( .A(n45670), .B(n45669), .Z(n53383) );
  NOR U58541 ( .A(n53374), .B(n53383), .Z(n49179) );
  IV U58542 ( .A(n45671), .Z(n45672) );
  NOR U58543 ( .A(n45673), .B(n45672), .Z(n45674) );
  IV U58544 ( .A(n45674), .Z(n46031) );
  IV U58545 ( .A(n45675), .Z(n45676) );
  NOR U58546 ( .A(n45676), .B(n46027), .Z(n49485) );
  IV U58547 ( .A(n45677), .Z(n45678) );
  NOR U58548 ( .A(n45678), .B(n46027), .Z(n49198) );
  IV U58549 ( .A(n45679), .Z(n45684) );
  IV U58550 ( .A(n45680), .Z(n45681) );
  NOR U58551 ( .A(n45684), .B(n45681), .Z(n49195) );
  IV U58552 ( .A(n45682), .Z(n45683) );
  NOR U58553 ( .A(n45684), .B(n45683), .Z(n49206) );
  IV U58554 ( .A(n45685), .Z(n45687) );
  NOR U58555 ( .A(n45687), .B(n45686), .Z(n45688) );
  IV U58556 ( .A(n45688), .Z(n46018) );
  IV U58557 ( .A(n45689), .Z(n45690) );
  NOR U58558 ( .A(n46016), .B(n45690), .Z(n49481) );
  IV U58559 ( .A(n45691), .Z(n45692) );
  NOR U58560 ( .A(n46004), .B(n45692), .Z(n45693) );
  IV U58561 ( .A(n45693), .Z(n49225) );
  IV U58562 ( .A(n45694), .Z(n45696) );
  IV U58563 ( .A(n45695), .Z(n45702) );
  NOR U58564 ( .A(n45696), .B(n45702), .Z(n49222) );
  IV U58565 ( .A(n45697), .Z(n45700) );
  IV U58566 ( .A(n45698), .Z(n45699) );
  NOR U58567 ( .A(n45700), .B(n45699), .Z(n49235) );
  IV U58568 ( .A(n45701), .Z(n45703) );
  NOR U58569 ( .A(n45703), .B(n45702), .Z(n49227) );
  NOR U58570 ( .A(n49235), .B(n49227), .Z(n45704) );
  IV U58571 ( .A(n45704), .Z(n46001) );
  IV U58572 ( .A(n45705), .Z(n45706) );
  NOR U58573 ( .A(n45706), .B(n45714), .Z(n49240) );
  IV U58574 ( .A(n45707), .Z(n45709) );
  NOR U58575 ( .A(n45709), .B(n45708), .Z(n49238) );
  NOR U58576 ( .A(n49240), .B(n49238), .Z(n46000) );
  IV U58577 ( .A(n45710), .Z(n45712) );
  NOR U58578 ( .A(n45712), .B(n45711), .Z(n49467) );
  IV U58579 ( .A(n45713), .Z(n45715) );
  NOR U58580 ( .A(n45715), .B(n45714), .Z(n49471) );
  NOR U58581 ( .A(n49467), .B(n49471), .Z(n45999) );
  IV U58582 ( .A(n45716), .Z(n45718) );
  NOR U58583 ( .A(n45718), .B(n45717), .Z(n45997) );
  IV U58584 ( .A(n45997), .Z(n45985) );
  IV U58585 ( .A(n45719), .Z(n45721) );
  NOR U58586 ( .A(n45721), .B(n45720), .Z(n49462) );
  IV U58587 ( .A(n45722), .Z(n45723) );
  NOR U58588 ( .A(n45975), .B(n45723), .Z(n49459) );
  IV U58589 ( .A(n45724), .Z(n45725) );
  NOR U58590 ( .A(n45725), .B(n45727), .Z(n49446) );
  IV U58591 ( .A(n45726), .Z(n45728) );
  NOR U58592 ( .A(n45728), .B(n45727), .Z(n49249) );
  IV U58593 ( .A(n45729), .Z(n45730) );
  NOR U58594 ( .A(n45730), .B(n45733), .Z(n49443) );
  NOR U58595 ( .A(n49249), .B(n49443), .Z(n45731) );
  IV U58596 ( .A(n45731), .Z(n45963) );
  IV U58597 ( .A(n45732), .Z(n45734) );
  NOR U58598 ( .A(n45734), .B(n45733), .Z(n45735) );
  IV U58599 ( .A(n45735), .Z(n49248) );
  IV U58600 ( .A(n45736), .Z(n45738) );
  NOR U58601 ( .A(n45738), .B(n45737), .Z(n49440) );
  IV U58602 ( .A(n45739), .Z(n49256) );
  NOR U58603 ( .A(n45740), .B(n49256), .Z(n45743) );
  IV U58604 ( .A(n45741), .Z(n45742) );
  NOR U58605 ( .A(n45746), .B(n45742), .Z(n49265) );
  NOR U58606 ( .A(n45743), .B(n49265), .Z(n45954) );
  IV U58607 ( .A(n45744), .Z(n45745) );
  NOR U58608 ( .A(n45746), .B(n45745), .Z(n49262) );
  IV U58609 ( .A(n45747), .Z(n45748) );
  NOR U58610 ( .A(n45748), .B(n45931), .Z(n45749) );
  IV U58611 ( .A(n45749), .Z(n49285) );
  IV U58612 ( .A(n45750), .Z(n45752) );
  NOR U58613 ( .A(n45752), .B(n45751), .Z(n45927) );
  IV U58614 ( .A(n45927), .Z(n45920) );
  IV U58615 ( .A(n45753), .Z(n45754) );
  NOR U58616 ( .A(n45754), .B(n45901), .Z(n49308) );
  IV U58617 ( .A(n45755), .Z(n45756) );
  NOR U58618 ( .A(n45757), .B(n45756), .Z(n53132) );
  IV U58619 ( .A(n45758), .Z(n45759) );
  NOR U58620 ( .A(n45760), .B(n45759), .Z(n53255) );
  NOR U58621 ( .A(n53132), .B(n53255), .Z(n49307) );
  IV U58622 ( .A(n45761), .Z(n45763) );
  NOR U58623 ( .A(n45763), .B(n45762), .Z(n45764) );
  IV U58624 ( .A(n45764), .Z(n45895) );
  IV U58625 ( .A(n45765), .Z(n49405) );
  IV U58626 ( .A(n45766), .Z(n45768) );
  NOR U58627 ( .A(n45768), .B(n45767), .Z(n49321) );
  IV U58628 ( .A(n45769), .Z(n45772) );
  NOR U58629 ( .A(n45770), .B(n45875), .Z(n45771) );
  IV U58630 ( .A(n45771), .Z(n45878) );
  NOR U58631 ( .A(n45772), .B(n45878), .Z(n49324) );
  NOR U58632 ( .A(n49321), .B(n49324), .Z(n45880) );
  IV U58633 ( .A(n45773), .Z(n45779) );
  IV U58634 ( .A(n45774), .Z(n45775) );
  NOR U58635 ( .A(n45779), .B(n45775), .Z(n49327) );
  NOR U58636 ( .A(n45777), .B(n45776), .Z(n49338) );
  IV U58637 ( .A(n45778), .Z(n45780) );
  NOR U58638 ( .A(n45780), .B(n45779), .Z(n49333) );
  NOR U58639 ( .A(n49338), .B(n49333), .Z(n45873) );
  IV U58640 ( .A(n45781), .Z(n45782) );
  NOR U58641 ( .A(n45783), .B(n45782), .Z(n45855) );
  IV U58642 ( .A(n45855), .Z(n45849) );
  IV U58643 ( .A(n45784), .Z(n45841) );
  IV U58644 ( .A(n45785), .Z(n45786) );
  NOR U58645 ( .A(n45841), .B(n45786), .Z(n49349) );
  IV U58646 ( .A(n45787), .Z(n45790) );
  NOR U58647 ( .A(n45788), .B(n45797), .Z(n45789) );
  IV U58648 ( .A(n45789), .Z(n45837) );
  NOR U58649 ( .A(n45790), .B(n45837), .Z(n45791) );
  IV U58650 ( .A(n45791), .Z(n49389) );
  IV U58651 ( .A(n45792), .Z(n45793) );
  NOR U58652 ( .A(n45794), .B(n45793), .Z(n49370) );
  IV U58653 ( .A(n45795), .Z(n45796) );
  NOR U58654 ( .A(n45797), .B(n45796), .Z(n49385) );
  NOR U58655 ( .A(n49370), .B(n49385), .Z(n45798) );
  IV U58656 ( .A(n45798), .Z(n45835) );
  IV U58657 ( .A(n45799), .Z(n45806) );
  IV U58658 ( .A(n45800), .Z(n45801) );
  NOR U58659 ( .A(n45806), .B(n45801), .Z(n49372) );
  NOR U58660 ( .A(n45803), .B(n45802), .Z(n45808) );
  IV U58661 ( .A(n45804), .Z(n45805) );
  NOR U58662 ( .A(n45806), .B(n45805), .Z(n45807) );
  NOR U58663 ( .A(n45808), .B(n45807), .Z(n49358) );
  IV U58664 ( .A(n45809), .Z(n45810) );
  NOR U58665 ( .A(n45810), .B(n45815), .Z(n49361) );
  IV U58666 ( .A(n45811), .Z(n45813) );
  NOR U58667 ( .A(n45813), .B(n45812), .Z(n49366) );
  NOR U58668 ( .A(n49361), .B(n49366), .Z(n45833) );
  IV U58669 ( .A(n45814), .Z(n45816) );
  NOR U58670 ( .A(n45816), .B(n45815), .Z(n45830) );
  IV U58671 ( .A(n45822), .Z(n45823) );
  NOR U58672 ( .A(n45824), .B(n45823), .Z(n49364) );
  IV U58673 ( .A(n45825), .Z(n45827) );
  NOR U58674 ( .A(n45827), .B(n45826), .Z(n49363) );
  NOR U58675 ( .A(n49364), .B(n49363), .Z(n45828) );
  XOR U58676 ( .A(n49365), .B(n45828), .Z(n45829) );
  NOR U58677 ( .A(n45830), .B(n45829), .Z(n49362) );
  IV U58678 ( .A(n45830), .Z(n45832) );
  XOR U58679 ( .A(n49364), .B(n49365), .Z(n45831) );
  NOR U58680 ( .A(n45832), .B(n45831), .Z(n49360) );
  NOR U58681 ( .A(n49362), .B(n49360), .Z(n49367) );
  XOR U58682 ( .A(n45833), .B(n49367), .Z(n49359) );
  XOR U58683 ( .A(n49358), .B(n49359), .Z(n45834) );
  IV U58684 ( .A(n45834), .Z(n49374) );
  XOR U58685 ( .A(n49372), .B(n49374), .Z(n49386) );
  XOR U58686 ( .A(n45835), .B(n49386), .Z(n49388) );
  XOR U58687 ( .A(n49389), .B(n49388), .Z(n49353) );
  IV U58688 ( .A(n45836), .Z(n45838) );
  NOR U58689 ( .A(n45838), .B(n45837), .Z(n49392) );
  IV U58690 ( .A(n45839), .Z(n45840) );
  NOR U58691 ( .A(n45841), .B(n45840), .Z(n49352) );
  IV U58692 ( .A(n45842), .Z(n45843) );
  NOR U58693 ( .A(n45844), .B(n45843), .Z(n49356) );
  NOR U58694 ( .A(n49352), .B(n49356), .Z(n45845) );
  IV U58695 ( .A(n45845), .Z(n45846) );
  NOR U58696 ( .A(n49392), .B(n45846), .Z(n45847) );
  XOR U58697 ( .A(n49353), .B(n45847), .Z(n49351) );
  XOR U58698 ( .A(n49349), .B(n49351), .Z(n45848) );
  NOR U58699 ( .A(n45849), .B(n45848), .Z(n53200) );
  IV U58700 ( .A(n45850), .Z(n45851) );
  NOR U58701 ( .A(n45852), .B(n45851), .Z(n49346) );
  NOR U58702 ( .A(n49349), .B(n49346), .Z(n45853) );
  XOR U58703 ( .A(n49351), .B(n45853), .Z(n45854) );
  NOR U58704 ( .A(n45855), .B(n45854), .Z(n45856) );
  NOR U58705 ( .A(n53200), .B(n45856), .Z(n49397) );
  IV U58706 ( .A(n45857), .Z(n45858) );
  NOR U58707 ( .A(n45859), .B(n45858), .Z(n49396) );
  NOR U58708 ( .A(n45861), .B(n45860), .Z(n49400) );
  NOR U58709 ( .A(n49396), .B(n49400), .Z(n45862) );
  XOR U58710 ( .A(n49397), .B(n45862), .Z(n49345) );
  IV U58711 ( .A(n45863), .Z(n45864) );
  NOR U58712 ( .A(n45865), .B(n45864), .Z(n45872) );
  IV U58713 ( .A(n45872), .Z(n45866) );
  NOR U58714 ( .A(n49345), .B(n45866), .Z(n49337) );
  IV U58715 ( .A(n45867), .Z(n45868) );
  NOR U58716 ( .A(n45869), .B(n45868), .Z(n49341) );
  NOR U58717 ( .A(n49343), .B(n49341), .Z(n45870) );
  XOR U58718 ( .A(n45870), .B(n49345), .Z(n45871) );
  NOR U58719 ( .A(n45872), .B(n45871), .Z(n49340) );
  NOR U58720 ( .A(n49337), .B(n49340), .Z(n49334) );
  XOR U58721 ( .A(n45873), .B(n49334), .Z(n49329) );
  XOR U58722 ( .A(n49327), .B(n49329), .Z(n53148) );
  IV U58723 ( .A(n45874), .Z(n45876) );
  NOR U58724 ( .A(n45876), .B(n45875), .Z(n53153) );
  IV U58725 ( .A(n45877), .Z(n45879) );
  NOR U58726 ( .A(n45879), .B(n45878), .Z(n53147) );
  NOR U58727 ( .A(n53153), .B(n53147), .Z(n49330) );
  XOR U58728 ( .A(n53148), .B(n49330), .Z(n49322) );
  XOR U58729 ( .A(n45880), .B(n49322), .Z(n49319) );
  IV U58730 ( .A(n45881), .Z(n45882) );
  NOR U58731 ( .A(n45883), .B(n45882), .Z(n49318) );
  NOR U58732 ( .A(n45885), .B(n45884), .Z(n49315) );
  NOR U58733 ( .A(n49318), .B(n49315), .Z(n45886) );
  XOR U58734 ( .A(n49319), .B(n45886), .Z(n49404) );
  XOR U58735 ( .A(n49405), .B(n49404), .Z(n45893) );
  NOR U58736 ( .A(n45895), .B(n45893), .Z(n53243) );
  IV U58737 ( .A(n45887), .Z(n45888) );
  NOR U58738 ( .A(n45889), .B(n45888), .Z(n49312) );
  IV U58739 ( .A(n45890), .Z(n45892) );
  IV U58740 ( .A(n45891), .Z(n49408) );
  NOR U58741 ( .A(n45892), .B(n49408), .Z(n45894) );
  XOR U58742 ( .A(n45894), .B(n45893), .Z(n49313) );
  IV U58743 ( .A(n49313), .Z(n45896) );
  XOR U58744 ( .A(n49312), .B(n45896), .Z(n45898) );
  NOR U58745 ( .A(n45896), .B(n45895), .Z(n45897) );
  NOR U58746 ( .A(n45898), .B(n45897), .Z(n45899) );
  NOR U58747 ( .A(n53243), .B(n45899), .Z(n49306) );
  XOR U58748 ( .A(n49307), .B(n49306), .Z(n49309) );
  XOR U58749 ( .A(n49308), .B(n49309), .Z(n49302) );
  IV U58750 ( .A(n45900), .Z(n45902) );
  NOR U58751 ( .A(n45902), .B(n45901), .Z(n49300) );
  XOR U58752 ( .A(n49302), .B(n49300), .Z(n49304) );
  IV U58753 ( .A(n45903), .Z(n45904) );
  NOR U58754 ( .A(n45905), .B(n45904), .Z(n49303) );
  IV U58755 ( .A(n45906), .Z(n45908) );
  NOR U58756 ( .A(n45908), .B(n45907), .Z(n49294) );
  NOR U58757 ( .A(n49303), .B(n49294), .Z(n45909) );
  XOR U58758 ( .A(n49304), .B(n45909), .Z(n49291) );
  IV U58759 ( .A(n45910), .Z(n45912) );
  NOR U58760 ( .A(n45912), .B(n45911), .Z(n49296) );
  IV U58761 ( .A(n45913), .Z(n45914) );
  NOR U58762 ( .A(n45915), .B(n45914), .Z(n49292) );
  NOR U58763 ( .A(n49296), .B(n49292), .Z(n45916) );
  XOR U58764 ( .A(n49291), .B(n45916), .Z(n49425) );
  NOR U58765 ( .A(n45917), .B(n49287), .Z(n49424) );
  NOR U58766 ( .A(n49424), .B(n49421), .Z(n45918) );
  XOR U58767 ( .A(n49425), .B(n45918), .Z(n45923) );
  IV U58768 ( .A(n45923), .Z(n45919) );
  NOR U58769 ( .A(n45920), .B(n45919), .Z(n53113) );
  IV U58770 ( .A(n45924), .Z(n45922) );
  XOR U58771 ( .A(n49424), .B(n49425), .Z(n45921) );
  NOR U58772 ( .A(n45922), .B(n45921), .Z(n53112) );
  NOR U58773 ( .A(n45924), .B(n45923), .Z(n45925) );
  NOR U58774 ( .A(n53112), .B(n45925), .Z(n45926) );
  NOR U58775 ( .A(n45927), .B(n45926), .Z(n45928) );
  NOR U58776 ( .A(n53113), .B(n45928), .Z(n49280) );
  XOR U58777 ( .A(n49285), .B(n49280), .Z(n49278) );
  IV U58778 ( .A(n45929), .Z(n45930) );
  NOR U58779 ( .A(n45931), .B(n45930), .Z(n49276) );
  XOR U58780 ( .A(n49278), .B(n49276), .Z(n49274) );
  IV U58781 ( .A(n45932), .Z(n49281) );
  NOR U58782 ( .A(n49281), .B(n45933), .Z(n45938) );
  NOR U58783 ( .A(n45935), .B(n45934), .Z(n49273) );
  NOR U58784 ( .A(n49273), .B(n49271), .Z(n45936) );
  IV U58785 ( .A(n45936), .Z(n45937) );
  NOR U58786 ( .A(n45938), .B(n45937), .Z(n45939) );
  XOR U58787 ( .A(n49274), .B(n45939), .Z(n45946) );
  IV U58788 ( .A(n45946), .Z(n45945) );
  IV U58789 ( .A(n45940), .Z(n45943) );
  IV U58790 ( .A(n45941), .Z(n45942) );
  NOR U58791 ( .A(n45943), .B(n45942), .Z(n45947) );
  IV U58792 ( .A(n45947), .Z(n45944) );
  NOR U58793 ( .A(n45945), .B(n45944), .Z(n53272) );
  NOR U58794 ( .A(n45947), .B(n45946), .Z(n49270) );
  IV U58795 ( .A(n45948), .Z(n45951) );
  IV U58796 ( .A(n45949), .Z(n45950) );
  NOR U58797 ( .A(n45951), .B(n45950), .Z(n49268) );
  XOR U58798 ( .A(n49270), .B(n49268), .Z(n45952) );
  NOR U58799 ( .A(n53272), .B(n45952), .Z(n45953) );
  IV U58800 ( .A(n45953), .Z(n49264) );
  XOR U58801 ( .A(n49262), .B(n49264), .Z(n49267) );
  XOR U58802 ( .A(n45954), .B(n49267), .Z(n45955) );
  IV U58803 ( .A(n45955), .Z(n49442) );
  XOR U58804 ( .A(n49440), .B(n49442), .Z(n49253) );
  IV U58805 ( .A(n45956), .Z(n45958) );
  NOR U58806 ( .A(n45958), .B(n45957), .Z(n49439) );
  IV U58807 ( .A(n45959), .Z(n45961) );
  NOR U58808 ( .A(n45961), .B(n45960), .Z(n49252) );
  NOR U58809 ( .A(n49439), .B(n49252), .Z(n45962) );
  XOR U58810 ( .A(n49253), .B(n45962), .Z(n49247) );
  XOR U58811 ( .A(n49248), .B(n49247), .Z(n49445) );
  XOR U58812 ( .A(n45963), .B(n49445), .Z(n49448) );
  XOR U58813 ( .A(n49446), .B(n49448), .Z(n49450) );
  IV U58814 ( .A(n45964), .Z(n45968) );
  NOR U58815 ( .A(n45966), .B(n45965), .Z(n45967) );
  IV U58816 ( .A(n45967), .Z(n45971) );
  NOR U58817 ( .A(n45968), .B(n45971), .Z(n45969) );
  IV U58818 ( .A(n45969), .Z(n49449) );
  XOR U58819 ( .A(n49450), .B(n49449), .Z(n49455) );
  IV U58820 ( .A(n45970), .Z(n45972) );
  NOR U58821 ( .A(n45972), .B(n45971), .Z(n49454) );
  XOR U58822 ( .A(n49455), .B(n49454), .Z(n53056) );
  IV U58823 ( .A(n45973), .Z(n45974) );
  NOR U58824 ( .A(n45975), .B(n45974), .Z(n45980) );
  IV U58825 ( .A(n45976), .Z(n45978) );
  NOR U58826 ( .A(n45978), .B(n45977), .Z(n45979) );
  NOR U58827 ( .A(n45980), .B(n45979), .Z(n53058) );
  XOR U58828 ( .A(n53056), .B(n53058), .Z(n49461) );
  XOR U58829 ( .A(n49459), .B(n49461), .Z(n49463) );
  XOR U58830 ( .A(n49462), .B(n49463), .Z(n49245) );
  IV U58831 ( .A(n45981), .Z(n45991) );
  IV U58832 ( .A(n45982), .Z(n45983) );
  NOR U58833 ( .A(n45991), .B(n45983), .Z(n49243) );
  XOR U58834 ( .A(n49245), .B(n49243), .Z(n45984) );
  NOR U58835 ( .A(n45985), .B(n45984), .Z(n53314) );
  IV U58836 ( .A(n45986), .Z(n45987) );
  NOR U58837 ( .A(n45988), .B(n45987), .Z(n45993) );
  IV U58838 ( .A(n45989), .Z(n45990) );
  NOR U58839 ( .A(n45991), .B(n45990), .Z(n45992) );
  NOR U58840 ( .A(n45993), .B(n45992), .Z(n49246) );
  IV U58841 ( .A(n49246), .Z(n45994) );
  NOR U58842 ( .A(n49243), .B(n45994), .Z(n45995) );
  XOR U58843 ( .A(n49245), .B(n45995), .Z(n45996) );
  NOR U58844 ( .A(n45997), .B(n45996), .Z(n45998) );
  NOR U58845 ( .A(n53314), .B(n45998), .Z(n49468) );
  XOR U58846 ( .A(n45999), .B(n49468), .Z(n49242) );
  XOR U58847 ( .A(n46000), .B(n49242), .Z(n49230) );
  IV U58848 ( .A(n49230), .Z(n49232) );
  XOR U58849 ( .A(n49231), .B(n49232), .Z(n49229) );
  XOR U58850 ( .A(n46001), .B(n49229), .Z(n49224) );
  XOR U58851 ( .A(n49222), .B(n49224), .Z(n49477) );
  XOR U58852 ( .A(n49225), .B(n49477), .Z(n49217) );
  IV U58853 ( .A(n46002), .Z(n46003) );
  NOR U58854 ( .A(n46004), .B(n46003), .Z(n49218) );
  IV U58855 ( .A(n46005), .Z(n46007) );
  IV U58856 ( .A(n46006), .Z(n46010) );
  NOR U58857 ( .A(n46007), .B(n46010), .Z(n49475) );
  NOR U58858 ( .A(n49218), .B(n49475), .Z(n46008) );
  XOR U58859 ( .A(n49217), .B(n46008), .Z(n49480) );
  IV U58860 ( .A(n46009), .Z(n46011) );
  NOR U58861 ( .A(n46011), .B(n46010), .Z(n49478) );
  XOR U58862 ( .A(n49480), .B(n49478), .Z(n49483) );
  XOR U58863 ( .A(n49481), .B(n49483), .Z(n49216) );
  NOR U58864 ( .A(n46018), .B(n49216), .Z(n53023) );
  IV U58865 ( .A(n46012), .Z(n46013) );
  NOR U58866 ( .A(n46013), .B(n46023), .Z(n49211) );
  IV U58867 ( .A(n46014), .Z(n46015) );
  NOR U58868 ( .A(n46016), .B(n46015), .Z(n46017) );
  IV U58869 ( .A(n46017), .Z(n49215) );
  XOR U58870 ( .A(n49216), .B(n49215), .Z(n49212) );
  XOR U58871 ( .A(n49211), .B(n49212), .Z(n46020) );
  NOR U58872 ( .A(n49212), .B(n46018), .Z(n46019) );
  NOR U58873 ( .A(n46020), .B(n46019), .Z(n46021) );
  NOR U58874 ( .A(n53023), .B(n46021), .Z(n49203) );
  IV U58875 ( .A(n46022), .Z(n46024) );
  NOR U58876 ( .A(n46024), .B(n46023), .Z(n46025) );
  IV U58877 ( .A(n46025), .Z(n49204) );
  XOR U58878 ( .A(n49203), .B(n49204), .Z(n49207) );
  XOR U58879 ( .A(n49206), .B(n49207), .Z(n49196) );
  XOR U58880 ( .A(n49195), .B(n49196), .Z(n49200) );
  XOR U58881 ( .A(n49198), .B(n49200), .Z(n49487) );
  XOR U58882 ( .A(n49485), .B(n49487), .Z(n49489) );
  NOR U58883 ( .A(n46031), .B(n49489), .Z(n53009) );
  IV U58884 ( .A(n46026), .Z(n46028) );
  NOR U58885 ( .A(n46028), .B(n46027), .Z(n49488) );
  XOR U58886 ( .A(n49488), .B(n49489), .Z(n49194) );
  IV U58887 ( .A(n46029), .Z(n46030) );
  NOR U58888 ( .A(n46038), .B(n46030), .Z(n46032) );
  IV U58889 ( .A(n46032), .Z(n49193) );
  XOR U58890 ( .A(n49194), .B(n49193), .Z(n46034) );
  NOR U58891 ( .A(n46032), .B(n46031), .Z(n46033) );
  NOR U58892 ( .A(n46034), .B(n46033), .Z(n46035) );
  NOR U58893 ( .A(n53009), .B(n46035), .Z(n46036) );
  IV U58894 ( .A(n46036), .Z(n49192) );
  IV U58895 ( .A(n46037), .Z(n46039) );
  NOR U58896 ( .A(n46039), .B(n46038), .Z(n49190) );
  IV U58897 ( .A(n46040), .Z(n49182) );
  NOR U58898 ( .A(n49182), .B(n46041), .Z(n46042) );
  NOR U58899 ( .A(n49190), .B(n46042), .Z(n46043) );
  XOR U58900 ( .A(n49192), .B(n46043), .Z(n49176) );
  IV U58901 ( .A(n46044), .Z(n46046) );
  NOR U58902 ( .A(n46046), .B(n46045), .Z(n46055) );
  IV U58903 ( .A(n46055), .Z(n49178) );
  NOR U58904 ( .A(n49176), .B(n49178), .Z(n46057) );
  NOR U58905 ( .A(n46048), .B(n46047), .Z(n46051) );
  IV U58906 ( .A(n46051), .Z(n46050) );
  XOR U58907 ( .A(n49190), .B(n49192), .Z(n46049) );
  NOR U58908 ( .A(n46050), .B(n46049), .Z(n52989) );
  NOR U58909 ( .A(n49176), .B(n46051), .Z(n46052) );
  NOR U58910 ( .A(n52989), .B(n46052), .Z(n46053) );
  IV U58911 ( .A(n46053), .Z(n46054) );
  NOR U58912 ( .A(n46055), .B(n46054), .Z(n46056) );
  NOR U58913 ( .A(n46057), .B(n46056), .Z(n53376) );
  XOR U58914 ( .A(n49179), .B(n53376), .Z(n49172) );
  IV U58915 ( .A(n46058), .Z(n46059) );
  NOR U58916 ( .A(n46060), .B(n46059), .Z(n49174) );
  IV U58917 ( .A(n46061), .Z(n46063) );
  NOR U58918 ( .A(n46063), .B(n46062), .Z(n49171) );
  NOR U58919 ( .A(n49174), .B(n49171), .Z(n46064) );
  XOR U58920 ( .A(n49172), .B(n46064), .Z(n49169) );
  XOR U58921 ( .A(n46065), .B(n49169), .Z(n49160) );
  XOR U58922 ( .A(n49159), .B(n49160), .Z(n49162) );
  IV U58923 ( .A(n46066), .Z(n46067) );
  NOR U58924 ( .A(n46068), .B(n46067), .Z(n49161) );
  IV U58925 ( .A(n46069), .Z(n46071) );
  NOR U58926 ( .A(n46071), .B(n46070), .Z(n49164) );
  NOR U58927 ( .A(n49161), .B(n49164), .Z(n46072) );
  XOR U58928 ( .A(n49162), .B(n46072), .Z(n49500) );
  XOR U58929 ( .A(n49499), .B(n49500), .Z(n53390) );
  XOR U58930 ( .A(n49502), .B(n53390), .Z(n49508) );
  IV U58931 ( .A(n49508), .Z(n49506) );
  IV U58932 ( .A(n46073), .Z(n46075) );
  NOR U58933 ( .A(n46075), .B(n46074), .Z(n49507) );
  XOR U58934 ( .A(n49506), .B(n49507), .Z(n49155) );
  XOR U58935 ( .A(n46076), .B(n49155), .Z(n46089) );
  IV U58936 ( .A(n46089), .Z(n46085) );
  IV U58937 ( .A(n46077), .Z(n46079) );
  NOR U58938 ( .A(n46079), .B(n46078), .Z(n46086) );
  IV U58939 ( .A(n46080), .Z(n46082) );
  NOR U58940 ( .A(n46082), .B(n46081), .Z(n46088) );
  NOR U58941 ( .A(n46086), .B(n46088), .Z(n46083) );
  IV U58942 ( .A(n46083), .Z(n46084) );
  NOR U58943 ( .A(n46085), .B(n46084), .Z(n46092) );
  IV U58944 ( .A(n46086), .Z(n46087) );
  NOR U58945 ( .A(n46087), .B(n49155), .Z(n52966) );
  IV U58946 ( .A(n46088), .Z(n46090) );
  NOR U58947 ( .A(n46090), .B(n46089), .Z(n52961) );
  NOR U58948 ( .A(n52966), .B(n52961), .Z(n46091) );
  IV U58949 ( .A(n46091), .Z(n49517) );
  NOR U58950 ( .A(n46092), .B(n49517), .Z(n49148) );
  XOR U58951 ( .A(n49149), .B(n49148), .Z(n49152) );
  IV U58952 ( .A(n46093), .Z(n46094) );
  NOR U58953 ( .A(n46095), .B(n46094), .Z(n49150) );
  XOR U58954 ( .A(n49152), .B(n49150), .Z(n49146) );
  XOR U58955 ( .A(n49147), .B(n49146), .Z(n49133) );
  IV U58956 ( .A(n46096), .Z(n46098) );
  NOR U58957 ( .A(n46098), .B(n46097), .Z(n46102) );
  IV U58958 ( .A(n46099), .Z(n46101) );
  NOR U58959 ( .A(n46101), .B(n46100), .Z(n49132) );
  NOR U58960 ( .A(n46102), .B(n49132), .Z(n46103) );
  XOR U58961 ( .A(n49133), .B(n46103), .Z(n49131) );
  IV U58962 ( .A(n46104), .Z(n46105) );
  NOR U58963 ( .A(n46106), .B(n46105), .Z(n49129) );
  IV U58964 ( .A(n46107), .Z(n46109) );
  NOR U58965 ( .A(n46109), .B(n46108), .Z(n49127) );
  NOR U58966 ( .A(n49129), .B(n49127), .Z(n46110) );
  XOR U58967 ( .A(n49131), .B(n46110), .Z(n46111) );
  NOR U58968 ( .A(n46112), .B(n46111), .Z(n46115) );
  IV U58969 ( .A(n46112), .Z(n46114) );
  XOR U58970 ( .A(n49129), .B(n49131), .Z(n46113) );
  NOR U58971 ( .A(n46114), .B(n46113), .Z(n53420) );
  NOR U58972 ( .A(n46115), .B(n53420), .Z(n49124) );
  NOR U58973 ( .A(n46117), .B(n46116), .Z(n46118) );
  IV U58974 ( .A(n46118), .Z(n49126) );
  XOR U58975 ( .A(n49124), .B(n49126), .Z(n49120) );
  XOR U58976 ( .A(n49118), .B(n49120), .Z(n49123) );
  NOR U58977 ( .A(n46119), .B(n49123), .Z(n52932) );
  IV U58978 ( .A(n46120), .Z(n46124) );
  NOR U58979 ( .A(n46121), .B(n46127), .Z(n46122) );
  IV U58980 ( .A(n46122), .Z(n46123) );
  NOR U58981 ( .A(n46124), .B(n46123), .Z(n49121) );
  XOR U58982 ( .A(n49123), .B(n49121), .Z(n49528) );
  IV U58983 ( .A(n46125), .Z(n46126) );
  NOR U58984 ( .A(n46127), .B(n46126), .Z(n46128) );
  IV U58985 ( .A(n46128), .Z(n49527) );
  XOR U58986 ( .A(n49528), .B(n49527), .Z(n46129) );
  NOR U58987 ( .A(n46130), .B(n46129), .Z(n46131) );
  NOR U58988 ( .A(n52932), .B(n46131), .Z(n49116) );
  IV U58989 ( .A(n46132), .Z(n46134) );
  NOR U58990 ( .A(n46134), .B(n46133), .Z(n49523) );
  IV U58991 ( .A(n46135), .Z(n46136) );
  NOR U58992 ( .A(n46136), .B(n46140), .Z(n49115) );
  NOR U58993 ( .A(n49523), .B(n49115), .Z(n46137) );
  XOR U58994 ( .A(n49116), .B(n46137), .Z(n49114) );
  IV U58995 ( .A(n46138), .Z(n46139) );
  NOR U58996 ( .A(n46140), .B(n46139), .Z(n49112) );
  IV U58997 ( .A(n46141), .Z(n46144) );
  IV U58998 ( .A(n46142), .Z(n46143) );
  NOR U58999 ( .A(n46144), .B(n46143), .Z(n49110) );
  NOR U59000 ( .A(n49112), .B(n49110), .Z(n46145) );
  XOR U59001 ( .A(n49114), .B(n46145), .Z(n49104) );
  XOR U59002 ( .A(n49105), .B(n49104), .Z(n49540) );
  IV U59003 ( .A(n46146), .Z(n46148) );
  NOR U59004 ( .A(n46148), .B(n46147), .Z(n49106) );
  XOR U59005 ( .A(n49540), .B(n49106), .Z(n46149) );
  XOR U59006 ( .A(n46150), .B(n46149), .Z(n49542) );
  XOR U59007 ( .A(n46151), .B(n49542), .Z(n49100) );
  XOR U59008 ( .A(n46152), .B(n49100), .Z(n49561) );
  XOR U59009 ( .A(n49560), .B(n49561), .Z(n46163) );
  IV U59010 ( .A(n46155), .Z(n46153) );
  NOR U59011 ( .A(n46169), .B(n46153), .Z(n46160) );
  IV U59012 ( .A(n46154), .Z(n46157) );
  XOR U59013 ( .A(n46155), .B(n46169), .Z(n46156) );
  NOR U59014 ( .A(n46157), .B(n46156), .Z(n46162) );
  NOR U59015 ( .A(n46160), .B(n46162), .Z(n46158) );
  IV U59016 ( .A(n46158), .Z(n46159) );
  NOR U59017 ( .A(n46163), .B(n46159), .Z(n46167) );
  IV U59018 ( .A(n46160), .Z(n46161) );
  NOR U59019 ( .A(n49561), .B(n46161), .Z(n49562) );
  IV U59020 ( .A(n46162), .Z(n46165) );
  IV U59021 ( .A(n46163), .Z(n46164) );
  NOR U59022 ( .A(n46165), .B(n46164), .Z(n49567) );
  NOR U59023 ( .A(n49562), .B(n49567), .Z(n52917) );
  IV U59024 ( .A(n52917), .Z(n46166) );
  NOR U59025 ( .A(n46167), .B(n46166), .Z(n49565) );
  IV U59026 ( .A(n46168), .Z(n46170) );
  NOR U59027 ( .A(n46170), .B(n46169), .Z(n49564) );
  NOR U59028 ( .A(n46172), .B(n46171), .Z(n49569) );
  NOR U59029 ( .A(n49564), .B(n49569), .Z(n46173) );
  XOR U59030 ( .A(n49565), .B(n46173), .Z(n49577) );
  IV U59031 ( .A(n46174), .Z(n46176) );
  IV U59032 ( .A(n46175), .Z(n46181) );
  NOR U59033 ( .A(n46176), .B(n46181), .Z(n49575) );
  XOR U59034 ( .A(n49577), .B(n49575), .Z(n49585) );
  IV U59035 ( .A(n46177), .Z(n46178) );
  NOR U59036 ( .A(n46179), .B(n46178), .Z(n49584) );
  IV U59037 ( .A(n46180), .Z(n46182) );
  NOR U59038 ( .A(n46182), .B(n46181), .Z(n49578) );
  NOR U59039 ( .A(n49584), .B(n49578), .Z(n46183) );
  XOR U59040 ( .A(n49585), .B(n46183), .Z(n49096) );
  XOR U59041 ( .A(n46184), .B(n49096), .Z(n49091) );
  XOR U59042 ( .A(n49090), .B(n49091), .Z(n49094) );
  XOR U59043 ( .A(n49093), .B(n49094), .Z(n49087) );
  XOR U59044 ( .A(n46185), .B(n49087), .Z(n49081) );
  XOR U59045 ( .A(n49079), .B(n49081), .Z(n49082) );
  XOR U59046 ( .A(n49083), .B(n49082), .Z(n49073) );
  IV U59047 ( .A(n46186), .Z(n46187) );
  NOR U59048 ( .A(n46188), .B(n46187), .Z(n49075) );
  IV U59049 ( .A(n46189), .Z(n46190) );
  NOR U59050 ( .A(n46191), .B(n46190), .Z(n49072) );
  NOR U59051 ( .A(n49075), .B(n49072), .Z(n46192) );
  XOR U59052 ( .A(n49073), .B(n46192), .Z(n49595) );
  XOR U59053 ( .A(n49594), .B(n49595), .Z(n49601) );
  XOR U59054 ( .A(n49597), .B(n49601), .Z(n49070) );
  XOR U59055 ( .A(n46193), .B(n49070), .Z(n49068) );
  XOR U59056 ( .A(n49066), .B(n49068), .Z(n49608) );
  IV U59057 ( .A(n46194), .Z(n46196) );
  NOR U59058 ( .A(n46196), .B(n46195), .Z(n46197) );
  IV U59059 ( .A(n46197), .Z(n49605) );
  XOR U59060 ( .A(n49608), .B(n49605), .Z(n49613) );
  IV U59061 ( .A(n46198), .Z(n46199) );
  NOR U59062 ( .A(n46199), .B(n46201), .Z(n49614) );
  IV U59063 ( .A(n46200), .Z(n46202) );
  NOR U59064 ( .A(n46202), .B(n46201), .Z(n49606) );
  NOR U59065 ( .A(n49614), .B(n49606), .Z(n46203) );
  XOR U59066 ( .A(n49613), .B(n46203), .Z(n49612) );
  IV U59067 ( .A(n46204), .Z(n46205) );
  NOR U59068 ( .A(n46206), .B(n46205), .Z(n46212) );
  IV U59069 ( .A(n46212), .Z(n46207) );
  NOR U59070 ( .A(n49612), .B(n46207), .Z(n49065) );
  IV U59071 ( .A(n46208), .Z(n46209) );
  NOR U59072 ( .A(n46210), .B(n46209), .Z(n49610) );
  XOR U59073 ( .A(n49610), .B(n49612), .Z(n46223) );
  IV U59074 ( .A(n46223), .Z(n46211) );
  NOR U59075 ( .A(n46212), .B(n46211), .Z(n46213) );
  NOR U59076 ( .A(n49065), .B(n46213), .Z(n46214) );
  NOR U59077 ( .A(n46215), .B(n46214), .Z(n46217) );
  IV U59078 ( .A(n46215), .Z(n46216) );
  NOR U59079 ( .A(n46223), .B(n46216), .Z(n53540) );
  NOR U59080 ( .A(n46217), .B(n53540), .Z(n49061) );
  IV U59081 ( .A(n46233), .Z(n46218) );
  NOR U59082 ( .A(n46232), .B(n46218), .Z(n46228) );
  IV U59083 ( .A(n46228), .Z(n49063) );
  NOR U59084 ( .A(n49061), .B(n49063), .Z(n46230) );
  IV U59085 ( .A(n46219), .Z(n46221) );
  NOR U59086 ( .A(n46221), .B(n46220), .Z(n46224) );
  IV U59087 ( .A(n46224), .Z(n46222) );
  NOR U59088 ( .A(n46223), .B(n46222), .Z(n52864) );
  NOR U59089 ( .A(n49061), .B(n46224), .Z(n46225) );
  NOR U59090 ( .A(n52864), .B(n46225), .Z(n46226) );
  IV U59091 ( .A(n46226), .Z(n46227) );
  NOR U59092 ( .A(n46228), .B(n46227), .Z(n46229) );
  NOR U59093 ( .A(n46230), .B(n46229), .Z(n49058) );
  IV U59094 ( .A(n46231), .Z(n46238) );
  XOR U59095 ( .A(n46233), .B(n46232), .Z(n46234) );
  NOR U59096 ( .A(n46235), .B(n46234), .Z(n46236) );
  IV U59097 ( .A(n46236), .Z(n46237) );
  NOR U59098 ( .A(n46238), .B(n46237), .Z(n49056) );
  XOR U59099 ( .A(n49058), .B(n49056), .Z(n49059) );
  XOR U59100 ( .A(n49060), .B(n49059), .Z(n49054) );
  NOR U59101 ( .A(n46240), .B(n46239), .Z(n52846) );
  NOR U59102 ( .A(n52846), .B(n53545), .Z(n49055) );
  XOR U59103 ( .A(n49054), .B(n49055), .Z(n49047) );
  XOR U59104 ( .A(n49046), .B(n49047), .Z(n49051) );
  XOR U59105 ( .A(n49049), .B(n49051), .Z(n49042) );
  XOR U59106 ( .A(n49040), .B(n49042), .Z(n49043) );
  NOR U59107 ( .A(n46248), .B(n49043), .Z(n53557) );
  IV U59108 ( .A(n46241), .Z(n46242) );
  NOR U59109 ( .A(n46243), .B(n46242), .Z(n49622) );
  IV U59110 ( .A(n46244), .Z(n46245) );
  NOR U59111 ( .A(n46246), .B(n46245), .Z(n46247) );
  IV U59112 ( .A(n46247), .Z(n49044) );
  XOR U59113 ( .A(n49044), .B(n49043), .Z(n49623) );
  XOR U59114 ( .A(n49622), .B(n49623), .Z(n46250) );
  NOR U59115 ( .A(n49623), .B(n46248), .Z(n46249) );
  NOR U59116 ( .A(n46250), .B(n46249), .Z(n46251) );
  NOR U59117 ( .A(n53557), .B(n46251), .Z(n49627) );
  XOR U59118 ( .A(n49626), .B(n49627), .Z(n49633) );
  IV U59119 ( .A(n46252), .Z(n46253) );
  NOR U59120 ( .A(n46254), .B(n46253), .Z(n52827) );
  IV U59121 ( .A(n46255), .Z(n46257) );
  NOR U59122 ( .A(n46257), .B(n46256), .Z(n52834) );
  NOR U59123 ( .A(n52827), .B(n52834), .Z(n49634) );
  XOR U59124 ( .A(n49633), .B(n49634), .Z(n49038) );
  XOR U59125 ( .A(n49037), .B(n49038), .Z(n49641) );
  XOR U59126 ( .A(n49639), .B(n49641), .Z(n49646) );
  XOR U59127 ( .A(n46258), .B(n49646), .Z(n49649) );
  XOR U59128 ( .A(n49650), .B(n49649), .Z(n49035) );
  XOR U59129 ( .A(n49034), .B(n49035), .Z(n49029) );
  XOR U59130 ( .A(n49028), .B(n49029), .Z(n49032) );
  XOR U59131 ( .A(n46259), .B(n49032), .Z(n49659) );
  XOR U59132 ( .A(n46260), .B(n49659), .Z(n46263) );
  IV U59133 ( .A(n46263), .Z(n46261) );
  NOR U59134 ( .A(n46262), .B(n46261), .Z(n53580) );
  NOR U59135 ( .A(n46264), .B(n46263), .Z(n49665) );
  IV U59136 ( .A(n46265), .Z(n46266) );
  NOR U59137 ( .A(n46267), .B(n46266), .Z(n49663) );
  XOR U59138 ( .A(n49665), .B(n49663), .Z(n46268) );
  NOR U59139 ( .A(n53580), .B(n46268), .Z(n46269) );
  IV U59140 ( .A(n46269), .Z(n49670) );
  XOR U59141 ( .A(n49661), .B(n49670), .Z(n49017) );
  XOR U59142 ( .A(n46270), .B(n49017), .Z(n49010) );
  XOR U59143 ( .A(n46271), .B(n49010), .Z(n49674) );
  XOR U59144 ( .A(n49672), .B(n49674), .Z(n49676) );
  XOR U59145 ( .A(n49675), .B(n49676), .Z(n49690) );
  XOR U59146 ( .A(n46272), .B(n49690), .Z(n49000) );
  XOR U59147 ( .A(n46273), .B(n49000), .Z(n49694) );
  XOR U59148 ( .A(n46274), .B(n49694), .Z(n48994) );
  XOR U59149 ( .A(n46275), .B(n48994), .Z(n48991) );
  IV U59150 ( .A(n46276), .Z(n46278) );
  NOR U59151 ( .A(n46278), .B(n46277), .Z(n48988) );
  NOR U59152 ( .A(n48990), .B(n48988), .Z(n46279) );
  XOR U59153 ( .A(n48991), .B(n46279), .Z(n46293) );
  IV U59154 ( .A(n46293), .Z(n46286) );
  IV U59155 ( .A(n46280), .Z(n46281) );
  NOR U59156 ( .A(n46282), .B(n46281), .Z(n46283) );
  IV U59157 ( .A(n46283), .Z(n46284) );
  NOR U59158 ( .A(n46289), .B(n46284), .Z(n46296) );
  IV U59159 ( .A(n46296), .Z(n46285) );
  NOR U59160 ( .A(n46286), .B(n46285), .Z(n52753) );
  XOR U59161 ( .A(n48990), .B(n48991), .Z(n46291) );
  IV U59162 ( .A(n46287), .Z(n46288) );
  NOR U59163 ( .A(n46289), .B(n46288), .Z(n46292) );
  IV U59164 ( .A(n46292), .Z(n46290) );
  NOR U59165 ( .A(n46291), .B(n46290), .Z(n52750) );
  NOR U59166 ( .A(n46293), .B(n46292), .Z(n46294) );
  NOR U59167 ( .A(n52750), .B(n46294), .Z(n46295) );
  NOR U59168 ( .A(n46296), .B(n46295), .Z(n46297) );
  NOR U59169 ( .A(n52753), .B(n46297), .Z(n46298) );
  IV U59170 ( .A(n46298), .Z(n49701) );
  IV U59171 ( .A(n46299), .Z(n46300) );
  NOR U59172 ( .A(n46301), .B(n46300), .Z(n49699) );
  XOR U59173 ( .A(n49701), .B(n49699), .Z(n48983) );
  XOR U59174 ( .A(n48982), .B(n48983), .Z(n48987) );
  IV U59175 ( .A(n46302), .Z(n46304) );
  NOR U59176 ( .A(n46304), .B(n46303), .Z(n48985) );
  XOR U59177 ( .A(n48987), .B(n48985), .Z(n49705) );
  NOR U59178 ( .A(n46306), .B(n46305), .Z(n46311) );
  IV U59179 ( .A(n46306), .Z(n46308) );
  NOR U59180 ( .A(n46308), .B(n46307), .Z(n48980) );
  NOR U59181 ( .A(n46309), .B(n48980), .Z(n46310) );
  NOR U59182 ( .A(n46311), .B(n46310), .Z(n46312) );
  XOR U59183 ( .A(n49705), .B(n46312), .Z(n49710) );
  IV U59184 ( .A(n46313), .Z(n46314) );
  NOR U59185 ( .A(n49706), .B(n46314), .Z(n46315) );
  IV U59186 ( .A(n46315), .Z(n49709) );
  XOR U59187 ( .A(n49710), .B(n49709), .Z(n48978) );
  IV U59188 ( .A(n46316), .Z(n46317) );
  NOR U59189 ( .A(n46318), .B(n46317), .Z(n53643) );
  NOR U59190 ( .A(n46320), .B(n46319), .Z(n52732) );
  NOR U59191 ( .A(n53643), .B(n52732), .Z(n48979) );
  XOR U59192 ( .A(n48978), .B(n48979), .Z(n49720) );
  XOR U59193 ( .A(n49718), .B(n49720), .Z(n48976) );
  XOR U59194 ( .A(n48975), .B(n48976), .Z(n49729) );
  XOR U59195 ( .A(n46321), .B(n49729), .Z(n48964) );
  IV U59196 ( .A(n46322), .Z(n46324) );
  NOR U59197 ( .A(n46324), .B(n46323), .Z(n48970) );
  NOR U59198 ( .A(n48963), .B(n48970), .Z(n46325) );
  XOR U59199 ( .A(n48964), .B(n46325), .Z(n49746) );
  IV U59200 ( .A(n46326), .Z(n46329) );
  IV U59201 ( .A(n46327), .Z(n46328) );
  NOR U59202 ( .A(n46329), .B(n46328), .Z(n48966) );
  IV U59203 ( .A(n46330), .Z(n46336) );
  IV U59204 ( .A(n46331), .Z(n46332) );
  NOR U59205 ( .A(n46336), .B(n46332), .Z(n49745) );
  NOR U59206 ( .A(n48966), .B(n49745), .Z(n46333) );
  XOR U59207 ( .A(n49746), .B(n46333), .Z(n49739) );
  IV U59208 ( .A(n46334), .Z(n46335) );
  NOR U59209 ( .A(n46336), .B(n46335), .Z(n49742) );
  IV U59210 ( .A(n46337), .Z(n46338) );
  NOR U59211 ( .A(n46339), .B(n46338), .Z(n49740) );
  NOR U59212 ( .A(n49742), .B(n49740), .Z(n46340) );
  XOR U59213 ( .A(n49739), .B(n46340), .Z(n49752) );
  IV U59214 ( .A(n46341), .Z(n46343) );
  NOR U59215 ( .A(n46343), .B(n46342), .Z(n49751) );
  IV U59216 ( .A(n46344), .Z(n46346) );
  NOR U59217 ( .A(n46346), .B(n46345), .Z(n49749) );
  NOR U59218 ( .A(n49751), .B(n49749), .Z(n46347) );
  XOR U59219 ( .A(n49752), .B(n46347), .Z(n46348) );
  XOR U59220 ( .A(n46349), .B(n46348), .Z(n48949) );
  XOR U59221 ( .A(n46350), .B(n48949), .Z(n49759) );
  IV U59222 ( .A(n46351), .Z(n46353) );
  NOR U59223 ( .A(n46353), .B(n46352), .Z(n49758) );
  IV U59224 ( .A(n46354), .Z(n46356) );
  NOR U59225 ( .A(n46356), .B(n46355), .Z(n48943) );
  NOR U59226 ( .A(n49758), .B(n48943), .Z(n46357) );
  XOR U59227 ( .A(n49759), .B(n46357), .Z(n48941) );
  XOR U59228 ( .A(n46358), .B(n48941), .Z(n48938) );
  XOR U59229 ( .A(n48937), .B(n48938), .Z(n46367) );
  IV U59230 ( .A(n46359), .Z(n46360) );
  NOR U59231 ( .A(n46361), .B(n46360), .Z(n46370) );
  NOR U59232 ( .A(n46363), .B(n46362), .Z(n46366) );
  NOR U59233 ( .A(n46370), .B(n46366), .Z(n46364) );
  IV U59234 ( .A(n46364), .Z(n46365) );
  NOR U59235 ( .A(n46367), .B(n46365), .Z(n46373) );
  IV U59236 ( .A(n46366), .Z(n46369) );
  IV U59237 ( .A(n46367), .Z(n46368) );
  NOR U59238 ( .A(n46369), .B(n46368), .Z(n52710) );
  IV U59239 ( .A(n46370), .Z(n46371) );
  NOR U59240 ( .A(n48938), .B(n46371), .Z(n52712) );
  NOR U59241 ( .A(n52710), .B(n52712), .Z(n46372) );
  IV U59242 ( .A(n46372), .Z(n48939) );
  NOR U59243 ( .A(n46373), .B(n48939), .Z(n48932) );
  XOR U59244 ( .A(n48934), .B(n48932), .Z(n48935) );
  XOR U59245 ( .A(n48936), .B(n48935), .Z(n48930) );
  IV U59246 ( .A(n46374), .Z(n46375) );
  NOR U59247 ( .A(n46376), .B(n46375), .Z(n52701) );
  IV U59248 ( .A(n46377), .Z(n46379) );
  NOR U59249 ( .A(n46379), .B(n46378), .Z(n52696) );
  NOR U59250 ( .A(n52701), .B(n52696), .Z(n48931) );
  XOR U59251 ( .A(n48930), .B(n48931), .Z(n48925) );
  XOR U59252 ( .A(n48924), .B(n48925), .Z(n48928) );
  XOR U59253 ( .A(n48927), .B(n48928), .Z(n48923) );
  XOR U59254 ( .A(n46380), .B(n48923), .Z(n48913) );
  IV U59255 ( .A(n46381), .Z(n46383) );
  NOR U59256 ( .A(n46383), .B(n46382), .Z(n48912) );
  IV U59257 ( .A(n46384), .Z(n46385) );
  NOR U59258 ( .A(n46386), .B(n46385), .Z(n48917) );
  NOR U59259 ( .A(n48912), .B(n48917), .Z(n46387) );
  XOR U59260 ( .A(n48913), .B(n46387), .Z(n49769) );
  XOR U59261 ( .A(n49768), .B(n49769), .Z(n49772) );
  XOR U59262 ( .A(n49771), .B(n49772), .Z(n49776) );
  XOR U59263 ( .A(n49775), .B(n49776), .Z(n48909) );
  NOR U59264 ( .A(n46392), .B(n48909), .Z(n55865) );
  IV U59265 ( .A(n46388), .Z(n46391) );
  IV U59266 ( .A(n46389), .Z(n46390) );
  NOR U59267 ( .A(n46391), .B(n46390), .Z(n48908) );
  IV U59268 ( .A(n48909), .Z(n46393) );
  XOR U59269 ( .A(n48908), .B(n46393), .Z(n46395) );
  NOR U59270 ( .A(n46393), .B(n46392), .Z(n46394) );
  NOR U59271 ( .A(n46395), .B(n46394), .Z(n48905) );
  NOR U59272 ( .A(n55865), .B(n48905), .Z(n49782) );
  IV U59273 ( .A(n46396), .Z(n46398) );
  NOR U59274 ( .A(n46398), .B(n46397), .Z(n48904) );
  IV U59275 ( .A(n46399), .Z(n46403) );
  NOR U59276 ( .A(n46401), .B(n46400), .Z(n46402) );
  IV U59277 ( .A(n46402), .Z(n46406) );
  NOR U59278 ( .A(n46403), .B(n46406), .Z(n49783) );
  NOR U59279 ( .A(n48904), .B(n49783), .Z(n46404) );
  XOR U59280 ( .A(n49782), .B(n46404), .Z(n48903) );
  IV U59281 ( .A(n46405), .Z(n46407) );
  NOR U59282 ( .A(n46407), .B(n46406), .Z(n48901) );
  XOR U59283 ( .A(n48903), .B(n48901), .Z(n49799) );
  XOR U59284 ( .A(n49798), .B(n49799), .Z(n49807) );
  XOR U59285 ( .A(n49806), .B(n49807), .Z(n49815) );
  XOR U59286 ( .A(n46408), .B(n49815), .Z(n49818) );
  XOR U59287 ( .A(n46409), .B(n49818), .Z(n48894) );
  XOR U59288 ( .A(n48892), .B(n48894), .Z(n49830) );
  XOR U59289 ( .A(n48889), .B(n49830), .Z(n46417) );
  IV U59290 ( .A(n46410), .Z(n46413) );
  NOR U59291 ( .A(n46411), .B(n46419), .Z(n46412) );
  IV U59292 ( .A(n46412), .Z(n46424) );
  NOR U59293 ( .A(n46413), .B(n46424), .Z(n46414) );
  IV U59294 ( .A(n46414), .Z(n46415) );
  NOR U59295 ( .A(n46423), .B(n46415), .Z(n46428) );
  IV U59296 ( .A(n46428), .Z(n46416) );
  NOR U59297 ( .A(n46417), .B(n46416), .Z(n53738) );
  IV U59298 ( .A(n46418), .Z(n46420) );
  NOR U59299 ( .A(n46420), .B(n46419), .Z(n49829) );
  NOR U59300 ( .A(n48889), .B(n49829), .Z(n46421) );
  IV U59301 ( .A(n46421), .Z(n46422) );
  XOR U59302 ( .A(n46422), .B(n49830), .Z(n49833) );
  IV U59303 ( .A(n46423), .Z(n46425) );
  NOR U59304 ( .A(n46425), .B(n46424), .Z(n46426) );
  IV U59305 ( .A(n46426), .Z(n49832) );
  XOR U59306 ( .A(n49833), .B(n49832), .Z(n46427) );
  NOR U59307 ( .A(n46428), .B(n46427), .Z(n46429) );
  NOR U59308 ( .A(n53738), .B(n46429), .Z(n48886) );
  IV U59309 ( .A(n46430), .Z(n46432) );
  NOR U59310 ( .A(n46432), .B(n46431), .Z(n46433) );
  IV U59311 ( .A(n46433), .Z(n48887) );
  XOR U59312 ( .A(n48886), .B(n48887), .Z(n49838) );
  XOR U59313 ( .A(n49836), .B(n49838), .Z(n49841) );
  XOR U59314 ( .A(n46434), .B(n49841), .Z(n48878) );
  IV U59315 ( .A(n46435), .Z(n46436) );
  NOR U59316 ( .A(n46437), .B(n46436), .Z(n48880) );
  IV U59317 ( .A(n46438), .Z(n46439) );
  NOR U59318 ( .A(n46440), .B(n46439), .Z(n48877) );
  NOR U59319 ( .A(n48880), .B(n48877), .Z(n46441) );
  XOR U59320 ( .A(n48878), .B(n46441), .Z(n49847) );
  XOR U59321 ( .A(n49846), .B(n49847), .Z(n48875) );
  XOR U59322 ( .A(n46442), .B(n48875), .Z(n49854) );
  XOR U59323 ( .A(n49852), .B(n49854), .Z(n46443) );
  XOR U59324 ( .A(n46444), .B(n46443), .Z(n48863) );
  IV U59325 ( .A(n46445), .Z(n46448) );
  IV U59326 ( .A(n46446), .Z(n46447) );
  NOR U59327 ( .A(n46448), .B(n46447), .Z(n48861) );
  IV U59328 ( .A(n48861), .Z(n48862) );
  XOR U59329 ( .A(n48863), .B(n48862), .Z(n49859) );
  IV U59330 ( .A(n46449), .Z(n46450) );
  NOR U59331 ( .A(n46457), .B(n46450), .Z(n48865) );
  IV U59332 ( .A(n46451), .Z(n46453) );
  NOR U59333 ( .A(n46453), .B(n46452), .Z(n49860) );
  NOR U59334 ( .A(n48865), .B(n49860), .Z(n46454) );
  XOR U59335 ( .A(n49859), .B(n46454), .Z(n48851) );
  IV U59336 ( .A(n46455), .Z(n46456) );
  NOR U59337 ( .A(n46457), .B(n46456), .Z(n48849) );
  XOR U59338 ( .A(n48851), .B(n48849), .Z(n48853) );
  XOR U59339 ( .A(n46458), .B(n48853), .Z(n48846) );
  XOR U59340 ( .A(n48844), .B(n48846), .Z(n48839) );
  XOR U59341 ( .A(n48838), .B(n48839), .Z(n48842) );
  XOR U59342 ( .A(n48841), .B(n48842), .Z(n48832) );
  IV U59343 ( .A(n46459), .Z(n46461) );
  NOR U59344 ( .A(n46461), .B(n46460), .Z(n46466) );
  IV U59345 ( .A(n46462), .Z(n46463) );
  NOR U59346 ( .A(n46464), .B(n46463), .Z(n46465) );
  NOR U59347 ( .A(n46466), .B(n46465), .Z(n48833) );
  XOR U59348 ( .A(n48832), .B(n48833), .Z(n48834) );
  XOR U59349 ( .A(n48835), .B(n48834), .Z(n53783) );
  XOR U59350 ( .A(n53784), .B(n53783), .Z(n46467) );
  XOR U59351 ( .A(n46468), .B(n46467), .Z(n49876) );
  IV U59352 ( .A(n46469), .Z(n46471) );
  NOR U59353 ( .A(n46471), .B(n46470), .Z(n49872) );
  IV U59354 ( .A(n46472), .Z(n46473) );
  NOR U59355 ( .A(n46474), .B(n46473), .Z(n49874) );
  NOR U59356 ( .A(n49872), .B(n49874), .Z(n46475) );
  XOR U59357 ( .A(n49876), .B(n46475), .Z(n49877) );
  XOR U59358 ( .A(n49878), .B(n49877), .Z(n49891) );
  IV U59359 ( .A(n49891), .Z(n46483) );
  IV U59360 ( .A(n46476), .Z(n46477) );
  NOR U59361 ( .A(n46478), .B(n46477), .Z(n49890) );
  IV U59362 ( .A(n46479), .Z(n46481) );
  NOR U59363 ( .A(n46481), .B(n46480), .Z(n49879) );
  NOR U59364 ( .A(n49890), .B(n49879), .Z(n46482) );
  XOR U59365 ( .A(n46483), .B(n46482), .Z(n49885) );
  IV U59366 ( .A(n46484), .Z(n46486) );
  NOR U59367 ( .A(n46486), .B(n46485), .Z(n49883) );
  XOR U59368 ( .A(n49885), .B(n49883), .Z(n49888) );
  XOR U59369 ( .A(n49887), .B(n49888), .Z(n49900) );
  XOR U59370 ( .A(n49898), .B(n49900), .Z(n49902) );
  XOR U59371 ( .A(n46487), .B(n49902), .Z(n48798) );
  XOR U59372 ( .A(n46488), .B(n48798), .Z(n48795) );
  IV U59373 ( .A(n46489), .Z(n46490) );
  NOR U59374 ( .A(n46491), .B(n46490), .Z(n48794) );
  IV U59375 ( .A(n46492), .Z(n46494) );
  NOR U59376 ( .A(n46494), .B(n46493), .Z(n48792) );
  NOR U59377 ( .A(n48794), .B(n48792), .Z(n46495) );
  XOR U59378 ( .A(n48795), .B(n46495), .Z(n46496) );
  NOR U59379 ( .A(n46497), .B(n46496), .Z(n46500) );
  XOR U59380 ( .A(n48794), .B(n48795), .Z(n46499) );
  IV U59381 ( .A(n46497), .Z(n46498) );
  NOR U59382 ( .A(n46499), .B(n46498), .Z(n52570) );
  NOR U59383 ( .A(n46500), .B(n52570), .Z(n48789) );
  XOR U59384 ( .A(n48791), .B(n48789), .Z(n49921) );
  IV U59385 ( .A(n46501), .Z(n46502) );
  NOR U59386 ( .A(n46503), .B(n46502), .Z(n49919) );
  XOR U59387 ( .A(n49921), .B(n49919), .Z(n49924) );
  IV U59388 ( .A(n46504), .Z(n46505) );
  NOR U59389 ( .A(n46505), .B(n46507), .Z(n49922) );
  XOR U59390 ( .A(n49924), .B(n49922), .Z(n48786) );
  IV U59391 ( .A(n46506), .Z(n46508) );
  NOR U59392 ( .A(n46508), .B(n46507), .Z(n48784) );
  XOR U59393 ( .A(n48786), .B(n48784), .Z(n48782) );
  XOR U59394 ( .A(n48783), .B(n48782), .Z(n46509) );
  XOR U59395 ( .A(n46510), .B(n46509), .Z(n49929) );
  IV U59396 ( .A(n46511), .Z(n46513) );
  NOR U59397 ( .A(n46513), .B(n46512), .Z(n49927) );
  XOR U59398 ( .A(n49929), .B(n49927), .Z(n49932) );
  XOR U59399 ( .A(n49930), .B(n49932), .Z(n49937) );
  XOR U59400 ( .A(n49934), .B(n49937), .Z(n46514) );
  NOR U59401 ( .A(n46515), .B(n46514), .Z(n53842) );
  IV U59402 ( .A(n46516), .Z(n46518) );
  NOR U59403 ( .A(n46518), .B(n46517), .Z(n49936) );
  NOR U59404 ( .A(n49934), .B(n49936), .Z(n46519) );
  XOR U59405 ( .A(n46519), .B(n49937), .Z(n49942) );
  NOR U59406 ( .A(n46520), .B(n49942), .Z(n46521) );
  NOR U59407 ( .A(n53842), .B(n46521), .Z(n49945) );
  NOR U59408 ( .A(n46523), .B(n46522), .Z(n49941) );
  IV U59409 ( .A(n46524), .Z(n46526) );
  IV U59410 ( .A(n46525), .Z(n46532) );
  NOR U59411 ( .A(n46526), .B(n46532), .Z(n49946) );
  NOR U59412 ( .A(n49941), .B(n49946), .Z(n46527) );
  XOR U59413 ( .A(n49945), .B(n46527), .Z(n53850) );
  IV U59414 ( .A(n46528), .Z(n46529) );
  NOR U59415 ( .A(n46530), .B(n46529), .Z(n53849) );
  IV U59416 ( .A(n46531), .Z(n46533) );
  NOR U59417 ( .A(n46533), .B(n46532), .Z(n53854) );
  NOR U59418 ( .A(n53849), .B(n53854), .Z(n48777) );
  XOR U59419 ( .A(n53850), .B(n48777), .Z(n49953) );
  XOR U59420 ( .A(n49954), .B(n49953), .Z(n49965) );
  IV U59421 ( .A(n46534), .Z(n46536) );
  NOR U59422 ( .A(n46536), .B(n46535), .Z(n49964) );
  NOR U59423 ( .A(n49952), .B(n49964), .Z(n53871) );
  XOR U59424 ( .A(n49965), .B(n53871), .Z(n49961) );
  XOR U59425 ( .A(n49960), .B(n49961), .Z(n52535) );
  XOR U59426 ( .A(n48775), .B(n52535), .Z(n48768) );
  NOR U59427 ( .A(n46537), .B(n48772), .Z(n46541) );
  IV U59428 ( .A(n46538), .Z(n46540) );
  NOR U59429 ( .A(n46540), .B(n46539), .Z(n48767) );
  NOR U59430 ( .A(n46541), .B(n48767), .Z(n46542) );
  XOR U59431 ( .A(n48768), .B(n46542), .Z(n49982) );
  XOR U59432 ( .A(n48765), .B(n49982), .Z(n46543) );
  XOR U59433 ( .A(n46544), .B(n46543), .Z(n48750) );
  XOR U59434 ( .A(n46545), .B(n48750), .Z(n48745) );
  XOR U59435 ( .A(n46546), .B(n48745), .Z(n48741) );
  IV U59436 ( .A(n46547), .Z(n46549) );
  NOR U59437 ( .A(n46549), .B(n46548), .Z(n46550) );
  IV U59438 ( .A(n46550), .Z(n48740) );
  XOR U59439 ( .A(n48741), .B(n48740), .Z(n46551) );
  XOR U59440 ( .A(n46552), .B(n46551), .Z(n48728) );
  IV U59441 ( .A(n46553), .Z(n46560) );
  IV U59442 ( .A(n46554), .Z(n46562) );
  NOR U59443 ( .A(n46555), .B(n46562), .Z(n46556) );
  IV U59444 ( .A(n46556), .Z(n46557) );
  NOR U59445 ( .A(n46558), .B(n46557), .Z(n46559) );
  IV U59446 ( .A(n46559), .Z(n46565) );
  NOR U59447 ( .A(n46560), .B(n46565), .Z(n48719) );
  IV U59448 ( .A(n46561), .Z(n46563) );
  NOR U59449 ( .A(n46563), .B(n46562), .Z(n48727) );
  IV U59450 ( .A(n46564), .Z(n46566) );
  NOR U59451 ( .A(n46566), .B(n46565), .Z(n48729) );
  XOR U59452 ( .A(n48727), .B(n48729), .Z(n46567) );
  NOR U59453 ( .A(n48719), .B(n46567), .Z(n46568) );
  XOR U59454 ( .A(n48728), .B(n46568), .Z(n48722) );
  XOR U59455 ( .A(n48721), .B(n48722), .Z(n49988) );
  IV U59456 ( .A(n46569), .Z(n46571) );
  NOR U59457 ( .A(n46571), .B(n46570), .Z(n49985) );
  NOR U59458 ( .A(n49992), .B(n49990), .Z(n46572) );
  NOR U59459 ( .A(n49985), .B(n46572), .Z(n46573) );
  XOR U59460 ( .A(n49988), .B(n46573), .Z(n49998) );
  XOR U59461 ( .A(n49994), .B(n49998), .Z(n46578) );
  IV U59462 ( .A(n46574), .Z(n46576) );
  IV U59463 ( .A(n46575), .Z(n46586) );
  NOR U59464 ( .A(n46576), .B(n46586), .Z(n46583) );
  IV U59465 ( .A(n46583), .Z(n46577) );
  NOR U59466 ( .A(n46578), .B(n46577), .Z(n50008) );
  NOR U59467 ( .A(n46580), .B(n46579), .Z(n49996) );
  NOR U59468 ( .A(n49994), .B(n49996), .Z(n46581) );
  XOR U59469 ( .A(n49998), .B(n46581), .Z(n46582) );
  NOR U59470 ( .A(n46583), .B(n46582), .Z(n46584) );
  NOR U59471 ( .A(n50008), .B(n46584), .Z(n50000) );
  IV U59472 ( .A(n46585), .Z(n46589) );
  NOR U59473 ( .A(n46587), .B(n46586), .Z(n46588) );
  IV U59474 ( .A(n46588), .Z(n46594) );
  NOR U59475 ( .A(n46589), .B(n46594), .Z(n50001) );
  XOR U59476 ( .A(n50000), .B(n50001), .Z(n50012) );
  IV U59477 ( .A(n46590), .Z(n46591) );
  NOR U59478 ( .A(n46592), .B(n46591), .Z(n50023) );
  IV U59479 ( .A(n46593), .Z(n46595) );
  NOR U59480 ( .A(n46595), .B(n46594), .Z(n50013) );
  NOR U59481 ( .A(n50023), .B(n50013), .Z(n46596) );
  XOR U59482 ( .A(n50012), .B(n46596), .Z(n50045) );
  IV U59483 ( .A(n46597), .Z(n46598) );
  NOR U59484 ( .A(n46598), .B(n48714), .Z(n50020) );
  XOR U59485 ( .A(n50045), .B(n50020), .Z(n50038) );
  XOR U59486 ( .A(n46599), .B(n50038), .Z(n50055) );
  XOR U59487 ( .A(n50053), .B(n50055), .Z(n50057) );
  XOR U59488 ( .A(n48706), .B(n50057), .Z(n48700) );
  NOR U59489 ( .A(n46601), .B(n46600), .Z(n48703) );
  IV U59490 ( .A(n46602), .Z(n46604) );
  IV U59491 ( .A(n46603), .Z(n46608) );
  NOR U59492 ( .A(n46604), .B(n46608), .Z(n48701) );
  NOR U59493 ( .A(n48703), .B(n48701), .Z(n46605) );
  XOR U59494 ( .A(n48700), .B(n46605), .Z(n50064) );
  IV U59495 ( .A(n46606), .Z(n46607) );
  NOR U59496 ( .A(n46608), .B(n46607), .Z(n48698) );
  XOR U59497 ( .A(n50064), .B(n48698), .Z(n48696) );
  XOR U59498 ( .A(n46609), .B(n48696), .Z(n50067) );
  XOR U59499 ( .A(n50065), .B(n50067), .Z(n50069) );
  XOR U59500 ( .A(n50068), .B(n50069), .Z(n48690) );
  XOR U59501 ( .A(n48691), .B(n48690), .Z(n48687) );
  IV U59502 ( .A(n46610), .Z(n46612) );
  NOR U59503 ( .A(n46612), .B(n46611), .Z(n48692) );
  IV U59504 ( .A(n46613), .Z(n46614) );
  NOR U59505 ( .A(n46615), .B(n46614), .Z(n48686) );
  NOR U59506 ( .A(n48692), .B(n48686), .Z(n46616) );
  XOR U59507 ( .A(n48687), .B(n46616), .Z(n50077) );
  XOR U59508 ( .A(n50074), .B(n50077), .Z(n50085) );
  XOR U59509 ( .A(n46617), .B(n50085), .Z(n50083) );
  XOR U59510 ( .A(n50082), .B(n50083), .Z(n48679) );
  IV U59511 ( .A(n46618), .Z(n46619) );
  NOR U59512 ( .A(n46620), .B(n46619), .Z(n48683) );
  IV U59513 ( .A(n46621), .Z(n46622) );
  NOR U59514 ( .A(n46626), .B(n46622), .Z(n48680) );
  NOR U59515 ( .A(n48683), .B(n48680), .Z(n46623) );
  XOR U59516 ( .A(n48679), .B(n46623), .Z(n48673) );
  IV U59517 ( .A(n46624), .Z(n46625) );
  NOR U59518 ( .A(n46626), .B(n46625), .Z(n48671) );
  XOR U59519 ( .A(n48673), .B(n48671), .Z(n48676) );
  XOR U59520 ( .A(n48674), .B(n48676), .Z(n50092) );
  XOR U59521 ( .A(n50090), .B(n50092), .Z(n46635) );
  IV U59522 ( .A(n46627), .Z(n46629) );
  NOR U59523 ( .A(n46629), .B(n46628), .Z(n46630) );
  IV U59524 ( .A(n46630), .Z(n46637) );
  NOR U59525 ( .A(n46635), .B(n46637), .Z(n50102) );
  IV U59526 ( .A(n46631), .Z(n46632) );
  NOR U59527 ( .A(n48665), .B(n46632), .Z(n48661) );
  IV U59528 ( .A(n46633), .Z(n46634) );
  NOR U59529 ( .A(n46634), .B(n48665), .Z(n46636) );
  XOR U59530 ( .A(n46636), .B(n46635), .Z(n48662) );
  IV U59531 ( .A(n48662), .Z(n46638) );
  XOR U59532 ( .A(n48661), .B(n46638), .Z(n46640) );
  NOR U59533 ( .A(n46638), .B(n46637), .Z(n46639) );
  NOR U59534 ( .A(n46640), .B(n46639), .Z(n46641) );
  NOR U59535 ( .A(n50102), .B(n46641), .Z(n48655) );
  XOR U59536 ( .A(n48657), .B(n48655), .Z(n48658) );
  IV U59537 ( .A(n46642), .Z(n46643) );
  NOR U59538 ( .A(n46644), .B(n46643), .Z(n46649) );
  IV U59539 ( .A(n46645), .Z(n46647) );
  NOR U59540 ( .A(n46647), .B(n46646), .Z(n46648) );
  NOR U59541 ( .A(n46649), .B(n46648), .Z(n48659) );
  XOR U59542 ( .A(n48658), .B(n48659), .Z(n48653) );
  XOR U59543 ( .A(n46650), .B(n48653), .Z(n50106) );
  XOR U59544 ( .A(n50104), .B(n50106), .Z(n50113) );
  IV U59545 ( .A(n46651), .Z(n46652) );
  NOR U59546 ( .A(n46653), .B(n46652), .Z(n50111) );
  XOR U59547 ( .A(n50113), .B(n50111), .Z(n50115) );
  XOR U59548 ( .A(n50114), .B(n50115), .Z(n50124) );
  IV U59549 ( .A(n46654), .Z(n46655) );
  NOR U59550 ( .A(n46656), .B(n46655), .Z(n48649) );
  IV U59551 ( .A(n46657), .Z(n46659) );
  NOR U59552 ( .A(n46659), .B(n46658), .Z(n50122) );
  NOR U59553 ( .A(n48649), .B(n50122), .Z(n46660) );
  XOR U59554 ( .A(n50124), .B(n46660), .Z(n46671) );
  IV U59555 ( .A(n46671), .Z(n50121) );
  IV U59556 ( .A(n46661), .Z(n46662) );
  NOR U59557 ( .A(n46663), .B(n46662), .Z(n46664) );
  IV U59558 ( .A(n46664), .Z(n46672) );
  NOR U59559 ( .A(n50121), .B(n46672), .Z(n52411) );
  IV U59560 ( .A(n46665), .Z(n46666) );
  NOR U59561 ( .A(n46667), .B(n46666), .Z(n48641) );
  IV U59562 ( .A(n46668), .Z(n46670) );
  NOR U59563 ( .A(n46670), .B(n46669), .Z(n50119) );
  XOR U59564 ( .A(n50119), .B(n46671), .Z(n48642) );
  XOR U59565 ( .A(n48641), .B(n48642), .Z(n46674) );
  NOR U59566 ( .A(n48642), .B(n46672), .Z(n46673) );
  NOR U59567 ( .A(n46674), .B(n46673), .Z(n46675) );
  NOR U59568 ( .A(n52411), .B(n46675), .Z(n48645) );
  IV U59569 ( .A(n46676), .Z(n46678) );
  NOR U59570 ( .A(n46678), .B(n46677), .Z(n52402) );
  IV U59571 ( .A(n46679), .Z(n46680) );
  NOR U59572 ( .A(n46681), .B(n46680), .Z(n54001) );
  NOR U59573 ( .A(n52402), .B(n54001), .Z(n48646) );
  XOR U59574 ( .A(n48645), .B(n48646), .Z(n50132) );
  XOR U59575 ( .A(n46682), .B(n50132), .Z(n50135) );
  XOR U59576 ( .A(n46683), .B(n50135), .Z(n48631) );
  XOR U59577 ( .A(n46684), .B(n48631), .Z(n50138) );
  XOR U59578 ( .A(n46685), .B(n50138), .Z(n50141) );
  IV U59579 ( .A(n46686), .Z(n46687) );
  NOR U59580 ( .A(n46688), .B(n46687), .Z(n50140) );
  IV U59581 ( .A(n46689), .Z(n46691) );
  NOR U59582 ( .A(n46691), .B(n46690), .Z(n46692) );
  NOR U59583 ( .A(n50140), .B(n46692), .Z(n50150) );
  XOR U59584 ( .A(n50141), .B(n50150), .Z(n50152) );
  XOR U59585 ( .A(n46693), .B(n50152), .Z(n48626) );
  IV U59586 ( .A(n46694), .Z(n46696) );
  NOR U59587 ( .A(n46696), .B(n46695), .Z(n46703) );
  IV U59588 ( .A(n46703), .Z(n46697) );
  NOR U59589 ( .A(n48626), .B(n46697), .Z(n52389) );
  NOR U59590 ( .A(n46706), .B(n52389), .Z(n46698) );
  IV U59591 ( .A(n46698), .Z(n46705) );
  IV U59592 ( .A(n46699), .Z(n46700) );
  NOR U59593 ( .A(n46701), .B(n46700), .Z(n46702) );
  IV U59594 ( .A(n46702), .Z(n48625) );
  XOR U59595 ( .A(n48625), .B(n48626), .Z(n48620) );
  NOR U59596 ( .A(n46703), .B(n48620), .Z(n46704) );
  NOR U59597 ( .A(n46705), .B(n46704), .Z(n46709) );
  IV U59598 ( .A(n46706), .Z(n46707) );
  NOR U59599 ( .A(n48620), .B(n46707), .Z(n46708) );
  NOR U59600 ( .A(n46709), .B(n46708), .Z(n48614) );
  XOR U59601 ( .A(n48612), .B(n48614), .Z(n48616) );
  XOR U59602 ( .A(n48615), .B(n48616), .Z(n50167) );
  XOR U59603 ( .A(n46710), .B(n50167), .Z(n48606) );
  XOR U59604 ( .A(n46711), .B(n48606), .Z(n50169) );
  XOR U59605 ( .A(n46712), .B(n50169), .Z(n48600) );
  XOR U59606 ( .A(n48598), .B(n48600), .Z(n50174) );
  XOR U59607 ( .A(n46713), .B(n50174), .Z(n52357) );
  XOR U59608 ( .A(n50179), .B(n52357), .Z(n48591) );
  IV U59609 ( .A(n46714), .Z(n46716) );
  NOR U59610 ( .A(n46716), .B(n46715), .Z(n50180) );
  NOR U59611 ( .A(n46718), .B(n46717), .Z(n48590) );
  NOR U59612 ( .A(n50180), .B(n48590), .Z(n46719) );
  XOR U59613 ( .A(n48591), .B(n46719), .Z(n48589) );
  IV U59614 ( .A(n46720), .Z(n46722) );
  NOR U59615 ( .A(n46722), .B(n46721), .Z(n48587) );
  XOR U59616 ( .A(n48589), .B(n48587), .Z(n48595) );
  XOR U59617 ( .A(n48594), .B(n48595), .Z(n50191) );
  XOR U59618 ( .A(n46723), .B(n50191), .Z(n50195) );
  XOR U59619 ( .A(n50193), .B(n50195), .Z(n50198) );
  IV U59620 ( .A(n46724), .Z(n46726) );
  NOR U59621 ( .A(n46726), .B(n46725), .Z(n50196) );
  XOR U59622 ( .A(n50198), .B(n50196), .Z(n48583) );
  IV U59623 ( .A(n46727), .Z(n46728) );
  NOR U59624 ( .A(n46729), .B(n46728), .Z(n48585) );
  IV U59625 ( .A(n46730), .Z(n46731) );
  NOR U59626 ( .A(n46732), .B(n46731), .Z(n48582) );
  NOR U59627 ( .A(n48585), .B(n48582), .Z(n46733) );
  XOR U59628 ( .A(n48583), .B(n46733), .Z(n48576) );
  IV U59629 ( .A(n46734), .Z(n46735) );
  NOR U59630 ( .A(n46736), .B(n46735), .Z(n48579) );
  IV U59631 ( .A(n46737), .Z(n46738) );
  NOR U59632 ( .A(n46739), .B(n46738), .Z(n48577) );
  NOR U59633 ( .A(n48579), .B(n48577), .Z(n46740) );
  XOR U59634 ( .A(n48576), .B(n46740), .Z(n50202) );
  XOR U59635 ( .A(n50203), .B(n50202), .Z(n50205) );
  NOR U59636 ( .A(n46742), .B(n46741), .Z(n48574) );
  IV U59637 ( .A(n46743), .Z(n46749) );
  IV U59638 ( .A(n46744), .Z(n46745) );
  NOR U59639 ( .A(n46749), .B(n46745), .Z(n50204) );
  NOR U59640 ( .A(n48574), .B(n50204), .Z(n46746) );
  XOR U59641 ( .A(n50205), .B(n46746), .Z(n48573) );
  IV U59642 ( .A(n46747), .Z(n46748) );
  NOR U59643 ( .A(n46749), .B(n46748), .Z(n48571) );
  XOR U59644 ( .A(n48573), .B(n48571), .Z(n46750) );
  NOR U59645 ( .A(n46751), .B(n46750), .Z(n52307) );
  IV U59646 ( .A(n46752), .Z(n46753) );
  NOR U59647 ( .A(n46754), .B(n46753), .Z(n48565) );
  NOR U59648 ( .A(n48565), .B(n48571), .Z(n46755) );
  XOR U59649 ( .A(n48573), .B(n46755), .Z(n48562) );
  NOR U59650 ( .A(n46756), .B(n48562), .Z(n46757) );
  NOR U59651 ( .A(n52307), .B(n46757), .Z(n48568) );
  XOR U59652 ( .A(n48570), .B(n48568), .Z(n48560) );
  NOR U59653 ( .A(n46759), .B(n46758), .Z(n48561) );
  IV U59654 ( .A(n46760), .Z(n46762) );
  IV U59655 ( .A(n46761), .Z(n46769) );
  NOR U59656 ( .A(n46762), .B(n46769), .Z(n48558) );
  NOR U59657 ( .A(n48561), .B(n48558), .Z(n46763) );
  XOR U59658 ( .A(n48560), .B(n46763), .Z(n48551) );
  IV U59659 ( .A(n46764), .Z(n46765) );
  NOR U59660 ( .A(n46766), .B(n46765), .Z(n48552) );
  IV U59661 ( .A(n46767), .Z(n46768) );
  NOR U59662 ( .A(n46769), .B(n46768), .Z(n48555) );
  NOR U59663 ( .A(n48552), .B(n48555), .Z(n46770) );
  XOR U59664 ( .A(n48551), .B(n46770), .Z(n50217) );
  XOR U59665 ( .A(n46771), .B(n50217), .Z(n50224) );
  IV U59666 ( .A(n46772), .Z(n46773) );
  NOR U59667 ( .A(n46774), .B(n46773), .Z(n50216) );
  IV U59668 ( .A(n46775), .Z(n46776) );
  NOR U59669 ( .A(n46777), .B(n46776), .Z(n50223) );
  NOR U59670 ( .A(n50216), .B(n50223), .Z(n46778) );
  XOR U59671 ( .A(n50224), .B(n46778), .Z(n46779) );
  IV U59672 ( .A(n46779), .Z(n50222) );
  XOR U59673 ( .A(n50220), .B(n50222), .Z(n48541) );
  XOR U59674 ( .A(n46780), .B(n48541), .Z(n48535) );
  XOR U59675 ( .A(n48534), .B(n48535), .Z(n48529) );
  IV U59676 ( .A(n46781), .Z(n46782) );
  NOR U59677 ( .A(n46783), .B(n46782), .Z(n48532) );
  NOR U59678 ( .A(n46785), .B(n46784), .Z(n48528) );
  NOR U59679 ( .A(n48532), .B(n48528), .Z(n46786) );
  XOR U59680 ( .A(n48529), .B(n46786), .Z(n48527) );
  IV U59681 ( .A(n46787), .Z(n46788) );
  NOR U59682 ( .A(n46789), .B(n46788), .Z(n48525) );
  XOR U59683 ( .A(n48527), .B(n48525), .Z(n48521) );
  XOR U59684 ( .A(n48519), .B(n48521), .Z(n48517) );
  XOR U59685 ( .A(n48516), .B(n48517), .Z(n48512) );
  IV U59686 ( .A(n46790), .Z(n46791) );
  NOR U59687 ( .A(n46792), .B(n46791), .Z(n48514) );
  IV U59688 ( .A(n46793), .Z(n46795) );
  NOR U59689 ( .A(n46795), .B(n46794), .Z(n48511) );
  NOR U59690 ( .A(n48514), .B(n48511), .Z(n46796) );
  XOR U59691 ( .A(n48512), .B(n46796), .Z(n48501) );
  XOR U59692 ( .A(n48502), .B(n48501), .Z(n48505) );
  IV U59693 ( .A(n46797), .Z(n46799) );
  NOR U59694 ( .A(n46799), .B(n46798), .Z(n46800) );
  IV U59695 ( .A(n46800), .Z(n48504) );
  XOR U59696 ( .A(n48505), .B(n48504), .Z(n50232) );
  IV U59697 ( .A(n46801), .Z(n48498) );
  NOR U59698 ( .A(n46802), .B(n48498), .Z(n46806) );
  IV U59699 ( .A(n46803), .Z(n46805) );
  NOR U59700 ( .A(n46805), .B(n46804), .Z(n50231) );
  NOR U59701 ( .A(n46806), .B(n50231), .Z(n46807) );
  XOR U59702 ( .A(n50232), .B(n46807), .Z(n50239) );
  XOR U59703 ( .A(n50235), .B(n50239), .Z(n48496) );
  XOR U59704 ( .A(n46808), .B(n48496), .Z(n48493) );
  XOR U59705 ( .A(n48492), .B(n48493), .Z(n48484) );
  IV U59706 ( .A(n46809), .Z(n46810) );
  NOR U59707 ( .A(n46811), .B(n46810), .Z(n48490) );
  IV U59708 ( .A(n46812), .Z(n46814) );
  NOR U59709 ( .A(n46814), .B(n46813), .Z(n48485) );
  NOR U59710 ( .A(n48490), .B(n48485), .Z(n46815) );
  XOR U59711 ( .A(n48484), .B(n46815), .Z(n48483) );
  IV U59712 ( .A(n46816), .Z(n46818) );
  NOR U59713 ( .A(n46818), .B(n46817), .Z(n48481) );
  XOR U59714 ( .A(n48483), .B(n48481), .Z(n50243) );
  XOR U59715 ( .A(n50242), .B(n50243), .Z(n50246) );
  XOR U59716 ( .A(n50245), .B(n50246), .Z(n48476) );
  XOR U59717 ( .A(n48475), .B(n48476), .Z(n50251) );
  XOR U59718 ( .A(n48478), .B(n50251), .Z(n48474) );
  XOR U59719 ( .A(n48472), .B(n48474), .Z(n48470) );
  XOR U59720 ( .A(n46819), .B(n48470), .Z(n48466) );
  XOR U59721 ( .A(n46820), .B(n48466), .Z(n50254) );
  XOR U59722 ( .A(n50253), .B(n50254), .Z(n52201) );
  XOR U59723 ( .A(n46821), .B(n52201), .Z(n52193) );
  XOR U59724 ( .A(n48462), .B(n52193), .Z(n46831) );
  IV U59725 ( .A(n46822), .Z(n46823) );
  NOR U59726 ( .A(n46824), .B(n46823), .Z(n46834) );
  IV U59727 ( .A(n46825), .Z(n46827) );
  NOR U59728 ( .A(n46827), .B(n46826), .Z(n46830) );
  NOR U59729 ( .A(n46834), .B(n46830), .Z(n46828) );
  IV U59730 ( .A(n46828), .Z(n46829) );
  NOR U59731 ( .A(n46831), .B(n46829), .Z(n46837) );
  IV U59732 ( .A(n46830), .Z(n46833) );
  IV U59733 ( .A(n46831), .Z(n46832) );
  NOR U59734 ( .A(n46833), .B(n46832), .Z(n52187) );
  IV U59735 ( .A(n46834), .Z(n46835) );
  NOR U59736 ( .A(n46835), .B(n52193), .Z(n52189) );
  NOR U59737 ( .A(n52187), .B(n52189), .Z(n46836) );
  IV U59738 ( .A(n46836), .Z(n48464) );
  NOR U59739 ( .A(n46837), .B(n48464), .Z(n48456) );
  IV U59740 ( .A(n46838), .Z(n46839) );
  NOR U59741 ( .A(n46840), .B(n46839), .Z(n46841) );
  IV U59742 ( .A(n46841), .Z(n48458) );
  XOR U59743 ( .A(n48456), .B(n48458), .Z(n48461) );
  XOR U59744 ( .A(n48459), .B(n48461), .Z(n50266) );
  XOR U59745 ( .A(n50264), .B(n50266), .Z(n50268) );
  XOR U59746 ( .A(n50267), .B(n50268), .Z(n48454) );
  XOR U59747 ( .A(n48453), .B(n48454), .Z(n50278) );
  XOR U59748 ( .A(n50276), .B(n50278), .Z(n50282) );
  XOR U59749 ( .A(n50279), .B(n50282), .Z(n46842) );
  NOR U59750 ( .A(n46843), .B(n46842), .Z(n52169) );
  IV U59751 ( .A(n46844), .Z(n46845) );
  NOR U59752 ( .A(n46846), .B(n46845), .Z(n50281) );
  NOR U59753 ( .A(n50281), .B(n50279), .Z(n46847) );
  XOR U59754 ( .A(n46847), .B(n50282), .Z(n48445) );
  NOR U59755 ( .A(n46848), .B(n48445), .Z(n46849) );
  NOR U59756 ( .A(n52169), .B(n46849), .Z(n48436) );
  NOR U59757 ( .A(n46850), .B(n48447), .Z(n46854) );
  IV U59758 ( .A(n46851), .Z(n48438) );
  NOR U59759 ( .A(n46852), .B(n48438), .Z(n46853) );
  NOR U59760 ( .A(n46854), .B(n46853), .Z(n46855) );
  XOR U59761 ( .A(n48436), .B(n46855), .Z(n48432) );
  IV U59762 ( .A(n46856), .Z(n46858) );
  NOR U59763 ( .A(n46858), .B(n46857), .Z(n48428) );
  IV U59764 ( .A(n46859), .Z(n46861) );
  NOR U59765 ( .A(n46861), .B(n46860), .Z(n48430) );
  NOR U59766 ( .A(n48428), .B(n48430), .Z(n46862) );
  XOR U59767 ( .A(n48432), .B(n46862), .Z(n46863) );
  NOR U59768 ( .A(n46864), .B(n46863), .Z(n46867) );
  IV U59769 ( .A(n46864), .Z(n46866) );
  XOR U59770 ( .A(n48428), .B(n48432), .Z(n46865) );
  NOR U59771 ( .A(n46866), .B(n46865), .Z(n52149) );
  NOR U59772 ( .A(n46867), .B(n52149), .Z(n50289) );
  IV U59773 ( .A(n46868), .Z(n46870) );
  NOR U59774 ( .A(n46870), .B(n46869), .Z(n46871) );
  IV U59775 ( .A(n46871), .Z(n50290) );
  XOR U59776 ( .A(n50289), .B(n50290), .Z(n48422) );
  XOR U59777 ( .A(n46872), .B(n48422), .Z(n48412) );
  IV U59778 ( .A(n46873), .Z(n46874) );
  NOR U59779 ( .A(n46875), .B(n46874), .Z(n48415) );
  IV U59780 ( .A(n46876), .Z(n46877) );
  NOR U59781 ( .A(n46878), .B(n46877), .Z(n48413) );
  NOR U59782 ( .A(n48415), .B(n48413), .Z(n46879) );
  XOR U59783 ( .A(n48412), .B(n46879), .Z(n50302) );
  XOR U59784 ( .A(n50293), .B(n50302), .Z(n50297) );
  XOR U59785 ( .A(n50295), .B(n50297), .Z(n46886) );
  NOR U59786 ( .A(n46890), .B(n46886), .Z(n50315) );
  IV U59787 ( .A(n46880), .Z(n46882) );
  NOR U59788 ( .A(n46882), .B(n46881), .Z(n48402) );
  IV U59789 ( .A(n46883), .Z(n50303) );
  NOR U59790 ( .A(n50303), .B(n46884), .Z(n46888) );
  IV U59791 ( .A(n46888), .Z(n46885) );
  NOR U59792 ( .A(n46885), .B(n50302), .Z(n48409) );
  IV U59793 ( .A(n46886), .Z(n46887) );
  NOR U59794 ( .A(n46888), .B(n46887), .Z(n46889) );
  NOR U59795 ( .A(n48409), .B(n46889), .Z(n48403) );
  XOR U59796 ( .A(n48402), .B(n48403), .Z(n46892) );
  NOR U59797 ( .A(n48403), .B(n46890), .Z(n46891) );
  NOR U59798 ( .A(n46892), .B(n46891), .Z(n46893) );
  NOR U59799 ( .A(n50315), .B(n46893), .Z(n46894) );
  IV U59800 ( .A(n46894), .Z(n54197) );
  XOR U59801 ( .A(n46895), .B(n54197), .Z(n48397) );
  IV U59802 ( .A(n46896), .Z(n46898) );
  NOR U59803 ( .A(n46898), .B(n46897), .Z(n48396) );
  NOR U59804 ( .A(n46899), .B(n48396), .Z(n46900) );
  XOR U59805 ( .A(n48397), .B(n46900), .Z(n50321) );
  XOR U59806 ( .A(n50317), .B(n50321), .Z(n46905) );
  IV U59807 ( .A(n46901), .Z(n46914) );
  IV U59808 ( .A(n46902), .Z(n46903) );
  NOR U59809 ( .A(n46914), .B(n46903), .Z(n46910) );
  IV U59810 ( .A(n46910), .Z(n46904) );
  NOR U59811 ( .A(n46905), .B(n46904), .Z(n52122) );
  NOR U59812 ( .A(n46907), .B(n46906), .Z(n50319) );
  NOR U59813 ( .A(n50317), .B(n50319), .Z(n46908) );
  XOR U59814 ( .A(n50321), .B(n46908), .Z(n46909) );
  NOR U59815 ( .A(n46910), .B(n46909), .Z(n46911) );
  NOR U59816 ( .A(n52122), .B(n46911), .Z(n46912) );
  IV U59817 ( .A(n46912), .Z(n50325) );
  IV U59818 ( .A(n46913), .Z(n46915) );
  NOR U59819 ( .A(n46915), .B(n46914), .Z(n50323) );
  XOR U59820 ( .A(n50325), .B(n50323), .Z(n48395) );
  IV U59821 ( .A(n48395), .Z(n46922) );
  IV U59822 ( .A(n46916), .Z(n46917) );
  NOR U59823 ( .A(n46920), .B(n46917), .Z(n48390) );
  IV U59824 ( .A(n46918), .Z(n46919) );
  NOR U59825 ( .A(n46920), .B(n46919), .Z(n48393) );
  NOR U59826 ( .A(n48390), .B(n48393), .Z(n46921) );
  XOR U59827 ( .A(n46922), .B(n46921), .Z(n50332) );
  XOR U59828 ( .A(n50330), .B(n50332), .Z(n50327) );
  XOR U59829 ( .A(n50328), .B(n50327), .Z(n48384) );
  IV U59830 ( .A(n46923), .Z(n46927) );
  IV U59831 ( .A(n46924), .Z(n48386) );
  NOR U59832 ( .A(n46925), .B(n48386), .Z(n46926) );
  IV U59833 ( .A(n46926), .Z(n46943) );
  NOR U59834 ( .A(n46927), .B(n46943), .Z(n46936) );
  IV U59835 ( .A(n46936), .Z(n46928) );
  NOR U59836 ( .A(n48384), .B(n46928), .Z(n46938) );
  NOR U59837 ( .A(n46930), .B(n46929), .Z(n46932) );
  IV U59838 ( .A(n46932), .Z(n46931) );
  NOR U59839 ( .A(n46931), .B(n50327), .Z(n52103) );
  NOR U59840 ( .A(n48384), .B(n46932), .Z(n46933) );
  NOR U59841 ( .A(n52103), .B(n46933), .Z(n46934) );
  IV U59842 ( .A(n46934), .Z(n46935) );
  NOR U59843 ( .A(n46936), .B(n46935), .Z(n46937) );
  NOR U59844 ( .A(n46938), .B(n46937), .Z(n48381) );
  IV U59845 ( .A(n46939), .Z(n46940) );
  NOR U59846 ( .A(n48386), .B(n46940), .Z(n48380) );
  IV U59847 ( .A(n46941), .Z(n46942) );
  NOR U59848 ( .A(n46943), .B(n46942), .Z(n46944) );
  NOR U59849 ( .A(n48380), .B(n46944), .Z(n46945) );
  XOR U59850 ( .A(n48381), .B(n46945), .Z(n48372) );
  IV U59851 ( .A(n46946), .Z(n46947) );
  NOR U59852 ( .A(n46950), .B(n46947), .Z(n48375) );
  IV U59853 ( .A(n46948), .Z(n46949) );
  NOR U59854 ( .A(n46950), .B(n46949), .Z(n48377) );
  NOR U59855 ( .A(n48377), .B(n48373), .Z(n46951) );
  IV U59856 ( .A(n46951), .Z(n46952) );
  NOR U59857 ( .A(n48375), .B(n46952), .Z(n46953) );
  XOR U59858 ( .A(n48372), .B(n46953), .Z(n48369) );
  IV U59859 ( .A(n46954), .Z(n46957) );
  IV U59860 ( .A(n46955), .Z(n46956) );
  NOR U59861 ( .A(n46957), .B(n46956), .Z(n48367) );
  XOR U59862 ( .A(n48369), .B(n48367), .Z(n48366) );
  IV U59863 ( .A(n46958), .Z(n46961) );
  IV U59864 ( .A(n46959), .Z(n46960) );
  NOR U59865 ( .A(n46961), .B(n46960), .Z(n48364) );
  XOR U59866 ( .A(n48366), .B(n48364), .Z(n48357) );
  IV U59867 ( .A(n46962), .Z(n46963) );
  NOR U59868 ( .A(n46964), .B(n46963), .Z(n48362) );
  IV U59869 ( .A(n46965), .Z(n46967) );
  NOR U59870 ( .A(n46967), .B(n46966), .Z(n48356) );
  NOR U59871 ( .A(n48362), .B(n48356), .Z(n46968) );
  XOR U59872 ( .A(n48357), .B(n46968), .Z(n48352) );
  IV U59873 ( .A(n46969), .Z(n46971) );
  NOR U59874 ( .A(n46971), .B(n46970), .Z(n48359) );
  IV U59875 ( .A(n46972), .Z(n46974) );
  NOR U59876 ( .A(n46974), .B(n46973), .Z(n48351) );
  NOR U59877 ( .A(n48359), .B(n48351), .Z(n46975) );
  XOR U59878 ( .A(n48352), .B(n46975), .Z(n50345) );
  IV U59879 ( .A(n46976), .Z(n46977) );
  NOR U59880 ( .A(n46978), .B(n46977), .Z(n48349) );
  IV U59881 ( .A(n46979), .Z(n46981) );
  NOR U59882 ( .A(n46981), .B(n46980), .Z(n50344) );
  NOR U59883 ( .A(n48349), .B(n50344), .Z(n46982) );
  XOR U59884 ( .A(n50345), .B(n46982), .Z(n48347) );
  XOR U59885 ( .A(n46983), .B(n48347), .Z(n48339) );
  XOR U59886 ( .A(n48340), .B(n48339), .Z(n48342) );
  IV U59887 ( .A(n46984), .Z(n46986) );
  NOR U59888 ( .A(n46986), .B(n46985), .Z(n48341) );
  IV U59889 ( .A(n46987), .Z(n46989) );
  NOR U59890 ( .A(n46989), .B(n46988), .Z(n50351) );
  NOR U59891 ( .A(n48341), .B(n50351), .Z(n46990) );
  XOR U59892 ( .A(n48342), .B(n46990), .Z(n50356) );
  XOR U59893 ( .A(n50354), .B(n50356), .Z(n48330) );
  XOR U59894 ( .A(n46991), .B(n48330), .Z(n50364) );
  XOR U59895 ( .A(n50362), .B(n50364), .Z(n50359) );
  IV U59896 ( .A(n46992), .Z(n46994) );
  NOR U59897 ( .A(n46994), .B(n46993), .Z(n48327) );
  NOR U59898 ( .A(n50358), .B(n48327), .Z(n46995) );
  XOR U59899 ( .A(n50359), .B(n46995), .Z(n50371) );
  IV U59900 ( .A(n46996), .Z(n46998) );
  NOR U59901 ( .A(n46998), .B(n46997), .Z(n50372) );
  NOR U59902 ( .A(n50374), .B(n50372), .Z(n46999) );
  XOR U59903 ( .A(n50371), .B(n46999), .Z(n50381) );
  IV U59904 ( .A(n47000), .Z(n47001) );
  NOR U59905 ( .A(n47002), .B(n47001), .Z(n50369) );
  IV U59906 ( .A(n47003), .Z(n47005) );
  NOR U59907 ( .A(n47005), .B(n47004), .Z(n50380) );
  NOR U59908 ( .A(n50369), .B(n50380), .Z(n47006) );
  XOR U59909 ( .A(n50381), .B(n47006), .Z(n47007) );
  IV U59910 ( .A(n47007), .Z(n50389) );
  IV U59911 ( .A(n47008), .Z(n47010) );
  NOR U59912 ( .A(n47010), .B(n47009), .Z(n50385) );
  XOR U59913 ( .A(n50389), .B(n50385), .Z(n47011) );
  XOR U59914 ( .A(n47012), .B(n47011), .Z(n48319) );
  XOR U59915 ( .A(n48320), .B(n48319), .Z(n48322) );
  IV U59916 ( .A(n47013), .Z(n47015) );
  NOR U59917 ( .A(n47015), .B(n47014), .Z(n48321) );
  IV U59918 ( .A(n47016), .Z(n47017) );
  NOR U59919 ( .A(n47018), .B(n47017), .Z(n48317) );
  NOR U59920 ( .A(n48321), .B(n48317), .Z(n47019) );
  XOR U59921 ( .A(n48322), .B(n47019), .Z(n48314) );
  XOR U59922 ( .A(n47020), .B(n48314), .Z(n50400) );
  XOR U59923 ( .A(n50398), .B(n50400), .Z(n50404) );
  XOR U59924 ( .A(n47021), .B(n50404), .Z(n48307) );
  XOR U59925 ( .A(n48306), .B(n48307), .Z(n48304) );
  IV U59926 ( .A(n47022), .Z(n47024) );
  NOR U59927 ( .A(n47024), .B(n47023), .Z(n48308) );
  IV U59928 ( .A(n47025), .Z(n47027) );
  NOR U59929 ( .A(n47027), .B(n47026), .Z(n48303) );
  NOR U59930 ( .A(n48308), .B(n48303), .Z(n47028) );
  XOR U59931 ( .A(n48304), .B(n47028), .Z(n48301) );
  XOR U59932 ( .A(n48300), .B(n48301), .Z(n48298) );
  XOR U59933 ( .A(n48295), .B(n48298), .Z(n50408) );
  XOR U59934 ( .A(n47029), .B(n50408), .Z(n50415) );
  XOR U59935 ( .A(n50413), .B(n50415), .Z(n50419) );
  IV U59936 ( .A(n47030), .Z(n47032) );
  NOR U59937 ( .A(n47032), .B(n47031), .Z(n50416) );
  NOR U59938 ( .A(n47034), .B(n47033), .Z(n50418) );
  NOR U59939 ( .A(n50416), .B(n50418), .Z(n47035) );
  XOR U59940 ( .A(n50419), .B(n47035), .Z(n48291) );
  XOR U59941 ( .A(n48293), .B(n48291), .Z(n50427) );
  IV U59942 ( .A(n47036), .Z(n47039) );
  IV U59943 ( .A(n47037), .Z(n47038) );
  NOR U59944 ( .A(n47039), .B(n47038), .Z(n50425) );
  XOR U59945 ( .A(n50427), .B(n50425), .Z(n50442) );
  IV U59946 ( .A(n47040), .Z(n47041) );
  NOR U59947 ( .A(n47042), .B(n47041), .Z(n50428) );
  IV U59948 ( .A(n47043), .Z(n47045) );
  NOR U59949 ( .A(n47045), .B(n47044), .Z(n50441) );
  NOR U59950 ( .A(n50428), .B(n50441), .Z(n47046) );
  XOR U59951 ( .A(n50442), .B(n47046), .Z(n48287) );
  IV U59952 ( .A(n47047), .Z(n47049) );
  NOR U59953 ( .A(n47049), .B(n47048), .Z(n50446) );
  NOR U59954 ( .A(n47050), .B(n48288), .Z(n47051) );
  NOR U59955 ( .A(n50446), .B(n47051), .Z(n47052) );
  XOR U59956 ( .A(n48287), .B(n47052), .Z(n50459) );
  IV U59957 ( .A(n47053), .Z(n47055) );
  IV U59958 ( .A(n47054), .Z(n47057) );
  NOR U59959 ( .A(n47055), .B(n47057), .Z(n50457) );
  XOR U59960 ( .A(n50459), .B(n50457), .Z(n50462) );
  IV U59961 ( .A(n47056), .Z(n47058) );
  NOR U59962 ( .A(n47058), .B(n47057), .Z(n50460) );
  XOR U59963 ( .A(n50462), .B(n50460), .Z(n50478) );
  NOR U59964 ( .A(n48283), .B(n47059), .Z(n47063) );
  IV U59965 ( .A(n47060), .Z(n47062) );
  IV U59966 ( .A(n47061), .Z(n47073) );
  NOR U59967 ( .A(n47062), .B(n47073), .Z(n50476) );
  NOR U59968 ( .A(n47063), .B(n50476), .Z(n47064) );
  XOR U59969 ( .A(n50478), .B(n47064), .Z(n48276) );
  IV U59970 ( .A(n47065), .Z(n47066) );
  NOR U59971 ( .A(n47067), .B(n47066), .Z(n50481) );
  IV U59972 ( .A(n47068), .Z(n47069) );
  NOR U59973 ( .A(n47070), .B(n47069), .Z(n48278) );
  IV U59974 ( .A(n47071), .Z(n47072) );
  NOR U59975 ( .A(n47073), .B(n47072), .Z(n48279) );
  XOR U59976 ( .A(n48278), .B(n48279), .Z(n47074) );
  NOR U59977 ( .A(n50481), .B(n47074), .Z(n47075) );
  XOR U59978 ( .A(n48276), .B(n47075), .Z(n50485) );
  XOR U59979 ( .A(n50484), .B(n50485), .Z(n54335) );
  IV U59980 ( .A(n47076), .Z(n47081) );
  IV U59981 ( .A(n47077), .Z(n47078) );
  NOR U59982 ( .A(n47081), .B(n47078), .Z(n54334) );
  IV U59983 ( .A(n47079), .Z(n47080) );
  NOR U59984 ( .A(n47081), .B(n47080), .Z(n54328) );
  NOR U59985 ( .A(n54334), .B(n54328), .Z(n50489) );
  XOR U59986 ( .A(n54335), .B(n50489), .Z(n47089) );
  IV U59987 ( .A(n47089), .Z(n47082) );
  NOR U59988 ( .A(n47083), .B(n47082), .Z(n50488) );
  IV U59989 ( .A(n47084), .Z(n47086) );
  NOR U59990 ( .A(n47086), .B(n47085), .Z(n47090) );
  IV U59991 ( .A(n47090), .Z(n47088) );
  XOR U59992 ( .A(n54328), .B(n54335), .Z(n47087) );
  NOR U59993 ( .A(n47088), .B(n47087), .Z(n50492) );
  NOR U59994 ( .A(n47090), .B(n47089), .Z(n47091) );
  NOR U59995 ( .A(n50492), .B(n47091), .Z(n47092) );
  NOR U59996 ( .A(n47093), .B(n47092), .Z(n47094) );
  NOR U59997 ( .A(n50488), .B(n47094), .Z(n48272) );
  IV U59998 ( .A(n47095), .Z(n47097) );
  NOR U59999 ( .A(n47097), .B(n47096), .Z(n50500) );
  IV U60000 ( .A(n47098), .Z(n48273) );
  NOR U60001 ( .A(n47099), .B(n48273), .Z(n47100) );
  NOR U60002 ( .A(n50500), .B(n47100), .Z(n47101) );
  XOR U60003 ( .A(n48272), .B(n47101), .Z(n51986) );
  IV U60004 ( .A(n47102), .Z(n47103) );
  NOR U60005 ( .A(n47104), .B(n47103), .Z(n51984) );
  IV U60006 ( .A(n47105), .Z(n47106) );
  NOR U60007 ( .A(n47107), .B(n47106), .Z(n54342) );
  NOR U60008 ( .A(n51984), .B(n54342), .Z(n50513) );
  XOR U60009 ( .A(n51986), .B(n50513), .Z(n48268) );
  XOR U60010 ( .A(n48270), .B(n48268), .Z(n51981) );
  IV U60011 ( .A(n47108), .Z(n47109) );
  NOR U60012 ( .A(n47110), .B(n47109), .Z(n51978) );
  IV U60013 ( .A(n47111), .Z(n47112) );
  NOR U60014 ( .A(n47113), .B(n47112), .Z(n54346) );
  NOR U60015 ( .A(n51978), .B(n54346), .Z(n50518) );
  XOR U60016 ( .A(n51981), .B(n50518), .Z(n48262) );
  XOR U60017 ( .A(n47114), .B(n48262), .Z(n48267) );
  XOR U60018 ( .A(n47115), .B(n48267), .Z(n47116) );
  IV U60019 ( .A(n47116), .Z(n50527) );
  XOR U60020 ( .A(n50526), .B(n50527), .Z(n50530) );
  XOR U60021 ( .A(n50529), .B(n50530), .Z(n54355) );
  XOR U60022 ( .A(n48259), .B(n54355), .Z(n47117) );
  IV U60023 ( .A(n47117), .Z(n50536) );
  IV U60024 ( .A(n47118), .Z(n47124) );
  IV U60025 ( .A(n47119), .Z(n47120) );
  NOR U60026 ( .A(n47124), .B(n47120), .Z(n50534) );
  XOR U60027 ( .A(n50536), .B(n50534), .Z(n48256) );
  IV U60028 ( .A(n47121), .Z(n47122) );
  NOR U60029 ( .A(n47123), .B(n47122), .Z(n48252) );
  NOR U60030 ( .A(n47125), .B(n47124), .Z(n47126) );
  IV U60031 ( .A(n47126), .Z(n48255) );
  NOR U60032 ( .A(n48255), .B(n47127), .Z(n47128) );
  NOR U60033 ( .A(n48252), .B(n47128), .Z(n47129) );
  XOR U60034 ( .A(n48256), .B(n47129), .Z(n48250) );
  XOR U60035 ( .A(n48251), .B(n48250), .Z(n50545) );
  XOR U60036 ( .A(n50544), .B(n50545), .Z(n48248) );
  IV U60037 ( .A(n47130), .Z(n47131) );
  NOR U60038 ( .A(n47132), .B(n47131), .Z(n48247) );
  IV U60039 ( .A(n47133), .Z(n47135) );
  NOR U60040 ( .A(n47135), .B(n47134), .Z(n48242) );
  NOR U60041 ( .A(n48247), .B(n48242), .Z(n47136) );
  XOR U60042 ( .A(n48248), .B(n47136), .Z(n48234) );
  IV U60043 ( .A(n47137), .Z(n47139) );
  NOR U60044 ( .A(n47139), .B(n47138), .Z(n48244) );
  NOR U60045 ( .A(n47140), .B(n48235), .Z(n47141) );
  NOR U60046 ( .A(n48244), .B(n47141), .Z(n47142) );
  XOR U60047 ( .A(n48234), .B(n47142), .Z(n50561) );
  XOR U60048 ( .A(n47143), .B(n50561), .Z(n48230) );
  XOR U60049 ( .A(n47144), .B(n48230), .Z(n48226) );
  XOR U60050 ( .A(n48224), .B(n48226), .Z(n50570) );
  IV U60051 ( .A(n47145), .Z(n47147) );
  NOR U60052 ( .A(n47147), .B(n47146), .Z(n48227) );
  IV U60053 ( .A(n47148), .Z(n47150) );
  IV U60054 ( .A(n47149), .Z(n47154) );
  NOR U60055 ( .A(n47150), .B(n47154), .Z(n50569) );
  NOR U60056 ( .A(n48227), .B(n50569), .Z(n47151) );
  XOR U60057 ( .A(n50570), .B(n47151), .Z(n50566) );
  IV U60058 ( .A(n47152), .Z(n47153) );
  NOR U60059 ( .A(n47154), .B(n47153), .Z(n50567) );
  IV U60060 ( .A(n47155), .Z(n47156) );
  NOR U60061 ( .A(n47159), .B(n47156), .Z(n50573) );
  NOR U60062 ( .A(n50567), .B(n50573), .Z(n47157) );
  XOR U60063 ( .A(n50566), .B(n47157), .Z(n50580) );
  IV U60064 ( .A(n47158), .Z(n47160) );
  NOR U60065 ( .A(n47160), .B(n47159), .Z(n50578) );
  XOR U60066 ( .A(n50580), .B(n50578), .Z(n48223) );
  IV U60067 ( .A(n47161), .Z(n47163) );
  NOR U60068 ( .A(n47163), .B(n47162), .Z(n48221) );
  XOR U60069 ( .A(n48223), .B(n48221), .Z(n48220) );
  IV U60070 ( .A(n47164), .Z(n47173) );
  IV U60071 ( .A(n47165), .Z(n47166) );
  NOR U60072 ( .A(n47173), .B(n47166), .Z(n47167) );
  IV U60073 ( .A(n47167), .Z(n48219) );
  XOR U60074 ( .A(n48220), .B(n48219), .Z(n48214) );
  IV U60075 ( .A(n47168), .Z(n47170) );
  NOR U60076 ( .A(n47170), .B(n47169), .Z(n48213) );
  IV U60077 ( .A(n47171), .Z(n47172) );
  NOR U60078 ( .A(n47173), .B(n47172), .Z(n50590) );
  NOR U60079 ( .A(n48213), .B(n50590), .Z(n47174) );
  XOR U60080 ( .A(n48214), .B(n47174), .Z(n48218) );
  XOR U60081 ( .A(n48216), .B(n48218), .Z(n50597) );
  XOR U60082 ( .A(n50595), .B(n50597), .Z(n50600) );
  XOR U60083 ( .A(n50598), .B(n50600), .Z(n50607) );
  XOR U60084 ( .A(n47175), .B(n50607), .Z(n51898) );
  XOR U60085 ( .A(n51893), .B(n51898), .Z(n47176) );
  XOR U60086 ( .A(n47177), .B(n47176), .Z(n50621) );
  XOR U60087 ( .A(n47178), .B(n50621), .Z(n50617) );
  NOR U60088 ( .A(n47186), .B(n50617), .Z(n54429) );
  IV U60089 ( .A(n47179), .Z(n47180) );
  NOR U60090 ( .A(n47181), .B(n47180), .Z(n48205) );
  IV U60091 ( .A(n47182), .Z(n47184) );
  NOR U60092 ( .A(n47184), .B(n47183), .Z(n47185) );
  IV U60093 ( .A(n47185), .Z(n50618) );
  XOR U60094 ( .A(n50618), .B(n50617), .Z(n48206) );
  XOR U60095 ( .A(n48205), .B(n48206), .Z(n47188) );
  NOR U60096 ( .A(n48206), .B(n47186), .Z(n47187) );
  NOR U60097 ( .A(n47188), .B(n47187), .Z(n47189) );
  NOR U60098 ( .A(n54429), .B(n47189), .Z(n48203) );
  IV U60099 ( .A(n47190), .Z(n47192) );
  NOR U60100 ( .A(n47192), .B(n47191), .Z(n48209) );
  IV U60101 ( .A(n47193), .Z(n47194) );
  NOR U60102 ( .A(n47195), .B(n47194), .Z(n48202) );
  NOR U60103 ( .A(n48209), .B(n48202), .Z(n47196) );
  XOR U60104 ( .A(n48203), .B(n47196), .Z(n48196) );
  XOR U60105 ( .A(n48195), .B(n48196), .Z(n50627) );
  XOR U60106 ( .A(n48198), .B(n50627), .Z(n50630) );
  XOR U60107 ( .A(n47197), .B(n50630), .Z(n48191) );
  XOR U60108 ( .A(n47198), .B(n48191), .Z(n50633) );
  XOR U60109 ( .A(n50632), .B(n50633), .Z(n48182) );
  XOR U60110 ( .A(n47199), .B(n48182), .Z(n48173) );
  XOR U60111 ( .A(n48174), .B(n48173), .Z(n48176) );
  XOR U60112 ( .A(n47207), .B(n48176), .Z(n47203) );
  IV U60113 ( .A(n47200), .Z(n47201) );
  NOR U60114 ( .A(n47201), .B(n47214), .Z(n47210) );
  IV U60115 ( .A(n47210), .Z(n47202) );
  NOR U60116 ( .A(n47203), .B(n47202), .Z(n51864) );
  IV U60117 ( .A(n47204), .Z(n47206) );
  NOR U60118 ( .A(n47206), .B(n47205), .Z(n48171) );
  NOR U60119 ( .A(n47207), .B(n48171), .Z(n47208) );
  XOR U60120 ( .A(n48176), .B(n47208), .Z(n47209) );
  NOR U60121 ( .A(n47210), .B(n47209), .Z(n47211) );
  NOR U60122 ( .A(n51864), .B(n47211), .Z(n48164) );
  IV U60123 ( .A(n47212), .Z(n47213) );
  NOR U60124 ( .A(n47214), .B(n47213), .Z(n48167) );
  IV U60125 ( .A(n47215), .Z(n47224) );
  IV U60126 ( .A(n47216), .Z(n47217) );
  NOR U60127 ( .A(n47224), .B(n47217), .Z(n48165) );
  NOR U60128 ( .A(n48167), .B(n48165), .Z(n47218) );
  XOR U60129 ( .A(n48164), .B(n47218), .Z(n48162) );
  IV U60130 ( .A(n47219), .Z(n47221) );
  NOR U60131 ( .A(n47221), .B(n47220), .Z(n48155) );
  IV U60132 ( .A(n47222), .Z(n47223) );
  NOR U60133 ( .A(n47224), .B(n47223), .Z(n48160) );
  NOR U60134 ( .A(n48155), .B(n48160), .Z(n47225) );
  XOR U60135 ( .A(n48162), .B(n47225), .Z(n48157) );
  XOR U60136 ( .A(n48159), .B(n48157), .Z(n50657) );
  IV U60137 ( .A(n47226), .Z(n47227) );
  NOR U60138 ( .A(n47228), .B(n47227), .Z(n50649) );
  NOR U60139 ( .A(n50658), .B(n50649), .Z(n47229) );
  XOR U60140 ( .A(n50657), .B(n47229), .Z(n50653) );
  XOR U60141 ( .A(n47230), .B(n50653), .Z(n48154) );
  XOR U60142 ( .A(n47231), .B(n48154), .Z(n47253) );
  IV U60143 ( .A(n47253), .Z(n48149) );
  IV U60144 ( .A(n47232), .Z(n47233) );
  NOR U60145 ( .A(n47233), .B(n47241), .Z(n47234) );
  IV U60146 ( .A(n47234), .Z(n47235) );
  NOR U60147 ( .A(n47236), .B(n47235), .Z(n47237) );
  IV U60148 ( .A(n47237), .Z(n47254) );
  NOR U60149 ( .A(n48149), .B(n47254), .Z(n51830) );
  IV U60150 ( .A(n47238), .Z(n47240) );
  NOR U60151 ( .A(n47240), .B(n47239), .Z(n48143) );
  NOR U60152 ( .A(n47242), .B(n47241), .Z(n47243) );
  IV U60153 ( .A(n47243), .Z(n47252) );
  IV U60154 ( .A(n47244), .Z(n47245) );
  NOR U60155 ( .A(n47246), .B(n47245), .Z(n47247) );
  IV U60156 ( .A(n47247), .Z(n47249) );
  NOR U60157 ( .A(n47249), .B(n47248), .Z(n47250) );
  IV U60158 ( .A(n47250), .Z(n47251) );
  NOR U60159 ( .A(n47252), .B(n47251), .Z(n48147) );
  XOR U60160 ( .A(n47253), .B(n48147), .Z(n48144) );
  XOR U60161 ( .A(n48143), .B(n48144), .Z(n47256) );
  NOR U60162 ( .A(n48144), .B(n47254), .Z(n47255) );
  NOR U60163 ( .A(n47256), .B(n47255), .Z(n47257) );
  NOR U60164 ( .A(n51830), .B(n47257), .Z(n48138) );
  XOR U60165 ( .A(n48139), .B(n48138), .Z(n50664) );
  NOR U60166 ( .A(n47259), .B(n47258), .Z(n48140) );
  IV U60167 ( .A(n47260), .Z(n47262) );
  NOR U60168 ( .A(n47262), .B(n47261), .Z(n50662) );
  NOR U60169 ( .A(n48140), .B(n50662), .Z(n47263) );
  XOR U60170 ( .A(n50664), .B(n47263), .Z(n50668) );
  XOR U60171 ( .A(n50669), .B(n50668), .Z(n50673) );
  IV U60172 ( .A(n47264), .Z(n47265) );
  NOR U60173 ( .A(n47266), .B(n47265), .Z(n50670) );
  IV U60174 ( .A(n47267), .Z(n47269) );
  NOR U60175 ( .A(n47269), .B(n47268), .Z(n50674) );
  NOR U60176 ( .A(n50670), .B(n50674), .Z(n47270) );
  XOR U60177 ( .A(n50673), .B(n47270), .Z(n48134) );
  IV U60178 ( .A(n47271), .Z(n47273) );
  NOR U60179 ( .A(n47273), .B(n47272), .Z(n48132) );
  XOR U60180 ( .A(n48134), .B(n48132), .Z(n48136) );
  XOR U60181 ( .A(n48135), .B(n48136), .Z(n50682) );
  IV U60182 ( .A(n47274), .Z(n47275) );
  NOR U60183 ( .A(n47276), .B(n47275), .Z(n50679) );
  IV U60184 ( .A(n47277), .Z(n47279) );
  NOR U60185 ( .A(n47279), .B(n47278), .Z(n50683) );
  NOR U60186 ( .A(n50679), .B(n50683), .Z(n47280) );
  XOR U60187 ( .A(n50682), .B(n47280), .Z(n48123) );
  XOR U60188 ( .A(n47281), .B(n48123), .Z(n48121) );
  XOR U60189 ( .A(n48117), .B(n48121), .Z(n50693) );
  IV U60190 ( .A(n47282), .Z(n47284) );
  NOR U60191 ( .A(n47284), .B(n47283), .Z(n48119) );
  IV U60192 ( .A(n47285), .Z(n47287) );
  NOR U60193 ( .A(n47287), .B(n47286), .Z(n50692) );
  NOR U60194 ( .A(n48119), .B(n50692), .Z(n47288) );
  XOR U60195 ( .A(n50693), .B(n47288), .Z(n48114) );
  IV U60196 ( .A(n47289), .Z(n47291) );
  NOR U60197 ( .A(n47291), .B(n47290), .Z(n48115) );
  IV U60198 ( .A(n47297), .Z(n47292) );
  NOR U60199 ( .A(n47292), .B(n47296), .Z(n50699) );
  NOR U60200 ( .A(n48115), .B(n50699), .Z(n47293) );
  XOR U60201 ( .A(n48114), .B(n47293), .Z(n50716) );
  IV U60202 ( .A(n47294), .Z(n47295) );
  NOR U60203 ( .A(n47295), .B(n47296), .Z(n50715) );
  XOR U60204 ( .A(n47297), .B(n47296), .Z(n47300) );
  IV U60205 ( .A(n47298), .Z(n47299) );
  NOR U60206 ( .A(n47300), .B(n47299), .Z(n48112) );
  NOR U60207 ( .A(n50715), .B(n48112), .Z(n47301) );
  XOR U60208 ( .A(n50716), .B(n47301), .Z(n47302) );
  IV U60209 ( .A(n47302), .Z(n50714) );
  IV U60210 ( .A(n47303), .Z(n47305) );
  NOR U60211 ( .A(n47305), .B(n47304), .Z(n50712) );
  XOR U60212 ( .A(n50714), .B(n50712), .Z(n48107) );
  XOR U60213 ( .A(n48106), .B(n48107), .Z(n48111) );
  XOR U60214 ( .A(n48109), .B(n48111), .Z(n47306) );
  NOR U60215 ( .A(n47307), .B(n47306), .Z(n51777) );
  IV U60216 ( .A(n47308), .Z(n47309) );
  NOR U60217 ( .A(n47310), .B(n47309), .Z(n48104) );
  NOR U60218 ( .A(n48104), .B(n48109), .Z(n47311) );
  XOR U60219 ( .A(n47311), .B(n48111), .Z(n47316) );
  NOR U60220 ( .A(n47312), .B(n47316), .Z(n47313) );
  NOR U60221 ( .A(n51777), .B(n47313), .Z(n47314) );
  NOR U60222 ( .A(n47315), .B(n47314), .Z(n47319) );
  IV U60223 ( .A(n47315), .Z(n47318) );
  IV U60224 ( .A(n47316), .Z(n47317) );
  NOR U60225 ( .A(n47318), .B(n47317), .Z(n48103) );
  NOR U60226 ( .A(n47319), .B(n48103), .Z(n48095) );
  IV U60227 ( .A(n47320), .Z(n47321) );
  NOR U60228 ( .A(n47322), .B(n47321), .Z(n48100) );
  IV U60229 ( .A(n47323), .Z(n47324) );
  NOR U60230 ( .A(n47325), .B(n47324), .Z(n48098) );
  NOR U60231 ( .A(n48100), .B(n48098), .Z(n47326) );
  XOR U60232 ( .A(n48095), .B(n47326), .Z(n50723) );
  XOR U60233 ( .A(n47327), .B(n50723), .Z(n50725) );
  XOR U60234 ( .A(n50726), .B(n50725), .Z(n50735) );
  XOR U60235 ( .A(n47328), .B(n50735), .Z(n50731) );
  XOR U60236 ( .A(n47329), .B(n50731), .Z(n50742) );
  XOR U60237 ( .A(n50741), .B(n50742), .Z(n48089) );
  XOR U60238 ( .A(n47330), .B(n48089), .Z(n48084) );
  NOR U60239 ( .A(n47331), .B(n50747), .Z(n47335) );
  IV U60240 ( .A(n47332), .Z(n47334) );
  IV U60241 ( .A(n47333), .Z(n47338) );
  NOR U60242 ( .A(n47334), .B(n47338), .Z(n48085) );
  NOR U60243 ( .A(n47335), .B(n48085), .Z(n47336) );
  XOR U60244 ( .A(n48084), .B(n47336), .Z(n48079) );
  IV U60245 ( .A(n47337), .Z(n47339) );
  NOR U60246 ( .A(n47339), .B(n47338), .Z(n47340) );
  IV U60247 ( .A(n47340), .Z(n48078) );
  XOR U60248 ( .A(n48079), .B(n48078), .Z(n50760) );
  NOR U60249 ( .A(n48075), .B(n47341), .Z(n47345) );
  IV U60250 ( .A(n47342), .Z(n47344) );
  NOR U60251 ( .A(n47344), .B(n47343), .Z(n50759) );
  NOR U60252 ( .A(n47345), .B(n50759), .Z(n47346) );
  XOR U60253 ( .A(n50760), .B(n47346), .Z(n50758) );
  XOR U60254 ( .A(n50756), .B(n50758), .Z(n51729) );
  XOR U60255 ( .A(n50764), .B(n51729), .Z(n48072) );
  IV U60256 ( .A(n47347), .Z(n47349) );
  NOR U60257 ( .A(n47349), .B(n47348), .Z(n50765) );
  IV U60258 ( .A(n47350), .Z(n47352) );
  NOR U60259 ( .A(n47352), .B(n47351), .Z(n48071) );
  NOR U60260 ( .A(n50765), .B(n48071), .Z(n47353) );
  XOR U60261 ( .A(n48072), .B(n47353), .Z(n48067) );
  IV U60262 ( .A(n47354), .Z(n47356) );
  NOR U60263 ( .A(n47356), .B(n47355), .Z(n48065) );
  XOR U60264 ( .A(n48067), .B(n48065), .Z(n48069) );
  XOR U60265 ( .A(n48068), .B(n48069), .Z(n48058) );
  XOR U60266 ( .A(n48056), .B(n48058), .Z(n48063) );
  XOR U60267 ( .A(n48059), .B(n48063), .Z(n47357) );
  NOR U60268 ( .A(n47358), .B(n47357), .Z(n51706) );
  IV U60269 ( .A(n47359), .Z(n47360) );
  NOR U60270 ( .A(n47361), .B(n47360), .Z(n48062) );
  NOR U60271 ( .A(n48059), .B(n48062), .Z(n47362) );
  XOR U60272 ( .A(n47362), .B(n48063), .Z(n50774) );
  NOR U60273 ( .A(n47363), .B(n50774), .Z(n47364) );
  NOR U60274 ( .A(n51706), .B(n47364), .Z(n50789) );
  IV U60275 ( .A(n47365), .Z(n47367) );
  NOR U60276 ( .A(n47367), .B(n47366), .Z(n50773) );
  IV U60277 ( .A(n47368), .Z(n47369) );
  NOR U60278 ( .A(n47370), .B(n47369), .Z(n50788) );
  NOR U60279 ( .A(n50773), .B(n50788), .Z(n47371) );
  XOR U60280 ( .A(n50789), .B(n47371), .Z(n50779) );
  IV U60281 ( .A(n47372), .Z(n47373) );
  NOR U60282 ( .A(n50783), .B(n47373), .Z(n47376) );
  NOR U60283 ( .A(n47374), .B(n48046), .Z(n47375) );
  NOR U60284 ( .A(n47376), .B(n47375), .Z(n47377) );
  XOR U60285 ( .A(n50779), .B(n47377), .Z(n48034) );
  IV U60286 ( .A(n47378), .Z(n48042) );
  NOR U60287 ( .A(n47379), .B(n48042), .Z(n48035) );
  IV U60288 ( .A(n47380), .Z(n47382) );
  NOR U60289 ( .A(n47382), .B(n47381), .Z(n48038) );
  NOR U60290 ( .A(n48035), .B(n48038), .Z(n47383) );
  XOR U60291 ( .A(n48034), .B(n47383), .Z(n50798) );
  XOR U60292 ( .A(n47384), .B(n50798), .Z(n50796) );
  XOR U60293 ( .A(n50795), .B(n50796), .Z(n48030) );
  XOR U60294 ( .A(n48028), .B(n48030), .Z(n51670) );
  XOR U60295 ( .A(n51671), .B(n51670), .Z(n47385) );
  IV U60296 ( .A(n47385), .Z(n50809) );
  IV U60297 ( .A(n47386), .Z(n47387) );
  NOR U60298 ( .A(n47387), .B(n50810), .Z(n50803) );
  XOR U60299 ( .A(n50809), .B(n50803), .Z(n51660) );
  NOR U60300 ( .A(n47388), .B(n50808), .Z(n47389) );
  NOR U60301 ( .A(n47389), .B(n50810), .Z(n47390) );
  XOR U60302 ( .A(n51660), .B(n47390), .Z(n51642) );
  IV U60303 ( .A(n51642), .Z(n50818) );
  IV U60304 ( .A(n47391), .Z(n47392) );
  NOR U60305 ( .A(n47393), .B(n47392), .Z(n51641) );
  IV U60306 ( .A(n47394), .Z(n47395) );
  NOR U60307 ( .A(n47396), .B(n47395), .Z(n54616) );
  NOR U60308 ( .A(n51641), .B(n54616), .Z(n50819) );
  XOR U60309 ( .A(n50818), .B(n50819), .Z(n54623) );
  XOR U60310 ( .A(n50821), .B(n54623), .Z(n50839) );
  IV U60311 ( .A(n50839), .Z(n47402) );
  IV U60312 ( .A(n50837), .Z(n47397) );
  NOR U60313 ( .A(n47398), .B(n47397), .Z(n50835) );
  NOR U60314 ( .A(n47399), .B(n50830), .Z(n47400) );
  NOR U60315 ( .A(n50835), .B(n47400), .Z(n47401) );
  XOR U60316 ( .A(n47402), .B(n47401), .Z(n50856) );
  XOR U60317 ( .A(n47403), .B(n50856), .Z(n50860) );
  NOR U60318 ( .A(n47405), .B(n47404), .Z(n50854) );
  IV U60319 ( .A(n47406), .Z(n47408) );
  IV U60320 ( .A(n47407), .Z(n47411) );
  NOR U60321 ( .A(n47408), .B(n47411), .Z(n50858) );
  NOR U60322 ( .A(n50854), .B(n50858), .Z(n47409) );
  XOR U60323 ( .A(n50860), .B(n47409), .Z(n48013) );
  IV U60324 ( .A(n47410), .Z(n47412) );
  NOR U60325 ( .A(n47412), .B(n47411), .Z(n48012) );
  IV U60326 ( .A(n47413), .Z(n47414) );
  NOR U60327 ( .A(n47415), .B(n47414), .Z(n48015) );
  NOR U60328 ( .A(n48012), .B(n48015), .Z(n47416) );
  XOR U60329 ( .A(n48013), .B(n47416), .Z(n51622) );
  XOR U60330 ( .A(n51623), .B(n51622), .Z(n48005) );
  IV U60331 ( .A(n47417), .Z(n47419) );
  NOR U60332 ( .A(n47419), .B(n47418), .Z(n48004) );
  IV U60333 ( .A(n47420), .Z(n47421) );
  NOR U60334 ( .A(n47422), .B(n47421), .Z(n50867) );
  NOR U60335 ( .A(n48004), .B(n50867), .Z(n47423) );
  XOR U60336 ( .A(n48005), .B(n47423), .Z(n48000) );
  NOR U60337 ( .A(n47429), .B(n48000), .Z(n51610) );
  IV U60338 ( .A(n47424), .Z(n47426) );
  NOR U60339 ( .A(n47426), .B(n47425), .Z(n47996) );
  NOR U60340 ( .A(n47427), .B(n48001), .Z(n47428) );
  XOR U60341 ( .A(n47428), .B(n48000), .Z(n47997) );
  IV U60342 ( .A(n47997), .Z(n47430) );
  XOR U60343 ( .A(n47996), .B(n47430), .Z(n47432) );
  NOR U60344 ( .A(n47430), .B(n47429), .Z(n47431) );
  NOR U60345 ( .A(n47432), .B(n47431), .Z(n47433) );
  NOR U60346 ( .A(n51610), .B(n47433), .Z(n47994) );
  XOR U60347 ( .A(n50879), .B(n47994), .Z(n50889) );
  IV U60348 ( .A(n47434), .Z(n47436) );
  NOR U60349 ( .A(n47436), .B(n47435), .Z(n47993) );
  NOR U60350 ( .A(n47438), .B(n47437), .Z(n50888) );
  NOR U60351 ( .A(n47993), .B(n50888), .Z(n47439) );
  XOR U60352 ( .A(n50889), .B(n47439), .Z(n50887) );
  IV U60353 ( .A(n47440), .Z(n47442) );
  NOR U60354 ( .A(n47442), .B(n47441), .Z(n50885) );
  XOR U60355 ( .A(n50887), .B(n50885), .Z(n50895) );
  XOR U60356 ( .A(n50893), .B(n50895), .Z(n50903) );
  XOR U60357 ( .A(n47443), .B(n50903), .Z(n50900) );
  XOR U60358 ( .A(n50899), .B(n50900), .Z(n47986) );
  NOR U60359 ( .A(n47445), .B(n47444), .Z(n47990) );
  IV U60360 ( .A(n47446), .Z(n47448) );
  IV U60361 ( .A(n47447), .Z(n47455) );
  NOR U60362 ( .A(n47448), .B(n47455), .Z(n47987) );
  NOR U60363 ( .A(n47990), .B(n47987), .Z(n47449) );
  XOR U60364 ( .A(n47986), .B(n47449), .Z(n50908) );
  IV U60365 ( .A(n47450), .Z(n47451) );
  NOR U60366 ( .A(n47452), .B(n47451), .Z(n47983) );
  IV U60367 ( .A(n47453), .Z(n47454) );
  NOR U60368 ( .A(n47455), .B(n47454), .Z(n50907) );
  NOR U60369 ( .A(n47983), .B(n50907), .Z(n47456) );
  XOR U60370 ( .A(n50908), .B(n47456), .Z(n47978) );
  IV U60371 ( .A(n47457), .Z(n47459) );
  NOR U60372 ( .A(n47459), .B(n47458), .Z(n50906) );
  NOR U60373 ( .A(n47460), .B(n47980), .Z(n47461) );
  NOR U60374 ( .A(n50906), .B(n47461), .Z(n47462) );
  XOR U60375 ( .A(n47978), .B(n47462), .Z(n50919) );
  IV U60376 ( .A(n47463), .Z(n47465) );
  NOR U60377 ( .A(n47465), .B(n47464), .Z(n50914) );
  IV U60378 ( .A(n47466), .Z(n47468) );
  NOR U60379 ( .A(n47468), .B(n47467), .Z(n50917) );
  NOR U60380 ( .A(n50914), .B(n50917), .Z(n47469) );
  XOR U60381 ( .A(n50919), .B(n47469), .Z(n50921) );
  IV U60382 ( .A(n47470), .Z(n47472) );
  NOR U60383 ( .A(n47472), .B(n47471), .Z(n50920) );
  NOR U60384 ( .A(n47474), .B(n47473), .Z(n50924) );
  NOR U60385 ( .A(n50920), .B(n50924), .Z(n47475) );
  XOR U60386 ( .A(n50921), .B(n47475), .Z(n50931) );
  IV U60387 ( .A(n47476), .Z(n47477) );
  NOR U60388 ( .A(n47477), .B(n47481), .Z(n50929) );
  XOR U60389 ( .A(n50931), .B(n50929), .Z(n47975) );
  XOR U60390 ( .A(n47974), .B(n47975), .Z(n47973) );
  NOR U60391 ( .A(n47478), .B(n47973), .Z(n47971) );
  IV U60392 ( .A(n47479), .Z(n47480) );
  NOR U60393 ( .A(n47481), .B(n47480), .Z(n47482) );
  IV U60394 ( .A(n47482), .Z(n47972) );
  XOR U60395 ( .A(n47973), .B(n47972), .Z(n47964) );
  NOR U60396 ( .A(n47483), .B(n47964), .Z(n47484) );
  NOR U60397 ( .A(n47971), .B(n47484), .Z(n47491) );
  IV U60398 ( .A(n47485), .Z(n47487) );
  NOR U60399 ( .A(n47487), .B(n47486), .Z(n47963) );
  NOR U60400 ( .A(n47489), .B(n47488), .Z(n47967) );
  NOR U60401 ( .A(n47963), .B(n47967), .Z(n47490) );
  XOR U60402 ( .A(n47491), .B(n47490), .Z(n50944) );
  XOR U60403 ( .A(n50944), .B(n50942), .Z(n50946) );
  XOR U60404 ( .A(n50945), .B(n50946), .Z(n50952) );
  XOR U60405 ( .A(n50951), .B(n50952), .Z(n47961) );
  XOR U60406 ( .A(n47960), .B(n47961), .Z(n50963) );
  IV U60407 ( .A(n47492), .Z(n47497) );
  NOR U60408 ( .A(n47494), .B(n47493), .Z(n47495) );
  IV U60409 ( .A(n47495), .Z(n47496) );
  NOR U60410 ( .A(n47497), .B(n47496), .Z(n50961) );
  XOR U60411 ( .A(n50963), .B(n50961), .Z(n50965) );
  IV U60412 ( .A(n47498), .Z(n47499) );
  NOR U60413 ( .A(n47500), .B(n47499), .Z(n50964) );
  IV U60414 ( .A(n47501), .Z(n47503) );
  NOR U60415 ( .A(n47503), .B(n47502), .Z(n47958) );
  NOR U60416 ( .A(n50964), .B(n47958), .Z(n47504) );
  XOR U60417 ( .A(n50965), .B(n47504), .Z(n47509) );
  IV U60418 ( .A(n47509), .Z(n47951) );
  NOR U60419 ( .A(n47510), .B(n47951), .Z(n54680) );
  NOR U60420 ( .A(n47519), .B(n47505), .Z(n47954) );
  IV U60421 ( .A(n47506), .Z(n47507) );
  NOR U60422 ( .A(n47508), .B(n47507), .Z(n47950) );
  XOR U60423 ( .A(n47950), .B(n47509), .Z(n47955) );
  XOR U60424 ( .A(n47954), .B(n47955), .Z(n47512) );
  NOR U60425 ( .A(n47955), .B(n47510), .Z(n47511) );
  NOR U60426 ( .A(n47512), .B(n47511), .Z(n47513) );
  NOR U60427 ( .A(n54680), .B(n47513), .Z(n47948) );
  IV U60428 ( .A(n47514), .Z(n47517) );
  IV U60429 ( .A(n47515), .Z(n47516) );
  NOR U60430 ( .A(n47517), .B(n47516), .Z(n47947) );
  IV U60431 ( .A(n47518), .Z(n47522) );
  NOR U60432 ( .A(n47520), .B(n47519), .Z(n47521) );
  IV U60433 ( .A(n47521), .Z(n47528) );
  NOR U60434 ( .A(n47522), .B(n47528), .Z(n50971) );
  NOR U60435 ( .A(n47947), .B(n50971), .Z(n47523) );
  XOR U60436 ( .A(n47948), .B(n47523), .Z(n50976) );
  IV U60437 ( .A(n47524), .Z(n47525) );
  NOR U60438 ( .A(n47535), .B(n47525), .Z(n47531) );
  IV U60439 ( .A(n47531), .Z(n47526) );
  NOR U60440 ( .A(n50976), .B(n47526), .Z(n54697) );
  IV U60441 ( .A(n47527), .Z(n47529) );
  NOR U60442 ( .A(n47529), .B(n47528), .Z(n47530) );
  IV U60443 ( .A(n47530), .Z(n50975) );
  XOR U60444 ( .A(n50975), .B(n50976), .Z(n47945) );
  NOR U60445 ( .A(n47531), .B(n47945), .Z(n47532) );
  NOR U60446 ( .A(n54697), .B(n47532), .Z(n47537) );
  IV U60447 ( .A(n47533), .Z(n47534) );
  NOR U60448 ( .A(n47535), .B(n47534), .Z(n50978) );
  NOR U60449 ( .A(n47944), .B(n50978), .Z(n47536) );
  XOR U60450 ( .A(n47537), .B(n47536), .Z(n50989) );
  IV U60451 ( .A(n50989), .Z(n47545) );
  IV U60452 ( .A(n47538), .Z(n47540) );
  NOR U60453 ( .A(n47540), .B(n47539), .Z(n50987) );
  IV U60454 ( .A(n47541), .Z(n47543) );
  NOR U60455 ( .A(n47543), .B(n47542), .Z(n50985) );
  NOR U60456 ( .A(n50987), .B(n50985), .Z(n47544) );
  XOR U60457 ( .A(n47545), .B(n47544), .Z(n50982) );
  IV U60458 ( .A(n47548), .Z(n47546) );
  NOR U60459 ( .A(n47547), .B(n47546), .Z(n47554) );
  IV U60460 ( .A(n47547), .Z(n47549) );
  NOR U60461 ( .A(n47549), .B(n47548), .Z(n50981) );
  XOR U60462 ( .A(n47551), .B(n47550), .Z(n47552) );
  NOR U60463 ( .A(n50981), .B(n47552), .Z(n47553) );
  NOR U60464 ( .A(n47554), .B(n47553), .Z(n47555) );
  XOR U60465 ( .A(n50982), .B(n47555), .Z(n47942) );
  IV U60466 ( .A(n47942), .Z(n51000) );
  IV U60467 ( .A(n47556), .Z(n47557) );
  NOR U60468 ( .A(n47558), .B(n47557), .Z(n47941) );
  NOR U60469 ( .A(n47559), .B(n47938), .Z(n47560) );
  NOR U60470 ( .A(n47941), .B(n47560), .Z(n47561) );
  XOR U60471 ( .A(n51000), .B(n47561), .Z(n47574) );
  IV U60472 ( .A(n47562), .Z(n47564) );
  NOR U60473 ( .A(n47564), .B(n47563), .Z(n47565) );
  IV U60474 ( .A(n47565), .Z(n47578) );
  NOR U60475 ( .A(n47574), .B(n47578), .Z(n54726) );
  IV U60476 ( .A(n47566), .Z(n47567) );
  NOR U60477 ( .A(n47568), .B(n47567), .Z(n51014) );
  IV U60478 ( .A(n47569), .Z(n47571) );
  NOR U60479 ( .A(n47571), .B(n47570), .Z(n47576) );
  IV U60480 ( .A(n47576), .Z(n47573) );
  XOR U60481 ( .A(n47941), .B(n47942), .Z(n47572) );
  NOR U60482 ( .A(n47573), .B(n47572), .Z(n54723) );
  IV U60483 ( .A(n47574), .Z(n47575) );
  NOR U60484 ( .A(n47576), .B(n47575), .Z(n47577) );
  NOR U60485 ( .A(n54723), .B(n47577), .Z(n51015) );
  XOR U60486 ( .A(n51014), .B(n51015), .Z(n47580) );
  NOR U60487 ( .A(n51015), .B(n47578), .Z(n47579) );
  NOR U60488 ( .A(n47580), .B(n47579), .Z(n47581) );
  NOR U60489 ( .A(n54726), .B(n47581), .Z(n51018) );
  XOR U60490 ( .A(n51020), .B(n51018), .Z(n47933) );
  XOR U60491 ( .A(n47932), .B(n47933), .Z(n47930) );
  XOR U60492 ( .A(n47931), .B(n47930), .Z(n47922) );
  XOR U60493 ( .A(n47921), .B(n47922), .Z(n51537) );
  IV U60494 ( .A(n47582), .Z(n47583) );
  NOR U60495 ( .A(n47584), .B(n47583), .Z(n47926) );
  IV U60496 ( .A(n47585), .Z(n47586) );
  NOR U60497 ( .A(n47591), .B(n47586), .Z(n47925) );
  NOR U60498 ( .A(n47926), .B(n47925), .Z(n51539) );
  XOR U60499 ( .A(n51537), .B(n51539), .Z(n47919) );
  XOR U60500 ( .A(n47915), .B(n47919), .Z(n47587) );
  NOR U60501 ( .A(n47588), .B(n47587), .Z(n51535) );
  IV U60502 ( .A(n47589), .Z(n47590) );
  NOR U60503 ( .A(n47591), .B(n47590), .Z(n47917) );
  NOR U60504 ( .A(n47915), .B(n47917), .Z(n47592) );
  XOR U60505 ( .A(n47592), .B(n47919), .Z(n51027) );
  NOR U60506 ( .A(n47593), .B(n51027), .Z(n47594) );
  NOR U60507 ( .A(n51535), .B(n47594), .Z(n47911) );
  XOR U60508 ( .A(n47595), .B(n47911), .Z(n51032) );
  XOR U60509 ( .A(n51030), .B(n51032), .Z(n51037) );
  IV U60510 ( .A(n47596), .Z(n47597) );
  NOR U60511 ( .A(n47598), .B(n47597), .Z(n51033) );
  XOR U60512 ( .A(n51037), .B(n51033), .Z(n47909) );
  IV U60513 ( .A(n47599), .Z(n47600) );
  NOR U60514 ( .A(n47601), .B(n47600), .Z(n51036) );
  NOR U60515 ( .A(n47602), .B(n47601), .Z(n47603) );
  IV U60516 ( .A(n47603), .Z(n47607) );
  NOR U60517 ( .A(n47604), .B(n47607), .Z(n47907) );
  NOR U60518 ( .A(n51036), .B(n47907), .Z(n47605) );
  XOR U60519 ( .A(n47909), .B(n47605), .Z(n51041) );
  IV U60520 ( .A(n47606), .Z(n47608) );
  NOR U60521 ( .A(n47608), .B(n47607), .Z(n47609) );
  IV U60522 ( .A(n47609), .Z(n47610) );
  NOR U60523 ( .A(n47611), .B(n47610), .Z(n47612) );
  IV U60524 ( .A(n47612), .Z(n51042) );
  XOR U60525 ( .A(n51041), .B(n51042), .Z(n47905) );
  NOR U60526 ( .A(n47620), .B(n47905), .Z(n51521) );
  IV U60527 ( .A(n47613), .Z(n47615) );
  NOR U60528 ( .A(n47615), .B(n47614), .Z(n47897) );
  IV U60529 ( .A(n47616), .Z(n47618) );
  NOR U60530 ( .A(n47618), .B(n47617), .Z(n47619) );
  IV U60531 ( .A(n47619), .Z(n47906) );
  XOR U60532 ( .A(n47906), .B(n47905), .Z(n47898) );
  XOR U60533 ( .A(n47897), .B(n47898), .Z(n47622) );
  NOR U60534 ( .A(n47898), .B(n47620), .Z(n47621) );
  NOR U60535 ( .A(n47622), .B(n47621), .Z(n47623) );
  NOR U60536 ( .A(n51521), .B(n47623), .Z(n47889) );
  IV U60537 ( .A(n47624), .Z(n47626) );
  NOR U60538 ( .A(n47626), .B(n47625), .Z(n47901) );
  IV U60539 ( .A(n47627), .Z(n47628) );
  NOR U60540 ( .A(n47628), .B(n47630), .Z(n47888) );
  IV U60541 ( .A(n47629), .Z(n47631) );
  NOR U60542 ( .A(n47631), .B(n47630), .Z(n47895) );
  NOR U60543 ( .A(n47888), .B(n47895), .Z(n47632) );
  IV U60544 ( .A(n47632), .Z(n47633) );
  NOR U60545 ( .A(n47901), .B(n47633), .Z(n47634) );
  XOR U60546 ( .A(n47889), .B(n47634), .Z(n47893) );
  XOR U60547 ( .A(n47635), .B(n47893), .Z(n47636) );
  IV U60548 ( .A(n47636), .Z(n51053) );
  XOR U60549 ( .A(n51052), .B(n51053), .Z(n51056) );
  XOR U60550 ( .A(n51055), .B(n51056), .Z(n47876) );
  XOR U60551 ( .A(n47637), .B(n47876), .Z(n47877) );
  XOR U60552 ( .A(n47878), .B(n47877), .Z(n51067) );
  XOR U60553 ( .A(n51066), .B(n51067), .Z(n51069) );
  NOR U60554 ( .A(n47645), .B(n51069), .Z(n51493) );
  IV U60555 ( .A(n47638), .Z(n47640) );
  NOR U60556 ( .A(n47640), .B(n47639), .Z(n47870) );
  IV U60557 ( .A(n47641), .Z(n47643) );
  NOR U60558 ( .A(n47643), .B(n47642), .Z(n47644) );
  IV U60559 ( .A(n47644), .Z(n51070) );
  XOR U60560 ( .A(n51070), .B(n51069), .Z(n47871) );
  XOR U60561 ( .A(n47870), .B(n47871), .Z(n47647) );
  NOR U60562 ( .A(n47871), .B(n47645), .Z(n47646) );
  NOR U60563 ( .A(n47647), .B(n47646), .Z(n47648) );
  NOR U60564 ( .A(n51493), .B(n47648), .Z(n47649) );
  IV U60565 ( .A(n47649), .Z(n47868) );
  XOR U60566 ( .A(n47867), .B(n47868), .Z(n47863) );
  XOR U60567 ( .A(n47650), .B(n47863), .Z(n47861) );
  XOR U60568 ( .A(n47859), .B(n47861), .Z(n47854) );
  XOR U60569 ( .A(n47853), .B(n47854), .Z(n47858) );
  IV U60570 ( .A(n47651), .Z(n47653) );
  IV U60571 ( .A(n47652), .Z(n47657) );
  NOR U60572 ( .A(n47653), .B(n47657), .Z(n47856) );
  XOR U60573 ( .A(n47858), .B(n47856), .Z(n51078) );
  IV U60574 ( .A(n47654), .Z(n47655) );
  NOR U60575 ( .A(n47662), .B(n47655), .Z(n47851) );
  IV U60576 ( .A(n47656), .Z(n47658) );
  NOR U60577 ( .A(n47658), .B(n47657), .Z(n51076) );
  NOR U60578 ( .A(n47851), .B(n51076), .Z(n47659) );
  XOR U60579 ( .A(n51078), .B(n47659), .Z(n47847) );
  IV U60580 ( .A(n47660), .Z(n47661) );
  NOR U60581 ( .A(n47662), .B(n47661), .Z(n51089) );
  IV U60582 ( .A(n47663), .Z(n47665) );
  NOR U60583 ( .A(n47665), .B(n47664), .Z(n47848) );
  NOR U60584 ( .A(n51089), .B(n47848), .Z(n47666) );
  XOR U60585 ( .A(n47847), .B(n47666), .Z(n47845) );
  XOR U60586 ( .A(n47846), .B(n47845), .Z(n47842) );
  IV U60587 ( .A(n47667), .Z(n47669) );
  NOR U60588 ( .A(n47669), .B(n47668), .Z(n54823) );
  NOR U60589 ( .A(n51465), .B(n54823), .Z(n47840) );
  XOR U60590 ( .A(n47842), .B(n47840), .Z(n54826) );
  XOR U60591 ( .A(n47838), .B(n54826), .Z(n47836) );
  XOR U60592 ( .A(n47835), .B(n47836), .Z(n51099) );
  NOR U60593 ( .A(n47671), .B(n47670), .Z(n47832) );
  IV U60594 ( .A(n47672), .Z(n47674) );
  NOR U60595 ( .A(n47674), .B(n47673), .Z(n51097) );
  NOR U60596 ( .A(n47832), .B(n51097), .Z(n47675) );
  XOR U60597 ( .A(n51099), .B(n47675), .Z(n51095) );
  XOR U60598 ( .A(n51096), .B(n51095), .Z(n51440) );
  IV U60599 ( .A(n47676), .Z(n47677) );
  NOR U60600 ( .A(n47678), .B(n47677), .Z(n51444) );
  IV U60601 ( .A(n47679), .Z(n47681) );
  NOR U60602 ( .A(n47681), .B(n47680), .Z(n51439) );
  NOR U60603 ( .A(n51444), .B(n51439), .Z(n51102) );
  XOR U60604 ( .A(n51440), .B(n51102), .Z(n47682) );
  IV U60605 ( .A(n47682), .Z(n51111) );
  XOR U60606 ( .A(n51103), .B(n51111), .Z(n51108) );
  XOR U60607 ( .A(n47683), .B(n51108), .Z(n51122) );
  XOR U60608 ( .A(n47684), .B(n51122), .Z(n47831) );
  XOR U60609 ( .A(n47829), .B(n47831), .Z(n47828) );
  XOR U60610 ( .A(n47826), .B(n47828), .Z(n51138) );
  XOR U60611 ( .A(n51136), .B(n51138), .Z(n47814) );
  XOR U60612 ( .A(n47685), .B(n47814), .Z(n51411) );
  XOR U60613 ( .A(n47813), .B(n51411), .Z(n47686) );
  IV U60614 ( .A(n47686), .Z(n47809) );
  IV U60615 ( .A(n47687), .Z(n47689) );
  NOR U60616 ( .A(n47689), .B(n47688), .Z(n47807) );
  XOR U60617 ( .A(n47809), .B(n47807), .Z(n47811) );
  XOR U60618 ( .A(n47810), .B(n47811), .Z(n47803) );
  XOR U60619 ( .A(n47802), .B(n47803), .Z(n47805) );
  XOR U60620 ( .A(n47806), .B(n47805), .Z(n47794) );
  IV U60621 ( .A(n47690), .Z(n47691) );
  NOR U60622 ( .A(n47692), .B(n47691), .Z(n47793) );
  IV U60623 ( .A(n47693), .Z(n47695) );
  NOR U60624 ( .A(n47695), .B(n47694), .Z(n47799) );
  NOR U60625 ( .A(n47793), .B(n47799), .Z(n47696) );
  XOR U60626 ( .A(n47794), .B(n47696), .Z(n47798) );
  XOR U60627 ( .A(n47796), .B(n47798), .Z(n51147) );
  XOR U60628 ( .A(n51146), .B(n51147), .Z(n51150) );
  XOR U60629 ( .A(n51149), .B(n51150), .Z(n47698) );
  NOR U60630 ( .A(n47697), .B(n47698), .Z(n54839) );
  IV U60631 ( .A(n47698), .Z(n47699) );
  NOR U60632 ( .A(n47700), .B(n47699), .Z(n51159) );
  IV U60633 ( .A(n47701), .Z(n47702) );
  NOR U60634 ( .A(n47707), .B(n47702), .Z(n51157) );
  XOR U60635 ( .A(n51159), .B(n51157), .Z(n47703) );
  NOR U60636 ( .A(n54839), .B(n47703), .Z(n47704) );
  IV U60637 ( .A(n47704), .Z(n51164) );
  IV U60638 ( .A(n47705), .Z(n47706) );
  NOR U60639 ( .A(n47707), .B(n47706), .Z(n51163) );
  IV U60640 ( .A(n47708), .Z(n47709) );
  NOR U60641 ( .A(n47710), .B(n47709), .Z(n51154) );
  NOR U60642 ( .A(n51163), .B(n51154), .Z(n47711) );
  XOR U60643 ( .A(n51164), .B(n47711), .Z(n47712) );
  NOR U60644 ( .A(n47713), .B(n47712), .Z(n47716) );
  IV U60645 ( .A(n47713), .Z(n47715) );
  XOR U60646 ( .A(n51163), .B(n51164), .Z(n47714) );
  NOR U60647 ( .A(n47715), .B(n47714), .Z(n54846) );
  NOR U60648 ( .A(n47716), .B(n54846), .Z(n47786) );
  XOR U60649 ( .A(n47717), .B(n47786), .Z(n51181) );
  XOR U60650 ( .A(n47718), .B(n51181), .Z(n47719) );
  IV U60651 ( .A(n47719), .Z(n51177) );
  XOR U60652 ( .A(n51176), .B(n51177), .Z(n51186) );
  XOR U60653 ( .A(n51185), .B(n51186), .Z(n47720) );
  NOR U60654 ( .A(n47721), .B(n47720), .Z(n51360) );
  IV U60655 ( .A(n47722), .Z(n47724) );
  NOR U60656 ( .A(n47724), .B(n47723), .Z(n51183) );
  NOR U60657 ( .A(n51185), .B(n51183), .Z(n47725) );
  XOR U60658 ( .A(n47725), .B(n51186), .Z(n51196) );
  NOR U60659 ( .A(n47726), .B(n51196), .Z(n47727) );
  NOR U60660 ( .A(n51360), .B(n47727), .Z(n51189) );
  XOR U60661 ( .A(n47728), .B(n51189), .Z(n47782) );
  XOR U60662 ( .A(n47729), .B(n47782), .Z(n47776) );
  XOR U60663 ( .A(n47730), .B(n47776), .Z(n51256) );
  NOR U60664 ( .A(n47732), .B(n47731), .Z(n47747) );
  NOR U60665 ( .A(n47747), .B(n47733), .Z(n47742) );
  IV U60666 ( .A(n47742), .Z(n47734) );
  NOR U60667 ( .A(n47759), .B(n47734), .Z(n47744) );
  XOR U60668 ( .A(n47747), .B(n47735), .Z(n51222) );
  IV U60669 ( .A(n47736), .Z(n47738) );
  NOR U60670 ( .A(n47738), .B(n47737), .Z(n51223) );
  IV U60671 ( .A(n51223), .Z(n47739) );
  NOR U60672 ( .A(n51222), .B(n47739), .Z(n47751) );
  IV U60673 ( .A(n47751), .Z(n47740) );
  NOR U60674 ( .A(n47741), .B(n47740), .Z(n51218) );
  IV U60675 ( .A(n51218), .Z(n47743) );
  XOR U60676 ( .A(n47759), .B(n47742), .Z(n51216) );
  NOR U60677 ( .A(n47743), .B(n51216), .Z(n47763) );
  NOR U60678 ( .A(n47744), .B(n47763), .Z(n47745) );
  XOR U60679 ( .A(n47746), .B(n47745), .Z(n51214) );
  NOR U60680 ( .A(n47748), .B(n47747), .Z(n47749) );
  XOR U60681 ( .A(n47750), .B(n47749), .Z(n51221) );
  NOR U60682 ( .A(n47751), .B(n51221), .Z(n47752) );
  NOR U60683 ( .A(n51218), .B(n47752), .Z(n51301) );
  IV U60684 ( .A(n51301), .Z(n51299) );
  IV U60685 ( .A(n47753), .Z(n47755) );
  NOR U60686 ( .A(n47755), .B(n47754), .Z(n47756) );
  IV U60687 ( .A(n47756), .Z(n51234) );
  NOR U60688 ( .A(n51222), .B(n51234), .Z(n51302) );
  IV U60689 ( .A(n51302), .Z(n47757) );
  NOR U60690 ( .A(n51299), .B(n47757), .Z(n51217) );
  IV U60691 ( .A(n51217), .Z(n47758) );
  NOR U60692 ( .A(n47759), .B(n47758), .Z(n51215) );
  IV U60693 ( .A(n51215), .Z(n47760) );
  NOR U60694 ( .A(n51214), .B(n47760), .Z(n51212) );
  IV U60695 ( .A(n51212), .Z(n47762) );
  XOR U60696 ( .A(n51210), .B(n51207), .Z(n47761) );
  NOR U60697 ( .A(n47762), .B(n47761), .Z(n51251) );
  IV U60698 ( .A(n51251), .Z(n47769) );
  IV U60699 ( .A(n47763), .Z(n47764) );
  NOR U60700 ( .A(n47765), .B(n47764), .Z(n51208) );
  IV U60701 ( .A(n51208), .Z(n47766) );
  NOR U60702 ( .A(n51210), .B(n47766), .Z(n47771) );
  XOR U60703 ( .A(n47768), .B(n47767), .Z(n47772) );
  XOR U60704 ( .A(n47771), .B(n47772), .Z(n51262) );
  NOR U60705 ( .A(n47769), .B(n51262), .Z(n51253) );
  IV U60706 ( .A(n51253), .Z(n47770) );
  NOR U60707 ( .A(n51256), .B(n47770), .Z(n51205) );
  IV U60708 ( .A(n51205), .Z(n51200) );
  IV U60709 ( .A(n47771), .Z(n47773) );
  NOR U60710 ( .A(n47773), .B(n47772), .Z(n51254) );
  IV U60711 ( .A(n51254), .Z(n47774) );
  NOR U60712 ( .A(n51256), .B(n47774), .Z(n54874) );
  IV U60713 ( .A(n47775), .Z(n47777) );
  IV U60714 ( .A(n47776), .Z(n51202) );
  NOR U60715 ( .A(n47777), .B(n51202), .Z(n54868) );
  IV U60716 ( .A(n47778), .Z(n47779) );
  NOR U60717 ( .A(n47782), .B(n47779), .Z(n51352) );
  IV U60718 ( .A(n47780), .Z(n47781) );
  NOR U60719 ( .A(n47782), .B(n47781), .Z(n54861) );
  IV U60720 ( .A(n47783), .Z(n47784) );
  NOR U60721 ( .A(n51181), .B(n47784), .Z(n51366) );
  IV U60722 ( .A(n51366), .Z(n51368) );
  IV U60723 ( .A(n47785), .Z(n47787) );
  IV U60724 ( .A(n47786), .Z(n51169) );
  NOR U60725 ( .A(n47787), .B(n51169), .Z(n51378) );
  IV U60726 ( .A(n47788), .Z(n47789) );
  NOR U60727 ( .A(n47789), .B(n51169), .Z(n47790) );
  IV U60728 ( .A(n47790), .Z(n47791) );
  NOR U60729 ( .A(n47792), .B(n47791), .Z(n51374) );
  NOR U60730 ( .A(n51378), .B(n51374), .Z(n51175) );
  IV U60731 ( .A(n47793), .Z(n47795) );
  IV U60732 ( .A(n47794), .Z(n47801) );
  NOR U60733 ( .A(n47795), .B(n47801), .Z(n51390) );
  IV U60734 ( .A(n47796), .Z(n47797) );
  NOR U60735 ( .A(n47798), .B(n47797), .Z(n51389) );
  NOR U60736 ( .A(n51390), .B(n51389), .Z(n51145) );
  IV U60737 ( .A(n47799), .Z(n47800) );
  NOR U60738 ( .A(n47801), .B(n47800), .Z(n51395) );
  IV U60739 ( .A(n47802), .Z(n47804) );
  NOR U60740 ( .A(n47804), .B(n47803), .Z(n51400) );
  NOR U60741 ( .A(n47806), .B(n47805), .Z(n51393) );
  NOR U60742 ( .A(n51400), .B(n51393), .Z(n51144) );
  IV U60743 ( .A(n47807), .Z(n47808) );
  NOR U60744 ( .A(n47809), .B(n47808), .Z(n51406) );
  IV U60745 ( .A(n47810), .Z(n47812) );
  NOR U60746 ( .A(n47812), .B(n47811), .Z(n51403) );
  NOR U60747 ( .A(n51406), .B(n51403), .Z(n51143) );
  NOR U60748 ( .A(n47813), .B(n51411), .Z(n51142) );
  NOR U60749 ( .A(n47815), .B(n47814), .Z(n47816) );
  IV U60750 ( .A(n47816), .Z(n51140) );
  NOR U60751 ( .A(n51140), .B(n47817), .Z(n47818) );
  IV U60752 ( .A(n47818), .Z(n47825) );
  XOR U60753 ( .A(n47820), .B(n47819), .Z(n47821) );
  NOR U60754 ( .A(n47822), .B(n47821), .Z(n47823) );
  IV U60755 ( .A(n47823), .Z(n47824) );
  NOR U60756 ( .A(n47825), .B(n47824), .Z(n51417) );
  IV U60757 ( .A(n47826), .Z(n47827) );
  NOR U60758 ( .A(n47828), .B(n47827), .Z(n51132) );
  IV U60759 ( .A(n47829), .Z(n47830) );
  NOR U60760 ( .A(n47831), .B(n47830), .Z(n51129) );
  IV U60761 ( .A(n51129), .Z(n51121) );
  IV U60762 ( .A(n47832), .Z(n47833) );
  NOR U60763 ( .A(n47833), .B(n47836), .Z(n47834) );
  IV U60764 ( .A(n47834), .Z(n51462) );
  IV U60765 ( .A(n47835), .Z(n47837) );
  NOR U60766 ( .A(n47837), .B(n47836), .Z(n51458) );
  IV U60767 ( .A(n47842), .Z(n51466) );
  NOR U60768 ( .A(n47840), .B(n51466), .Z(n47839) );
  NOR U60769 ( .A(n47839), .B(n47838), .Z(n47844) );
  IV U60770 ( .A(n47840), .Z(n47841) );
  NOR U60771 ( .A(n47842), .B(n47841), .Z(n47843) );
  NOR U60772 ( .A(n47844), .B(n47843), .Z(n51094) );
  NOR U60773 ( .A(n47846), .B(n47845), .Z(n54818) );
  IV U60774 ( .A(n47847), .Z(n51091) );
  IV U60775 ( .A(n47848), .Z(n47849) );
  NOR U60776 ( .A(n51091), .B(n47849), .Z(n54815) );
  NOR U60777 ( .A(n54818), .B(n54815), .Z(n47850) );
  IV U60778 ( .A(n47850), .Z(n51093) );
  IV U60779 ( .A(n47851), .Z(n47852) );
  NOR U60780 ( .A(n47852), .B(n47858), .Z(n51086) );
  IV U60781 ( .A(n51086), .Z(n51075) );
  IV U60782 ( .A(n47853), .Z(n47855) );
  NOR U60783 ( .A(n47855), .B(n47854), .Z(n51475) );
  IV U60784 ( .A(n47856), .Z(n47857) );
  NOR U60785 ( .A(n47858), .B(n47857), .Z(n51473) );
  NOR U60786 ( .A(n51475), .B(n51473), .Z(n51074) );
  IV U60787 ( .A(n47859), .Z(n47860) );
  NOR U60788 ( .A(n47861), .B(n47860), .Z(n51478) );
  IV U60789 ( .A(n47862), .Z(n47864) );
  NOR U60790 ( .A(n47864), .B(n47863), .Z(n51485) );
  NOR U60791 ( .A(n51478), .B(n51485), .Z(n51073) );
  IV U60792 ( .A(n47865), .Z(n47866) );
  NOR U60793 ( .A(n47866), .B(n47868), .Z(n51484) );
  IV U60794 ( .A(n47867), .Z(n47869) );
  NOR U60795 ( .A(n47869), .B(n47868), .Z(n51490) );
  IV U60796 ( .A(n47870), .Z(n47873) );
  IV U60797 ( .A(n47871), .Z(n47872) );
  NOR U60798 ( .A(n47873), .B(n47872), .Z(n51496) );
  IV U60799 ( .A(n47874), .Z(n47875) );
  NOR U60800 ( .A(n47876), .B(n47875), .Z(n54800) );
  IV U60801 ( .A(n47877), .Z(n54804) );
  NOR U60802 ( .A(n54804), .B(n47878), .Z(n51064) );
  IV U60803 ( .A(n47879), .Z(n47882) );
  NOR U60804 ( .A(n47880), .B(n51053), .Z(n47881) );
  IV U60805 ( .A(n47881), .Z(n47884) );
  NOR U60806 ( .A(n47882), .B(n47884), .Z(n51060) );
  IV U60807 ( .A(n47883), .Z(n47885) );
  NOR U60808 ( .A(n47885), .B(n47884), .Z(n51504) );
  IV U60809 ( .A(n47886), .Z(n47887) );
  NOR U60810 ( .A(n47893), .B(n47887), .Z(n54773) );
  IV U60811 ( .A(n47888), .Z(n47890) );
  IV U60812 ( .A(n47889), .Z(n47902) );
  NOR U60813 ( .A(n47890), .B(n47902), .Z(n51513) );
  NOR U60814 ( .A(n54773), .B(n51513), .Z(n51051) );
  IV U60815 ( .A(n47891), .Z(n47892) );
  NOR U60816 ( .A(n47893), .B(n47892), .Z(n47894) );
  IV U60817 ( .A(n47894), .Z(n51512) );
  IV U60818 ( .A(n47895), .Z(n47896) );
  NOR U60819 ( .A(n47896), .B(n47902), .Z(n51515) );
  IV U60820 ( .A(n47897), .Z(n47900) );
  IV U60821 ( .A(n47898), .Z(n47899) );
  NOR U60822 ( .A(n47900), .B(n47899), .Z(n51518) );
  IV U60823 ( .A(n47901), .Z(n47903) );
  NOR U60824 ( .A(n47903), .B(n47902), .Z(n54768) );
  NOR U60825 ( .A(n51518), .B(n54768), .Z(n47904) );
  IV U60826 ( .A(n47904), .Z(n51049) );
  NOR U60827 ( .A(n47906), .B(n47905), .Z(n51046) );
  IV U60828 ( .A(n51046), .Z(n51040) );
  IV U60829 ( .A(n47907), .Z(n47908) );
  NOR U60830 ( .A(n47909), .B(n47908), .Z(n54762) );
  IV U60831 ( .A(n47910), .Z(n47913) );
  IV U60832 ( .A(n47911), .Z(n47912) );
  NOR U60833 ( .A(n47913), .B(n47912), .Z(n47914) );
  IV U60834 ( .A(n47914), .Z(n51534) );
  IV U60835 ( .A(n47915), .Z(n47916) );
  NOR U60836 ( .A(n47919), .B(n47916), .Z(n54745) );
  IV U60837 ( .A(n47917), .Z(n47918) );
  NOR U60838 ( .A(n47919), .B(n47918), .Z(n54743) );
  XOR U60839 ( .A(n54745), .B(n54743), .Z(n47920) );
  NOR U60840 ( .A(n51535), .B(n47920), .Z(n51025) );
  NOR U60841 ( .A(n47921), .B(n47922), .Z(n47929) );
  IV U60842 ( .A(n47921), .Z(n47924) );
  IV U60843 ( .A(n47922), .Z(n47923) );
  NOR U60844 ( .A(n47924), .B(n47923), .Z(n51546) );
  XOR U60845 ( .A(n47926), .B(n47925), .Z(n47927) );
  NOR U60846 ( .A(n51546), .B(n47927), .Z(n47928) );
  NOR U60847 ( .A(n47929), .B(n47928), .Z(n51024) );
  NOR U60848 ( .A(n47931), .B(n47930), .Z(n51544) );
  IV U60849 ( .A(n47932), .Z(n47934) );
  NOR U60850 ( .A(n47934), .B(n47933), .Z(n47935) );
  IV U60851 ( .A(n47935), .Z(n51549) );
  NOR U60852 ( .A(n54723), .B(n54726), .Z(n47936) );
  IV U60853 ( .A(n47936), .Z(n51013) );
  IV U60854 ( .A(n47937), .Z(n47940) );
  NOR U60855 ( .A(n47938), .B(n47942), .Z(n47939) );
  IV U60856 ( .A(n47939), .Z(n51010) );
  NOR U60857 ( .A(n47940), .B(n51010), .Z(n51005) );
  IV U60858 ( .A(n47941), .Z(n47943) );
  NOR U60859 ( .A(n47943), .B(n47942), .Z(n51002) );
  IV U60860 ( .A(n51002), .Z(n50995) );
  IV U60861 ( .A(n47944), .Z(n47946) );
  IV U60862 ( .A(n47945), .Z(n50979) );
  NOR U60863 ( .A(n47946), .B(n50979), .Z(n51552) );
  IV U60864 ( .A(n47947), .Z(n47949) );
  IV U60865 ( .A(n47948), .Z(n50972) );
  NOR U60866 ( .A(n47949), .B(n50972), .Z(n54687) );
  IV U60867 ( .A(n47950), .Z(n47952) );
  NOR U60868 ( .A(n47952), .B(n47951), .Z(n54676) );
  NOR U60869 ( .A(n54676), .B(n54680), .Z(n47953) );
  IV U60870 ( .A(n47953), .Z(n50970) );
  IV U60871 ( .A(n47954), .Z(n47957) );
  IV U60872 ( .A(n47955), .Z(n47956) );
  NOR U60873 ( .A(n47957), .B(n47956), .Z(n51555) );
  IV U60874 ( .A(n47958), .Z(n47959) );
  NOR U60875 ( .A(n47959), .B(n50965), .Z(n54673) );
  IV U60876 ( .A(n47960), .Z(n47962) );
  NOR U60877 ( .A(n47962), .B(n47961), .Z(n50959) );
  IV U60878 ( .A(n50959), .Z(n50950) );
  IV U60879 ( .A(n47963), .Z(n47965) );
  IV U60880 ( .A(n47964), .Z(n47968) );
  NOR U60881 ( .A(n47965), .B(n47968), .Z(n47966) );
  IV U60882 ( .A(n47966), .Z(n51569) );
  IV U60883 ( .A(n47967), .Z(n47969) );
  NOR U60884 ( .A(n47969), .B(n47968), .Z(n47970) );
  IV U60885 ( .A(n47970), .Z(n51568) );
  IV U60886 ( .A(n47971), .Z(n54667) );
  NOR U60887 ( .A(n47973), .B(n47972), .Z(n50936) );
  IV U60888 ( .A(n47974), .Z(n47976) );
  NOR U60889 ( .A(n47976), .B(n47975), .Z(n50933) );
  IV U60890 ( .A(n50933), .Z(n50928) );
  IV U60891 ( .A(n47977), .Z(n47982) );
  IV U60892 ( .A(n47978), .Z(n47979) );
  NOR U60893 ( .A(n47980), .B(n47979), .Z(n47981) );
  IV U60894 ( .A(n47981), .Z(n50912) );
  NOR U60895 ( .A(n47982), .B(n50912), .Z(n51583) );
  IV U60896 ( .A(n47983), .Z(n47984) );
  NOR U60897 ( .A(n50908), .B(n47984), .Z(n51586) );
  IV U60898 ( .A(n50907), .Z(n47985) );
  NOR U60899 ( .A(n50908), .B(n47985), .Z(n54648) );
  IV U60900 ( .A(n47986), .Z(n47991) );
  IV U60901 ( .A(n47987), .Z(n47988) );
  NOR U60902 ( .A(n47991), .B(n47988), .Z(n54650) );
  XOR U60903 ( .A(n54648), .B(n54650), .Z(n47989) );
  NOR U60904 ( .A(n51586), .B(n47989), .Z(n50904) );
  IV U60905 ( .A(n47990), .Z(n47992) );
  NOR U60906 ( .A(n47992), .B(n47991), .Z(n54638) );
  IV U60907 ( .A(n47993), .Z(n47995) );
  IV U60908 ( .A(n47994), .Z(n50880) );
  NOR U60909 ( .A(n47995), .B(n50880), .Z(n50883) );
  IV U60910 ( .A(n50883), .Z(n50878) );
  IV U60911 ( .A(n47996), .Z(n47998) );
  NOR U60912 ( .A(n47998), .B(n47997), .Z(n51605) );
  IV U60913 ( .A(n47999), .Z(n48003) );
  NOR U60914 ( .A(n48001), .B(n48000), .Z(n48002) );
  IV U60915 ( .A(n48002), .Z(n50871) );
  NOR U60916 ( .A(n48003), .B(n50871), .Z(n51608) );
  NOR U60917 ( .A(n51610), .B(n51608), .Z(n50875) );
  IV U60918 ( .A(n48004), .Z(n48006) );
  IV U60919 ( .A(n48005), .Z(n50868) );
  NOR U60920 ( .A(n48006), .B(n50868), .Z(n50864) );
  IV U60921 ( .A(n48007), .Z(n48008) );
  NOR U60922 ( .A(n48008), .B(n51622), .Z(n50862) );
  IV U60923 ( .A(n48009), .Z(n48011) );
  NOR U60924 ( .A(n48012), .B(n48013), .Z(n48010) );
  NOR U60925 ( .A(n48011), .B(n48010), .Z(n48020) );
  IV U60926 ( .A(n48012), .Z(n48014) );
  IV U60927 ( .A(n48013), .Z(n48016) );
  NOR U60928 ( .A(n48014), .B(n48016), .Z(n51630) );
  IV U60929 ( .A(n48015), .Z(n48017) );
  NOR U60930 ( .A(n48017), .B(n48016), .Z(n51626) );
  NOR U60931 ( .A(n51630), .B(n51626), .Z(n48018) );
  IV U60932 ( .A(n48018), .Z(n48019) );
  NOR U60933 ( .A(n48020), .B(n48019), .Z(n48021) );
  IV U60934 ( .A(n48021), .Z(n50861) );
  IV U60935 ( .A(n48022), .Z(n48025) );
  NOR U60936 ( .A(n50856), .B(n48023), .Z(n48024) );
  IV U60937 ( .A(n48024), .Z(n50852) );
  NOR U60938 ( .A(n48025), .B(n50852), .Z(n50846) );
  IV U60939 ( .A(n48030), .Z(n54595) );
  NOR U60940 ( .A(n48028), .B(n54595), .Z(n48026) );
  NOR U60941 ( .A(n48027), .B(n48026), .Z(n48032) );
  IV U60942 ( .A(n48028), .Z(n48029) );
  NOR U60943 ( .A(n48030), .B(n48029), .Z(n48031) );
  NOR U60944 ( .A(n48032), .B(n48031), .Z(n50802) );
  IV U60945 ( .A(n48033), .Z(n48037) );
  IV U60946 ( .A(n48034), .Z(n48041) );
  XOR U60947 ( .A(n48035), .B(n48041), .Z(n48036) );
  NOR U60948 ( .A(n48037), .B(n48036), .Z(n51679) );
  IV U60949 ( .A(n48038), .Z(n48039) );
  NOR U60950 ( .A(n48039), .B(n48041), .Z(n51686) );
  IV U60951 ( .A(n48040), .Z(n48044) );
  NOR U60952 ( .A(n48042), .B(n48041), .Z(n48043) );
  IV U60953 ( .A(n48043), .Z(n48050) );
  NOR U60954 ( .A(n48044), .B(n48050), .Z(n51688) );
  NOR U60955 ( .A(n51686), .B(n51688), .Z(n50794) );
  IV U60956 ( .A(n48045), .Z(n48048) );
  NOR U60957 ( .A(n50779), .B(n48046), .Z(n48047) );
  IV U60958 ( .A(n48047), .Z(n48054) );
  NOR U60959 ( .A(n48048), .B(n48054), .Z(n51695) );
  IV U60960 ( .A(n48049), .Z(n48051) );
  NOR U60961 ( .A(n48051), .B(n48050), .Z(n51692) );
  NOR U60962 ( .A(n51695), .B(n51692), .Z(n48052) );
  IV U60963 ( .A(n48052), .Z(n50793) );
  IV U60964 ( .A(n48053), .Z(n48055) );
  NOR U60965 ( .A(n48055), .B(n48054), .Z(n51697) );
  IV U60966 ( .A(n48056), .Z(n48057) );
  NOR U60967 ( .A(n48058), .B(n48057), .Z(n51717) );
  IV U60968 ( .A(n48059), .Z(n48060) );
  NOR U60969 ( .A(n48060), .B(n48063), .Z(n51714) );
  NOR U60970 ( .A(n51717), .B(n51714), .Z(n48061) );
  IV U60971 ( .A(n48061), .Z(n50772) );
  IV U60972 ( .A(n48062), .Z(n48064) );
  NOR U60973 ( .A(n48064), .B(n48063), .Z(n51712) );
  IV U60974 ( .A(n48065), .Z(n48066) );
  NOR U60975 ( .A(n48067), .B(n48066), .Z(n51721) );
  IV U60976 ( .A(n48068), .Z(n48070) );
  NOR U60977 ( .A(n48070), .B(n48069), .Z(n51719) );
  NOR U60978 ( .A(n51721), .B(n51719), .Z(n55156) );
  IV U60979 ( .A(n48071), .Z(n48073) );
  IV U60980 ( .A(n48072), .Z(n50766) );
  NOR U60981 ( .A(n48073), .B(n50766), .Z(n58056) );
  IV U60982 ( .A(n48074), .Z(n48077) );
  NOR U60983 ( .A(n48075), .B(n48079), .Z(n48076) );
  IV U60984 ( .A(n48076), .Z(n48081) );
  NOR U60985 ( .A(n48077), .B(n48081), .Z(n51735) );
  NOR U60986 ( .A(n48079), .B(n48078), .Z(n54575) );
  IV U60987 ( .A(n48080), .Z(n48082) );
  NOR U60988 ( .A(n48082), .B(n48081), .Z(n51739) );
  NOR U60989 ( .A(n54575), .B(n51739), .Z(n48083) );
  IV U60990 ( .A(n48083), .Z(n50755) );
  IV U60991 ( .A(n48084), .Z(n50748) );
  IV U60992 ( .A(n48085), .Z(n48086) );
  NOR U60993 ( .A(n50748), .B(n48086), .Z(n54578) );
  IV U60994 ( .A(n48087), .Z(n48088) );
  NOR U60995 ( .A(n48088), .B(n48089), .Z(n54549) );
  NOR U60996 ( .A(n48090), .B(n48089), .Z(n48091) );
  IV U60997 ( .A(n48091), .Z(n48092) );
  NOR U60998 ( .A(n48093), .B(n48092), .Z(n51742) );
  IV U60999 ( .A(n48094), .Z(n48097) );
  IV U61000 ( .A(n48095), .Z(n48101) );
  XOR U61001 ( .A(n48100), .B(n48101), .Z(n48096) );
  NOR U61002 ( .A(n48097), .B(n48096), .Z(n51764) );
  IV U61003 ( .A(n48098), .Z(n48099) );
  NOR U61004 ( .A(n48099), .B(n48101), .Z(n51768) );
  IV U61005 ( .A(n48100), .Z(n48102) );
  NOR U61006 ( .A(n48102), .B(n48101), .Z(n51770) );
  NOR U61007 ( .A(n51768), .B(n51770), .Z(n50721) );
  IV U61008 ( .A(n48103), .Z(n51773) );
  IV U61009 ( .A(n48104), .Z(n48105) );
  NOR U61010 ( .A(n48105), .B(n48111), .Z(n51774) );
  IV U61011 ( .A(n48106), .Z(n48108) );
  NOR U61012 ( .A(n48108), .B(n48107), .Z(n57916) );
  IV U61013 ( .A(n48109), .Z(n48110) );
  NOR U61014 ( .A(n48111), .B(n48110), .Z(n57919) );
  NOR U61015 ( .A(n57916), .B(n57919), .Z(n51782) );
  IV U61016 ( .A(n51782), .Z(n50719) );
  IV U61017 ( .A(n48112), .Z(n48113) );
  NOR U61018 ( .A(n48113), .B(n50716), .Z(n50703) );
  IV U61019 ( .A(n48114), .Z(n50701) );
  IV U61020 ( .A(n48115), .Z(n48116) );
  NOR U61021 ( .A(n50701), .B(n48116), .Z(n54508) );
  IV U61022 ( .A(n48117), .Z(n48118) );
  NOR U61023 ( .A(n48121), .B(n48118), .Z(n51796) );
  IV U61024 ( .A(n48119), .Z(n48120) );
  NOR U61025 ( .A(n48121), .B(n48120), .Z(n51791) );
  NOR U61026 ( .A(n51796), .B(n51791), .Z(n50696) );
  IV U61027 ( .A(n48122), .Z(n48127) );
  IV U61028 ( .A(n48123), .Z(n48124) );
  NOR U61029 ( .A(n48125), .B(n48124), .Z(n48126) );
  IV U61030 ( .A(n48126), .Z(n48129) );
  NOR U61031 ( .A(n48127), .B(n48129), .Z(n51794) );
  IV U61032 ( .A(n48128), .Z(n48130) );
  NOR U61033 ( .A(n48130), .B(n48129), .Z(n54501) );
  IV U61034 ( .A(n50683), .Z(n48131) );
  NOR U61035 ( .A(n50682), .B(n48131), .Z(n51804) );
  IV U61036 ( .A(n48132), .Z(n48133) );
  NOR U61037 ( .A(n48134), .B(n48133), .Z(n51814) );
  IV U61038 ( .A(n48135), .Z(n48137) );
  NOR U61039 ( .A(n48137), .B(n48136), .Z(n51807) );
  NOR U61040 ( .A(n51814), .B(n51807), .Z(n50678) );
  IV U61041 ( .A(n48138), .Z(n48141) );
  NOR U61042 ( .A(n48139), .B(n48141), .Z(n51824) );
  IV U61043 ( .A(n48140), .Z(n48142) );
  NOR U61044 ( .A(n48142), .B(n48141), .Z(n51821) );
  NOR U61045 ( .A(n51824), .B(n51821), .Z(n50667) );
  IV U61046 ( .A(n48143), .Z(n48146) );
  IV U61047 ( .A(n48144), .Z(n48145) );
  NOR U61048 ( .A(n48146), .B(n48145), .Z(n51826) );
  IV U61049 ( .A(n48147), .Z(n48148) );
  NOR U61050 ( .A(n48149), .B(n48148), .Z(n54487) );
  IV U61051 ( .A(n48150), .Z(n48151) );
  NOR U61052 ( .A(n48154), .B(n48151), .Z(n51833) );
  IV U61053 ( .A(n48152), .Z(n48153) );
  NOR U61054 ( .A(n48154), .B(n48153), .Z(n51839) );
  IV U61055 ( .A(n48155), .Z(n48156) );
  NOR U61056 ( .A(n48162), .B(n48156), .Z(n54476) );
  IV U61057 ( .A(n48157), .Z(n48158) );
  NOR U61058 ( .A(n48159), .B(n48158), .Z(n54478) );
  NOR U61059 ( .A(n54476), .B(n54478), .Z(n50647) );
  IV U61060 ( .A(n48160), .Z(n48161) );
  NOR U61061 ( .A(n48162), .B(n48161), .Z(n48163) );
  IV U61062 ( .A(n48163), .Z(n51854) );
  IV U61063 ( .A(n48164), .Z(n48169) );
  IV U61064 ( .A(n48165), .Z(n48166) );
  NOR U61065 ( .A(n48169), .B(n48166), .Z(n51851) );
  IV U61066 ( .A(n48167), .Z(n48168) );
  NOR U61067 ( .A(n48169), .B(n48168), .Z(n51857) );
  NOR U61068 ( .A(n51864), .B(n51857), .Z(n48170) );
  IV U61069 ( .A(n48170), .Z(n50645) );
  IV U61070 ( .A(n48171), .Z(n48172) );
  NOR U61071 ( .A(n48172), .B(n48176), .Z(n51863) );
  IV U61072 ( .A(n51863), .Z(n51860) );
  IV U61073 ( .A(n48173), .Z(n51876) );
  NOR U61074 ( .A(n51876), .B(n48174), .Z(n48180) );
  IV U61075 ( .A(n48175), .Z(n48179) );
  NOR U61076 ( .A(n48177), .B(n48176), .Z(n48178) );
  IV U61077 ( .A(n48178), .Z(n50641) );
  NOR U61078 ( .A(n48179), .B(n50641), .Z(n51869) );
  NOR U61079 ( .A(n48180), .B(n51869), .Z(n50644) );
  IV U61080 ( .A(n48181), .Z(n48183) );
  NOR U61081 ( .A(n48183), .B(n48182), .Z(n51879) );
  IV U61082 ( .A(n48184), .Z(n48187) );
  NOR U61083 ( .A(n48185), .B(n50633), .Z(n48186) );
  IV U61084 ( .A(n48186), .Z(n48189) );
  NOR U61085 ( .A(n48187), .B(n48189), .Z(n54459) );
  IV U61086 ( .A(n48188), .Z(n48190) );
  NOR U61087 ( .A(n48190), .B(n48189), .Z(n54456) );
  IV U61088 ( .A(n48191), .Z(n50637) );
  IV U61089 ( .A(n48192), .Z(n48193) );
  NOR U61090 ( .A(n50637), .B(n48193), .Z(n48194) );
  IV U61091 ( .A(n48194), .Z(n54451) );
  IV U61092 ( .A(n48195), .Z(n48197) );
  NOR U61093 ( .A(n48197), .B(n48196), .Z(n48201) );
  IV U61094 ( .A(n48198), .Z(n48199) );
  NOR U61095 ( .A(n48199), .B(n50627), .Z(n48200) );
  NOR U61096 ( .A(n48201), .B(n48200), .Z(n54440) );
  IV U61097 ( .A(n48202), .Z(n48204) );
  IV U61098 ( .A(n48203), .Z(n48210) );
  NOR U61099 ( .A(n48204), .B(n48210), .Z(n54436) );
  IV U61100 ( .A(n48205), .Z(n48208) );
  IV U61101 ( .A(n48206), .Z(n48207) );
  NOR U61102 ( .A(n48208), .B(n48207), .Z(n54433) );
  IV U61103 ( .A(n48209), .Z(n48211) );
  NOR U61104 ( .A(n48211), .B(n48210), .Z(n51883) );
  NOR U61105 ( .A(n54433), .B(n51883), .Z(n48212) );
  IV U61106 ( .A(n48212), .Z(n50624) );
  IV U61107 ( .A(n48213), .Z(n48215) );
  IV U61108 ( .A(n48214), .Z(n50592) );
  NOR U61109 ( .A(n48215), .B(n50592), .Z(n51915) );
  IV U61110 ( .A(n48216), .Z(n48217) );
  NOR U61111 ( .A(n48218), .B(n48217), .Z(n54414) );
  NOR U61112 ( .A(n51915), .B(n54414), .Z(n50594) );
  NOR U61113 ( .A(n48220), .B(n48219), .Z(n50585) );
  IV U61114 ( .A(n48221), .Z(n48222) );
  NOR U61115 ( .A(n48223), .B(n48222), .Z(n50582) );
  IV U61116 ( .A(n50582), .Z(n50577) );
  IV U61117 ( .A(n48224), .Z(n48225) );
  NOR U61118 ( .A(n48226), .B(n48225), .Z(n51930) );
  IV U61119 ( .A(n48227), .Z(n48228) );
  NOR U61120 ( .A(n48228), .B(n50570), .Z(n51928) );
  NOR U61121 ( .A(n51930), .B(n51928), .Z(n50565) );
  IV U61122 ( .A(n48229), .Z(n48232) );
  IV U61123 ( .A(n48230), .Z(n48231) );
  NOR U61124 ( .A(n48232), .B(n48231), .Z(n54393) );
  IV U61125 ( .A(n48233), .Z(n48237) );
  IV U61126 ( .A(n48234), .Z(n48245) );
  NOR U61127 ( .A(n48235), .B(n48245), .Z(n48236) );
  IV U61128 ( .A(n48236), .Z(n48240) );
  NOR U61129 ( .A(n48237), .B(n48240), .Z(n48238) );
  IV U61130 ( .A(n48238), .Z(n51937) );
  IV U61131 ( .A(n48239), .Z(n48241) );
  NOR U61132 ( .A(n48241), .B(n48240), .Z(n51933) );
  IV U61133 ( .A(n48242), .Z(n48243) );
  NOR U61134 ( .A(n48243), .B(n48248), .Z(n51944) );
  IV U61135 ( .A(n48244), .Z(n48246) );
  NOR U61136 ( .A(n48246), .B(n48245), .Z(n51940) );
  NOR U61137 ( .A(n51944), .B(n51940), .Z(n50555) );
  IV U61138 ( .A(n48247), .Z(n48249) );
  NOR U61139 ( .A(n48249), .B(n48248), .Z(n50553) );
  IV U61140 ( .A(n50553), .Z(n50543) );
  IV U61141 ( .A(n48250), .Z(n51948) );
  NOR U61142 ( .A(n48251), .B(n51948), .Z(n50542) );
  IV U61143 ( .A(n48252), .Z(n48253) );
  NOR U61144 ( .A(n48253), .B(n48256), .Z(n51951) );
  IV U61145 ( .A(n48254), .Z(n48258) );
  NOR U61146 ( .A(n48256), .B(n48255), .Z(n48257) );
  IV U61147 ( .A(n48257), .Z(n50538) );
  NOR U61148 ( .A(n48258), .B(n50538), .Z(n51954) );
  NOR U61149 ( .A(n48259), .B(n54355), .Z(n50533) );
  IV U61150 ( .A(n48260), .Z(n48261) );
  NOR U61151 ( .A(n48267), .B(n48261), .Z(n51968) );
  IV U61152 ( .A(n48262), .Z(n50521) );
  IV U61153 ( .A(n48263), .Z(n48264) );
  NOR U61154 ( .A(n50521), .B(n48264), .Z(n51974) );
  NOR U61155 ( .A(n51968), .B(n51974), .Z(n50525) );
  IV U61156 ( .A(n48265), .Z(n48266) );
  NOR U61157 ( .A(n48267), .B(n48266), .Z(n51966) );
  IV U61158 ( .A(n48268), .Z(n48269) );
  NOR U61159 ( .A(n48270), .B(n48269), .Z(n50516) );
  IV U61160 ( .A(n50516), .Z(n50512) );
  IV U61161 ( .A(n48271), .Z(n48275) );
  IV U61162 ( .A(n48272), .Z(n50501) );
  NOR U61163 ( .A(n48273), .B(n50501), .Z(n48274) );
  IV U61164 ( .A(n48274), .Z(n50497) );
  NOR U61165 ( .A(n48275), .B(n50497), .Z(n50507) );
  IV U61166 ( .A(n48276), .Z(n50483) );
  IV U61167 ( .A(n48279), .Z(n48277) );
  NOR U61168 ( .A(n50483), .B(n48277), .Z(n54321) );
  IV U61169 ( .A(n48278), .Z(n48281) );
  XOR U61170 ( .A(n50483), .B(n48279), .Z(n48280) );
  NOR U61171 ( .A(n48281), .B(n48280), .Z(n52001) );
  NOR U61172 ( .A(n54321), .B(n52001), .Z(n50480) );
  IV U61173 ( .A(n48282), .Z(n48285) );
  NOR U61174 ( .A(n48283), .B(n50459), .Z(n48284) );
  IV U61175 ( .A(n48284), .Z(n50466) );
  NOR U61176 ( .A(n48285), .B(n50466), .Z(n50469) );
  IV U61177 ( .A(n48286), .Z(n48290) );
  IV U61178 ( .A(n48287), .Z(n50448) );
  NOR U61179 ( .A(n50448), .B(n48288), .Z(n48289) );
  IV U61180 ( .A(n48289), .Z(n50454) );
  NOR U61181 ( .A(n48290), .B(n50454), .Z(n50451) );
  IV U61182 ( .A(n50451), .Z(n50440) );
  IV U61183 ( .A(n48291), .Z(n48292) );
  NOR U61184 ( .A(n48293), .B(n48292), .Z(n48294) );
  IV U61185 ( .A(n48294), .Z(n54289) );
  IV U61186 ( .A(n48295), .Z(n48296) );
  NOR U61187 ( .A(n48296), .B(n48298), .Z(n54277) );
  IV U61188 ( .A(n48297), .Z(n48299) );
  NOR U61189 ( .A(n48299), .B(n48298), .Z(n52021) );
  NOR U61190 ( .A(n54277), .B(n52021), .Z(n50412) );
  IV U61191 ( .A(n48300), .Z(n48302) );
  NOR U61192 ( .A(n48302), .B(n48301), .Z(n54278) );
  IV U61193 ( .A(n48303), .Z(n48305) );
  IV U61194 ( .A(n48304), .Z(n48309) );
  NOR U61195 ( .A(n48305), .B(n48309), .Z(n54274) );
  NOR U61196 ( .A(n48307), .B(n48306), .Z(n52028) );
  IV U61197 ( .A(n48308), .Z(n48310) );
  NOR U61198 ( .A(n48310), .B(n48309), .Z(n54271) );
  NOR U61199 ( .A(n52028), .B(n54271), .Z(n48311) );
  IV U61200 ( .A(n48311), .Z(n50406) );
  IV U61201 ( .A(n48312), .Z(n48313) );
  NOR U61202 ( .A(n48313), .B(n50404), .Z(n52024) );
  IV U61203 ( .A(n48314), .Z(n50397) );
  IV U61204 ( .A(n48315), .Z(n48316) );
  NOR U61205 ( .A(n50397), .B(n48316), .Z(n54258) );
  IV U61206 ( .A(n48317), .Z(n48318) );
  NOR U61207 ( .A(n48318), .B(n48322), .Z(n52036) );
  IV U61208 ( .A(n48319), .Z(n52044) );
  NOR U61209 ( .A(n48320), .B(n52044), .Z(n48324) );
  IV U61210 ( .A(n48321), .Z(n48323) );
  NOR U61211 ( .A(n48323), .B(n48322), .Z(n52040) );
  NOR U61212 ( .A(n48324), .B(n52040), .Z(n50394) );
  IV U61213 ( .A(n48325), .Z(n48326) );
  NOR U61214 ( .A(n50389), .B(n48326), .Z(n50392) );
  IV U61215 ( .A(n50392), .Z(n50384) );
  IV U61216 ( .A(n48327), .Z(n48328) );
  NOR U61217 ( .A(n50364), .B(n48328), .Z(n52065) );
  IV U61218 ( .A(n48329), .Z(n48331) );
  NOR U61219 ( .A(n48331), .B(n48330), .Z(n52067) );
  IV U61220 ( .A(n48332), .Z(n48335) );
  NOR U61221 ( .A(n48333), .B(n50356), .Z(n48334) );
  IV U61222 ( .A(n48334), .Z(n48337) );
  NOR U61223 ( .A(n48335), .B(n48337), .Z(n52073) );
  IV U61224 ( .A(n48336), .Z(n48338) );
  NOR U61225 ( .A(n48338), .B(n48337), .Z(n52070) );
  NOR U61226 ( .A(n48340), .B(n48339), .Z(n48345) );
  IV U61227 ( .A(n48341), .Z(n48343) );
  IV U61228 ( .A(n48342), .Z(n50353) );
  NOR U61229 ( .A(n48343), .B(n50353), .Z(n48344) );
  NOR U61230 ( .A(n48345), .B(n48344), .Z(n57576) );
  IV U61231 ( .A(n48346), .Z(n48348) );
  IV U61232 ( .A(n48347), .Z(n50348) );
  NOR U61233 ( .A(n48348), .B(n50348), .Z(n54239) );
  IV U61234 ( .A(n48349), .Z(n48350) );
  NOR U61235 ( .A(n48350), .B(n50345), .Z(n48355) );
  IV U61236 ( .A(n48351), .Z(n48353) );
  IV U61237 ( .A(n48352), .Z(n48361) );
  NOR U61238 ( .A(n48353), .B(n48361), .Z(n48354) );
  NOR U61239 ( .A(n48355), .B(n48354), .Z(n52089) );
  IV U61240 ( .A(n52089), .Z(n50343) );
  IV U61241 ( .A(n48356), .Z(n48358) );
  NOR U61242 ( .A(n48358), .B(n48357), .Z(n54229) );
  IV U61243 ( .A(n48359), .Z(n48360) );
  NOR U61244 ( .A(n48361), .B(n48360), .Z(n52091) );
  NOR U61245 ( .A(n54229), .B(n52091), .Z(n50342) );
  IV U61246 ( .A(n48362), .Z(n48363) );
  NOR U61247 ( .A(n48363), .B(n48366), .Z(n54232) );
  IV U61248 ( .A(n48364), .Z(n48365) );
  NOR U61249 ( .A(n48366), .B(n48365), .Z(n52095) );
  IV U61250 ( .A(n48367), .Z(n48368) );
  NOR U61251 ( .A(n48369), .B(n48368), .Z(n54226) );
  NOR U61252 ( .A(n52095), .B(n54226), .Z(n48370) );
  IV U61253 ( .A(n48370), .Z(n48371) );
  NOR U61254 ( .A(n54232), .B(n48371), .Z(n50341) );
  IV U61255 ( .A(n48372), .Z(n48379) );
  IV U61256 ( .A(n48373), .Z(n48374) );
  NOR U61257 ( .A(n48379), .B(n48374), .Z(n54223) );
  IV U61258 ( .A(n48375), .Z(n48376) );
  NOR U61259 ( .A(n48379), .B(n48376), .Z(n52100) );
  IV U61260 ( .A(n48377), .Z(n48378) );
  NOR U61261 ( .A(n48379), .B(n48378), .Z(n52097) );
  IV U61262 ( .A(n48380), .Z(n48382) );
  NOR U61263 ( .A(n48382), .B(n48381), .Z(n52111) );
  IV U61264 ( .A(n48383), .Z(n48389) );
  IV U61265 ( .A(n48384), .Z(n48385) );
  NOR U61266 ( .A(n48386), .B(n48385), .Z(n48387) );
  IV U61267 ( .A(n48387), .Z(n48388) );
  NOR U61268 ( .A(n48389), .B(n48388), .Z(n52106) );
  IV U61269 ( .A(n48390), .Z(n48391) );
  NOR U61270 ( .A(n48391), .B(n48395), .Z(n48392) );
  IV U61271 ( .A(n48392), .Z(n52119) );
  IV U61272 ( .A(n48393), .Z(n48394) );
  NOR U61273 ( .A(n48395), .B(n48394), .Z(n54215) );
  IV U61274 ( .A(n48396), .Z(n48399) );
  IV U61275 ( .A(n48397), .Z(n48398) );
  NOR U61276 ( .A(n48399), .B(n48398), .Z(n52129) );
  IV U61277 ( .A(n52129), .Z(n52126) );
  NOR U61278 ( .A(n48400), .B(n54197), .Z(n48401) );
  IV U61279 ( .A(n48401), .Z(n54203) );
  IV U61280 ( .A(n48402), .Z(n48405) );
  IV U61281 ( .A(n48403), .Z(n48404) );
  NOR U61282 ( .A(n48405), .B(n48404), .Z(n54178) );
  IV U61283 ( .A(n48406), .Z(n48407) );
  NOR U61284 ( .A(n48407), .B(n54197), .Z(n54193) );
  NOR U61285 ( .A(n54178), .B(n54193), .Z(n48408) );
  IV U61286 ( .A(n48408), .Z(n50316) );
  IV U61287 ( .A(n48409), .Z(n48410) );
  NOR U61288 ( .A(n48411), .B(n48410), .Z(n50313) );
  IV U61289 ( .A(n50313), .Z(n50300) );
  IV U61290 ( .A(n48412), .Z(n48417) );
  IV U61291 ( .A(n48413), .Z(n48414) );
  NOR U61292 ( .A(n48417), .B(n48414), .Z(n54160) );
  IV U61293 ( .A(n48415), .Z(n48416) );
  NOR U61294 ( .A(n48417), .B(n48416), .Z(n54163) );
  IV U61295 ( .A(n48418), .Z(n48419) );
  NOR U61296 ( .A(n48419), .B(n48422), .Z(n54155) );
  NOR U61297 ( .A(n54163), .B(n54155), .Z(n48420) );
  IV U61298 ( .A(n48420), .Z(n50292) );
  IV U61299 ( .A(n48421), .Z(n48425) );
  NOR U61300 ( .A(n48423), .B(n48422), .Z(n48424) );
  IV U61301 ( .A(n48424), .Z(n52139) );
  NOR U61302 ( .A(n48425), .B(n52139), .Z(n52137) );
  IV U61303 ( .A(n48426), .Z(n48427) );
  NOR U61304 ( .A(n48427), .B(n52139), .Z(n54148) );
  IV U61305 ( .A(n48428), .Z(n48429) );
  NOR U61306 ( .A(n48432), .B(n48429), .Z(n52154) );
  IV U61307 ( .A(n48430), .Z(n48431) );
  NOR U61308 ( .A(n48432), .B(n48431), .Z(n52146) );
  XOR U61309 ( .A(n52154), .B(n52146), .Z(n48433) );
  NOR U61310 ( .A(n52149), .B(n48433), .Z(n48434) );
  IV U61311 ( .A(n48434), .Z(n50288) );
  IV U61312 ( .A(n48435), .Z(n48440) );
  IV U61313 ( .A(n48436), .Z(n48437) );
  NOR U61314 ( .A(n48438), .B(n48437), .Z(n48439) );
  IV U61315 ( .A(n48439), .Z(n48442) );
  NOR U61316 ( .A(n48440), .B(n48442), .Z(n52151) );
  IV U61317 ( .A(n48441), .Z(n48443) );
  NOR U61318 ( .A(n48443), .B(n48442), .Z(n52162) );
  IV U61319 ( .A(n48444), .Z(n48449) );
  IV U61320 ( .A(n48445), .Z(n48446) );
  NOR U61321 ( .A(n48447), .B(n48446), .Z(n48448) );
  IV U61322 ( .A(n48448), .Z(n48451) );
  NOR U61323 ( .A(n48449), .B(n48451), .Z(n52159) );
  IV U61324 ( .A(n48450), .Z(n48452) );
  NOR U61325 ( .A(n48452), .B(n48451), .Z(n52167) );
  NOR U61326 ( .A(n52169), .B(n52167), .Z(n50286) );
  IV U61327 ( .A(n48453), .Z(n48455) );
  NOR U61328 ( .A(n48455), .B(n48454), .Z(n50272) );
  IV U61329 ( .A(n48456), .Z(n48457) );
  NOR U61330 ( .A(n48458), .B(n48457), .Z(n54116) );
  IV U61331 ( .A(n48459), .Z(n48460) );
  NOR U61332 ( .A(n48461), .B(n48460), .Z(n54121) );
  NOR U61333 ( .A(n54116), .B(n54121), .Z(n50263) );
  NOR U61334 ( .A(n48462), .B(n52193), .Z(n48463) );
  NOR U61335 ( .A(n48464), .B(n48463), .Z(n50262) );
  NOR U61336 ( .A(n48465), .B(n52201), .Z(n50261) );
  IV U61337 ( .A(n48466), .Z(n50258) );
  IV U61338 ( .A(n48467), .Z(n48468) );
  NOR U61339 ( .A(n50258), .B(n48468), .Z(n52217) );
  IV U61340 ( .A(n48469), .Z(n48471) );
  NOR U61341 ( .A(n48471), .B(n48470), .Z(n52214) );
  IV U61342 ( .A(n48472), .Z(n48473) );
  NOR U61343 ( .A(n48474), .B(n48473), .Z(n52222) );
  IV U61344 ( .A(n48475), .Z(n48477) );
  NOR U61345 ( .A(n48477), .B(n48476), .Z(n52232) );
  IV U61346 ( .A(n48478), .Z(n48479) );
  NOR U61347 ( .A(n48479), .B(n50251), .Z(n52230) );
  NOR U61348 ( .A(n52232), .B(n52230), .Z(n48480) );
  IV U61349 ( .A(n48480), .Z(n50249) );
  IV U61350 ( .A(n48481), .Z(n48482) );
  NOR U61351 ( .A(n48483), .B(n48482), .Z(n48489) );
  IV U61352 ( .A(n48484), .Z(n48487) );
  IV U61353 ( .A(n48485), .Z(n48486) );
  NOR U61354 ( .A(n48487), .B(n48486), .Z(n48488) );
  NOR U61355 ( .A(n48489), .B(n48488), .Z(n52245) );
  IV U61356 ( .A(n48490), .Z(n48491) );
  NOR U61357 ( .A(n48493), .B(n48491), .Z(n52241) );
  NOR U61358 ( .A(n48493), .B(n48492), .Z(n52248) );
  IV U61359 ( .A(n48494), .Z(n48495) );
  NOR U61360 ( .A(n48496), .B(n48495), .Z(n52250) );
  NOR U61361 ( .A(n52248), .B(n52250), .Z(n50241) );
  IV U61362 ( .A(n48497), .Z(n48500) );
  NOR U61363 ( .A(n48498), .B(n48505), .Z(n48499) );
  IV U61364 ( .A(n48499), .Z(n48508) );
  NOR U61365 ( .A(n48500), .B(n48508), .Z(n54103) );
  IV U61366 ( .A(n48501), .Z(n48503) );
  NOR U61367 ( .A(n48503), .B(n48502), .Z(n54096) );
  NOR U61368 ( .A(n48505), .B(n48504), .Z(n52260) );
  NOR U61369 ( .A(n54096), .B(n52260), .Z(n48506) );
  XOR U61370 ( .A(n54103), .B(n48506), .Z(n50230) );
  IV U61371 ( .A(n48507), .Z(n48509) );
  NOR U61372 ( .A(n48509), .B(n48508), .Z(n48510) );
  IV U61373 ( .A(n48510), .Z(n52258) );
  IV U61374 ( .A(n48511), .Z(n48513) );
  NOR U61375 ( .A(n48513), .B(n48512), .Z(n52263) );
  IV U61376 ( .A(n48514), .Z(n48515) );
  NOR U61377 ( .A(n48515), .B(n48517), .Z(n54093) );
  IV U61378 ( .A(n48516), .Z(n48518) );
  NOR U61379 ( .A(n48518), .B(n48517), .Z(n54089) );
  IV U61380 ( .A(n48519), .Z(n48520) );
  NOR U61381 ( .A(n48521), .B(n48520), .Z(n52265) );
  NOR U61382 ( .A(n54089), .B(n52265), .Z(n48522) );
  IV U61383 ( .A(n48522), .Z(n48523) );
  NOR U61384 ( .A(n54093), .B(n48523), .Z(n48524) );
  IV U61385 ( .A(n48524), .Z(n50228) );
  IV U61386 ( .A(n48525), .Z(n48526) );
  NOR U61387 ( .A(n48527), .B(n48526), .Z(n52270) );
  IV U61388 ( .A(n48528), .Z(n48531) );
  IV U61389 ( .A(n48529), .Z(n48530) );
  NOR U61390 ( .A(n48531), .B(n48530), .Z(n52267) );
  IV U61391 ( .A(n48532), .Z(n48533) );
  NOR U61392 ( .A(n48535), .B(n48533), .Z(n54084) );
  NOR U61393 ( .A(n48535), .B(n48534), .Z(n54081) );
  IV U61394 ( .A(n48536), .Z(n48539) );
  NOR U61395 ( .A(n50222), .B(n48537), .Z(n48538) );
  IV U61396 ( .A(n48538), .Z(n48544) );
  NOR U61397 ( .A(n48539), .B(n48544), .Z(n52280) );
  IV U61398 ( .A(n48540), .Z(n48542) );
  NOR U61399 ( .A(n48542), .B(n48541), .Z(n52275) );
  IV U61400 ( .A(n48543), .Z(n48545) );
  NOR U61401 ( .A(n48545), .B(n48544), .Z(n52277) );
  IV U61402 ( .A(n48546), .Z(n48549) );
  NOR U61403 ( .A(n48547), .B(n50217), .Z(n48548) );
  IV U61404 ( .A(n48548), .Z(n50214) );
  NOR U61405 ( .A(n48549), .B(n50214), .Z(n48550) );
  IV U61406 ( .A(n48550), .Z(n52290) );
  IV U61407 ( .A(n48551), .Z(n48557) );
  IV U61408 ( .A(n48552), .Z(n48553) );
  NOR U61409 ( .A(n48557), .B(n48553), .Z(n48554) );
  IV U61410 ( .A(n48554), .Z(n52292) );
  IV U61411 ( .A(n48555), .Z(n48556) );
  NOR U61412 ( .A(n48557), .B(n48556), .Z(n52293) );
  IV U61413 ( .A(n48558), .Z(n48559) );
  NOR U61414 ( .A(n48560), .B(n48559), .Z(n52299) );
  IV U61415 ( .A(n48561), .Z(n48564) );
  IV U61416 ( .A(n48562), .Z(n48563) );
  NOR U61417 ( .A(n48564), .B(n48563), .Z(n52296) );
  IV U61418 ( .A(n48565), .Z(n48566) );
  NOR U61419 ( .A(n48573), .B(n48566), .Z(n52309) );
  NOR U61420 ( .A(n52307), .B(n52309), .Z(n48567) );
  IV U61421 ( .A(n48567), .Z(n50211) );
  IV U61422 ( .A(n48568), .Z(n48569) );
  NOR U61423 ( .A(n48570), .B(n48569), .Z(n52304) );
  IV U61424 ( .A(n48571), .Z(n48572) );
  NOR U61425 ( .A(n48573), .B(n48572), .Z(n52310) );
  IV U61426 ( .A(n48574), .Z(n48575) );
  NOR U61427 ( .A(n48575), .B(n50202), .Z(n52316) );
  IV U61428 ( .A(n48576), .Z(n48581) );
  IV U61429 ( .A(n48577), .Z(n48578) );
  NOR U61430 ( .A(n48581), .B(n48578), .Z(n52323) );
  NOR U61431 ( .A(n52316), .B(n52323), .Z(n50201) );
  IV U61432 ( .A(n48579), .Z(n48580) );
  NOR U61433 ( .A(n48581), .B(n48580), .Z(n52320) );
  IV U61434 ( .A(n48582), .Z(n48584) );
  NOR U61435 ( .A(n48584), .B(n48583), .Z(n52331) );
  IV U61436 ( .A(n48585), .Z(n48586) );
  NOR U61437 ( .A(n48586), .B(n50198), .Z(n52328) );
  IV U61438 ( .A(n48587), .Z(n48588) );
  NOR U61439 ( .A(n48589), .B(n48588), .Z(n52346) );
  IV U61440 ( .A(n48590), .Z(n48593) );
  IV U61441 ( .A(n48591), .Z(n48592) );
  NOR U61442 ( .A(n48593), .B(n48592), .Z(n52350) );
  NOR U61443 ( .A(n52346), .B(n52350), .Z(n50186) );
  IV U61444 ( .A(n48594), .Z(n48596) );
  NOR U61445 ( .A(n48596), .B(n48595), .Z(n48597) );
  IV U61446 ( .A(n48597), .Z(n52345) );
  IV U61447 ( .A(n48598), .Z(n48599) );
  NOR U61448 ( .A(n48600), .B(n48599), .Z(n52370) );
  IV U61449 ( .A(n48601), .Z(n48602) );
  NOR U61450 ( .A(n50174), .B(n48602), .Z(n52367) );
  NOR U61451 ( .A(n52370), .B(n52367), .Z(n50178) );
  IV U61452 ( .A(n48603), .Z(n48604) );
  NOR U61453 ( .A(n48604), .B(n48606), .Z(n52372) );
  IV U61454 ( .A(n48605), .Z(n48607) );
  NOR U61455 ( .A(n48607), .B(n48606), .Z(n52383) );
  IV U61456 ( .A(n48608), .Z(n48611) );
  NOR U61457 ( .A(n48614), .B(n48609), .Z(n48610) );
  IV U61458 ( .A(n48610), .Z(n50164) );
  NOR U61459 ( .A(n48611), .B(n50164), .Z(n54061) );
  IV U61460 ( .A(n48612), .Z(n48613) );
  NOR U61461 ( .A(n48614), .B(n48613), .Z(n52386) );
  IV U61462 ( .A(n48615), .Z(n48617) );
  NOR U61463 ( .A(n48617), .B(n48616), .Z(n54057) );
  NOR U61464 ( .A(n52386), .B(n54057), .Z(n48618) );
  IV U61465 ( .A(n48618), .Z(n50162) );
  IV U61466 ( .A(n48619), .Z(n48624) );
  IV U61467 ( .A(n48620), .Z(n48621) );
  NOR U61468 ( .A(n48622), .B(n48621), .Z(n48623) );
  IV U61469 ( .A(n48623), .Z(n50159) );
  NOR U61470 ( .A(n48624), .B(n50159), .Z(n54053) );
  NOR U61471 ( .A(n48626), .B(n48625), .Z(n54045) );
  IV U61472 ( .A(n48627), .Z(n48628) );
  NOR U61473 ( .A(n48628), .B(n50152), .Z(n50156) );
  IV U61474 ( .A(n50156), .Z(n50146) );
  IV U61475 ( .A(n48629), .Z(n48630) );
  NOR U61476 ( .A(n48630), .B(n50138), .Z(n52395) );
  IV U61477 ( .A(n48631), .Z(n48636) );
  IV U61478 ( .A(n48632), .Z(n48633) );
  NOR U61479 ( .A(n48636), .B(n48633), .Z(n52392) );
  IV U61480 ( .A(n48634), .Z(n48635) );
  NOR U61481 ( .A(n48636), .B(n48635), .Z(n54012) );
  IV U61482 ( .A(n48637), .Z(n48640) );
  NOR U61483 ( .A(n48638), .B(n50132), .Z(n48639) );
  IV U61484 ( .A(n48639), .Z(n50129) );
  NOR U61485 ( .A(n48640), .B(n50129), .Z(n53998) );
  IV U61486 ( .A(n48641), .Z(n48644) );
  IV U61487 ( .A(n48642), .Z(n48643) );
  NOR U61488 ( .A(n48644), .B(n48643), .Z(n52399) );
  IV U61489 ( .A(n48645), .Z(n52403) );
  NOR U61490 ( .A(n48646), .B(n52403), .Z(n48647) );
  NOR U61491 ( .A(n52399), .B(n48647), .Z(n48648) );
  IV U61492 ( .A(n48648), .Z(n50127) );
  IV U61493 ( .A(n48649), .Z(n48650) );
  NOR U61494 ( .A(n48650), .B(n50124), .Z(n48651) );
  IV U61495 ( .A(n48651), .Z(n52417) );
  IV U61496 ( .A(n48652), .Z(n48654) );
  IV U61497 ( .A(n48653), .Z(n50108) );
  NOR U61498 ( .A(n48654), .B(n50108), .Z(n52424) );
  IV U61499 ( .A(n48655), .Z(n48656) );
  NOR U61500 ( .A(n48657), .B(n48656), .Z(n52427) );
  NOR U61501 ( .A(n48659), .B(n48658), .Z(n53986) );
  NOR U61502 ( .A(n52427), .B(n53986), .Z(n48660) );
  IV U61503 ( .A(n48660), .Z(n50103) );
  IV U61504 ( .A(n48661), .Z(n48663) );
  NOR U61505 ( .A(n48663), .B(n48662), .Z(n50098) );
  IV U61506 ( .A(n48664), .Z(n48670) );
  NOR U61507 ( .A(n48665), .B(n50092), .Z(n48666) );
  IV U61508 ( .A(n48666), .Z(n48667) );
  NOR U61509 ( .A(n48668), .B(n48667), .Z(n48669) );
  IV U61510 ( .A(n48669), .Z(n50094) );
  NOR U61511 ( .A(n48670), .B(n50094), .Z(n52429) );
  IV U61512 ( .A(n48671), .Z(n48672) );
  NOR U61513 ( .A(n48673), .B(n48672), .Z(n48678) );
  IV U61514 ( .A(n48674), .Z(n48675) );
  NOR U61515 ( .A(n48676), .B(n48675), .Z(n48677) );
  NOR U61516 ( .A(n48678), .B(n48677), .Z(n52443) );
  IV U61517 ( .A(n48679), .Z(n48682) );
  IV U61518 ( .A(n48680), .Z(n48681) );
  NOR U61519 ( .A(n48682), .B(n48681), .Z(n52439) );
  IV U61520 ( .A(n48683), .Z(n48684) );
  NOR U61521 ( .A(n50083), .B(n48684), .Z(n48685) );
  IV U61522 ( .A(n48685), .Z(n52446) );
  IV U61523 ( .A(n48686), .Z(n48688) );
  IV U61524 ( .A(n48687), .Z(n48693) );
  NOR U61525 ( .A(n48688), .B(n48693), .Z(n48689) );
  IV U61526 ( .A(n48689), .Z(n52460) );
  NOR U61527 ( .A(n48691), .B(n48690), .Z(n53967) );
  IV U61528 ( .A(n48692), .Z(n48694) );
  NOR U61529 ( .A(n48694), .B(n48693), .Z(n52465) );
  NOR U61530 ( .A(n53967), .B(n52465), .Z(n50073) );
  IV U61531 ( .A(n48695), .Z(n48697) );
  NOR U61532 ( .A(n48697), .B(n48696), .Z(n52473) );
  IV U61533 ( .A(n48698), .Z(n48699) );
  NOR U61534 ( .A(n50064), .B(n48699), .Z(n53959) );
  IV U61535 ( .A(n48700), .Z(n48704) );
  IV U61536 ( .A(n48701), .Z(n48702) );
  NOR U61537 ( .A(n48704), .B(n48702), .Z(n52476) );
  NOR U61538 ( .A(n53959), .B(n52476), .Z(n50060) );
  IV U61539 ( .A(n48703), .Z(n48705) );
  NOR U61540 ( .A(n48705), .B(n48704), .Z(n52478) );
  NOR U61541 ( .A(n48706), .B(n50057), .Z(n48707) );
  IV U61542 ( .A(n48707), .Z(n48708) );
  NOR U61543 ( .A(n48709), .B(n48708), .Z(n53947) );
  IV U61544 ( .A(n48710), .Z(n48711) );
  NOR U61545 ( .A(n50038), .B(n48711), .Z(n48712) );
  IV U61546 ( .A(n48712), .Z(n48717) );
  NOR U61547 ( .A(n48714), .B(n48713), .Z(n48715) );
  IV U61548 ( .A(n48715), .Z(n48716) );
  NOR U61549 ( .A(n48717), .B(n48716), .Z(n48718) );
  IV U61550 ( .A(n48718), .Z(n53933) );
  IV U61551 ( .A(n48719), .Z(n48720) );
  NOR U61552 ( .A(n48728), .B(n48720), .Z(n48725) );
  IV U61553 ( .A(n48721), .Z(n48723) );
  IV U61554 ( .A(n48722), .Z(n49986) );
  NOR U61555 ( .A(n48723), .B(n49986), .Z(n48724) );
  NOR U61556 ( .A(n48725), .B(n48724), .Z(n53912) );
  IV U61557 ( .A(n48727), .Z(n48726) );
  NOR U61558 ( .A(n48728), .B(n48726), .Z(n48733) );
  XOR U61559 ( .A(n48728), .B(n48727), .Z(n48731) );
  IV U61560 ( .A(n48729), .Z(n48730) );
  NOR U61561 ( .A(n48731), .B(n48730), .Z(n48732) );
  NOR U61562 ( .A(n48733), .B(n48732), .Z(n53909) );
  IV U61563 ( .A(n48734), .Z(n48735) );
  NOR U61564 ( .A(n48741), .B(n48735), .Z(n53899) );
  IV U61565 ( .A(n48736), .Z(n48737) );
  NOR U61566 ( .A(n48737), .B(n48745), .Z(n52502) );
  IV U61567 ( .A(n48738), .Z(n48739) );
  NOR U61568 ( .A(n48741), .B(n48739), .Z(n53902) );
  NOR U61569 ( .A(n48741), .B(n48740), .Z(n52500) );
  NOR U61570 ( .A(n53902), .B(n52500), .Z(n48742) );
  IV U61571 ( .A(n48742), .Z(n48743) );
  NOR U61572 ( .A(n52502), .B(n48743), .Z(n48744) );
  IV U61573 ( .A(n48744), .Z(n49984) );
  NOR U61574 ( .A(n48746), .B(n48745), .Z(n48747) );
  IV U61575 ( .A(n48747), .Z(n52509) );
  NOR U61576 ( .A(n52509), .B(n48748), .Z(n49983) );
  IV U61577 ( .A(n48749), .Z(n48753) );
  IV U61578 ( .A(n48750), .Z(n48759) );
  NOR U61579 ( .A(n48759), .B(n48751), .Z(n48752) );
  IV U61580 ( .A(n48752), .Z(n48755) );
  NOR U61581 ( .A(n48753), .B(n48755), .Z(n52505) );
  IV U61582 ( .A(n48754), .Z(n48756) );
  NOR U61583 ( .A(n48756), .B(n48755), .Z(n52518) );
  IV U61584 ( .A(n48757), .Z(n48761) );
  NOR U61585 ( .A(n48759), .B(n48758), .Z(n48760) );
  IV U61586 ( .A(n48760), .Z(n48763) );
  NOR U61587 ( .A(n48761), .B(n48763), .Z(n52515) );
  IV U61588 ( .A(n48762), .Z(n48764) );
  NOR U61589 ( .A(n48764), .B(n48763), .Z(n52524) );
  IV U61590 ( .A(n48765), .Z(n48766) );
  NOR U61591 ( .A(n49982), .B(n48766), .Z(n52528) );
  IV U61592 ( .A(n48767), .Z(n48769) );
  IV U61593 ( .A(n48768), .Z(n48771) );
  NOR U61594 ( .A(n48769), .B(n48771), .Z(n52532) );
  NOR U61595 ( .A(n52528), .B(n52532), .Z(n49979) );
  IV U61596 ( .A(n48770), .Z(n48774) );
  NOR U61597 ( .A(n48772), .B(n48771), .Z(n48773) );
  IV U61598 ( .A(n48773), .Z(n49973) );
  NOR U61599 ( .A(n48774), .B(n49973), .Z(n53887) );
  NOR U61600 ( .A(n48775), .B(n52535), .Z(n48776) );
  IV U61601 ( .A(n48776), .Z(n53879) );
  NOR U61602 ( .A(n53850), .B(n48777), .Z(n49949) );
  IV U61603 ( .A(n48778), .Z(n48779) );
  NOR U61604 ( .A(n48779), .B(n48782), .Z(n52556) );
  IV U61605 ( .A(n48780), .Z(n48781) );
  NOR U61606 ( .A(n48781), .B(n48782), .Z(n52559) );
  NOR U61607 ( .A(n48783), .B(n48782), .Z(n52564) );
  IV U61608 ( .A(n48784), .Z(n48785) );
  NOR U61609 ( .A(n48786), .B(n48785), .Z(n53836) );
  NOR U61610 ( .A(n52564), .B(n53836), .Z(n48787) );
  IV U61611 ( .A(n48787), .Z(n48788) );
  NOR U61612 ( .A(n52559), .B(n48788), .Z(n49926) );
  IV U61613 ( .A(n48789), .Z(n48790) );
  NOR U61614 ( .A(n48791), .B(n48790), .Z(n52567) );
  IV U61615 ( .A(n48792), .Z(n48793) );
  NOR U61616 ( .A(n48795), .B(n48793), .Z(n53813) );
  IV U61617 ( .A(n48794), .Z(n48796) );
  NOR U61618 ( .A(n48796), .B(n48795), .Z(n52573) );
  IV U61619 ( .A(n48797), .Z(n48803) );
  IV U61620 ( .A(n48798), .Z(n48800) );
  NOR U61621 ( .A(n48800), .B(n48799), .Z(n48801) );
  IV U61622 ( .A(n48801), .Z(n48802) );
  NOR U61623 ( .A(n48803), .B(n48802), .Z(n52580) );
  NOR U61624 ( .A(n52573), .B(n52580), .Z(n48804) );
  IV U61625 ( .A(n48804), .Z(n49918) );
  IV U61626 ( .A(n48805), .Z(n48817) );
  IV U61627 ( .A(n48806), .Z(n48807) );
  NOR U61628 ( .A(n48808), .B(n48807), .Z(n48812) );
  XOR U61629 ( .A(n49901), .B(n49902), .Z(n48822) );
  NOR U61630 ( .A(n48809), .B(n48822), .Z(n48810) );
  IV U61631 ( .A(n48810), .Z(n48811) );
  NOR U61632 ( .A(n48812), .B(n48811), .Z(n48813) );
  IV U61633 ( .A(n48813), .Z(n48814) );
  NOR U61634 ( .A(n48815), .B(n48814), .Z(n48816) );
  IV U61635 ( .A(n48816), .Z(n48819) );
  NOR U61636 ( .A(n48817), .B(n48819), .Z(n52579) );
  IV U61637 ( .A(n48818), .Z(n48820) );
  NOR U61638 ( .A(n48820), .B(n48819), .Z(n52591) );
  IV U61639 ( .A(n48821), .Z(n48823) );
  NOR U61640 ( .A(n48823), .B(n48822), .Z(n52588) );
  IV U61641 ( .A(n48824), .Z(n48827) );
  NOR U61642 ( .A(n48825), .B(n49902), .Z(n48826) );
  IV U61643 ( .A(n48826), .Z(n49915) );
  NOR U61644 ( .A(n48827), .B(n49915), .Z(n49906) );
  IV U61645 ( .A(n48828), .Z(n48829) );
  NOR U61646 ( .A(n48829), .B(n53783), .Z(n53780) );
  NOR U61647 ( .A(n53776), .B(n48830), .Z(n48831) );
  NOR U61648 ( .A(n53783), .B(n48831), .Z(n49871) );
  NOR U61649 ( .A(n48833), .B(n48832), .Z(n52622) );
  IV U61650 ( .A(n48834), .Z(n52619) );
  NOR U61651 ( .A(n48835), .B(n52619), .Z(n48836) );
  NOR U61652 ( .A(n52622), .B(n48836), .Z(n48837) );
  IV U61653 ( .A(n48837), .Z(n49870) );
  IV U61654 ( .A(n48838), .Z(n48840) );
  NOR U61655 ( .A(n48840), .B(n48839), .Z(n52628) );
  IV U61656 ( .A(n48841), .Z(n48843) );
  NOR U61657 ( .A(n48843), .B(n48842), .Z(n52626) );
  NOR U61658 ( .A(n52628), .B(n52626), .Z(n49869) );
  IV U61659 ( .A(n48844), .Z(n48845) );
  NOR U61660 ( .A(n48846), .B(n48845), .Z(n53766) );
  IV U61661 ( .A(n48847), .Z(n48848) );
  NOR U61662 ( .A(n48848), .B(n48853), .Z(n53759) );
  NOR U61663 ( .A(n53766), .B(n53759), .Z(n49868) );
  IV U61664 ( .A(n48849), .Z(n48850) );
  NOR U61665 ( .A(n48851), .B(n48850), .Z(n52635) );
  IV U61666 ( .A(n48852), .Z(n48859) );
  NOR U61667 ( .A(n48854), .B(n48853), .Z(n48855) );
  IV U61668 ( .A(n48855), .Z(n48856) );
  NOR U61669 ( .A(n48857), .B(n48856), .Z(n48858) );
  IV U61670 ( .A(n48858), .Z(n49866) );
  NOR U61671 ( .A(n48859), .B(n49866), .Z(n53755) );
  NOR U61672 ( .A(n52635), .B(n53755), .Z(n49864) );
  IV U61673 ( .A(n48863), .Z(n48860) );
  NOR U61674 ( .A(n48861), .B(n48860), .Z(n48867) );
  NOR U61675 ( .A(n48863), .B(n48862), .Z(n48864) );
  NOR U61676 ( .A(n48865), .B(n48864), .Z(n48866) );
  NOR U61677 ( .A(n48867), .B(n48866), .Z(n48868) );
  IV U61678 ( .A(n48868), .Z(n52636) );
  IV U61679 ( .A(n48869), .Z(n48870) );
  NOR U61680 ( .A(n48870), .B(n48875), .Z(n53752) );
  IV U61681 ( .A(n48871), .Z(n48872) );
  NOR U61682 ( .A(n49854), .B(n48872), .Z(n52638) );
  NOR U61683 ( .A(n53752), .B(n52638), .Z(n48873) );
  IV U61684 ( .A(n48873), .Z(n49858) );
  IV U61685 ( .A(n48874), .Z(n48876) );
  NOR U61686 ( .A(n48876), .B(n48875), .Z(n49851) );
  IV U61687 ( .A(n49851), .Z(n49845) );
  IV U61688 ( .A(n48877), .Z(n48879) );
  IV U61689 ( .A(n48878), .Z(n48881) );
  NOR U61690 ( .A(n48879), .B(n48881), .Z(n52651) );
  IV U61691 ( .A(n48880), .Z(n48882) );
  NOR U61692 ( .A(n48882), .B(n48881), .Z(n52648) );
  IV U61693 ( .A(n48883), .Z(n48884) );
  NOR U61694 ( .A(n48884), .B(n49841), .Z(n48885) );
  IV U61695 ( .A(n48885), .Z(n52656) );
  IV U61696 ( .A(n48886), .Z(n48888) );
  NOR U61697 ( .A(n48888), .B(n48887), .Z(n53744) );
  NOR U61698 ( .A(n53738), .B(n53744), .Z(n49835) );
  IV U61699 ( .A(n48889), .Z(n48890) );
  NOR U61700 ( .A(n48890), .B(n49830), .Z(n48891) );
  IV U61701 ( .A(n48891), .Z(n53726) );
  IV U61702 ( .A(n48892), .Z(n48893) );
  NOR U61703 ( .A(n48894), .B(n48893), .Z(n48895) );
  IV U61704 ( .A(n48895), .Z(n49824) );
  IV U61705 ( .A(n48896), .Z(n48900) );
  NOR U61706 ( .A(n48897), .B(n49799), .Z(n48898) );
  IV U61707 ( .A(n48898), .Z(n48899) );
  NOR U61708 ( .A(n48900), .B(n48899), .Z(n49789) );
  IV U61709 ( .A(n48901), .Z(n48902) );
  NOR U61710 ( .A(n48903), .B(n48902), .Z(n49792) );
  IV U61711 ( .A(n48904), .Z(n48906) );
  NOR U61712 ( .A(n48906), .B(n48905), .Z(n48907) );
  NOR U61713 ( .A(n55865), .B(n48907), .Z(n53712) );
  IV U61714 ( .A(n48908), .Z(n48910) );
  NOR U61715 ( .A(n48910), .B(n48909), .Z(n48911) );
  IV U61716 ( .A(n48911), .Z(n49778) );
  IV U61717 ( .A(n48912), .Z(n48914) );
  IV U61718 ( .A(n48913), .Z(n48919) );
  NOR U61719 ( .A(n48914), .B(n48919), .Z(n53693) );
  IV U61720 ( .A(n48915), .Z(n48916) );
  NOR U61721 ( .A(n48923), .B(n48916), .Z(n52686) );
  IV U61722 ( .A(n48917), .Z(n48918) );
  NOR U61723 ( .A(n48919), .B(n48918), .Z(n53690) );
  NOR U61724 ( .A(n52686), .B(n53690), .Z(n48920) );
  IV U61725 ( .A(n48920), .Z(n49767) );
  IV U61726 ( .A(n48921), .Z(n48922) );
  NOR U61727 ( .A(n48923), .B(n48922), .Z(n52685) );
  IV U61728 ( .A(n48924), .Z(n48926) );
  NOR U61729 ( .A(n48926), .B(n48925), .Z(n52694) );
  IV U61730 ( .A(n48927), .Z(n48929) );
  NOR U61731 ( .A(n48929), .B(n48928), .Z(n52691) );
  NOR U61732 ( .A(n52694), .B(n52691), .Z(n49766) );
  IV U61733 ( .A(n48930), .Z(n52697) );
  NOR U61734 ( .A(n48931), .B(n52697), .Z(n49765) );
  IV U61735 ( .A(n48932), .Z(n48933) );
  NOR U61736 ( .A(n48934), .B(n48933), .Z(n52707) );
  NOR U61737 ( .A(n48936), .B(n48935), .Z(n52704) );
  NOR U61738 ( .A(n52707), .B(n52704), .Z(n49764) );
  NOR U61739 ( .A(n48938), .B(n48937), .Z(n53682) );
  NOR U61740 ( .A(n48939), .B(n53682), .Z(n49763) );
  IV U61741 ( .A(n48940), .Z(n48942) );
  IV U61742 ( .A(n48941), .Z(n48946) );
  NOR U61743 ( .A(n48942), .B(n48946), .Z(n53685) );
  IV U61744 ( .A(n48943), .Z(n48944) );
  NOR U61745 ( .A(n48944), .B(n49759), .Z(n52716) );
  IV U61746 ( .A(n48945), .Z(n48947) );
  NOR U61747 ( .A(n48947), .B(n48946), .Z(n53679) );
  NOR U61748 ( .A(n52716), .B(n53679), .Z(n48948) );
  IV U61749 ( .A(n48948), .Z(n49762) );
  IV U61750 ( .A(n48949), .Z(n49756) );
  IV U61751 ( .A(n48950), .Z(n48951) );
  NOR U61752 ( .A(n49756), .B(n48951), .Z(n48952) );
  IV U61753 ( .A(n48952), .Z(n52726) );
  NOR U61754 ( .A(n48954), .B(n48953), .Z(n48955) );
  IV U61755 ( .A(n48955), .Z(n48961) );
  XOR U61756 ( .A(n49751), .B(n49752), .Z(n48958) );
  IV U61757 ( .A(n48956), .Z(n48957) );
  NOR U61758 ( .A(n48958), .B(n48957), .Z(n48959) );
  IV U61759 ( .A(n48959), .Z(n48960) );
  NOR U61760 ( .A(n48961), .B(n48960), .Z(n48962) );
  IV U61761 ( .A(n48962), .Z(n53673) );
  IV U61762 ( .A(n48963), .Z(n48965) );
  IV U61763 ( .A(n48964), .Z(n48972) );
  NOR U61764 ( .A(n48965), .B(n48972), .Z(n48969) );
  IV U61765 ( .A(n48966), .Z(n48967) );
  NOR U61766 ( .A(n48967), .B(n49746), .Z(n48968) );
  NOR U61767 ( .A(n48969), .B(n48968), .Z(n52729) );
  IV U61768 ( .A(n48970), .Z(n48971) );
  NOR U61769 ( .A(n48972), .B(n48971), .Z(n49737) );
  IV U61770 ( .A(n49737), .Z(n49727) );
  IV U61771 ( .A(n48973), .Z(n48974) );
  NOR U61772 ( .A(n48974), .B(n49729), .Z(n53649) );
  IV U61773 ( .A(n48975), .Z(n48977) );
  NOR U61774 ( .A(n48977), .B(n48976), .Z(n49724) );
  IV U61775 ( .A(n49724), .Z(n49717) );
  IV U61776 ( .A(n48978), .Z(n52734) );
  NOR U61777 ( .A(n48979), .B(n52734), .Z(n49721) );
  IV U61778 ( .A(n48980), .Z(n48981) );
  NOR U61779 ( .A(n48981), .B(n49705), .Z(n53628) );
  IV U61780 ( .A(n48982), .Z(n48984) );
  NOR U61781 ( .A(n48984), .B(n48983), .Z(n52745) );
  IV U61782 ( .A(n48985), .Z(n48986) );
  NOR U61783 ( .A(n48987), .B(n48986), .Z(n52741) );
  NOR U61784 ( .A(n52745), .B(n52741), .Z(n49703) );
  IV U61785 ( .A(n48988), .Z(n48989) );
  NOR U61786 ( .A(n48989), .B(n48991), .Z(n52761) );
  IV U61787 ( .A(n48990), .Z(n48992) );
  NOR U61788 ( .A(n48992), .B(n48991), .Z(n52758) );
  IV U61789 ( .A(n48993), .Z(n48995) );
  IV U61790 ( .A(n48994), .Z(n48997) );
  NOR U61791 ( .A(n48995), .B(n48997), .Z(n52767) );
  IV U61792 ( .A(n48996), .Z(n48998) );
  NOR U61793 ( .A(n48998), .B(n48997), .Z(n52764) );
  IV U61794 ( .A(n49695), .Z(n48999) );
  NOR U61795 ( .A(n49694), .B(n48999), .Z(n52779) );
  IV U61796 ( .A(n49000), .Z(n49005) );
  IV U61797 ( .A(n49001), .Z(n49002) );
  NOR U61798 ( .A(n49005), .B(n49002), .Z(n53614) );
  IV U61799 ( .A(n49003), .Z(n49004) );
  NOR U61800 ( .A(n49005), .B(n49004), .Z(n53618) );
  IV U61801 ( .A(n49006), .Z(n49009) );
  NOR U61802 ( .A(n49007), .B(n49676), .Z(n49008) );
  IV U61803 ( .A(n49008), .Z(n49686) );
  NOR U61804 ( .A(n49009), .B(n49686), .Z(n49680) );
  IV U61805 ( .A(n49010), .Z(n49015) );
  IV U61806 ( .A(n49011), .Z(n49012) );
  NOR U61807 ( .A(n49015), .B(n49012), .Z(n53591) );
  IV U61808 ( .A(n49013), .Z(n49014) );
  NOR U61809 ( .A(n49015), .B(n49014), .Z(n53586) );
  IV U61810 ( .A(n49016), .Z(n49018) );
  NOR U61811 ( .A(n49018), .B(n49017), .Z(n53583) );
  IV U61812 ( .A(n49019), .Z(n49022) );
  NOR U61813 ( .A(n49659), .B(n49020), .Z(n49021) );
  IV U61814 ( .A(n49021), .Z(n49024) );
  NOR U61815 ( .A(n49022), .B(n49024), .Z(n53574) );
  IV U61816 ( .A(n49023), .Z(n49025) );
  NOR U61817 ( .A(n49025), .B(n49024), .Z(n52799) );
  IV U61818 ( .A(n49026), .Z(n49027) );
  NOR U61819 ( .A(n49027), .B(n49032), .Z(n52796) );
  IV U61820 ( .A(n49028), .Z(n49030) );
  NOR U61821 ( .A(n49030), .B(n49029), .Z(n52806) );
  IV U61822 ( .A(n49031), .Z(n49033) );
  NOR U61823 ( .A(n49033), .B(n49032), .Z(n52803) );
  NOR U61824 ( .A(n52806), .B(n52803), .Z(n49656) );
  IV U61825 ( .A(n49034), .Z(n49036) );
  NOR U61826 ( .A(n49036), .B(n49035), .Z(n49654) );
  IV U61827 ( .A(n49654), .Z(n49648) );
  IV U61828 ( .A(n49037), .Z(n49039) );
  NOR U61829 ( .A(n49039), .B(n49038), .Z(n49637) );
  IV U61830 ( .A(n49637), .Z(n49632) );
  IV U61831 ( .A(n49040), .Z(n49041) );
  NOR U61832 ( .A(n49042), .B(n49041), .Z(n53553) );
  NOR U61833 ( .A(n49044), .B(n49043), .Z(n52843) );
  NOR U61834 ( .A(n53553), .B(n52843), .Z(n49045) );
  IV U61835 ( .A(n49045), .Z(n49621) );
  IV U61836 ( .A(n49046), .Z(n49048) );
  NOR U61837 ( .A(n49048), .B(n49047), .Z(n49053) );
  IV U61838 ( .A(n49049), .Z(n49050) );
  NOR U61839 ( .A(n49051), .B(n49050), .Z(n49052) );
  NOR U61840 ( .A(n49053), .B(n49052), .Z(n53550) );
  IV U61841 ( .A(n49054), .Z(n52847) );
  NOR U61842 ( .A(n49055), .B(n52847), .Z(n49620) );
  IV U61843 ( .A(n49056), .Z(n49057) );
  NOR U61844 ( .A(n49058), .B(n49057), .Z(n52853) );
  NOR U61845 ( .A(n49060), .B(n49059), .Z(n52858) );
  NOR U61846 ( .A(n52853), .B(n52858), .Z(n49619) );
  IV U61847 ( .A(n49061), .Z(n49062) );
  NOR U61848 ( .A(n49063), .B(n49062), .Z(n52851) );
  XOR U61849 ( .A(n53540), .B(n52864), .Z(n49064) );
  NOR U61850 ( .A(n52851), .B(n49064), .Z(n49618) );
  IV U61851 ( .A(n49065), .Z(n53538) );
  IV U61852 ( .A(n49066), .Z(n49067) );
  NOR U61853 ( .A(n49068), .B(n49067), .Z(n52872) );
  IV U61854 ( .A(n49069), .Z(n49071) );
  NOR U61855 ( .A(n49071), .B(n49070), .Z(n53530) );
  NOR U61856 ( .A(n52872), .B(n53530), .Z(n49603) );
  IV U61857 ( .A(n49072), .Z(n49074) );
  IV U61858 ( .A(n49073), .Z(n49076) );
  NOR U61859 ( .A(n49074), .B(n49076), .Z(n49591) );
  IV U61860 ( .A(n49075), .Z(n49077) );
  NOR U61861 ( .A(n49077), .B(n49076), .Z(n49078) );
  IV U61862 ( .A(n49078), .Z(n52885) );
  IV U61863 ( .A(n49079), .Z(n49080) );
  NOR U61864 ( .A(n49081), .B(n49080), .Z(n52891) );
  NOR U61865 ( .A(n49083), .B(n49082), .Z(n52882) );
  NOR U61866 ( .A(n52891), .B(n52882), .Z(n49084) );
  IV U61867 ( .A(n49084), .Z(n49589) );
  IV U61868 ( .A(n49085), .Z(n49086) );
  NOR U61869 ( .A(n49087), .B(n49086), .Z(n52888) );
  IV U61870 ( .A(n49088), .Z(n49089) );
  NOR U61871 ( .A(n49089), .B(n49094), .Z(n52896) );
  IV U61872 ( .A(n49090), .Z(n49092) );
  NOR U61873 ( .A(n49092), .B(n49091), .Z(n53497) );
  IV U61874 ( .A(n49093), .Z(n49095) );
  NOR U61875 ( .A(n49095), .B(n49094), .Z(n53489) );
  NOR U61876 ( .A(n53497), .B(n53489), .Z(n56048) );
  IV U61877 ( .A(n49096), .Z(n49583) );
  IV U61878 ( .A(n49097), .Z(n49098) );
  NOR U61879 ( .A(n49583), .B(n49098), .Z(n53499) );
  IV U61880 ( .A(n53499), .Z(n53496) );
  IV U61881 ( .A(n49099), .Z(n49101) );
  NOR U61882 ( .A(n49101), .B(n49100), .Z(n49558) );
  IV U61883 ( .A(n49558), .Z(n49548) );
  IV U61884 ( .A(n49102), .Z(n49103) );
  NOR U61885 ( .A(n49103), .B(n49540), .Z(n53456) );
  IV U61886 ( .A(n49104), .Z(n53452) );
  NOR U61887 ( .A(n49105), .B(n53452), .Z(n49108) );
  IV U61888 ( .A(n49106), .Z(n49107) );
  NOR U61889 ( .A(n49540), .B(n49107), .Z(n53459) );
  NOR U61890 ( .A(n49108), .B(n53459), .Z(n49109) );
  IV U61891 ( .A(n49109), .Z(n49538) );
  IV U61892 ( .A(n49110), .Z(n49111) );
  NOR U61893 ( .A(n49114), .B(n49111), .Z(n53436) );
  IV U61894 ( .A(n49112), .Z(n49113) );
  NOR U61895 ( .A(n49114), .B(n49113), .Z(n53439) );
  IV U61896 ( .A(n49115), .Z(n49117) );
  IV U61897 ( .A(n49116), .Z(n49524) );
  NOR U61898 ( .A(n49117), .B(n49524), .Z(n52926) );
  IV U61899 ( .A(n49118), .Z(n49119) );
  NOR U61900 ( .A(n49120), .B(n49119), .Z(n52935) );
  IV U61901 ( .A(n49121), .Z(n49122) );
  NOR U61902 ( .A(n49123), .B(n49122), .Z(n53425) );
  NOR U61903 ( .A(n52935), .B(n53425), .Z(n49522) );
  IV U61904 ( .A(n49124), .Z(n49125) );
  NOR U61905 ( .A(n49126), .B(n49125), .Z(n52938) );
  NOR U61906 ( .A(n53420), .B(n52938), .Z(n49521) );
  IV U61907 ( .A(n49127), .Z(n49128) );
  NOR U61908 ( .A(n49131), .B(n49128), .Z(n52942) );
  IV U61909 ( .A(n49129), .Z(n49130) );
  NOR U61910 ( .A(n49131), .B(n49130), .Z(n52950) );
  NOR U61911 ( .A(n52942), .B(n52950), .Z(n49520) );
  IV U61912 ( .A(n49132), .Z(n49135) );
  IV U61913 ( .A(n49133), .Z(n49134) );
  NOR U61914 ( .A(n49135), .B(n49134), .Z(n52946) );
  NOR U61915 ( .A(n49146), .B(n49136), .Z(n49137) );
  IV U61916 ( .A(n49137), .Z(n49145) );
  NOR U61917 ( .A(n49139), .B(n49138), .Z(n49140) );
  IV U61918 ( .A(n49140), .Z(n49141) );
  NOR U61919 ( .A(n49142), .B(n49141), .Z(n49143) );
  IV U61920 ( .A(n49143), .Z(n49144) );
  NOR U61921 ( .A(n49145), .B(n49144), .Z(n53411) );
  NOR U61922 ( .A(n49147), .B(n49146), .Z(n53408) );
  IV U61923 ( .A(n49148), .Z(n52958) );
  NOR U61924 ( .A(n49149), .B(n52958), .Z(n49153) );
  IV U61925 ( .A(n49150), .Z(n49151) );
  NOR U61926 ( .A(n49152), .B(n49151), .Z(n53404) );
  NOR U61927 ( .A(n49153), .B(n53404), .Z(n49518) );
  IV U61928 ( .A(n49154), .Z(n49158) );
  NOR U61929 ( .A(n49510), .B(n49155), .Z(n49156) );
  IV U61930 ( .A(n49156), .Z(n49157) );
  NOR U61931 ( .A(n49158), .B(n49157), .Z(n52963) );
  NOR U61932 ( .A(n49160), .B(n49159), .Z(n52975) );
  IV U61933 ( .A(n49161), .Z(n49163) );
  IV U61934 ( .A(n49162), .Z(n49165) );
  NOR U61935 ( .A(n49163), .B(n49165), .Z(n52973) );
  NOR U61936 ( .A(n52975), .B(n52973), .Z(n49498) );
  IV U61937 ( .A(n49164), .Z(n49166) );
  NOR U61938 ( .A(n49166), .B(n49165), .Z(n49167) );
  IV U61939 ( .A(n49167), .Z(n52971) );
  IV U61940 ( .A(n49168), .Z(n49170) );
  NOR U61941 ( .A(n49170), .B(n49169), .Z(n52981) );
  IV U61942 ( .A(n49171), .Z(n49173) );
  IV U61943 ( .A(n49172), .Z(n49495) );
  NOR U61944 ( .A(n49173), .B(n49495), .Z(n52986) );
  IV U61945 ( .A(n49174), .Z(n49175) );
  NOR U61946 ( .A(n49175), .B(n49495), .Z(n53380) );
  IV U61947 ( .A(n49176), .Z(n49177) );
  NOR U61948 ( .A(n49178), .B(n49177), .Z(n52993) );
  NOR U61949 ( .A(n49179), .B(n53376), .Z(n49180) );
  NOR U61950 ( .A(n52993), .B(n49180), .Z(n49181) );
  IV U61951 ( .A(n49181), .Z(n49493) );
  NOR U61952 ( .A(n49182), .B(n49192), .Z(n49183) );
  IV U61953 ( .A(n49183), .Z(n53003) );
  XOR U61954 ( .A(n49185), .B(n49184), .Z(n49186) );
  NOR U61955 ( .A(n49187), .B(n49186), .Z(n53001) );
  IV U61956 ( .A(n49188), .Z(n52997) );
  XOR U61957 ( .A(n53001), .B(n52997), .Z(n49189) );
  NOR U61958 ( .A(n53003), .B(n49189), .Z(n49492) );
  IV U61959 ( .A(n49190), .Z(n49191) );
  NOR U61960 ( .A(n49192), .B(n49191), .Z(n53006) );
  NOR U61961 ( .A(n49194), .B(n49193), .Z(n53012) );
  IV U61962 ( .A(n49195), .Z(n49197) );
  NOR U61963 ( .A(n49197), .B(n49196), .Z(n49202) );
  IV U61964 ( .A(n49198), .Z(n49199) );
  NOR U61965 ( .A(n49200), .B(n49199), .Z(n49201) );
  NOR U61966 ( .A(n49202), .B(n49201), .Z(n53021) );
  IV U61967 ( .A(n49203), .Z(n49205) );
  NOR U61968 ( .A(n49205), .B(n49204), .Z(n49210) );
  IV U61969 ( .A(n49206), .Z(n49208) );
  NOR U61970 ( .A(n49208), .B(n49207), .Z(n49209) );
  NOR U61971 ( .A(n49210), .B(n49209), .Z(n53030) );
  IV U61972 ( .A(n49211), .Z(n49214) );
  IV U61973 ( .A(n49212), .Z(n49213) );
  NOR U61974 ( .A(n49214), .B(n49213), .Z(n53026) );
  NOR U61975 ( .A(n49216), .B(n49215), .Z(n53031) );
  NOR U61976 ( .A(n53031), .B(n53023), .Z(n49484) );
  IV U61977 ( .A(n49217), .Z(n49220) );
  IV U61978 ( .A(n49218), .Z(n49219) );
  NOR U61979 ( .A(n49220), .B(n49219), .Z(n49221) );
  IV U61980 ( .A(n49221), .Z(n53336) );
  IV U61981 ( .A(n49222), .Z(n49223) );
  NOR U61982 ( .A(n49224), .B(n49223), .Z(n53036) );
  NOR U61983 ( .A(n49225), .B(n49477), .Z(n53034) );
  NOR U61984 ( .A(n53036), .B(n53034), .Z(n49226) );
  IV U61985 ( .A(n49226), .Z(n49474) );
  IV U61986 ( .A(n49227), .Z(n49228) );
  NOR U61987 ( .A(n49229), .B(n49228), .Z(n53039) );
  NOR U61988 ( .A(n49231), .B(n49230), .Z(n49237) );
  IV U61989 ( .A(n49231), .Z(n49233) );
  NOR U61990 ( .A(n49233), .B(n49232), .Z(n49234) );
  NOR U61991 ( .A(n49235), .B(n49234), .Z(n49236) );
  NOR U61992 ( .A(n49237), .B(n49236), .Z(n53045) );
  IV U61993 ( .A(n49238), .Z(n49239) );
  NOR U61994 ( .A(n49242), .B(n49239), .Z(n53042) );
  IV U61995 ( .A(n49240), .Z(n49241) );
  NOR U61996 ( .A(n49242), .B(n49241), .Z(n53322) );
  IV U61997 ( .A(n49243), .Z(n49244) );
  NOR U61998 ( .A(n49245), .B(n49244), .Z(n53302) );
  NOR U61999 ( .A(n49246), .B(n49245), .Z(n53311) );
  NOR U62000 ( .A(n53302), .B(n53311), .Z(n49466) );
  IV U62001 ( .A(n49247), .Z(n49251) );
  NOR U62002 ( .A(n49251), .B(n49248), .Z(n53288) );
  IV U62003 ( .A(n49249), .Z(n49250) );
  NOR U62004 ( .A(n49251), .B(n49250), .Z(n53292) );
  NOR U62005 ( .A(n53288), .B(n53292), .Z(n56424) );
  IV U62006 ( .A(n49252), .Z(n49254) );
  NOR U62007 ( .A(n49254), .B(n49253), .Z(n53285) );
  IV U62008 ( .A(n49255), .Z(n49258) );
  NOR U62009 ( .A(n49256), .B(n49264), .Z(n49257) );
  IV U62010 ( .A(n49257), .Z(n49260) );
  NOR U62011 ( .A(n49258), .B(n49260), .Z(n53278) );
  IV U62012 ( .A(n49259), .Z(n49261) );
  NOR U62013 ( .A(n49261), .B(n49260), .Z(n53075) );
  IV U62014 ( .A(n49262), .Z(n49263) );
  NOR U62015 ( .A(n49264), .B(n49263), .Z(n53082) );
  IV U62016 ( .A(n49265), .Z(n49266) );
  NOR U62017 ( .A(n49267), .B(n49266), .Z(n53079) );
  NOR U62018 ( .A(n53082), .B(n53079), .Z(n49438) );
  IV U62019 ( .A(n49268), .Z(n49269) );
  NOR U62020 ( .A(n49270), .B(n49269), .Z(n53084) );
  NOR U62021 ( .A(n53272), .B(n53084), .Z(n49437) );
  IV U62022 ( .A(n49271), .Z(n49272) );
  NOR U62023 ( .A(n49272), .B(n49274), .Z(n53090) );
  IV U62024 ( .A(n49273), .Z(n49275) );
  NOR U62025 ( .A(n49275), .B(n49274), .Z(n53088) );
  IV U62026 ( .A(n49276), .Z(n49277) );
  NOR U62027 ( .A(n49278), .B(n49277), .Z(n53101) );
  IV U62028 ( .A(n49279), .Z(n49283) );
  IV U62029 ( .A(n49280), .Z(n49284) );
  NOR U62030 ( .A(n49281), .B(n49284), .Z(n49282) );
  IV U62031 ( .A(n49282), .Z(n49433) );
  NOR U62032 ( .A(n49283), .B(n49433), .Z(n53099) );
  NOR U62033 ( .A(n53101), .B(n53099), .Z(n49436) );
  NOR U62034 ( .A(n49285), .B(n49284), .Z(n53104) );
  NOR U62035 ( .A(n53113), .B(n53104), .Z(n49431) );
  IV U62036 ( .A(n49286), .Z(n49290) );
  NOR U62037 ( .A(n49287), .B(n49425), .Z(n49288) );
  IV U62038 ( .A(n49288), .Z(n49289) );
  NOR U62039 ( .A(n49290), .B(n49289), .Z(n53267) );
  IV U62040 ( .A(n49291), .Z(n49298) );
  IV U62041 ( .A(n49292), .Z(n49293) );
  NOR U62042 ( .A(n49298), .B(n49293), .Z(n53264) );
  IV U62043 ( .A(n49294), .Z(n49295) );
  NOR U62044 ( .A(n49295), .B(n49304), .Z(n53123) );
  IV U62045 ( .A(n49296), .Z(n49297) );
  NOR U62046 ( .A(n49298), .B(n49297), .Z(n53261) );
  NOR U62047 ( .A(n53123), .B(n53261), .Z(n49299) );
  IV U62048 ( .A(n49299), .Z(n49420) );
  IV U62049 ( .A(n49300), .Z(n49301) );
  NOR U62050 ( .A(n49302), .B(n49301), .Z(n53129) );
  IV U62051 ( .A(n49303), .Z(n49305) );
  NOR U62052 ( .A(n49305), .B(n49304), .Z(n53127) );
  NOR U62053 ( .A(n53129), .B(n53127), .Z(n49419) );
  IV U62054 ( .A(n49306), .Z(n53133) );
  NOR U62055 ( .A(n49307), .B(n53133), .Z(n49311) );
  IV U62056 ( .A(n49308), .Z(n49310) );
  NOR U62057 ( .A(n49310), .B(n49309), .Z(n53258) );
  NOR U62058 ( .A(n49311), .B(n53258), .Z(n49418) );
  IV U62059 ( .A(n49312), .Z(n49314) );
  NOR U62060 ( .A(n49314), .B(n49313), .Z(n53240) );
  IV U62061 ( .A(n49315), .Z(n49316) );
  NOR U62062 ( .A(n49316), .B(n49319), .Z(n49317) );
  IV U62063 ( .A(n49317), .Z(n53140) );
  IV U62064 ( .A(n49318), .Z(n49320) );
  NOR U62065 ( .A(n49320), .B(n49319), .Z(n53218) );
  IV U62066 ( .A(n49321), .Z(n49323) );
  IV U62067 ( .A(n49322), .Z(n49326) );
  NOR U62068 ( .A(n49323), .B(n49326), .Z(n53141) );
  IV U62069 ( .A(n49324), .Z(n49325) );
  NOR U62070 ( .A(n49326), .B(n49325), .Z(n53144) );
  IV U62071 ( .A(n49327), .Z(n49328) );
  NOR U62072 ( .A(n49329), .B(n49328), .Z(n53156) );
  NOR U62073 ( .A(n49330), .B(n53148), .Z(n49331) );
  NOR U62074 ( .A(n53156), .B(n49331), .Z(n49332) );
  IV U62075 ( .A(n49332), .Z(n49403) );
  IV U62076 ( .A(n49333), .Z(n49336) );
  IV U62077 ( .A(n49334), .Z(n49335) );
  NOR U62078 ( .A(n49336), .B(n49335), .Z(n53162) );
  NOR U62079 ( .A(n49338), .B(n49337), .Z(n49339) );
  NOR U62080 ( .A(n49340), .B(n49339), .Z(n53159) );
  IV U62081 ( .A(n49341), .Z(n49342) );
  NOR U62082 ( .A(n49345), .B(n49342), .Z(n53210) );
  IV U62083 ( .A(n49343), .Z(n49344) );
  NOR U62084 ( .A(n49345), .B(n49344), .Z(n53165) );
  IV U62085 ( .A(n49346), .Z(n49347) );
  NOR U62086 ( .A(n49351), .B(n49347), .Z(n49348) );
  IV U62087 ( .A(n49348), .Z(n53172) );
  IV U62088 ( .A(n49349), .Z(n49350) );
  NOR U62089 ( .A(n49351), .B(n49350), .Z(n53197) );
  IV U62090 ( .A(n49352), .Z(n49354) );
  IV U62091 ( .A(n49353), .Z(n49394) );
  NOR U62092 ( .A(n49354), .B(n49394), .Z(n53173) );
  NOR U62093 ( .A(n53197), .B(n53173), .Z(n49355) );
  IV U62094 ( .A(n49355), .Z(n49395) );
  IV U62095 ( .A(n49356), .Z(n49357) );
  NOR U62096 ( .A(n49394), .B(n49357), .Z(n53178) );
  NOR U62097 ( .A(n49359), .B(n49358), .Z(n53187) );
  IV U62098 ( .A(n49366), .Z(n49369) );
  IV U62099 ( .A(n49367), .Z(n49368) );
  NOR U62100 ( .A(n49369), .B(n49368), .Z(n53186) );
  XOR U62101 ( .A(n53189), .B(n53186), .Z(n49375) );
  XOR U62102 ( .A(n53187), .B(n49375), .Z(n53182) );
  IV U62103 ( .A(n53182), .Z(n49378) );
  IV U62104 ( .A(n49370), .Z(n49371) );
  NOR U62105 ( .A(n49371), .B(n49386), .Z(n49382) );
  IV U62106 ( .A(n49382), .Z(n53183) );
  NOR U62107 ( .A(n49378), .B(n53183), .Z(n49384) );
  IV U62108 ( .A(n49372), .Z(n49373) );
  NOR U62109 ( .A(n49374), .B(n49373), .Z(n49377) );
  IV U62110 ( .A(n49377), .Z(n49376) );
  NOR U62111 ( .A(n49376), .B(n49375), .Z(n53184) );
  NOR U62112 ( .A(n49378), .B(n49377), .Z(n49379) );
  NOR U62113 ( .A(n53184), .B(n49379), .Z(n49380) );
  IV U62114 ( .A(n49380), .Z(n49381) );
  NOR U62115 ( .A(n49382), .B(n49381), .Z(n49383) );
  NOR U62116 ( .A(n49384), .B(n49383), .Z(n53193) );
  IV U62117 ( .A(n49385), .Z(n49387) );
  NOR U62118 ( .A(n49387), .B(n49386), .Z(n53190) );
  NOR U62119 ( .A(n49389), .B(n49388), .Z(n53192) );
  NOR U62120 ( .A(n53190), .B(n53192), .Z(n49390) );
  XOR U62121 ( .A(n53193), .B(n49390), .Z(n49391) );
  IV U62122 ( .A(n49391), .Z(n53177) );
  IV U62123 ( .A(n49392), .Z(n49393) );
  NOR U62124 ( .A(n49394), .B(n49393), .Z(n53175) );
  XOR U62125 ( .A(n53177), .B(n53175), .Z(n53180) );
  XOR U62126 ( .A(n53178), .B(n53180), .Z(n53198) );
  XOR U62127 ( .A(n49395), .B(n53198), .Z(n53202) );
  XOR U62128 ( .A(n53172), .B(n53202), .Z(n53168) );
  IV U62129 ( .A(n49396), .Z(n49398) );
  IV U62130 ( .A(n49397), .Z(n49401) );
  NOR U62131 ( .A(n49398), .B(n49401), .Z(n53169) );
  NOR U62132 ( .A(n53200), .B(n53169), .Z(n49399) );
  XOR U62133 ( .A(n53168), .B(n49399), .Z(n53206) );
  IV U62134 ( .A(n49400), .Z(n49402) );
  NOR U62135 ( .A(n49402), .B(n49401), .Z(n53204) );
  XOR U62136 ( .A(n53206), .B(n53204), .Z(n53166) );
  XOR U62137 ( .A(n53165), .B(n53166), .Z(n53212) );
  XOR U62138 ( .A(n53210), .B(n53212), .Z(n53161) );
  XOR U62139 ( .A(n53159), .B(n53161), .Z(n53163) );
  XOR U62140 ( .A(n53162), .B(n53163), .Z(n53157) );
  XOR U62141 ( .A(n49403), .B(n53157), .Z(n53146) );
  XOR U62142 ( .A(n53144), .B(n53146), .Z(n53142) );
  XOR U62143 ( .A(n53141), .B(n53142), .Z(n53219) );
  XOR U62144 ( .A(n53218), .B(n53219), .Z(n53139) );
  XOR U62145 ( .A(n53140), .B(n53139), .Z(n53224) );
  IV U62146 ( .A(n49404), .Z(n49407) );
  NOR U62147 ( .A(n49405), .B(n49407), .Z(n53228) );
  IV U62148 ( .A(n49406), .Z(n49413) );
  NOR U62149 ( .A(n49408), .B(n49407), .Z(n49409) );
  IV U62150 ( .A(n49409), .Z(n49410) );
  NOR U62151 ( .A(n49411), .B(n49410), .Z(n49412) );
  IV U62152 ( .A(n49412), .Z(n49416) );
  NOR U62153 ( .A(n49413), .B(n49416), .Z(n53225) );
  NOR U62154 ( .A(n53228), .B(n53225), .Z(n49414) );
  XOR U62155 ( .A(n53224), .B(n49414), .Z(n53138) );
  IV U62156 ( .A(n49415), .Z(n49417) );
  NOR U62157 ( .A(n49417), .B(n49416), .Z(n53136) );
  XOR U62158 ( .A(n53138), .B(n53136), .Z(n53244) );
  XOR U62159 ( .A(n53243), .B(n53244), .Z(n53241) );
  XOR U62160 ( .A(n53240), .B(n53241), .Z(n53259) );
  XOR U62161 ( .A(n49418), .B(n53259), .Z(n53126) );
  XOR U62162 ( .A(n49419), .B(n53126), .Z(n53263) );
  XOR U62163 ( .A(n49420), .B(n53263), .Z(n53266) );
  XOR U62164 ( .A(n53264), .B(n53266), .Z(n53268) );
  XOR U62165 ( .A(n53267), .B(n53268), .Z(n53122) );
  IV U62166 ( .A(n49421), .Z(n49422) );
  NOR U62167 ( .A(n49422), .B(n49425), .Z(n53118) );
  IV U62168 ( .A(n49423), .Z(n49429) );
  IV U62169 ( .A(n49424), .Z(n49426) );
  NOR U62170 ( .A(n49426), .B(n49425), .Z(n49427) );
  IV U62171 ( .A(n49427), .Z(n49428) );
  NOR U62172 ( .A(n49429), .B(n49428), .Z(n53120) );
  NOR U62173 ( .A(n53118), .B(n53120), .Z(n49430) );
  XOR U62174 ( .A(n53122), .B(n49430), .Z(n53111) );
  IV U62175 ( .A(n53111), .Z(n53109) );
  XOR U62176 ( .A(n53112), .B(n53109), .Z(n53106) );
  XOR U62177 ( .A(n49431), .B(n53106), .Z(n53095) );
  IV U62178 ( .A(n49432), .Z(n49434) );
  NOR U62179 ( .A(n49434), .B(n49433), .Z(n53096) );
  XOR U62180 ( .A(n53095), .B(n53096), .Z(n49435) );
  XOR U62181 ( .A(n49436), .B(n49435), .Z(n53273) );
  XOR U62182 ( .A(n53088), .B(n53273), .Z(n53092) );
  XOR U62183 ( .A(n53090), .B(n53092), .Z(n53085) );
  XOR U62184 ( .A(n49437), .B(n53085), .Z(n53078) );
  XOR U62185 ( .A(n49438), .B(n53078), .Z(n53077) );
  XOR U62186 ( .A(n53075), .B(n53077), .Z(n53277) );
  XOR U62187 ( .A(n53278), .B(n53277), .Z(n56417) );
  NOR U62188 ( .A(n49440), .B(n49439), .Z(n49441) );
  NOR U62189 ( .A(n49442), .B(n49441), .Z(n53280) );
  XOR U62190 ( .A(n56417), .B(n53280), .Z(n53286) );
  XOR U62191 ( .A(n53285), .B(n53286), .Z(n56425) );
  XOR U62192 ( .A(n56424), .B(n56425), .Z(n53070) );
  IV U62193 ( .A(n49443), .Z(n49444) );
  NOR U62194 ( .A(n49445), .B(n49444), .Z(n53072) );
  XOR U62195 ( .A(n53070), .B(n53072), .Z(n53065) );
  IV U62196 ( .A(n49446), .Z(n49447) );
  NOR U62197 ( .A(n49448), .B(n49447), .Z(n53069) );
  NOR U62198 ( .A(n49450), .B(n49449), .Z(n53064) );
  NOR U62199 ( .A(n53069), .B(n53064), .Z(n49451) );
  XOR U62200 ( .A(n53065), .B(n49451), .Z(n53063) );
  IV U62201 ( .A(n49455), .Z(n49453) );
  IV U62202 ( .A(n49454), .Z(n49452) );
  NOR U62203 ( .A(n49453), .B(n49452), .Z(n53061) );
  NOR U62204 ( .A(n49455), .B(n49454), .Z(n49456) );
  NOR U62205 ( .A(n49456), .B(n53058), .Z(n49457) );
  NOR U62206 ( .A(n53061), .B(n49457), .Z(n49458) );
  XOR U62207 ( .A(n53063), .B(n49458), .Z(n53054) );
  IV U62208 ( .A(n49459), .Z(n49460) );
  NOR U62209 ( .A(n49461), .B(n49460), .Z(n53297) );
  IV U62210 ( .A(n49462), .Z(n49464) );
  NOR U62211 ( .A(n49464), .B(n49463), .Z(n53053) );
  NOR U62212 ( .A(n53297), .B(n53053), .Z(n49465) );
  XOR U62213 ( .A(n53054), .B(n49465), .Z(n53313) );
  XOR U62214 ( .A(n49466), .B(n53313), .Z(n53051) );
  IV U62215 ( .A(n49467), .Z(n49469) );
  IV U62216 ( .A(n49468), .Z(n49472) );
  NOR U62217 ( .A(n49469), .B(n49472), .Z(n53050) );
  NOR U62218 ( .A(n53314), .B(n53050), .Z(n49470) );
  XOR U62219 ( .A(n53051), .B(n49470), .Z(n53321) );
  IV U62220 ( .A(n49471), .Z(n49473) );
  NOR U62221 ( .A(n49473), .B(n49472), .Z(n53319) );
  XOR U62222 ( .A(n53321), .B(n53319), .Z(n53323) );
  XOR U62223 ( .A(n53322), .B(n53323), .Z(n53043) );
  XOR U62224 ( .A(n53042), .B(n53043), .Z(n53047) );
  XOR U62225 ( .A(n53045), .B(n53047), .Z(n53040) );
  XOR U62226 ( .A(n53039), .B(n53040), .Z(n53037) );
  XOR U62227 ( .A(n49474), .B(n53037), .Z(n53337) );
  XOR U62228 ( .A(n53336), .B(n53337), .Z(n53348) );
  IV U62229 ( .A(n53348), .Z(n53345) );
  IV U62230 ( .A(n49475), .Z(n49476) );
  NOR U62231 ( .A(n49477), .B(n49476), .Z(n53347) );
  XOR U62232 ( .A(n53345), .B(n53347), .Z(n56472) );
  IV U62233 ( .A(n49478), .Z(n49479) );
  NOR U62234 ( .A(n49480), .B(n49479), .Z(n53346) );
  IV U62235 ( .A(n49481), .Z(n49482) );
  NOR U62236 ( .A(n49483), .B(n49482), .Z(n53338) );
  NOR U62237 ( .A(n53346), .B(n53338), .Z(n56469) );
  XOR U62238 ( .A(n56472), .B(n56469), .Z(n53024) );
  XOR U62239 ( .A(n49484), .B(n53024), .Z(n53027) );
  XOR U62240 ( .A(n53026), .B(n53027), .Z(n53029) );
  XOR U62241 ( .A(n53030), .B(n53029), .Z(n53016) );
  IV U62242 ( .A(n53016), .Z(n53020) );
  XOR U62243 ( .A(n53021), .B(n53020), .Z(n53368) );
  IV U62244 ( .A(n49485), .Z(n49486) );
  NOR U62245 ( .A(n49487), .B(n49486), .Z(n53017) );
  IV U62246 ( .A(n49488), .Z(n49490) );
  NOR U62247 ( .A(n49490), .B(n49489), .Z(n53367) );
  NOR U62248 ( .A(n53017), .B(n53367), .Z(n56132) );
  XOR U62249 ( .A(n53368), .B(n56132), .Z(n53010) );
  XOR U62250 ( .A(n53009), .B(n53010), .Z(n53013) );
  XOR U62251 ( .A(n53012), .B(n53013), .Z(n53007) );
  XOR U62252 ( .A(n53006), .B(n53007), .Z(n49491) );
  XOR U62253 ( .A(n49492), .B(n49491), .Z(n52991) );
  XOR U62254 ( .A(n52989), .B(n52991), .Z(n53375) );
  XOR U62255 ( .A(n49493), .B(n53375), .Z(n53382) );
  XOR U62256 ( .A(n53380), .B(n53382), .Z(n52987) );
  XOR U62257 ( .A(n52986), .B(n52987), .Z(n52980) );
  IV U62258 ( .A(n49494), .Z(n49496) );
  NOR U62259 ( .A(n49496), .B(n49495), .Z(n52978) );
  XOR U62260 ( .A(n52980), .B(n52978), .Z(n52982) );
  XOR U62261 ( .A(n52981), .B(n52982), .Z(n52976) );
  XOR U62262 ( .A(n52971), .B(n52976), .Z(n49497) );
  XOR U62263 ( .A(n49498), .B(n49497), .Z(n53391) );
  IV U62264 ( .A(n49499), .Z(n49501) );
  NOR U62265 ( .A(n49501), .B(n49500), .Z(n52969) );
  NOR U62266 ( .A(n49502), .B(n53390), .Z(n49503) );
  NOR U62267 ( .A(n52969), .B(n49503), .Z(n49504) );
  XOR U62268 ( .A(n53391), .B(n49504), .Z(n53396) );
  IV U62269 ( .A(n49507), .Z(n49505) );
  NOR U62270 ( .A(n49506), .B(n49505), .Z(n49516) );
  NOR U62271 ( .A(n49508), .B(n49507), .Z(n49514) );
  IV U62272 ( .A(n49509), .Z(n49511) );
  NOR U62273 ( .A(n49511), .B(n49510), .Z(n49512) );
  IV U62274 ( .A(n49512), .Z(n49513) );
  NOR U62275 ( .A(n49514), .B(n49513), .Z(n49515) );
  NOR U62276 ( .A(n49516), .B(n49515), .Z(n53398) );
  XOR U62277 ( .A(n53396), .B(n53398), .Z(n52965) );
  XOR U62278 ( .A(n52963), .B(n52965), .Z(n52967) );
  XOR U62279 ( .A(n49517), .B(n52967), .Z(n53406) );
  XOR U62280 ( .A(n49518), .B(n53406), .Z(n49519) );
  IV U62281 ( .A(n49519), .Z(n53409) );
  XOR U62282 ( .A(n53408), .B(n53409), .Z(n53413) );
  XOR U62283 ( .A(n53411), .B(n53413), .Z(n52948) );
  XOR U62284 ( .A(n52946), .B(n52948), .Z(n52943) );
  XOR U62285 ( .A(n49520), .B(n52943), .Z(n52937) );
  XOR U62286 ( .A(n49521), .B(n52937), .Z(n53426) );
  XOR U62287 ( .A(n49522), .B(n53426), .Z(n52929) );
  IV U62288 ( .A(n49523), .Z(n49525) );
  NOR U62289 ( .A(n49525), .B(n49524), .Z(n52930) );
  NOR U62290 ( .A(n52932), .B(n52930), .Z(n49526) );
  NOR U62291 ( .A(n52929), .B(n49526), .Z(n49537) );
  IV U62292 ( .A(n49526), .Z(n49535) );
  NOR U62293 ( .A(n49528), .B(n49527), .Z(n49531) );
  IV U62294 ( .A(n49531), .Z(n49530) );
  XOR U62295 ( .A(n52935), .B(n53426), .Z(n49529) );
  NOR U62296 ( .A(n49530), .B(n49529), .Z(n53433) );
  NOR U62297 ( .A(n52929), .B(n49531), .Z(n49532) );
  NOR U62298 ( .A(n53433), .B(n49532), .Z(n49533) );
  IV U62299 ( .A(n49533), .Z(n49534) );
  NOR U62300 ( .A(n49535), .B(n49534), .Z(n49536) );
  NOR U62301 ( .A(n49537), .B(n49536), .Z(n52928) );
  XOR U62302 ( .A(n52926), .B(n52928), .Z(n53451) );
  XOR U62303 ( .A(n53439), .B(n53451), .Z(n53437) );
  XOR U62304 ( .A(n53436), .B(n53437), .Z(n53460) );
  XOR U62305 ( .A(n49538), .B(n53460), .Z(n53458) );
  XOR U62306 ( .A(n53456), .B(n53458), .Z(n53469) );
  IV U62307 ( .A(n49539), .Z(n49541) );
  NOR U62308 ( .A(n49541), .B(n49540), .Z(n53467) );
  XOR U62309 ( .A(n53469), .B(n53467), .Z(n53471) );
  IV U62310 ( .A(n49542), .Z(n49549) );
  IV U62311 ( .A(n49543), .Z(n49544) );
  NOR U62312 ( .A(n49549), .B(n49544), .Z(n52924) );
  IV U62313 ( .A(n49550), .Z(n49545) );
  NOR U62314 ( .A(n49549), .B(n49545), .Z(n53470) );
  NOR U62315 ( .A(n52924), .B(n53470), .Z(n49546) );
  XOR U62316 ( .A(n53471), .B(n49546), .Z(n49555) );
  IV U62317 ( .A(n49555), .Z(n49547) );
  NOR U62318 ( .A(n49548), .B(n49547), .Z(n52923) );
  XOR U62319 ( .A(n49550), .B(n49549), .Z(n49553) );
  IV U62320 ( .A(n49551), .Z(n49552) );
  NOR U62321 ( .A(n49553), .B(n49552), .Z(n49556) );
  IV U62322 ( .A(n49556), .Z(n49554) );
  NOR U62323 ( .A(n49554), .B(n53471), .Z(n53480) );
  NOR U62324 ( .A(n49556), .B(n49555), .Z(n49557) );
  NOR U62325 ( .A(n53480), .B(n49557), .Z(n52918) );
  NOR U62326 ( .A(n49558), .B(n52918), .Z(n49559) );
  NOR U62327 ( .A(n52923), .B(n49559), .Z(n52915) );
  NOR U62328 ( .A(n49561), .B(n49560), .Z(n52919) );
  NOR U62329 ( .A(n52919), .B(n49562), .Z(n49563) );
  XOR U62330 ( .A(n52915), .B(n49563), .Z(n52914) );
  IV U62331 ( .A(n49564), .Z(n49566) );
  IV U62332 ( .A(n49565), .Z(n49570) );
  NOR U62333 ( .A(n49566), .B(n49570), .Z(n52912) );
  NOR U62334 ( .A(n49567), .B(n52912), .Z(n49568) );
  XOR U62335 ( .A(n52914), .B(n49568), .Z(n52909) );
  IV U62336 ( .A(n49569), .Z(n49571) );
  NOR U62337 ( .A(n49571), .B(n49570), .Z(n49572) );
  NOR U62338 ( .A(n52909), .B(n49572), .Z(n49574) );
  IV U62339 ( .A(n49572), .Z(n49573) );
  NOR U62340 ( .A(n52914), .B(n49573), .Z(n56055) );
  NOR U62341 ( .A(n49574), .B(n56055), .Z(n52904) );
  IV U62342 ( .A(n49575), .Z(n49576) );
  NOR U62343 ( .A(n49577), .B(n49576), .Z(n52908) );
  IV U62344 ( .A(n49578), .Z(n49579) );
  NOR U62345 ( .A(n49585), .B(n49579), .Z(n52905) );
  NOR U62346 ( .A(n52908), .B(n52905), .Z(n49580) );
  XOR U62347 ( .A(n52904), .B(n49580), .Z(n52903) );
  IV U62348 ( .A(n49581), .Z(n49582) );
  NOR U62349 ( .A(n49583), .B(n49582), .Z(n52899) );
  IV U62350 ( .A(n49584), .Z(n49586) );
  NOR U62351 ( .A(n49586), .B(n49585), .Z(n52901) );
  NOR U62352 ( .A(n52899), .B(n52901), .Z(n49587) );
  XOR U62353 ( .A(n52903), .B(n49587), .Z(n53498) );
  XOR U62354 ( .A(n53496), .B(n53498), .Z(n56044) );
  XOR U62355 ( .A(n56048), .B(n56044), .Z(n49588) );
  IV U62356 ( .A(n49588), .Z(n52898) );
  XOR U62357 ( .A(n52896), .B(n52898), .Z(n52890) );
  XOR U62358 ( .A(n52888), .B(n52890), .Z(n52892) );
  XOR U62359 ( .A(n49589), .B(n52892), .Z(n52884) );
  XOR U62360 ( .A(n52885), .B(n52884), .Z(n49590) );
  NOR U62361 ( .A(n49591), .B(n49590), .Z(n53513) );
  IV U62362 ( .A(n49591), .Z(n49593) );
  XOR U62363 ( .A(n52891), .B(n52892), .Z(n49592) );
  NOR U62364 ( .A(n49593), .B(n49592), .Z(n53510) );
  NOR U62365 ( .A(n53513), .B(n53510), .Z(n52879) );
  IV U62366 ( .A(n49594), .Z(n49596) );
  NOR U62367 ( .A(n49596), .B(n49595), .Z(n53511) );
  IV U62368 ( .A(n49597), .Z(n49598) );
  NOR U62369 ( .A(n49598), .B(n49601), .Z(n52878) );
  NOR U62370 ( .A(n53511), .B(n52878), .Z(n49599) );
  XOR U62371 ( .A(n52879), .B(n49599), .Z(n53517) );
  IV U62372 ( .A(n49600), .Z(n49602) );
  NOR U62373 ( .A(n49602), .B(n49601), .Z(n53515) );
  XOR U62374 ( .A(n53517), .B(n53515), .Z(n53531) );
  XOR U62375 ( .A(n49603), .B(n53531), .Z(n49604) );
  IV U62376 ( .A(n49604), .Z(n52875) );
  NOR U62377 ( .A(n49608), .B(n49605), .Z(n52874) );
  IV U62378 ( .A(n49606), .Z(n49607) );
  NOR U62379 ( .A(n49608), .B(n49607), .Z(n52869) );
  XOR U62380 ( .A(n52874), .B(n52869), .Z(n49609) );
  XOR U62381 ( .A(n52875), .B(n49609), .Z(n53535) );
  IV U62382 ( .A(n49610), .Z(n49611) );
  NOR U62383 ( .A(n49612), .B(n49611), .Z(n52867) );
  IV U62384 ( .A(n49613), .Z(n49616) );
  IV U62385 ( .A(n49614), .Z(n49615) );
  NOR U62386 ( .A(n49616), .B(n49615), .Z(n53534) );
  NOR U62387 ( .A(n52867), .B(n53534), .Z(n49617) );
  XOR U62388 ( .A(n53535), .B(n49617), .Z(n53537) );
  XOR U62389 ( .A(n53538), .B(n53537), .Z(n53541) );
  XOR U62390 ( .A(n49618), .B(n53541), .Z(n52859) );
  XOR U62391 ( .A(n49619), .B(n52859), .Z(n52848) );
  XOR U62392 ( .A(n49620), .B(n52848), .Z(n53551) );
  IV U62393 ( .A(n53551), .Z(n53549) );
  XOR U62394 ( .A(n53550), .B(n53549), .Z(n52844) );
  XOR U62395 ( .A(n49621), .B(n52844), .Z(n53559) );
  XOR U62396 ( .A(n53557), .B(n53559), .Z(n52840) );
  IV U62397 ( .A(n49622), .Z(n49625) );
  IV U62398 ( .A(n49623), .Z(n49624) );
  NOR U62399 ( .A(n49625), .B(n49624), .Z(n52839) );
  IV U62400 ( .A(n49626), .Z(n49629) );
  IV U62401 ( .A(n49627), .Z(n49628) );
  NOR U62402 ( .A(n49629), .B(n49628), .Z(n52832) );
  NOR U62403 ( .A(n52839), .B(n52832), .Z(n49630) );
  XOR U62404 ( .A(n52840), .B(n49630), .Z(n49635) );
  IV U62405 ( .A(n49635), .Z(n49631) );
  NOR U62406 ( .A(n49632), .B(n49631), .Z(n56699) );
  IV U62407 ( .A(n49633), .Z(n52829) );
  NOR U62408 ( .A(n49634), .B(n52829), .Z(n49636) );
  XOR U62409 ( .A(n49636), .B(n49635), .Z(n52824) );
  NOR U62410 ( .A(n49637), .B(n52824), .Z(n49638) );
  NOR U62411 ( .A(n56699), .B(n49638), .Z(n52819) );
  IV U62412 ( .A(n49639), .Z(n49640) );
  NOR U62413 ( .A(n49641), .B(n49640), .Z(n52823) );
  IV U62414 ( .A(n49642), .Z(n49643) );
  NOR U62415 ( .A(n49646), .B(n49643), .Z(n52820) );
  NOR U62416 ( .A(n52823), .B(n52820), .Z(n49644) );
  XOR U62417 ( .A(n52819), .B(n49644), .Z(n52818) );
  IV U62418 ( .A(n49645), .Z(n49647) );
  NOR U62419 ( .A(n49647), .B(n49646), .Z(n52816) );
  XOR U62420 ( .A(n52818), .B(n52816), .Z(n49651) );
  NOR U62421 ( .A(n49648), .B(n49651), .Z(n55993) );
  IV U62422 ( .A(n49649), .Z(n52810) );
  NOR U62423 ( .A(n49650), .B(n52810), .Z(n49652) );
  XOR U62424 ( .A(n49652), .B(n49651), .Z(n52807) );
  IV U62425 ( .A(n52807), .Z(n49653) );
  NOR U62426 ( .A(n49654), .B(n49653), .Z(n49655) );
  NOR U62427 ( .A(n55993), .B(n49655), .Z(n52802) );
  XOR U62428 ( .A(n49656), .B(n52802), .Z(n52798) );
  XOR U62429 ( .A(n52796), .B(n52798), .Z(n52800) );
  XOR U62430 ( .A(n52799), .B(n52800), .Z(n53575) );
  XOR U62431 ( .A(n53574), .B(n53575), .Z(n53581) );
  IV U62432 ( .A(n49657), .Z(n49658) );
  NOR U62433 ( .A(n49659), .B(n49658), .Z(n49660) );
  IV U62434 ( .A(n49660), .Z(n53577) );
  XOR U62435 ( .A(n53581), .B(n53577), .Z(n52788) );
  IV U62436 ( .A(n49661), .Z(n49662) );
  NOR U62437 ( .A(n49670), .B(n49662), .Z(n52789) );
  IV U62438 ( .A(n49663), .Z(n49664) );
  NOR U62439 ( .A(n49665), .B(n49664), .Z(n52793) );
  NOR U62440 ( .A(n53580), .B(n52793), .Z(n49666) );
  IV U62441 ( .A(n49666), .Z(n49667) );
  NOR U62442 ( .A(n52789), .B(n49667), .Z(n49668) );
  XOR U62443 ( .A(n52788), .B(n49668), .Z(n52787) );
  IV U62444 ( .A(n49669), .Z(n49671) );
  NOR U62445 ( .A(n49671), .B(n49670), .Z(n52785) );
  XOR U62446 ( .A(n52787), .B(n52785), .Z(n53585) );
  XOR U62447 ( .A(n53583), .B(n53585), .Z(n53588) );
  XOR U62448 ( .A(n53586), .B(n53588), .Z(n53593) );
  XOR U62449 ( .A(n53591), .B(n53593), .Z(n53603) );
  IV U62450 ( .A(n49672), .Z(n49673) );
  NOR U62451 ( .A(n49674), .B(n49673), .Z(n53594) );
  IV U62452 ( .A(n49675), .Z(n49677) );
  NOR U62453 ( .A(n49677), .B(n49676), .Z(n53602) );
  NOR U62454 ( .A(n53594), .B(n53602), .Z(n49678) );
  XOR U62455 ( .A(n53603), .B(n49678), .Z(n49679) );
  NOR U62456 ( .A(n49680), .B(n49679), .Z(n49683) );
  XOR U62457 ( .A(n53594), .B(n53603), .Z(n49682) );
  IV U62458 ( .A(n49680), .Z(n49681) );
  NOR U62459 ( .A(n49682), .B(n49681), .Z(n53610) );
  NOR U62460 ( .A(n49683), .B(n53610), .Z(n49684) );
  IV U62461 ( .A(n49684), .Z(n53608) );
  IV U62462 ( .A(n49685), .Z(n49687) );
  NOR U62463 ( .A(n49687), .B(n49686), .Z(n53606) );
  XOR U62464 ( .A(n53608), .B(n53606), .Z(n52784) );
  IV U62465 ( .A(n49688), .Z(n49689) );
  NOR U62466 ( .A(n49690), .B(n49689), .Z(n52782) );
  XOR U62467 ( .A(n52784), .B(n52782), .Z(n53619) );
  XOR U62468 ( .A(n53618), .B(n53619), .Z(n53615) );
  XOR U62469 ( .A(n53614), .B(n53615), .Z(n52780) );
  XOR U62470 ( .A(n52779), .B(n52780), .Z(n52773) );
  IV U62471 ( .A(n49691), .Z(n49692) );
  NOR U62472 ( .A(n49694), .B(n49692), .Z(n52772) );
  IV U62473 ( .A(n49693), .Z(n49697) );
  XOR U62474 ( .A(n49695), .B(n49694), .Z(n49696) );
  NOR U62475 ( .A(n49697), .B(n49696), .Z(n52776) );
  XOR U62476 ( .A(n52772), .B(n52776), .Z(n49698) );
  XOR U62477 ( .A(n52773), .B(n49698), .Z(n52765) );
  XOR U62478 ( .A(n52764), .B(n52765), .Z(n52768) );
  XOR U62479 ( .A(n52767), .B(n52768), .Z(n52759) );
  XOR U62480 ( .A(n52758), .B(n52759), .Z(n52762) );
  XOR U62481 ( .A(n52761), .B(n52762), .Z(n52751) );
  XOR U62482 ( .A(n52750), .B(n52751), .Z(n52754) );
  IV U62483 ( .A(n49699), .Z(n49700) );
  NOR U62484 ( .A(n49701), .B(n49700), .Z(n52748) );
  NOR U62485 ( .A(n52753), .B(n52748), .Z(n49702) );
  XOR U62486 ( .A(n52754), .B(n49702), .Z(n52742) );
  XOR U62487 ( .A(n49703), .B(n52742), .Z(n53630) );
  XOR U62488 ( .A(n53628), .B(n53630), .Z(n53633) );
  IV U62489 ( .A(n49704), .Z(n49708) );
  NOR U62490 ( .A(n49706), .B(n49705), .Z(n49707) );
  IV U62491 ( .A(n49707), .Z(n49712) );
  NOR U62492 ( .A(n49708), .B(n49712), .Z(n53631) );
  XOR U62493 ( .A(n53633), .B(n53631), .Z(n53641) );
  IV U62494 ( .A(n53641), .Z(n49715) );
  NOR U62495 ( .A(n49710), .B(n49709), .Z(n53640) );
  IV U62496 ( .A(n49711), .Z(n49713) );
  NOR U62497 ( .A(n49713), .B(n49712), .Z(n52739) );
  NOR U62498 ( .A(n53640), .B(n52739), .Z(n49714) );
  XOR U62499 ( .A(n49715), .B(n49714), .Z(n52733) );
  XOR U62500 ( .A(n49721), .B(n52733), .Z(n49716) );
  NOR U62501 ( .A(n49717), .B(n49716), .Z(n53653) );
  IV U62502 ( .A(n49718), .Z(n49719) );
  NOR U62503 ( .A(n49720), .B(n49719), .Z(n52730) );
  NOR U62504 ( .A(n49721), .B(n52730), .Z(n49722) );
  XOR U62505 ( .A(n52733), .B(n49722), .Z(n49723) );
  NOR U62506 ( .A(n49724), .B(n49723), .Z(n49725) );
  NOR U62507 ( .A(n53653), .B(n49725), .Z(n49726) );
  IV U62508 ( .A(n49726), .Z(n53651) );
  XOR U62509 ( .A(n53649), .B(n53651), .Z(n49732) );
  NOR U62510 ( .A(n49727), .B(n49732), .Z(n55909) );
  IV U62511 ( .A(n49728), .Z(n49730) );
  NOR U62512 ( .A(n49730), .B(n49729), .Z(n49734) );
  IV U62513 ( .A(n49734), .Z(n49731) );
  NOR U62514 ( .A(n53651), .B(n49731), .Z(n55924) );
  IV U62515 ( .A(n49732), .Z(n49733) );
  NOR U62516 ( .A(n49734), .B(n49733), .Z(n49735) );
  NOR U62517 ( .A(n55924), .B(n49735), .Z(n49736) );
  NOR U62518 ( .A(n49737), .B(n49736), .Z(n49738) );
  NOR U62519 ( .A(n55909), .B(n49738), .Z(n52727) );
  XOR U62520 ( .A(n52729), .B(n52727), .Z(n55898) );
  IV U62521 ( .A(n55898), .Z(n53657) );
  IV U62522 ( .A(n49739), .Z(n49744) );
  IV U62523 ( .A(n49740), .Z(n49741) );
  NOR U62524 ( .A(n49744), .B(n49741), .Z(n53659) );
  IV U62525 ( .A(n49742), .Z(n49743) );
  NOR U62526 ( .A(n49744), .B(n49743), .Z(n55911) );
  IV U62527 ( .A(n49745), .Z(n49747) );
  NOR U62528 ( .A(n49747), .B(n49746), .Z(n55900) );
  NOR U62529 ( .A(n55911), .B(n55900), .Z(n53658) );
  XOR U62530 ( .A(n53659), .B(n53658), .Z(n49748) );
  XOR U62531 ( .A(n53657), .B(n49748), .Z(n53666) );
  IV U62532 ( .A(n49749), .Z(n49750) );
  NOR U62533 ( .A(n49750), .B(n49752), .Z(n53665) );
  IV U62534 ( .A(n49751), .Z(n49753) );
  NOR U62535 ( .A(n49753), .B(n49752), .Z(n53662) );
  NOR U62536 ( .A(n53665), .B(n53662), .Z(n49754) );
  XOR U62537 ( .A(n53666), .B(n49754), .Z(n53672) );
  XOR U62538 ( .A(n53673), .B(n53672), .Z(n52725) );
  XOR U62539 ( .A(n52726), .B(n52725), .Z(n52718) );
  IV U62540 ( .A(n49755), .Z(n49757) );
  NOR U62541 ( .A(n49757), .B(n49756), .Z(n53669) );
  IV U62542 ( .A(n49758), .Z(n49760) );
  NOR U62543 ( .A(n49760), .B(n49759), .Z(n52715) );
  NOR U62544 ( .A(n53669), .B(n52715), .Z(n49761) );
  XOR U62545 ( .A(n52718), .B(n49761), .Z(n53686) );
  XOR U62546 ( .A(n49762), .B(n53686), .Z(n52714) );
  XOR U62547 ( .A(n53685), .B(n52714), .Z(n53683) );
  XOR U62548 ( .A(n49763), .B(n53683), .Z(n52705) );
  XOR U62549 ( .A(n49764), .B(n52705), .Z(n52698) );
  XOR U62550 ( .A(n49765), .B(n52698), .Z(n52693) );
  XOR U62551 ( .A(n49766), .B(n52693), .Z(n52684) );
  IV U62552 ( .A(n52684), .Z(n52682) );
  XOR U62553 ( .A(n52685), .B(n52682), .Z(n53691) );
  XOR U62554 ( .A(n49767), .B(n53691), .Z(n53695) );
  XOR U62555 ( .A(n53693), .B(n53695), .Z(n53700) );
  IV U62556 ( .A(n49768), .Z(n49770) );
  NOR U62557 ( .A(n49770), .B(n49769), .Z(n53696) );
  IV U62558 ( .A(n49771), .Z(n49773) );
  NOR U62559 ( .A(n49773), .B(n49772), .Z(n53699) );
  NOR U62560 ( .A(n53696), .B(n53699), .Z(n49774) );
  XOR U62561 ( .A(n53700), .B(n49774), .Z(n49779) );
  IV U62562 ( .A(n49779), .Z(n53707) );
  NOR U62563 ( .A(n49778), .B(n53707), .Z(n55869) );
  IV U62564 ( .A(n49775), .Z(n49777) );
  NOR U62565 ( .A(n49777), .B(n49776), .Z(n53706) );
  XOR U62566 ( .A(n53706), .B(n49779), .Z(n49781) );
  NOR U62567 ( .A(n49779), .B(n49778), .Z(n49780) );
  NOR U62568 ( .A(n49781), .B(n49780), .Z(n55867) );
  NOR U62569 ( .A(n55869), .B(n55867), .Z(n53710) );
  XOR U62570 ( .A(n53712), .B(n53710), .Z(n52679) );
  IV U62571 ( .A(n49782), .Z(n56857) );
  IV U62572 ( .A(n49783), .Z(n49784) );
  NOR U62573 ( .A(n56857), .B(n49784), .Z(n49785) );
  IV U62574 ( .A(n49785), .Z(n52678) );
  XOR U62575 ( .A(n52679), .B(n52678), .Z(n49788) );
  NOR U62576 ( .A(n49792), .B(n49788), .Z(n49786) );
  IV U62577 ( .A(n49786), .Z(n49787) );
  NOR U62578 ( .A(n49789), .B(n49787), .Z(n49795) );
  IV U62579 ( .A(n49788), .Z(n49791) );
  IV U62580 ( .A(n49789), .Z(n49790) );
  NOR U62581 ( .A(n49791), .B(n49790), .Z(n53714) );
  IV U62582 ( .A(n49792), .Z(n49793) );
  NOR U62583 ( .A(n49793), .B(n52679), .Z(n52680) );
  NOR U62584 ( .A(n53714), .B(n52680), .Z(n55864) );
  IV U62585 ( .A(n55864), .Z(n49794) );
  NOR U62586 ( .A(n49795), .B(n49794), .Z(n49796) );
  IV U62587 ( .A(n49796), .Z(n52677) );
  IV U62588 ( .A(n49797), .Z(n49803) );
  IV U62589 ( .A(n49798), .Z(n49800) );
  NOR U62590 ( .A(n49800), .B(n49799), .Z(n49801) );
  IV U62591 ( .A(n49801), .Z(n49802) );
  NOR U62592 ( .A(n49803), .B(n49802), .Z(n52675) );
  XOR U62593 ( .A(n52677), .B(n52675), .Z(n53719) );
  IV U62594 ( .A(n49804), .Z(n49805) );
  NOR U62595 ( .A(n49805), .B(n49807), .Z(n53717) );
  IV U62596 ( .A(n49806), .Z(n49808) );
  NOR U62597 ( .A(n49808), .B(n49807), .Z(n52673) );
  IV U62598 ( .A(n49809), .Z(n49810) );
  NOR U62599 ( .A(n49810), .B(n49815), .Z(n52671) );
  NOR U62600 ( .A(n52673), .B(n52671), .Z(n49811) );
  IV U62601 ( .A(n49811), .Z(n49812) );
  NOR U62602 ( .A(n53717), .B(n49812), .Z(n49813) );
  XOR U62603 ( .A(n53719), .B(n49813), .Z(n52663) );
  IV U62604 ( .A(n49814), .Z(n49816) );
  NOR U62605 ( .A(n49816), .B(n49815), .Z(n49817) );
  IV U62606 ( .A(n49817), .Z(n52664) );
  XOR U62607 ( .A(n52663), .B(n52664), .Z(n52668) );
  NOR U62608 ( .A(n49824), .B(n52668), .Z(n56872) );
  IV U62609 ( .A(n49818), .Z(n49823) );
  IV U62610 ( .A(n49819), .Z(n49820) );
  NOR U62611 ( .A(n49823), .B(n49820), .Z(n52666) );
  XOR U62612 ( .A(n52668), .B(n52666), .Z(n52662) );
  IV U62613 ( .A(n49821), .Z(n49822) );
  NOR U62614 ( .A(n49823), .B(n49822), .Z(n49825) );
  IV U62615 ( .A(n49825), .Z(n52661) );
  XOR U62616 ( .A(n52662), .B(n52661), .Z(n49827) );
  NOR U62617 ( .A(n49825), .B(n49824), .Z(n49826) );
  NOR U62618 ( .A(n49827), .B(n49826), .Z(n49828) );
  NOR U62619 ( .A(n56872), .B(n49828), .Z(n53724) );
  XOR U62620 ( .A(n53726), .B(n53724), .Z(n53732) );
  IV U62621 ( .A(n49829), .Z(n49831) );
  NOR U62622 ( .A(n49831), .B(n49830), .Z(n53731) );
  NOR U62623 ( .A(n49833), .B(n49832), .Z(n52659) );
  NOR U62624 ( .A(n53731), .B(n52659), .Z(n49834) );
  XOR U62625 ( .A(n53732), .B(n49834), .Z(n53739) );
  XOR U62626 ( .A(n49835), .B(n53739), .Z(n53742) );
  XOR U62627 ( .A(n52656), .B(n53742), .Z(n49843) );
  IV U62628 ( .A(n49836), .Z(n49837) );
  NOR U62629 ( .A(n49838), .B(n49837), .Z(n53741) );
  IV U62630 ( .A(n49839), .Z(n49840) );
  NOR U62631 ( .A(n49841), .B(n49840), .Z(n52657) );
  NOR U62632 ( .A(n53741), .B(n52657), .Z(n49842) );
  XOR U62633 ( .A(n49843), .B(n49842), .Z(n52650) );
  XOR U62634 ( .A(n52648), .B(n52650), .Z(n52652) );
  XOR U62635 ( .A(n52651), .B(n52652), .Z(n49844) );
  NOR U62636 ( .A(n49845), .B(n49844), .Z(n53751) );
  IV U62637 ( .A(n49846), .Z(n49848) );
  NOR U62638 ( .A(n49848), .B(n49847), .Z(n52646) );
  NOR U62639 ( .A(n52651), .B(n52646), .Z(n49849) );
  XOR U62640 ( .A(n52652), .B(n49849), .Z(n49850) );
  NOR U62641 ( .A(n49851), .B(n49850), .Z(n53754) );
  NOR U62642 ( .A(n53751), .B(n53754), .Z(n52639) );
  NOR U62643 ( .A(n49852), .B(n49854), .Z(n52643) );
  IV U62644 ( .A(n49853), .Z(n49855) );
  NOR U62645 ( .A(n49855), .B(n49854), .Z(n52641) );
  NOR U62646 ( .A(n52643), .B(n52641), .Z(n49856) );
  XOR U62647 ( .A(n52639), .B(n49856), .Z(n49857) );
  XOR U62648 ( .A(n49858), .B(n49857), .Z(n52637) );
  XOR U62649 ( .A(n52636), .B(n52637), .Z(n52634) );
  IV U62650 ( .A(n49859), .Z(n49862) );
  IV U62651 ( .A(n49860), .Z(n49861) );
  NOR U62652 ( .A(n49862), .B(n49861), .Z(n52633) );
  XOR U62653 ( .A(n52634), .B(n52633), .Z(n49863) );
  XOR U62654 ( .A(n49864), .B(n49863), .Z(n53761) );
  IV U62655 ( .A(n49865), .Z(n49867) );
  NOR U62656 ( .A(n49867), .B(n49866), .Z(n52631) );
  XOR U62657 ( .A(n53761), .B(n52631), .Z(n53767) );
  XOR U62658 ( .A(n49868), .B(n53767), .Z(n52625) );
  XOR U62659 ( .A(n49869), .B(n52625), .Z(n52623) );
  XOR U62660 ( .A(n49870), .B(n52623), .Z(n53787) );
  XOR U62661 ( .A(n49871), .B(n53787), .Z(n53782) );
  XOR U62662 ( .A(n53780), .B(n53782), .Z(n52612) );
  IV U62663 ( .A(n49872), .Z(n49873) );
  NOR U62664 ( .A(n49876), .B(n49873), .Z(n52610) );
  XOR U62665 ( .A(n52612), .B(n52610), .Z(n52615) );
  IV U62666 ( .A(n49874), .Z(n49875) );
  NOR U62667 ( .A(n49876), .B(n49875), .Z(n52613) );
  XOR U62668 ( .A(n52615), .B(n52613), .Z(n53798) );
  IV U62669 ( .A(n49877), .Z(n52606) );
  NOR U62670 ( .A(n49878), .B(n52606), .Z(n49881) );
  IV U62671 ( .A(n49879), .Z(n49880) );
  NOR U62672 ( .A(n49891), .B(n49880), .Z(n53796) );
  NOR U62673 ( .A(n49881), .B(n53796), .Z(n49882) );
  XOR U62674 ( .A(n53798), .B(n49882), .Z(n49893) );
  IV U62675 ( .A(n49893), .Z(n53795) );
  IV U62676 ( .A(n49883), .Z(n49884) );
  NOR U62677 ( .A(n49885), .B(n49884), .Z(n49886) );
  IV U62678 ( .A(n49886), .Z(n49894) );
  NOR U62679 ( .A(n53795), .B(n49894), .Z(n56975) );
  IV U62680 ( .A(n49887), .Z(n49889) );
  NOR U62681 ( .A(n49889), .B(n49888), .Z(n53802) );
  IV U62682 ( .A(n49890), .Z(n49892) );
  NOR U62683 ( .A(n49892), .B(n49891), .Z(n53793) );
  XOR U62684 ( .A(n53793), .B(n49893), .Z(n53803) );
  XOR U62685 ( .A(n53802), .B(n53803), .Z(n49896) );
  NOR U62686 ( .A(n53803), .B(n49894), .Z(n49895) );
  NOR U62687 ( .A(n49896), .B(n49895), .Z(n49897) );
  NOR U62688 ( .A(n56975), .B(n49897), .Z(n49908) );
  IV U62689 ( .A(n49908), .Z(n52603) );
  IV U62690 ( .A(n49898), .Z(n49899) );
  NOR U62691 ( .A(n49900), .B(n49899), .Z(n52602) );
  IV U62692 ( .A(n49901), .Z(n49903) );
  NOR U62693 ( .A(n49903), .B(n49902), .Z(n49907) );
  NOR U62694 ( .A(n52602), .B(n49907), .Z(n49904) );
  XOR U62695 ( .A(n52603), .B(n49904), .Z(n49905) );
  NOR U62696 ( .A(n49906), .B(n49905), .Z(n49913) );
  IV U62697 ( .A(n49906), .Z(n49912) );
  XOR U62698 ( .A(n52602), .B(n49908), .Z(n49910) );
  IV U62699 ( .A(n49907), .Z(n52599) );
  NOR U62700 ( .A(n49908), .B(n52599), .Z(n49909) );
  NOR U62701 ( .A(n49910), .B(n49909), .Z(n49911) );
  NOR U62702 ( .A(n49912), .B(n49911), .Z(n52600) );
  NOR U62703 ( .A(n49913), .B(n52600), .Z(n52585) );
  IV U62704 ( .A(n49914), .Z(n49916) );
  NOR U62705 ( .A(n49916), .B(n49915), .Z(n49917) );
  IV U62706 ( .A(n49917), .Z(n52586) );
  XOR U62707 ( .A(n52585), .B(n52586), .Z(n52589) );
  XOR U62708 ( .A(n52588), .B(n52589), .Z(n52593) );
  XOR U62709 ( .A(n52591), .B(n52593), .Z(n52577) );
  XOR U62710 ( .A(n52579), .B(n52577), .Z(n52574) );
  XOR U62711 ( .A(n49918), .B(n52574), .Z(n52572) );
  XOR U62712 ( .A(n52570), .B(n52572), .Z(n53814) );
  XOR U62713 ( .A(n53813), .B(n53814), .Z(n52568) );
  XOR U62714 ( .A(n52567), .B(n52568), .Z(n53837) );
  IV U62715 ( .A(n49919), .Z(n49920) );
  NOR U62716 ( .A(n49921), .B(n49920), .Z(n53838) );
  IV U62717 ( .A(n49922), .Z(n49923) );
  NOR U62718 ( .A(n49924), .B(n49923), .Z(n53823) );
  NOR U62719 ( .A(n53838), .B(n53823), .Z(n49925) );
  XOR U62720 ( .A(n53837), .B(n49925), .Z(n52560) );
  XOR U62721 ( .A(n49926), .B(n52560), .Z(n52558) );
  XOR U62722 ( .A(n52556), .B(n52558), .Z(n52554) );
  IV U62723 ( .A(n49927), .Z(n49928) );
  NOR U62724 ( .A(n49929), .B(n49928), .Z(n52553) );
  IV U62725 ( .A(n49930), .Z(n49931) );
  NOR U62726 ( .A(n49932), .B(n49931), .Z(n52551) );
  NOR U62727 ( .A(n52553), .B(n52551), .Z(n49933) );
  XOR U62728 ( .A(n52554), .B(n49933), .Z(n52543) );
  IV U62729 ( .A(n49934), .Z(n49935) );
  NOR U62730 ( .A(n49935), .B(n49937), .Z(n52546) );
  IV U62731 ( .A(n49936), .Z(n49938) );
  NOR U62732 ( .A(n49938), .B(n49937), .Z(n52545) );
  XOR U62733 ( .A(n52546), .B(n52545), .Z(n49939) );
  NOR U62734 ( .A(n53842), .B(n49939), .Z(n49940) );
  XOR U62735 ( .A(n52543), .B(n49940), .Z(n53847) );
  IV U62736 ( .A(n49941), .Z(n49944) );
  IV U62737 ( .A(n49942), .Z(n49943) );
  NOR U62738 ( .A(n49944), .B(n49943), .Z(n53845) );
  XOR U62739 ( .A(n53847), .B(n53845), .Z(n53859) );
  IV U62740 ( .A(n49945), .Z(n49948) );
  IV U62741 ( .A(n49946), .Z(n49947) );
  NOR U62742 ( .A(n49948), .B(n49947), .Z(n53857) );
  XOR U62743 ( .A(n53859), .B(n53857), .Z(n52541) );
  XOR U62744 ( .A(n49949), .B(n52541), .Z(n53873) );
  IV U62745 ( .A(n53873), .Z(n49959) );
  IV U62746 ( .A(n49954), .Z(n49951) );
  IV U62747 ( .A(n49953), .Z(n49950) );
  NOR U62748 ( .A(n49951), .B(n49950), .Z(n52540) );
  IV U62749 ( .A(n49952), .Z(n49956) );
  NOR U62750 ( .A(n49954), .B(n49953), .Z(n49955) );
  NOR U62751 ( .A(n49956), .B(n49955), .Z(n49957) );
  NOR U62752 ( .A(n52540), .B(n49957), .Z(n49958) );
  XOR U62753 ( .A(n49959), .B(n49958), .Z(n49968) );
  IV U62754 ( .A(n49960), .Z(n49962) );
  NOR U62755 ( .A(n49962), .B(n49961), .Z(n49970) );
  IV U62756 ( .A(n49970), .Z(n49963) );
  NOR U62757 ( .A(n49968), .B(n49963), .Z(n57045) );
  IV U62758 ( .A(n49964), .Z(n49966) );
  IV U62759 ( .A(n49965), .Z(n53870) );
  NOR U62760 ( .A(n49966), .B(n53870), .Z(n49967) );
  XOR U62761 ( .A(n49968), .B(n49967), .Z(n52536) );
  IV U62762 ( .A(n52536), .Z(n49969) );
  NOR U62763 ( .A(n49970), .B(n49969), .Z(n49971) );
  NOR U62764 ( .A(n57045), .B(n49971), .Z(n52531) );
  XOR U62765 ( .A(n53879), .B(n52531), .Z(n53886) );
  IV U62766 ( .A(n49972), .Z(n49974) );
  NOR U62767 ( .A(n49974), .B(n49973), .Z(n53884) );
  XOR U62768 ( .A(n53886), .B(n53884), .Z(n53888) );
  XOR U62769 ( .A(n53887), .B(n53888), .Z(n52529) );
  IV U62770 ( .A(n49975), .Z(n49976) );
  NOR U62771 ( .A(n49982), .B(n49976), .Z(n49977) );
  IV U62772 ( .A(n49977), .Z(n52527) );
  XOR U62773 ( .A(n52529), .B(n52527), .Z(n49978) );
  XOR U62774 ( .A(n49979), .B(n49978), .Z(n52523) );
  IV U62775 ( .A(n49980), .Z(n49981) );
  NOR U62776 ( .A(n49982), .B(n49981), .Z(n52521) );
  XOR U62777 ( .A(n52523), .B(n52521), .Z(n52526) );
  XOR U62778 ( .A(n52524), .B(n52526), .Z(n52516) );
  XOR U62779 ( .A(n52515), .B(n52516), .Z(n52520) );
  XOR U62780 ( .A(n52518), .B(n52520), .Z(n52506) );
  XOR U62781 ( .A(n52505), .B(n52506), .Z(n52510) );
  XOR U62782 ( .A(n49983), .B(n52510), .Z(n53903) );
  XOR U62783 ( .A(n49984), .B(n53903), .Z(n53901) );
  XOR U62784 ( .A(n53899), .B(n53901), .Z(n53908) );
  XOR U62785 ( .A(n53909), .B(n53908), .Z(n53910) );
  XOR U62786 ( .A(n53912), .B(n53910), .Z(n53915) );
  IV U62787 ( .A(n49985), .Z(n49987) );
  NOR U62788 ( .A(n49987), .B(n49986), .Z(n53913) );
  XOR U62789 ( .A(n53915), .B(n53913), .Z(n52496) );
  IV U62790 ( .A(n49988), .Z(n49989) );
  NOR U62791 ( .A(n49990), .B(n49989), .Z(n49991) );
  IV U62792 ( .A(n49991), .Z(n52495) );
  NOR U62793 ( .A(n49992), .B(n52495), .Z(n49993) );
  XOR U62794 ( .A(n52496), .B(n49993), .Z(n53926) );
  IV U62795 ( .A(n49994), .Z(n49995) );
  NOR U62796 ( .A(n49998), .B(n49995), .Z(n52492) );
  IV U62797 ( .A(n49996), .Z(n49997) );
  NOR U62798 ( .A(n49998), .B(n49997), .Z(n53925) );
  NOR U62799 ( .A(n52492), .B(n53925), .Z(n49999) );
  XOR U62800 ( .A(n53926), .B(n49999), .Z(n50007) );
  IV U62801 ( .A(n50007), .Z(n50005) );
  IV U62802 ( .A(n50000), .Z(n50003) );
  IV U62803 ( .A(n50001), .Z(n50002) );
  NOR U62804 ( .A(n50003), .B(n50002), .Z(n50010) );
  IV U62805 ( .A(n50010), .Z(n50004) );
  NOR U62806 ( .A(n50005), .B(n50004), .Z(n55741) );
  IV U62807 ( .A(n50008), .Z(n50006) );
  NOR U62808 ( .A(n50006), .B(n53926), .Z(n55740) );
  NOR U62809 ( .A(n50008), .B(n50007), .Z(n50009) );
  NOR U62810 ( .A(n55740), .B(n50009), .Z(n50015) );
  NOR U62811 ( .A(n50010), .B(n50015), .Z(n50011) );
  NOR U62812 ( .A(n55741), .B(n50011), .Z(n50022) );
  IV U62813 ( .A(n50012), .Z(n50024) );
  IV U62814 ( .A(n50013), .Z(n50014) );
  NOR U62815 ( .A(n50024), .B(n50014), .Z(n50016) );
  NOR U62816 ( .A(n50022), .B(n50016), .Z(n50019) );
  IV U62817 ( .A(n50015), .Z(n50018) );
  IV U62818 ( .A(n50016), .Z(n50017) );
  NOR U62819 ( .A(n50018), .B(n50017), .Z(n57142) );
  NOR U62820 ( .A(n50019), .B(n57142), .Z(n53930) );
  IV U62821 ( .A(n50020), .Z(n50021) );
  NOR U62822 ( .A(n50045), .B(n50021), .Z(n50032) );
  IV U62823 ( .A(n50032), .Z(n53932) );
  NOR U62824 ( .A(n53930), .B(n53932), .Z(n50034) );
  IV U62825 ( .A(n50022), .Z(n50027) );
  IV U62826 ( .A(n50023), .Z(n50025) );
  NOR U62827 ( .A(n50025), .B(n50024), .Z(n50028) );
  IV U62828 ( .A(n50028), .Z(n50026) );
  NOR U62829 ( .A(n50027), .B(n50026), .Z(n52491) );
  NOR U62830 ( .A(n53930), .B(n50028), .Z(n50029) );
  NOR U62831 ( .A(n52491), .B(n50029), .Z(n50030) );
  IV U62832 ( .A(n50030), .Z(n50031) );
  NOR U62833 ( .A(n50032), .B(n50031), .Z(n50033) );
  NOR U62834 ( .A(n50034), .B(n50033), .Z(n53934) );
  IV U62835 ( .A(n50035), .Z(n50041) );
  IV U62836 ( .A(n50036), .Z(n50037) );
  NOR U62837 ( .A(n50038), .B(n50037), .Z(n50039) );
  IV U62838 ( .A(n50039), .Z(n50040) );
  NOR U62839 ( .A(n50041), .B(n50040), .Z(n50042) );
  IV U62840 ( .A(n50042), .Z(n52490) );
  XOR U62841 ( .A(n53934), .B(n52490), .Z(n50043) );
  XOR U62842 ( .A(n53933), .B(n50043), .Z(n52489) );
  IV U62843 ( .A(n50044), .Z(n50048) );
  NOR U62844 ( .A(n50046), .B(n50045), .Z(n50047) );
  IV U62845 ( .A(n50047), .Z(n50050) );
  NOR U62846 ( .A(n50048), .B(n50050), .Z(n52487) );
  XOR U62847 ( .A(n52489), .B(n52487), .Z(n53939) );
  IV U62848 ( .A(n50049), .Z(n50051) );
  NOR U62849 ( .A(n50051), .B(n50050), .Z(n50052) );
  IV U62850 ( .A(n50052), .Z(n53938) );
  XOR U62851 ( .A(n53939), .B(n53938), .Z(n52482) );
  IV U62852 ( .A(n50053), .Z(n50054) );
  NOR U62853 ( .A(n50055), .B(n50054), .Z(n52484) );
  IV U62854 ( .A(n50056), .Z(n50058) );
  NOR U62855 ( .A(n50058), .B(n50057), .Z(n52481) );
  NOR U62856 ( .A(n52484), .B(n52481), .Z(n50059) );
  XOR U62857 ( .A(n52482), .B(n50059), .Z(n53948) );
  XOR U62858 ( .A(n53947), .B(n53948), .Z(n52480) );
  XOR U62859 ( .A(n52478), .B(n52480), .Z(n53960) );
  XOR U62860 ( .A(n50060), .B(n53960), .Z(n50061) );
  IV U62861 ( .A(n50061), .Z(n52472) );
  IV U62862 ( .A(n50062), .Z(n50063) );
  NOR U62863 ( .A(n50064), .B(n50063), .Z(n52470) );
  XOR U62864 ( .A(n52472), .B(n52470), .Z(n52474) );
  XOR U62865 ( .A(n52473), .B(n52474), .Z(n53965) );
  IV U62866 ( .A(n50065), .Z(n50066) );
  NOR U62867 ( .A(n50067), .B(n50066), .Z(n52467) );
  IV U62868 ( .A(n50068), .Z(n50070) );
  NOR U62869 ( .A(n50070), .B(n50069), .Z(n53964) );
  NOR U62870 ( .A(n52467), .B(n53964), .Z(n50071) );
  XOR U62871 ( .A(n53965), .B(n50071), .Z(n50072) );
  XOR U62872 ( .A(n50073), .B(n50072), .Z(n52461) );
  XOR U62873 ( .A(n52460), .B(n52461), .Z(n52456) );
  IV U62874 ( .A(n50074), .Z(n50075) );
  NOR U62875 ( .A(n50075), .B(n50077), .Z(n52462) );
  IV U62876 ( .A(n50076), .Z(n50078) );
  NOR U62877 ( .A(n50078), .B(n50077), .Z(n52455) );
  NOR U62878 ( .A(n52462), .B(n52455), .Z(n50079) );
  XOR U62879 ( .A(n52456), .B(n50079), .Z(n52454) );
  IV U62880 ( .A(n50080), .Z(n50081) );
  NOR U62881 ( .A(n50081), .B(n50085), .Z(n52452) );
  XOR U62882 ( .A(n52454), .B(n52452), .Z(n52450) );
  XOR U62883 ( .A(n52446), .B(n52450), .Z(n50088) );
  NOR U62884 ( .A(n50083), .B(n50082), .Z(n52447) );
  IV U62885 ( .A(n50084), .Z(n50086) );
  NOR U62886 ( .A(n50086), .B(n50085), .Z(n52449) );
  NOR U62887 ( .A(n52447), .B(n52449), .Z(n50087) );
  XOR U62888 ( .A(n50088), .B(n50087), .Z(n52441) );
  XOR U62889 ( .A(n52439), .B(n52441), .Z(n52442) );
  XOR U62890 ( .A(n52443), .B(n52442), .Z(n50089) );
  IV U62891 ( .A(n50089), .Z(n52437) );
  XOR U62892 ( .A(n52429), .B(n52437), .Z(n52432) );
  IV U62893 ( .A(n50090), .Z(n50091) );
  NOR U62894 ( .A(n50092), .B(n50091), .Z(n52436) );
  IV U62895 ( .A(n50093), .Z(n50095) );
  NOR U62896 ( .A(n50095), .B(n50094), .Z(n52431) );
  NOR U62897 ( .A(n52436), .B(n52431), .Z(n50096) );
  XOR U62898 ( .A(n52432), .B(n50096), .Z(n50097) );
  NOR U62899 ( .A(n50098), .B(n50097), .Z(n50101) );
  IV U62900 ( .A(n50098), .Z(n50100) );
  XOR U62901 ( .A(n52436), .B(n52432), .Z(n50099) );
  NOR U62902 ( .A(n50100), .B(n50099), .Z(n53982) );
  NOR U62903 ( .A(n50101), .B(n53982), .Z(n53976) );
  IV U62904 ( .A(n50102), .Z(n53978) );
  XOR U62905 ( .A(n53976), .B(n53978), .Z(n53987) );
  XOR U62906 ( .A(n50103), .B(n53987), .Z(n53995) );
  XOR U62907 ( .A(n52424), .B(n53995), .Z(n52422) );
  IV U62908 ( .A(n50104), .Z(n50105) );
  NOR U62909 ( .A(n50106), .B(n50105), .Z(n52421) );
  IV U62910 ( .A(n50107), .Z(n50109) );
  NOR U62911 ( .A(n50109), .B(n50108), .Z(n53993) );
  NOR U62912 ( .A(n52421), .B(n53993), .Z(n50110) );
  XOR U62913 ( .A(n52422), .B(n50110), .Z(n52418) );
  IV U62914 ( .A(n50111), .Z(n50112) );
  NOR U62915 ( .A(n50113), .B(n50112), .Z(n50118) );
  IV U62916 ( .A(n50114), .Z(n50116) );
  NOR U62917 ( .A(n50116), .B(n50115), .Z(n50117) );
  NOR U62918 ( .A(n50118), .B(n50117), .Z(n52419) );
  XOR U62919 ( .A(n52418), .B(n52419), .Z(n52416) );
  XOR U62920 ( .A(n52417), .B(n52416), .Z(n52408) );
  IV U62921 ( .A(n50119), .Z(n50120) );
  NOR U62922 ( .A(n50121), .B(n50120), .Z(n50126) );
  IV U62923 ( .A(n50122), .Z(n50123) );
  NOR U62924 ( .A(n50124), .B(n50123), .Z(n50125) );
  NOR U62925 ( .A(n50126), .B(n50125), .Z(n52410) );
  XOR U62926 ( .A(n52408), .B(n52410), .Z(n52412) );
  XOR U62927 ( .A(n52411), .B(n52412), .Z(n52400) );
  XOR U62928 ( .A(n50127), .B(n52400), .Z(n54000) );
  XOR U62929 ( .A(n53998), .B(n54000), .Z(n54007) );
  IV U62930 ( .A(n50128), .Z(n50130) );
  NOR U62931 ( .A(n50130), .B(n50129), .Z(n54005) );
  XOR U62932 ( .A(n54007), .B(n54005), .Z(n54010) );
  IV U62933 ( .A(n50131), .Z(n50133) );
  NOR U62934 ( .A(n50133), .B(n50132), .Z(n54008) );
  XOR U62935 ( .A(n54010), .B(n54008), .Z(n54017) );
  IV U62936 ( .A(n50134), .Z(n50136) );
  NOR U62937 ( .A(n50136), .B(n50135), .Z(n54015) );
  XOR U62938 ( .A(n54017), .B(n54015), .Z(n54013) );
  XOR U62939 ( .A(n54012), .B(n54013), .Z(n52393) );
  XOR U62940 ( .A(n52392), .B(n52393), .Z(n52396) );
  XOR U62941 ( .A(n52395), .B(n52396), .Z(n54029) );
  IV U62942 ( .A(n54029), .Z(n50148) );
  IV U62943 ( .A(n50137), .Z(n50139) );
  NOR U62944 ( .A(n50139), .B(n50138), .Z(n50147) );
  IV U62945 ( .A(n50140), .Z(n50142) );
  IV U62946 ( .A(n50141), .Z(n50149) );
  NOR U62947 ( .A(n50142), .B(n50149), .Z(n50143) );
  NOR U62948 ( .A(n50147), .B(n50143), .Z(n50144) );
  XOR U62949 ( .A(n50148), .B(n50144), .Z(n50145) );
  NOR U62950 ( .A(n50146), .B(n50145), .Z(n55634) );
  IV U62951 ( .A(n50147), .Z(n54030) );
  XOR U62952 ( .A(n54030), .B(n50148), .Z(n54043) );
  NOR U62953 ( .A(n50150), .B(n50149), .Z(n54027) );
  IV U62954 ( .A(n50151), .Z(n50153) );
  NOR U62955 ( .A(n50153), .B(n50152), .Z(n54041) );
  NOR U62956 ( .A(n54027), .B(n54041), .Z(n50154) );
  XOR U62957 ( .A(n54043), .B(n50154), .Z(n50155) );
  NOR U62958 ( .A(n50156), .B(n50155), .Z(n50157) );
  NOR U62959 ( .A(n55634), .B(n50157), .Z(n54046) );
  XOR U62960 ( .A(n54045), .B(n54046), .Z(n52390) );
  IV U62961 ( .A(n50158), .Z(n50160) );
  NOR U62962 ( .A(n50160), .B(n50159), .Z(n54050) );
  NOR U62963 ( .A(n52389), .B(n54050), .Z(n50161) );
  XOR U62964 ( .A(n52390), .B(n50161), .Z(n54055) );
  XOR U62965 ( .A(n54053), .B(n54055), .Z(n54058) );
  XOR U62966 ( .A(n50162), .B(n54058), .Z(n54063) );
  XOR U62967 ( .A(n54061), .B(n54063), .Z(n54066) );
  IV U62968 ( .A(n50163), .Z(n50165) );
  NOR U62969 ( .A(n50165), .B(n50164), .Z(n54064) );
  XOR U62970 ( .A(n54066), .B(n54064), .Z(n52382) );
  IV U62971 ( .A(n50166), .Z(n50168) );
  NOR U62972 ( .A(n50168), .B(n50167), .Z(n52380) );
  XOR U62973 ( .A(n52382), .B(n52380), .Z(n52384) );
  XOR U62974 ( .A(n52383), .B(n52384), .Z(n52373) );
  XOR U62975 ( .A(n52372), .B(n52373), .Z(n52377) );
  IV U62976 ( .A(n50169), .Z(n50172) );
  IV U62977 ( .A(n50170), .Z(n50171) );
  NOR U62978 ( .A(n50172), .B(n50171), .Z(n52375) );
  XOR U62979 ( .A(n52377), .B(n52375), .Z(n52368) );
  IV U62980 ( .A(n50173), .Z(n50175) );
  NOR U62981 ( .A(n50175), .B(n50174), .Z(n50176) );
  IV U62982 ( .A(n50176), .Z(n52366) );
  XOR U62983 ( .A(n52368), .B(n52366), .Z(n50177) );
  XOR U62984 ( .A(n50178), .B(n50177), .Z(n52356) );
  IV U62985 ( .A(n52356), .Z(n50184) );
  NOR U62986 ( .A(n52357), .B(n50179), .Z(n50182) );
  IV U62987 ( .A(n50180), .Z(n50181) );
  NOR U62988 ( .A(n52357), .B(n50181), .Z(n52348) );
  NOR U62989 ( .A(n50182), .B(n52348), .Z(n50183) );
  XOR U62990 ( .A(n50184), .B(n50183), .Z(n52352) );
  XOR U62991 ( .A(n52345), .B(n52352), .Z(n50185) );
  XOR U62992 ( .A(n50186), .B(n50185), .Z(n52343) );
  IV U62993 ( .A(n50187), .Z(n50188) );
  NOR U62994 ( .A(n50188), .B(n50191), .Z(n52341) );
  XOR U62995 ( .A(n52343), .B(n52341), .Z(n52335) );
  IV U62996 ( .A(n50189), .Z(n50190) );
  NOR U62997 ( .A(n50191), .B(n50190), .Z(n50192) );
  IV U62998 ( .A(n50192), .Z(n52334) );
  XOR U62999 ( .A(n52335), .B(n52334), .Z(n52336) );
  IV U63000 ( .A(n50193), .Z(n50194) );
  NOR U63001 ( .A(n50195), .B(n50194), .Z(n50200) );
  IV U63002 ( .A(n50196), .Z(n50197) );
  NOR U63003 ( .A(n50198), .B(n50197), .Z(n50199) );
  NOR U63004 ( .A(n50200), .B(n50199), .Z(n52338) );
  XOR U63005 ( .A(n52336), .B(n52338), .Z(n52330) );
  XOR U63006 ( .A(n52328), .B(n52330), .Z(n52333) );
  XOR U63007 ( .A(n52331), .B(n52333), .Z(n52322) );
  XOR U63008 ( .A(n52320), .B(n52322), .Z(n52325) );
  XOR U63009 ( .A(n50201), .B(n52325), .Z(n50209) );
  NOR U63010 ( .A(n50203), .B(n50202), .Z(n52318) );
  IV U63011 ( .A(n50204), .Z(n50207) );
  IV U63012 ( .A(n50205), .Z(n50206) );
  NOR U63013 ( .A(n50207), .B(n50206), .Z(n52313) );
  NOR U63014 ( .A(n52318), .B(n52313), .Z(n50208) );
  XOR U63015 ( .A(n50209), .B(n50208), .Z(n52312) );
  XOR U63016 ( .A(n52310), .B(n52312), .Z(n52306) );
  XOR U63017 ( .A(n52304), .B(n52306), .Z(n50210) );
  XOR U63018 ( .A(n50211), .B(n50210), .Z(n52298) );
  XOR U63019 ( .A(n52296), .B(n52298), .Z(n52300) );
  XOR U63020 ( .A(n52299), .B(n52300), .Z(n52294) );
  XOR U63021 ( .A(n52293), .B(n52294), .Z(n52291) );
  XOR U63022 ( .A(n52292), .B(n52291), .Z(n50212) );
  XOR U63023 ( .A(n52290), .B(n50212), .Z(n54076) );
  IV U63024 ( .A(n50213), .Z(n50215) );
  NOR U63025 ( .A(n50215), .B(n50214), .Z(n54074) );
  XOR U63026 ( .A(n54076), .B(n54074), .Z(n54078) );
  IV U63027 ( .A(n50216), .Z(n50218) );
  NOR U63028 ( .A(n50218), .B(n50217), .Z(n50219) );
  IV U63029 ( .A(n50219), .Z(n54077) );
  XOR U63030 ( .A(n54078), .B(n54077), .Z(n52285) );
  IV U63031 ( .A(n50220), .Z(n50221) );
  NOR U63032 ( .A(n50222), .B(n50221), .Z(n52284) );
  IV U63033 ( .A(n50223), .Z(n50225) );
  NOR U63034 ( .A(n50225), .B(n50224), .Z(n52287) );
  NOR U63035 ( .A(n52284), .B(n52287), .Z(n50226) );
  XOR U63036 ( .A(n52285), .B(n50226), .Z(n52279) );
  XOR U63037 ( .A(n52277), .B(n52279), .Z(n52282) );
  XOR U63038 ( .A(n52275), .B(n52282), .Z(n50227) );
  XOR U63039 ( .A(n52280), .B(n50227), .Z(n54082) );
  XOR U63040 ( .A(n54081), .B(n54082), .Z(n54085) );
  XOR U63041 ( .A(n54084), .B(n54085), .Z(n52269) );
  XOR U63042 ( .A(n52267), .B(n52269), .Z(n52271) );
  XOR U63043 ( .A(n52270), .B(n52271), .Z(n54095) );
  XOR U63044 ( .A(n50228), .B(n54095), .Z(n54098) );
  XOR U63045 ( .A(n52263), .B(n54098), .Z(n52261) );
  XOR U63046 ( .A(n52258), .B(n52261), .Z(n50229) );
  XOR U63047 ( .A(n50230), .B(n50229), .Z(n54104) );
  IV U63048 ( .A(n50231), .Z(n50234) );
  IV U63049 ( .A(n50232), .Z(n50233) );
  NOR U63050 ( .A(n50234), .B(n50233), .Z(n54101) );
  XOR U63051 ( .A(n54104), .B(n54101), .Z(n52255) );
  IV U63052 ( .A(n50235), .Z(n50236) );
  NOR U63053 ( .A(n50239), .B(n50236), .Z(n52256) );
  IV U63054 ( .A(n50237), .Z(n50238) );
  NOR U63055 ( .A(n50239), .B(n50238), .Z(n52253) );
  NOR U63056 ( .A(n52256), .B(n52253), .Z(n50240) );
  XOR U63057 ( .A(n52255), .B(n50240), .Z(n52247) );
  XOR U63058 ( .A(n50241), .B(n52247), .Z(n52243) );
  XOR U63059 ( .A(n52241), .B(n52243), .Z(n52244) );
  XOR U63060 ( .A(n52245), .B(n52244), .Z(n52236) );
  IV U63061 ( .A(n50242), .Z(n50244) );
  NOR U63062 ( .A(n50244), .B(n50243), .Z(n52238) );
  IV U63063 ( .A(n50245), .Z(n50247) );
  NOR U63064 ( .A(n50247), .B(n50246), .Z(n52235) );
  NOR U63065 ( .A(n52238), .B(n52235), .Z(n50248) );
  XOR U63066 ( .A(n52236), .B(n50248), .Z(n52233) );
  XOR U63067 ( .A(n50249), .B(n52233), .Z(n52223) );
  XOR U63068 ( .A(n52222), .B(n52223), .Z(n52227) );
  IV U63069 ( .A(n50250), .Z(n50252) );
  NOR U63070 ( .A(n50252), .B(n50251), .Z(n52225) );
  XOR U63071 ( .A(n52227), .B(n52225), .Z(n52215) );
  XOR U63072 ( .A(n52214), .B(n52215), .Z(n52218) );
  XOR U63073 ( .A(n52217), .B(n52218), .Z(n52213) );
  IV U63074 ( .A(n52213), .Z(n50260) );
  IV U63075 ( .A(n50253), .Z(n50255) );
  NOR U63076 ( .A(n50255), .B(n50254), .Z(n52209) );
  IV U63077 ( .A(n50256), .Z(n50257) );
  NOR U63078 ( .A(n50258), .B(n50257), .Z(n52211) );
  NOR U63079 ( .A(n52209), .B(n52211), .Z(n50259) );
  XOR U63080 ( .A(n50260), .B(n50259), .Z(n52200) );
  XOR U63081 ( .A(n50261), .B(n52200), .Z(n52190) );
  XOR U63082 ( .A(n50262), .B(n52190), .Z(n54115) );
  XOR U63083 ( .A(n50263), .B(n54115), .Z(n52185) );
  IV U63084 ( .A(n50264), .Z(n50265) );
  NOR U63085 ( .A(n50266), .B(n50265), .Z(n52182) );
  IV U63086 ( .A(n50267), .Z(n50269) );
  NOR U63087 ( .A(n50269), .B(n50268), .Z(n52184) );
  NOR U63088 ( .A(n52182), .B(n52184), .Z(n50270) );
  XOR U63089 ( .A(n52185), .B(n50270), .Z(n50271) );
  NOR U63090 ( .A(n50272), .B(n50271), .Z(n50275) );
  IV U63091 ( .A(n50272), .Z(n50274) );
  XOR U63092 ( .A(n52182), .B(n52185), .Z(n50273) );
  NOR U63093 ( .A(n50274), .B(n50273), .Z(n52181) );
  NOR U63094 ( .A(n50275), .B(n52181), .Z(n52173) );
  IV U63095 ( .A(n50276), .Z(n50277) );
  NOR U63096 ( .A(n50278), .B(n50277), .Z(n52177) );
  IV U63097 ( .A(n50279), .Z(n50280) );
  NOR U63098 ( .A(n50282), .B(n50280), .Z(n52175) );
  IV U63099 ( .A(n50281), .Z(n50283) );
  NOR U63100 ( .A(n50283), .B(n50282), .Z(n52172) );
  NOR U63101 ( .A(n52175), .B(n52172), .Z(n50284) );
  XOR U63102 ( .A(n52177), .B(n50284), .Z(n50285) );
  XOR U63103 ( .A(n52173), .B(n50285), .Z(n52171) );
  XOR U63104 ( .A(n50286), .B(n52171), .Z(n50287) );
  IV U63105 ( .A(n50287), .Z(n52161) );
  XOR U63106 ( .A(n52159), .B(n52161), .Z(n52163) );
  XOR U63107 ( .A(n52162), .B(n52163), .Z(n52152) );
  XOR U63108 ( .A(n52151), .B(n52152), .Z(n52155) );
  XOR U63109 ( .A(n50288), .B(n52155), .Z(n54146) );
  IV U63110 ( .A(n50289), .Z(n50291) );
  NOR U63111 ( .A(n50291), .B(n50290), .Z(n54145) );
  XOR U63112 ( .A(n54146), .B(n54145), .Z(n54150) );
  XOR U63113 ( .A(n54148), .B(n54150), .Z(n52136) );
  XOR U63114 ( .A(n52137), .B(n52136), .Z(n54165) );
  XOR U63115 ( .A(n50292), .B(n54165), .Z(n54162) );
  XOR U63116 ( .A(n54160), .B(n54162), .Z(n54170) );
  IV U63117 ( .A(n50293), .Z(n50294) );
  NOR U63118 ( .A(n50302), .B(n50294), .Z(n54169) );
  IV U63119 ( .A(n50295), .Z(n50296) );
  NOR U63120 ( .A(n50297), .B(n50296), .Z(n54168) );
  NOR U63121 ( .A(n54169), .B(n54168), .Z(n50298) );
  XOR U63122 ( .A(n54170), .B(n50298), .Z(n50310) );
  IV U63123 ( .A(n50310), .Z(n50299) );
  NOR U63124 ( .A(n50300), .B(n50299), .Z(n54176) );
  XOR U63125 ( .A(n54169), .B(n54170), .Z(n50308) );
  IV U63126 ( .A(n50301), .Z(n50306) );
  NOR U63127 ( .A(n50303), .B(n50302), .Z(n50304) );
  IV U63128 ( .A(n50304), .Z(n50305) );
  NOR U63129 ( .A(n50306), .B(n50305), .Z(n50309) );
  IV U63130 ( .A(n50309), .Z(n50307) );
  NOR U63131 ( .A(n50308), .B(n50307), .Z(n54173) );
  NOR U63132 ( .A(n50310), .B(n50309), .Z(n50311) );
  NOR U63133 ( .A(n54173), .B(n50311), .Z(n50312) );
  NOR U63134 ( .A(n50313), .B(n50312), .Z(n50314) );
  NOR U63135 ( .A(n54176), .B(n50314), .Z(n54181) );
  IV U63136 ( .A(n50315), .Z(n54183) );
  XOR U63137 ( .A(n54181), .B(n54183), .Z(n54194) );
  XOR U63138 ( .A(n50316), .B(n54194), .Z(n54204) );
  XOR U63139 ( .A(n54203), .B(n54204), .Z(n52128) );
  XOR U63140 ( .A(n52126), .B(n52128), .Z(n54210) );
  IV U63141 ( .A(n50317), .Z(n50318) );
  NOR U63142 ( .A(n50321), .B(n50318), .Z(n52127) );
  IV U63143 ( .A(n50319), .Z(n50320) );
  NOR U63144 ( .A(n50321), .B(n50320), .Z(n54209) );
  NOR U63145 ( .A(n52127), .B(n54209), .Z(n50322) );
  XOR U63146 ( .A(n54210), .B(n50322), .Z(n52121) );
  IV U63147 ( .A(n50323), .Z(n50324) );
  NOR U63148 ( .A(n50325), .B(n50324), .Z(n54212) );
  NOR U63149 ( .A(n52122), .B(n54212), .Z(n50326) );
  XOR U63150 ( .A(n52121), .B(n50326), .Z(n54216) );
  XOR U63151 ( .A(n54215), .B(n54216), .Z(n52118) );
  XOR U63152 ( .A(n52119), .B(n52118), .Z(n52104) );
  NOR U63153 ( .A(n50328), .B(n50327), .Z(n52114) );
  NOR U63154 ( .A(n52103), .B(n52114), .Z(n50329) );
  NOR U63155 ( .A(n52104), .B(n50329), .Z(n50340) );
  IV U63156 ( .A(n50329), .Z(n50338) );
  IV U63157 ( .A(n50330), .Z(n50331) );
  NOR U63158 ( .A(n50332), .B(n50331), .Z(n50334) );
  IV U63159 ( .A(n50334), .Z(n50333) );
  NOR U63160 ( .A(n50333), .B(n52118), .Z(n55451) );
  NOR U63161 ( .A(n50334), .B(n52104), .Z(n50335) );
  NOR U63162 ( .A(n55451), .B(n50335), .Z(n50336) );
  IV U63163 ( .A(n50336), .Z(n50337) );
  NOR U63164 ( .A(n50338), .B(n50337), .Z(n50339) );
  NOR U63165 ( .A(n50340), .B(n50339), .Z(n52107) );
  XOR U63166 ( .A(n52106), .B(n52107), .Z(n52113) );
  XOR U63167 ( .A(n52111), .B(n52113), .Z(n52099) );
  XOR U63168 ( .A(n52097), .B(n52099), .Z(n52101) );
  XOR U63169 ( .A(n52100), .B(n52101), .Z(n54225) );
  XOR U63170 ( .A(n54223), .B(n54225), .Z(n54234) );
  XOR U63171 ( .A(n50341), .B(n54234), .Z(n52090) );
  XOR U63172 ( .A(n50342), .B(n52090), .Z(n52088) );
  XOR U63173 ( .A(n50343), .B(n52088), .Z(n52086) );
  IV U63174 ( .A(n50344), .Z(n50346) );
  NOR U63175 ( .A(n50346), .B(n50345), .Z(n52085) );
  IV U63176 ( .A(n50347), .Z(n50349) );
  NOR U63177 ( .A(n50349), .B(n50348), .Z(n52083) );
  NOR U63178 ( .A(n52085), .B(n52083), .Z(n50350) );
  XOR U63179 ( .A(n52086), .B(n50350), .Z(n54238) );
  IV U63180 ( .A(n54238), .Z(n54236) );
  XOR U63181 ( .A(n54239), .B(n54236), .Z(n57579) );
  XOR U63182 ( .A(n57576), .B(n57579), .Z(n52078) );
  IV U63183 ( .A(n50351), .Z(n50352) );
  NOR U63184 ( .A(n50353), .B(n50352), .Z(n52080) );
  IV U63185 ( .A(n50354), .Z(n50355) );
  NOR U63186 ( .A(n50356), .B(n50355), .Z(n52077) );
  NOR U63187 ( .A(n52080), .B(n52077), .Z(n50357) );
  XOR U63188 ( .A(n52078), .B(n50357), .Z(n52072) );
  XOR U63189 ( .A(n52070), .B(n52072), .Z(n52074) );
  XOR U63190 ( .A(n52073), .B(n52074), .Z(n52068) );
  XOR U63191 ( .A(n52067), .B(n52068), .Z(n54245) );
  XOR U63192 ( .A(n52065), .B(n54245), .Z(n50366) );
  IV U63193 ( .A(n50358), .Z(n50360) );
  NOR U63194 ( .A(n50360), .B(n50359), .Z(n50367) );
  IV U63195 ( .A(n50367), .Z(n50361) );
  NOR U63196 ( .A(n50366), .B(n50361), .Z(n55410) );
  IV U63197 ( .A(n50362), .Z(n50363) );
  NOR U63198 ( .A(n50364), .B(n50363), .Z(n50365) );
  IV U63199 ( .A(n50365), .Z(n54246) );
  XOR U63200 ( .A(n54246), .B(n50366), .Z(n54248) );
  NOR U63201 ( .A(n50367), .B(n54248), .Z(n50368) );
  NOR U63202 ( .A(n55410), .B(n50368), .Z(n52061) );
  IV U63203 ( .A(n50369), .Z(n50370) );
  NOR U63204 ( .A(n50370), .B(n50381), .Z(n52062) );
  IV U63205 ( .A(n50371), .Z(n50376) );
  IV U63206 ( .A(n50372), .Z(n50373) );
  NOR U63207 ( .A(n50376), .B(n50373), .Z(n54252) );
  IV U63208 ( .A(n50374), .Z(n50375) );
  NOR U63209 ( .A(n50376), .B(n50375), .Z(n54247) );
  NOR U63210 ( .A(n54252), .B(n54247), .Z(n50377) );
  IV U63211 ( .A(n50377), .Z(n50378) );
  NOR U63212 ( .A(n52062), .B(n50378), .Z(n50379) );
  XOR U63213 ( .A(n52061), .B(n50379), .Z(n52060) );
  IV U63214 ( .A(n50380), .Z(n50382) );
  NOR U63215 ( .A(n50382), .B(n50381), .Z(n52058) );
  XOR U63216 ( .A(n52060), .B(n52058), .Z(n50383) );
  NOR U63217 ( .A(n50384), .B(n50383), .Z(n55402) );
  IV U63218 ( .A(n50385), .Z(n50386) );
  NOR U63219 ( .A(n50389), .B(n50386), .Z(n52052) );
  IV U63220 ( .A(n50387), .Z(n50388) );
  NOR U63221 ( .A(n50389), .B(n50388), .Z(n52050) );
  NOR U63222 ( .A(n52050), .B(n52058), .Z(n50390) );
  XOR U63223 ( .A(n52060), .B(n50390), .Z(n52053) );
  XOR U63224 ( .A(n52052), .B(n52053), .Z(n50391) );
  NOR U63225 ( .A(n50392), .B(n50391), .Z(n50393) );
  NOR U63226 ( .A(n55402), .B(n50393), .Z(n52039) );
  XOR U63227 ( .A(n50394), .B(n52039), .Z(n52038) );
  XOR U63228 ( .A(n52036), .B(n52038), .Z(n54259) );
  XOR U63229 ( .A(n54258), .B(n54259), .Z(n54263) );
  IV U63230 ( .A(n54263), .Z(n50402) );
  IV U63231 ( .A(n50395), .Z(n50396) );
  NOR U63232 ( .A(n50397), .B(n50396), .Z(n52034) );
  IV U63233 ( .A(n50398), .Z(n50399) );
  NOR U63234 ( .A(n50400), .B(n50399), .Z(n54262) );
  NOR U63235 ( .A(n52034), .B(n54262), .Z(n50401) );
  XOR U63236 ( .A(n50402), .B(n50401), .Z(n52033) );
  IV U63237 ( .A(n50403), .Z(n50405) );
  NOR U63238 ( .A(n50405), .B(n50404), .Z(n52031) );
  XOR U63239 ( .A(n52033), .B(n52031), .Z(n52026) );
  XOR U63240 ( .A(n52024), .B(n52026), .Z(n54272) );
  XOR U63241 ( .A(n50406), .B(n54272), .Z(n54276) );
  XOR U63242 ( .A(n54274), .B(n54276), .Z(n54280) );
  XOR U63243 ( .A(n54278), .B(n54280), .Z(n52020) );
  IV U63244 ( .A(n50407), .Z(n50409) );
  NOR U63245 ( .A(n50409), .B(n50408), .Z(n50410) );
  IV U63246 ( .A(n50410), .Z(n52019) );
  XOR U63247 ( .A(n52020), .B(n52019), .Z(n50411) );
  XOR U63248 ( .A(n50412), .B(n50411), .Z(n54292) );
  IV U63249 ( .A(n54292), .Z(n50424) );
  IV U63250 ( .A(n50413), .Z(n50414) );
  NOR U63251 ( .A(n50415), .B(n50414), .Z(n54284) );
  IV U63252 ( .A(n50416), .Z(n50417) );
  NOR U63253 ( .A(n50417), .B(n50419), .Z(n52017) );
  IV U63254 ( .A(n50418), .Z(n50420) );
  NOR U63255 ( .A(n50420), .B(n50419), .Z(n54290) );
  NOR U63256 ( .A(n52017), .B(n54290), .Z(n50421) );
  IV U63257 ( .A(n50421), .Z(n50422) );
  NOR U63258 ( .A(n54284), .B(n50422), .Z(n50423) );
  XOR U63259 ( .A(n50424), .B(n50423), .Z(n54288) );
  XOR U63260 ( .A(n54289), .B(n54288), .Z(n50435) );
  IV U63261 ( .A(n50425), .Z(n50426) );
  NOR U63262 ( .A(n50427), .B(n50426), .Z(n50432) );
  IV U63263 ( .A(n50428), .Z(n50429) );
  NOR U63264 ( .A(n50429), .B(n50442), .Z(n50434) );
  NOR U63265 ( .A(n50432), .B(n50434), .Z(n50430) );
  IV U63266 ( .A(n50430), .Z(n50431) );
  NOR U63267 ( .A(n50435), .B(n50431), .Z(n50439) );
  IV U63268 ( .A(n50432), .Z(n50433) );
  NOR U63269 ( .A(n50433), .B(n54288), .Z(n54296) );
  IV U63270 ( .A(n50434), .Z(n50437) );
  IV U63271 ( .A(n50435), .Z(n50436) );
  NOR U63272 ( .A(n50437), .B(n50436), .Z(n54304) );
  NOR U63273 ( .A(n54296), .B(n54304), .Z(n50438) );
  IV U63274 ( .A(n50438), .Z(n54300) );
  NOR U63275 ( .A(n50439), .B(n54300), .Z(n50445) );
  IV U63276 ( .A(n50445), .Z(n52015) );
  NOR U63277 ( .A(n50440), .B(n52015), .Z(n57644) );
  IV U63278 ( .A(n50441), .Z(n50443) );
  NOR U63279 ( .A(n50443), .B(n50442), .Z(n50444) );
  IV U63280 ( .A(n50444), .Z(n52016) );
  XOR U63281 ( .A(n52016), .B(n50445), .Z(n54313) );
  IV U63282 ( .A(n50446), .Z(n50447) );
  NOR U63283 ( .A(n50448), .B(n50447), .Z(n50449) );
  IV U63284 ( .A(n50449), .Z(n54312) );
  XOR U63285 ( .A(n54313), .B(n54312), .Z(n50450) );
  NOR U63286 ( .A(n50451), .B(n50450), .Z(n50452) );
  NOR U63287 ( .A(n57644), .B(n50452), .Z(n52007) );
  IV U63288 ( .A(n50453), .Z(n50455) );
  NOR U63289 ( .A(n50455), .B(n50454), .Z(n50456) );
  IV U63290 ( .A(n50456), .Z(n52008) );
  XOR U63291 ( .A(n52007), .B(n52008), .Z(n52011) );
  IV U63292 ( .A(n50457), .Z(n50458) );
  NOR U63293 ( .A(n50459), .B(n50458), .Z(n52010) );
  IV U63294 ( .A(n50460), .Z(n50461) );
  NOR U63295 ( .A(n50462), .B(n50461), .Z(n52004) );
  NOR U63296 ( .A(n52010), .B(n52004), .Z(n50463) );
  XOR U63297 ( .A(n52011), .B(n50463), .Z(n50464) );
  NOR U63298 ( .A(n50469), .B(n50464), .Z(n50472) );
  IV U63299 ( .A(n50465), .Z(n50467) );
  NOR U63300 ( .A(n50467), .B(n50466), .Z(n50474) );
  IV U63301 ( .A(n50474), .Z(n50468) );
  NOR U63302 ( .A(n50472), .B(n50468), .Z(n54317) );
  IV U63303 ( .A(n50469), .Z(n50471) );
  XOR U63304 ( .A(n52010), .B(n52011), .Z(n50470) );
  NOR U63305 ( .A(n50471), .B(n50470), .Z(n55333) );
  NOR U63306 ( .A(n50472), .B(n55333), .Z(n50473) );
  NOR U63307 ( .A(n50474), .B(n50473), .Z(n50475) );
  NOR U63308 ( .A(n54317), .B(n50475), .Z(n54318) );
  IV U63309 ( .A(n50476), .Z(n50477) );
  NOR U63310 ( .A(n50478), .B(n50477), .Z(n50479) );
  IV U63311 ( .A(n50479), .Z(n54319) );
  XOR U63312 ( .A(n54318), .B(n54319), .Z(n54322) );
  XOR U63313 ( .A(n50480), .B(n54322), .Z(n51999) );
  IV U63314 ( .A(n50481), .Z(n50482) );
  NOR U63315 ( .A(n50483), .B(n50482), .Z(n51998) );
  IV U63316 ( .A(n50484), .Z(n50486) );
  NOR U63317 ( .A(n50486), .B(n50485), .Z(n54325) );
  NOR U63318 ( .A(n51998), .B(n54325), .Z(n50487) );
  XOR U63319 ( .A(n51999), .B(n50487), .Z(n54336) );
  IV U63320 ( .A(n50488), .Z(n50491) );
  NOR U63321 ( .A(n54336), .B(n50491), .Z(n51995) );
  NOR U63322 ( .A(n50489), .B(n54335), .Z(n50490) );
  XOR U63323 ( .A(n50490), .B(n54336), .Z(n51997) );
  IV U63324 ( .A(n50492), .Z(n51996) );
  XOR U63325 ( .A(n51997), .B(n51996), .Z(n50494) );
  NOR U63326 ( .A(n50492), .B(n50491), .Z(n50493) );
  NOR U63327 ( .A(n50494), .B(n50493), .Z(n50495) );
  NOR U63328 ( .A(n51995), .B(n50495), .Z(n50503) );
  IV U63329 ( .A(n50503), .Z(n51993) );
  IV U63330 ( .A(n50496), .Z(n50498) );
  NOR U63331 ( .A(n50498), .B(n50497), .Z(n50504) );
  IV U63332 ( .A(n50504), .Z(n50499) );
  NOR U63333 ( .A(n51993), .B(n50499), .Z(n55293) );
  IV U63334 ( .A(n50500), .Z(n50502) );
  NOR U63335 ( .A(n50502), .B(n50501), .Z(n51991) );
  XOR U63336 ( .A(n50503), .B(n51991), .Z(n50508) );
  NOR U63337 ( .A(n50504), .B(n50508), .Z(n50505) );
  NOR U63338 ( .A(n55293), .B(n50505), .Z(n50506) );
  NOR U63339 ( .A(n50507), .B(n50506), .Z(n50511) );
  IV U63340 ( .A(n50507), .Z(n50510) );
  IV U63341 ( .A(n50508), .Z(n50509) );
  NOR U63342 ( .A(n50510), .B(n50509), .Z(n51990) );
  NOR U63343 ( .A(n50511), .B(n51990), .Z(n50515) );
  IV U63344 ( .A(n50515), .Z(n51985) );
  NOR U63345 ( .A(n50512), .B(n51985), .Z(n54350) );
  NOR U63346 ( .A(n51986), .B(n50513), .Z(n50514) );
  XOR U63347 ( .A(n50515), .B(n50514), .Z(n51979) );
  NOR U63348 ( .A(n50516), .B(n51979), .Z(n50517) );
  NOR U63349 ( .A(n54350), .B(n50517), .Z(n51970) );
  NOR U63350 ( .A(n50518), .B(n51981), .Z(n50522) );
  IV U63351 ( .A(n50519), .Z(n50520) );
  NOR U63352 ( .A(n50521), .B(n50520), .Z(n51971) );
  NOR U63353 ( .A(n50522), .B(n51971), .Z(n50523) );
  XOR U63354 ( .A(n51970), .B(n50523), .Z(n51976) );
  XOR U63355 ( .A(n51966), .B(n51976), .Z(n50524) );
  XOR U63356 ( .A(n50525), .B(n50524), .Z(n51960) );
  IV U63357 ( .A(n50526), .Z(n50528) );
  NOR U63358 ( .A(n50528), .B(n50527), .Z(n51963) );
  IV U63359 ( .A(n50529), .Z(n50531) );
  NOR U63360 ( .A(n50531), .B(n50530), .Z(n51961) );
  NOR U63361 ( .A(n51963), .B(n51961), .Z(n50532) );
  XOR U63362 ( .A(n51960), .B(n50532), .Z(n54354) );
  XOR U63363 ( .A(n50533), .B(n54354), .Z(n54364) );
  IV U63364 ( .A(n50534), .Z(n50535) );
  NOR U63365 ( .A(n50536), .B(n50535), .Z(n51958) );
  IV U63366 ( .A(n50537), .Z(n50539) );
  NOR U63367 ( .A(n50539), .B(n50538), .Z(n54363) );
  NOR U63368 ( .A(n51958), .B(n54363), .Z(n50540) );
  XOR U63369 ( .A(n54364), .B(n50540), .Z(n50541) );
  IV U63370 ( .A(n50541), .Z(n51956) );
  XOR U63371 ( .A(n51954), .B(n51956), .Z(n51952) );
  XOR U63372 ( .A(n51951), .B(n51952), .Z(n50547) );
  XOR U63373 ( .A(n50542), .B(n50547), .Z(n51945) );
  NOR U63374 ( .A(n50543), .B(n51945), .Z(n54381) );
  IV U63375 ( .A(n50544), .Z(n50546) );
  NOR U63376 ( .A(n50546), .B(n50545), .Z(n50550) );
  IV U63377 ( .A(n50550), .Z(n50548) );
  NOR U63378 ( .A(n50548), .B(n50547), .Z(n54380) );
  IV U63379 ( .A(n51945), .Z(n50549) );
  NOR U63380 ( .A(n50550), .B(n50549), .Z(n50551) );
  NOR U63381 ( .A(n54380), .B(n50551), .Z(n50552) );
  NOR U63382 ( .A(n50553), .B(n50552), .Z(n50554) );
  NOR U63383 ( .A(n54381), .B(n50554), .Z(n51941) );
  XOR U63384 ( .A(n50555), .B(n51941), .Z(n51935) );
  XOR U63385 ( .A(n51933), .B(n51935), .Z(n51936) );
  XOR U63386 ( .A(n51937), .B(n51936), .Z(n54384) );
  IV U63387 ( .A(n50562), .Z(n50556) );
  NOR U63388 ( .A(n50561), .B(n50556), .Z(n54383) );
  IV U63389 ( .A(n50557), .Z(n50558) );
  NOR U63390 ( .A(n50561), .B(n50558), .Z(n54386) );
  NOR U63391 ( .A(n54383), .B(n54386), .Z(n50559) );
  XOR U63392 ( .A(n54384), .B(n50559), .Z(n54392) );
  IV U63393 ( .A(n50560), .Z(n50564) );
  XOR U63394 ( .A(n50562), .B(n50561), .Z(n50563) );
  NOR U63395 ( .A(n50564), .B(n50563), .Z(n54390) );
  XOR U63396 ( .A(n54392), .B(n54390), .Z(n54394) );
  XOR U63397 ( .A(n54393), .B(n54394), .Z(n51931) );
  XOR U63398 ( .A(n50565), .B(n51931), .Z(n51923) );
  IV U63399 ( .A(n50566), .Z(n50575) );
  IV U63400 ( .A(n50567), .Z(n50568) );
  NOR U63401 ( .A(n50575), .B(n50568), .Z(n51922) );
  IV U63402 ( .A(n50569), .Z(n50571) );
  NOR U63403 ( .A(n50571), .B(n50570), .Z(n51925) );
  NOR U63404 ( .A(n51922), .B(n51925), .Z(n50572) );
  XOR U63405 ( .A(n51923), .B(n50572), .Z(n51921) );
  IV U63406 ( .A(n50573), .Z(n50574) );
  NOR U63407 ( .A(n50575), .B(n50574), .Z(n51919) );
  XOR U63408 ( .A(n51921), .B(n51919), .Z(n50576) );
  NOR U63409 ( .A(n50577), .B(n50576), .Z(n55211) );
  IV U63410 ( .A(n50578), .Z(n50579) );
  NOR U63411 ( .A(n50580), .B(n50579), .Z(n51917) );
  NOR U63412 ( .A(n51917), .B(n51919), .Z(n50581) );
  XOR U63413 ( .A(n51921), .B(n50581), .Z(n50586) );
  NOR U63414 ( .A(n50582), .B(n50586), .Z(n50583) );
  NOR U63415 ( .A(n55211), .B(n50583), .Z(n50584) );
  NOR U63416 ( .A(n50585), .B(n50584), .Z(n50589) );
  IV U63417 ( .A(n50585), .Z(n50588) );
  IV U63418 ( .A(n50586), .Z(n50587) );
  NOR U63419 ( .A(n50588), .B(n50587), .Z(n54411) );
  NOR U63420 ( .A(n50589), .B(n54411), .Z(n54405) );
  IV U63421 ( .A(n50590), .Z(n50591) );
  NOR U63422 ( .A(n50592), .B(n50591), .Z(n50593) );
  IV U63423 ( .A(n50593), .Z(n54407) );
  XOR U63424 ( .A(n54405), .B(n54407), .Z(n54415) );
  XOR U63425 ( .A(n50594), .B(n54415), .Z(n54420) );
  IV U63426 ( .A(n50595), .Z(n50596) );
  NOR U63427 ( .A(n50597), .B(n50596), .Z(n51913) );
  IV U63428 ( .A(n50598), .Z(n50599) );
  NOR U63429 ( .A(n50600), .B(n50599), .Z(n54419) );
  NOR U63430 ( .A(n51913), .B(n54419), .Z(n50601) );
  XOR U63431 ( .A(n54420), .B(n50601), .Z(n51907) );
  IV U63432 ( .A(n50602), .Z(n50603) );
  NOR U63433 ( .A(n50603), .B(n51898), .Z(n51903) );
  IV U63434 ( .A(n50604), .Z(n50605) );
  NOR U63435 ( .A(n50605), .B(n50607), .Z(n51908) );
  IV U63436 ( .A(n50606), .Z(n50608) );
  NOR U63437 ( .A(n50608), .B(n50607), .Z(n51906) );
  XOR U63438 ( .A(n51908), .B(n51906), .Z(n50609) );
  NOR U63439 ( .A(n51903), .B(n50609), .Z(n50610) );
  XOR U63440 ( .A(n51907), .B(n50610), .Z(n50611) );
  IV U63441 ( .A(n50611), .Z(n51895) );
  NOR U63442 ( .A(n51897), .B(n50612), .Z(n50613) );
  NOR U63443 ( .A(n50613), .B(n51898), .Z(n50614) );
  XOR U63444 ( .A(n51895), .B(n50614), .Z(n51892) );
  IV U63445 ( .A(n50615), .Z(n50616) );
  NOR U63446 ( .A(n50621), .B(n50616), .Z(n51890) );
  XOR U63447 ( .A(n51892), .B(n51890), .Z(n51886) );
  NOR U63448 ( .A(n50618), .B(n50617), .Z(n51885) );
  IV U63449 ( .A(n50619), .Z(n50620) );
  NOR U63450 ( .A(n50621), .B(n50620), .Z(n51888) );
  NOR U63451 ( .A(n51885), .B(n51888), .Z(n50622) );
  XOR U63452 ( .A(n51886), .B(n50622), .Z(n54428) );
  IV U63453 ( .A(n54428), .Z(n54431) );
  XOR U63454 ( .A(n54429), .B(n54431), .Z(n50623) );
  XOR U63455 ( .A(n50624), .B(n50623), .Z(n54438) );
  XOR U63456 ( .A(n54436), .B(n54438), .Z(n54439) );
  XOR U63457 ( .A(n54440), .B(n54439), .Z(n50625) );
  IV U63458 ( .A(n50625), .Z(n54444) );
  IV U63459 ( .A(n50626), .Z(n50628) );
  NOR U63460 ( .A(n50628), .B(n50627), .Z(n54442) );
  XOR U63461 ( .A(n54444), .B(n54442), .Z(n54447) );
  IV U63462 ( .A(n50629), .Z(n50631) );
  NOR U63463 ( .A(n50631), .B(n50630), .Z(n54445) );
  XOR U63464 ( .A(n54447), .B(n54445), .Z(n54450) );
  XOR U63465 ( .A(n54451), .B(n54450), .Z(n54452) );
  IV U63466 ( .A(n50632), .Z(n50634) );
  NOR U63467 ( .A(n50634), .B(n50633), .Z(n50639) );
  IV U63468 ( .A(n50635), .Z(n50636) );
  NOR U63469 ( .A(n50637), .B(n50636), .Z(n50638) );
  NOR U63470 ( .A(n50639), .B(n50638), .Z(n54454) );
  XOR U63471 ( .A(n54452), .B(n54454), .Z(n54458) );
  XOR U63472 ( .A(n54456), .B(n54458), .Z(n54461) );
  XOR U63473 ( .A(n54459), .B(n54461), .Z(n51880) );
  XOR U63474 ( .A(n51879), .B(n51880), .Z(n51873) );
  IV U63475 ( .A(n50640), .Z(n50642) );
  NOR U63476 ( .A(n50642), .B(n50641), .Z(n51871) );
  XOR U63477 ( .A(n51873), .B(n51871), .Z(n50643) );
  XOR U63478 ( .A(n50644), .B(n50643), .Z(n51862) );
  XOR U63479 ( .A(n51860), .B(n51862), .Z(n51859) );
  XOR U63480 ( .A(n50645), .B(n51859), .Z(n51853) );
  XOR U63481 ( .A(n51851), .B(n51853), .Z(n54479) );
  XOR U63482 ( .A(n51854), .B(n54479), .Z(n50646) );
  XOR U63483 ( .A(n50647), .B(n50646), .Z(n51850) );
  IV U63484 ( .A(n50658), .Z(n50648) );
  NOR U63485 ( .A(n50648), .B(n50657), .Z(n51848) );
  IV U63486 ( .A(n50649), .Z(n50650) );
  NOR U63487 ( .A(n50650), .B(n50657), .Z(n51845) );
  NOR U63488 ( .A(n51848), .B(n51845), .Z(n50651) );
  XOR U63489 ( .A(n51850), .B(n50651), .Z(n50652) );
  IV U63490 ( .A(n50652), .Z(n51844) );
  IV U63491 ( .A(n50653), .Z(n50656) );
  IV U63492 ( .A(n50654), .Z(n50655) );
  NOR U63493 ( .A(n50656), .B(n50655), .Z(n51842) );
  XOR U63494 ( .A(n51844), .B(n51842), .Z(n51838) );
  XOR U63495 ( .A(n50658), .B(n50657), .Z(n50661) );
  IV U63496 ( .A(n50659), .Z(n50660) );
  NOR U63497 ( .A(n50661), .B(n50660), .Z(n51836) );
  XOR U63498 ( .A(n51838), .B(n51836), .Z(n51840) );
  XOR U63499 ( .A(n51839), .B(n51840), .Z(n51834) );
  XOR U63500 ( .A(n51833), .B(n51834), .Z(n54488) );
  XOR U63501 ( .A(n54487), .B(n54488), .Z(n51831) );
  XOR U63502 ( .A(n51830), .B(n51831), .Z(n51827) );
  XOR U63503 ( .A(n51826), .B(n51827), .Z(n51822) );
  IV U63504 ( .A(n50662), .Z(n50663) );
  NOR U63505 ( .A(n50664), .B(n50663), .Z(n50665) );
  IV U63506 ( .A(n50665), .Z(n51820) );
  XOR U63507 ( .A(n51822), .B(n51820), .Z(n50666) );
  XOR U63508 ( .A(n50667), .B(n50666), .Z(n51819) );
  IV U63509 ( .A(n50668), .Z(n50672) );
  NOR U63510 ( .A(n50670), .B(n50669), .Z(n50671) );
  NOR U63511 ( .A(n50672), .B(n50671), .Z(n51817) );
  XOR U63512 ( .A(n51819), .B(n51817), .Z(n51812) );
  IV U63513 ( .A(n50673), .Z(n50676) );
  IV U63514 ( .A(n50674), .Z(n50675) );
  NOR U63515 ( .A(n50676), .B(n50675), .Z(n51810) );
  XOR U63516 ( .A(n51812), .B(n51810), .Z(n50677) );
  XOR U63517 ( .A(n50678), .B(n50677), .Z(n51803) );
  XOR U63518 ( .A(n51804), .B(n51803), .Z(n51799) );
  IV U63519 ( .A(n50679), .Z(n50680) );
  NOR U63520 ( .A(n50680), .B(n50682), .Z(n51805) );
  IV U63521 ( .A(n50681), .Z(n50687) );
  XOR U63522 ( .A(n50683), .B(n50682), .Z(n50684) );
  NOR U63523 ( .A(n50685), .B(n50684), .Z(n50686) );
  IV U63524 ( .A(n50686), .Z(n50690) );
  NOR U63525 ( .A(n50687), .B(n50690), .Z(n51800) );
  NOR U63526 ( .A(n51805), .B(n51800), .Z(n50688) );
  XOR U63527 ( .A(n51799), .B(n50688), .Z(n54500) );
  IV U63528 ( .A(n50689), .Z(n50691) );
  NOR U63529 ( .A(n50691), .B(n50690), .Z(n54498) );
  XOR U63530 ( .A(n54500), .B(n54498), .Z(n54503) );
  XOR U63531 ( .A(n54501), .B(n54503), .Z(n51797) );
  XOR U63532 ( .A(n51794), .B(n51797), .Z(n51792) );
  IV U63533 ( .A(n50692), .Z(n50694) );
  NOR U63534 ( .A(n50694), .B(n50693), .Z(n51789) );
  XOR U63535 ( .A(n51792), .B(n51789), .Z(n50695) );
  XOR U63536 ( .A(n50696), .B(n50695), .Z(n50704) );
  XOR U63537 ( .A(n54508), .B(n50704), .Z(n50697) );
  NOR U63538 ( .A(n50703), .B(n50697), .Z(n50698) );
  IV U63539 ( .A(n50698), .Z(n50702) );
  IV U63540 ( .A(n50699), .Z(n50700) );
  NOR U63541 ( .A(n50701), .B(n50700), .Z(n50706) );
  NOR U63542 ( .A(n50702), .B(n50706), .Z(n50711) );
  IV U63543 ( .A(n50703), .Z(n50705) );
  IV U63544 ( .A(n50704), .Z(n54510) );
  NOR U63545 ( .A(n50705), .B(n54510), .Z(n50710) );
  IV U63546 ( .A(n50706), .Z(n50708) );
  XOR U63547 ( .A(n54510), .B(n54508), .Z(n50707) );
  NOR U63548 ( .A(n50708), .B(n50707), .Z(n50709) );
  NOR U63549 ( .A(n50710), .B(n50709), .Z(n57978) );
  IV U63550 ( .A(n57978), .Z(n54511) );
  NOR U63551 ( .A(n50711), .B(n54511), .Z(n51784) );
  IV U63552 ( .A(n50712), .Z(n50713) );
  NOR U63553 ( .A(n50714), .B(n50713), .Z(n51783) );
  IV U63554 ( .A(n50715), .Z(n50717) );
  NOR U63555 ( .A(n50717), .B(n50716), .Z(n51786) );
  NOR U63556 ( .A(n51783), .B(n51786), .Z(n50718) );
  XOR U63557 ( .A(n51784), .B(n50718), .Z(n57924) );
  XOR U63558 ( .A(n50719), .B(n57924), .Z(n51775) );
  XOR U63559 ( .A(n51774), .B(n51775), .Z(n51778) );
  XOR U63560 ( .A(n51777), .B(n51778), .Z(n51772) );
  XOR U63561 ( .A(n51773), .B(n51772), .Z(n50720) );
  XOR U63562 ( .A(n50721), .B(n50720), .Z(n54521) );
  IV U63563 ( .A(n50722), .Z(n50724) );
  NOR U63564 ( .A(n50724), .B(n50723), .Z(n54519) );
  XOR U63565 ( .A(n54521), .B(n54519), .Z(n51765) );
  XOR U63566 ( .A(n51764), .B(n51765), .Z(n54526) );
  IV U63567 ( .A(n50725), .Z(n51759) );
  NOR U63568 ( .A(n51759), .B(n50726), .Z(n50729) );
  IV U63569 ( .A(n50727), .Z(n50728) );
  NOR U63570 ( .A(n50728), .B(n50735), .Z(n54524) );
  NOR U63571 ( .A(n50729), .B(n54524), .Z(n50730) );
  XOR U63572 ( .A(n54526), .B(n50730), .Z(n51751) );
  IV U63573 ( .A(n50731), .Z(n50740) );
  IV U63574 ( .A(n50732), .Z(n50733) );
  NOR U63575 ( .A(n50740), .B(n50733), .Z(n54542) );
  IV U63576 ( .A(n50734), .Z(n50736) );
  NOR U63577 ( .A(n50736), .B(n50735), .Z(n51752) );
  NOR U63578 ( .A(n54542), .B(n51752), .Z(n50737) );
  XOR U63579 ( .A(n51751), .B(n50737), .Z(n51749) );
  IV U63580 ( .A(n50738), .Z(n50739) );
  NOR U63581 ( .A(n50740), .B(n50739), .Z(n51748) );
  IV U63582 ( .A(n50741), .Z(n50743) );
  NOR U63583 ( .A(n50743), .B(n50742), .Z(n51745) );
  NOR U63584 ( .A(n51748), .B(n51745), .Z(n50744) );
  XOR U63585 ( .A(n51749), .B(n50744), .Z(n50745) );
  IV U63586 ( .A(n50745), .Z(n51744) );
  XOR U63587 ( .A(n51742), .B(n51744), .Z(n54568) );
  XOR U63588 ( .A(n54549), .B(n54568), .Z(n54552) );
  IV U63589 ( .A(n50746), .Z(n50750) );
  NOR U63590 ( .A(n50748), .B(n50747), .Z(n50749) );
  IV U63591 ( .A(n50749), .Z(n50752) );
  NOR U63592 ( .A(n50750), .B(n50752), .Z(n54567) );
  IV U63593 ( .A(n50751), .Z(n50753) );
  NOR U63594 ( .A(n50753), .B(n50752), .Z(n54551) );
  XOR U63595 ( .A(n54567), .B(n54551), .Z(n50754) );
  XOR U63596 ( .A(n54552), .B(n50754), .Z(n54576) );
  XOR U63597 ( .A(n54578), .B(n54576), .Z(n51741) );
  XOR U63598 ( .A(n50755), .B(n51741), .Z(n51737) );
  XOR U63599 ( .A(n51735), .B(n51737), .Z(n54586) );
  IV U63600 ( .A(n50756), .Z(n50757) );
  NOR U63601 ( .A(n50758), .B(n50757), .Z(n54584) );
  IV U63602 ( .A(n50759), .Z(n50762) );
  IV U63603 ( .A(n50760), .Z(n50761) );
  NOR U63604 ( .A(n50762), .B(n50761), .Z(n54585) );
  NOR U63605 ( .A(n54584), .B(n54585), .Z(n50763) );
  XOR U63606 ( .A(n54586), .B(n50763), .Z(n51723) );
  NOR U63607 ( .A(n50764), .B(n51729), .Z(n50768) );
  IV U63608 ( .A(n50765), .Z(n50767) );
  NOR U63609 ( .A(n50767), .B(n50766), .Z(n51724) );
  NOR U63610 ( .A(n50768), .B(n51724), .Z(n50769) );
  XOR U63611 ( .A(n51723), .B(n50769), .Z(n58057) );
  XOR U63612 ( .A(n58056), .B(n58057), .Z(n55152) );
  XOR U63613 ( .A(n55156), .B(n55152), .Z(n50770) );
  IV U63614 ( .A(n50770), .Z(n51715) );
  XOR U63615 ( .A(n51712), .B(n51715), .Z(n50771) );
  XOR U63616 ( .A(n50772), .B(n50771), .Z(n51708) );
  XOR U63617 ( .A(n51706), .B(n51708), .Z(n51710) );
  IV U63618 ( .A(n50773), .Z(n50776) );
  IV U63619 ( .A(n50774), .Z(n50775) );
  NOR U63620 ( .A(n50776), .B(n50775), .Z(n50777) );
  IV U63621 ( .A(n50777), .Z(n51709) );
  XOR U63622 ( .A(n51710), .B(n51709), .Z(n51701) );
  NOR U63623 ( .A(n50779), .B(n50778), .Z(n50780) );
  IV U63624 ( .A(n50780), .Z(n50787) );
  XOR U63625 ( .A(n50782), .B(n50781), .Z(n50784) );
  NOR U63626 ( .A(n50784), .B(n50783), .Z(n50785) );
  IV U63627 ( .A(n50785), .Z(n50786) );
  NOR U63628 ( .A(n50787), .B(n50786), .Z(n51700) );
  IV U63629 ( .A(n50788), .Z(n50791) );
  IV U63630 ( .A(n50789), .Z(n50790) );
  NOR U63631 ( .A(n50791), .B(n50790), .Z(n51703) );
  NOR U63632 ( .A(n51700), .B(n51703), .Z(n50792) );
  XOR U63633 ( .A(n51701), .B(n50792), .Z(n51699) );
  XOR U63634 ( .A(n51697), .B(n51699), .Z(n51694) );
  XOR U63635 ( .A(n50793), .B(n51694), .Z(n51690) );
  XOR U63636 ( .A(n50794), .B(n51690), .Z(n51678) );
  IV U63637 ( .A(n51678), .Z(n51680) );
  XOR U63638 ( .A(n51679), .B(n51680), .Z(n51676) );
  NOR U63639 ( .A(n50796), .B(n50795), .Z(n51675) );
  IV U63640 ( .A(n50797), .Z(n50799) );
  NOR U63641 ( .A(n50799), .B(n50798), .Z(n51682) );
  NOR U63642 ( .A(n51675), .B(n51682), .Z(n50800) );
  XOR U63643 ( .A(n51676), .B(n50800), .Z(n50801) );
  IV U63644 ( .A(n50801), .Z(n54596) );
  XOR U63645 ( .A(n50802), .B(n54596), .Z(n51669) );
  IV U63646 ( .A(n50803), .Z(n50804) );
  NOR U63647 ( .A(n50809), .B(n50804), .Z(n51667) );
  IV U63648 ( .A(n50805), .Z(n50806) );
  NOR U63649 ( .A(n50806), .B(n51670), .Z(n50807) );
  NOR U63650 ( .A(n51667), .B(n50807), .Z(n50814) );
  IV U63651 ( .A(n50808), .Z(n50813) );
  NOR U63652 ( .A(n50810), .B(n50809), .Z(n50811) );
  IV U63653 ( .A(n50811), .Z(n50812) );
  NOR U63654 ( .A(n50813), .B(n50812), .Z(n51665) );
  XOR U63655 ( .A(n50814), .B(n51665), .Z(n50815) );
  XOR U63656 ( .A(n51669), .B(n50815), .Z(n50816) );
  IV U63657 ( .A(n50816), .Z(n51647) );
  IV U63658 ( .A(n50819), .Z(n50817) );
  NOR U63659 ( .A(n50818), .B(n50817), .Z(n50823) );
  NOR U63660 ( .A(n50819), .B(n51642), .Z(n50820) );
  NOR U63661 ( .A(n50821), .B(n50820), .Z(n50822) );
  NOR U63662 ( .A(n50823), .B(n50822), .Z(n50824) );
  XOR U63663 ( .A(n51647), .B(n50824), .Z(n50828) );
  IV U63664 ( .A(n50825), .Z(n50826) );
  NOR U63665 ( .A(n51660), .B(n50826), .Z(n50827) );
  XOR U63666 ( .A(n50828), .B(n50827), .Z(n54622) );
  IV U63667 ( .A(n50829), .Z(n50833) );
  NOR U63668 ( .A(n50830), .B(n50839), .Z(n50831) );
  IV U63669 ( .A(n50831), .Z(n50832) );
  NOR U63670 ( .A(n50833), .B(n50832), .Z(n50844) );
  IV U63671 ( .A(n50844), .Z(n50834) );
  NOR U63672 ( .A(n54622), .B(n50834), .Z(n55106) );
  NOR U63673 ( .A(n50836), .B(n50835), .Z(n50843) );
  NOR U63674 ( .A(n50838), .B(n50837), .Z(n50840) );
  NOR U63675 ( .A(n50840), .B(n50839), .Z(n50841) );
  IV U63676 ( .A(n50841), .Z(n50842) );
  NOR U63677 ( .A(n50843), .B(n50842), .Z(n54620) );
  IV U63678 ( .A(n54622), .Z(n54626) );
  XOR U63679 ( .A(n54620), .B(n54626), .Z(n50847) );
  NOR U63680 ( .A(n50844), .B(n50847), .Z(n50845) );
  NOR U63681 ( .A(n55106), .B(n50845), .Z(n51637) );
  NOR U63682 ( .A(n50846), .B(n51637), .Z(n50850) );
  IV U63683 ( .A(n50846), .Z(n50849) );
  IV U63684 ( .A(n50847), .Z(n50848) );
  NOR U63685 ( .A(n50849), .B(n50848), .Z(n55112) );
  NOR U63686 ( .A(n50850), .B(n55112), .Z(n51633) );
  IV U63687 ( .A(n50851), .Z(n50853) );
  NOR U63688 ( .A(n50853), .B(n50852), .Z(n51638) );
  IV U63689 ( .A(n50854), .Z(n50855) );
  NOR U63690 ( .A(n50856), .B(n50855), .Z(n51634) );
  NOR U63691 ( .A(n51638), .B(n51634), .Z(n50857) );
  XOR U63692 ( .A(n51633), .B(n50857), .Z(n51632) );
  IV U63693 ( .A(n50858), .Z(n50859) );
  NOR U63694 ( .A(n50860), .B(n50859), .Z(n51629) );
  XOR U63695 ( .A(n51632), .B(n51629), .Z(n51627) );
  XOR U63696 ( .A(n50861), .B(n51627), .Z(n50866) );
  XOR U63697 ( .A(n50862), .B(n50866), .Z(n51617) );
  IV U63698 ( .A(n51617), .Z(n50863) );
  NOR U63699 ( .A(n50864), .B(n50863), .Z(n51621) );
  IV U63700 ( .A(n50864), .Z(n50865) );
  NOR U63701 ( .A(n50866), .B(n50865), .Z(n51618) );
  NOR U63702 ( .A(n51621), .B(n51618), .Z(n50874) );
  IV U63703 ( .A(n50867), .Z(n50869) );
  NOR U63704 ( .A(n50869), .B(n50868), .Z(n51619) );
  IV U63705 ( .A(n50870), .Z(n50872) );
  NOR U63706 ( .A(n50872), .B(n50871), .Z(n51615) );
  NOR U63707 ( .A(n51619), .B(n51615), .Z(n50873) );
  XOR U63708 ( .A(n50874), .B(n50873), .Z(n51612) );
  XOR U63709 ( .A(n50875), .B(n51612), .Z(n50876) );
  IV U63710 ( .A(n50876), .Z(n51606) );
  XOR U63711 ( .A(n51605), .B(n51606), .Z(n50877) );
  NOR U63712 ( .A(n50878), .B(n50877), .Z(n58155) );
  IV U63713 ( .A(n50879), .Z(n50881) );
  NOR U63714 ( .A(n50881), .B(n50880), .Z(n51603) );
  NOR U63715 ( .A(n51605), .B(n51603), .Z(n50882) );
  XOR U63716 ( .A(n50882), .B(n51606), .Z(n51599) );
  NOR U63717 ( .A(n50883), .B(n51599), .Z(n50884) );
  NOR U63718 ( .A(n58155), .B(n50884), .Z(n51596) );
  IV U63719 ( .A(n50885), .Z(n50886) );
  NOR U63720 ( .A(n50887), .B(n50886), .Z(n51595) );
  IV U63721 ( .A(n50888), .Z(n50891) );
  IV U63722 ( .A(n50889), .Z(n50890) );
  NOR U63723 ( .A(n50891), .B(n50890), .Z(n51600) );
  NOR U63724 ( .A(n51595), .B(n51600), .Z(n50892) );
  XOR U63725 ( .A(n51596), .B(n50892), .Z(n54633) );
  IV U63726 ( .A(n50893), .Z(n50894) );
  NOR U63727 ( .A(n50895), .B(n50894), .Z(n51593) );
  IV U63728 ( .A(n50896), .Z(n50897) );
  NOR U63729 ( .A(n50897), .B(n50903), .Z(n54631) );
  NOR U63730 ( .A(n51593), .B(n54631), .Z(n50898) );
  XOR U63731 ( .A(n54633), .B(n50898), .Z(n54634) );
  NOR U63732 ( .A(n50900), .B(n50899), .Z(n58167) );
  IV U63733 ( .A(n50901), .Z(n50902) );
  NOR U63734 ( .A(n50903), .B(n50902), .Z(n58176) );
  NOR U63735 ( .A(n58167), .B(n58176), .Z(n54635) );
  XOR U63736 ( .A(n54634), .B(n54635), .Z(n54639) );
  XOR U63737 ( .A(n54638), .B(n54639), .Z(n54649) );
  XOR U63738 ( .A(n50904), .B(n54649), .Z(n50905) );
  IV U63739 ( .A(n50905), .Z(n51590) );
  IV U63740 ( .A(n50906), .Z(n50910) );
  XOR U63741 ( .A(n50908), .B(n50907), .Z(n50909) );
  NOR U63742 ( .A(n50910), .B(n50909), .Z(n51588) );
  XOR U63743 ( .A(n51590), .B(n51588), .Z(n51584) );
  XOR U63744 ( .A(n51583), .B(n51584), .Z(n54658) );
  IV U63745 ( .A(n50911), .Z(n50913) );
  NOR U63746 ( .A(n50913), .B(n50912), .Z(n54656) );
  XOR U63747 ( .A(n54658), .B(n54656), .Z(n51582) );
  IV U63748 ( .A(n50914), .Z(n50915) );
  NOR U63749 ( .A(n50919), .B(n50915), .Z(n50916) );
  IV U63750 ( .A(n50916), .Z(n51581) );
  XOR U63751 ( .A(n51582), .B(n51581), .Z(n51575) );
  IV U63752 ( .A(n50917), .Z(n50918) );
  NOR U63753 ( .A(n50919), .B(n50918), .Z(n51578) );
  IV U63754 ( .A(n50920), .Z(n50922) );
  IV U63755 ( .A(n50921), .Z(n50925) );
  NOR U63756 ( .A(n50922), .B(n50925), .Z(n51576) );
  NOR U63757 ( .A(n51578), .B(n51576), .Z(n50923) );
  XOR U63758 ( .A(n51575), .B(n50923), .Z(n51574) );
  IV U63759 ( .A(n50924), .Z(n50926) );
  NOR U63760 ( .A(n50926), .B(n50925), .Z(n51572) );
  XOR U63761 ( .A(n51574), .B(n51572), .Z(n50927) );
  NOR U63762 ( .A(n50928), .B(n50927), .Z(n51571) );
  IV U63763 ( .A(n50929), .Z(n50930) );
  NOR U63764 ( .A(n50931), .B(n50930), .Z(n51573) );
  NOR U63765 ( .A(n51573), .B(n51572), .Z(n50932) );
  XOR U63766 ( .A(n51574), .B(n50932), .Z(n50937) );
  NOR U63767 ( .A(n50933), .B(n50937), .Z(n50934) );
  NOR U63768 ( .A(n51571), .B(n50934), .Z(n50935) );
  NOR U63769 ( .A(n50936), .B(n50935), .Z(n50940) );
  IV U63770 ( .A(n50936), .Z(n50939) );
  IV U63771 ( .A(n50937), .Z(n50938) );
  NOR U63772 ( .A(n50939), .B(n50938), .Z(n55074) );
  NOR U63773 ( .A(n50940), .B(n55074), .Z(n51567) );
  XOR U63774 ( .A(n54667), .B(n51567), .Z(n51570) );
  XOR U63775 ( .A(n51568), .B(n51570), .Z(n50941) );
  XOR U63776 ( .A(n51569), .B(n50941), .Z(n51565) );
  IV U63777 ( .A(n50942), .Z(n50943) );
  NOR U63778 ( .A(n50944), .B(n50943), .Z(n51564) );
  IV U63779 ( .A(n50945), .Z(n50947) );
  NOR U63780 ( .A(n50947), .B(n50946), .Z(n51562) );
  NOR U63781 ( .A(n51564), .B(n51562), .Z(n50948) );
  XOR U63782 ( .A(n51565), .B(n50948), .Z(n50956) );
  IV U63783 ( .A(n50956), .Z(n50949) );
  NOR U63784 ( .A(n50950), .B(n50949), .Z(n51561) );
  IV U63785 ( .A(n50951), .Z(n50953) );
  NOR U63786 ( .A(n50953), .B(n50952), .Z(n50957) );
  IV U63787 ( .A(n50957), .Z(n50955) );
  XOR U63788 ( .A(n51564), .B(n51565), .Z(n50954) );
  NOR U63789 ( .A(n50955), .B(n50954), .Z(n58226) );
  NOR U63790 ( .A(n50957), .B(n50956), .Z(n50958) );
  NOR U63791 ( .A(n58226), .B(n50958), .Z(n51558) );
  NOR U63792 ( .A(n50959), .B(n51558), .Z(n50960) );
  NOR U63793 ( .A(n51561), .B(n50960), .Z(n50968) );
  IV U63794 ( .A(n50961), .Z(n50962) );
  NOR U63795 ( .A(n50963), .B(n50962), .Z(n51557) );
  IV U63796 ( .A(n50964), .Z(n50966) );
  NOR U63797 ( .A(n50966), .B(n50965), .Z(n54670) );
  NOR U63798 ( .A(n51557), .B(n54670), .Z(n50967) );
  XOR U63799 ( .A(n50968), .B(n50967), .Z(n54675) );
  XOR U63800 ( .A(n54673), .B(n54675), .Z(n54681) );
  XOR U63801 ( .A(n51555), .B(n54681), .Z(n50969) );
  XOR U63802 ( .A(n50970), .B(n50969), .Z(n54689) );
  XOR U63803 ( .A(n54687), .B(n54689), .Z(n54692) );
  IV U63804 ( .A(n50971), .Z(n50973) );
  NOR U63805 ( .A(n50973), .B(n50972), .Z(n50974) );
  IV U63806 ( .A(n50974), .Z(n54691) );
  XOR U63807 ( .A(n54692), .B(n54691), .Z(n54694) );
  NOR U63808 ( .A(n50976), .B(n50975), .Z(n54693) );
  NOR U63809 ( .A(n54697), .B(n54693), .Z(n50977) );
  XOR U63810 ( .A(n54694), .B(n50977), .Z(n54704) );
  IV U63811 ( .A(n50978), .Z(n50980) );
  NOR U63812 ( .A(n50980), .B(n50979), .Z(n54702) );
  XOR U63813 ( .A(n54704), .B(n54702), .Z(n51554) );
  XOR U63814 ( .A(n51552), .B(n51554), .Z(n54708) );
  IV U63815 ( .A(n50981), .Z(n50983) );
  NOR U63816 ( .A(n50983), .B(n50982), .Z(n50984) );
  IV U63817 ( .A(n50984), .Z(n50991) );
  NOR U63818 ( .A(n54708), .B(n50991), .Z(n58270) );
  IV U63819 ( .A(n50985), .Z(n50986) );
  NOR U63820 ( .A(n50989), .B(n50986), .Z(n54710) );
  IV U63821 ( .A(n50987), .Z(n50988) );
  NOR U63822 ( .A(n50989), .B(n50988), .Z(n50990) );
  IV U63823 ( .A(n50990), .Z(n54709) );
  XOR U63824 ( .A(n54709), .B(n54708), .Z(n54711) );
  XOR U63825 ( .A(n54710), .B(n54711), .Z(n50993) );
  NOR U63826 ( .A(n54711), .B(n50991), .Z(n50992) );
  NOR U63827 ( .A(n50993), .B(n50992), .Z(n50994) );
  NOR U63828 ( .A(n58270), .B(n50994), .Z(n51001) );
  IV U63829 ( .A(n51001), .Z(n54716) );
  NOR U63830 ( .A(n50995), .B(n54716), .Z(n58313) );
  NOR U63831 ( .A(n50997), .B(n50996), .Z(n50998) );
  IV U63832 ( .A(n50998), .Z(n50999) );
  NOR U63833 ( .A(n51000), .B(n50999), .Z(n54715) );
  XOR U63834 ( .A(n54715), .B(n51001), .Z(n51006) );
  NOR U63835 ( .A(n51002), .B(n51006), .Z(n51003) );
  NOR U63836 ( .A(n58313), .B(n51003), .Z(n51004) );
  NOR U63837 ( .A(n51005), .B(n51004), .Z(n51008) );
  IV U63838 ( .A(n51005), .Z(n51007) );
  IV U63839 ( .A(n51006), .Z(n54724) );
  NOR U63840 ( .A(n51007), .B(n54724), .Z(n58310) );
  NOR U63841 ( .A(n51008), .B(n58310), .Z(n54719) );
  IV U63842 ( .A(n51009), .Z(n51011) );
  NOR U63843 ( .A(n51011), .B(n51010), .Z(n51012) );
  IV U63844 ( .A(n51012), .Z(n54720) );
  XOR U63845 ( .A(n54719), .B(n54720), .Z(n54727) );
  XOR U63846 ( .A(n51013), .B(n54727), .Z(n54731) );
  XOR U63847 ( .A(n51549), .B(n54731), .Z(n51022) );
  IV U63848 ( .A(n51014), .Z(n51017) );
  IV U63849 ( .A(n51015), .Z(n51016) );
  NOR U63850 ( .A(n51017), .B(n51016), .Z(n54729) );
  IV U63851 ( .A(n51018), .Z(n51019) );
  NOR U63852 ( .A(n51020), .B(n51019), .Z(n51550) );
  NOR U63853 ( .A(n54729), .B(n51550), .Z(n51021) );
  XOR U63854 ( .A(n51022), .B(n51021), .Z(n51548) );
  XOR U63855 ( .A(n51544), .B(n51548), .Z(n51023) );
  XOR U63856 ( .A(n51024), .B(n51023), .Z(n54744) );
  IV U63857 ( .A(n54744), .Z(n51542) );
  XOR U63858 ( .A(n51025), .B(n51542), .Z(n54754) );
  IV U63859 ( .A(n51026), .Z(n51029) );
  IV U63860 ( .A(n51027), .Z(n51028) );
  NOR U63861 ( .A(n51029), .B(n51028), .Z(n54752) );
  XOR U63862 ( .A(n54754), .B(n54752), .Z(n51533) );
  XOR U63863 ( .A(n51534), .B(n51533), .Z(n51527) );
  IV U63864 ( .A(n51030), .Z(n51031) );
  NOR U63865 ( .A(n51032), .B(n51031), .Z(n51529) );
  IV U63866 ( .A(n51033), .Z(n51034) );
  NOR U63867 ( .A(n51037), .B(n51034), .Z(n51526) );
  NOR U63868 ( .A(n51529), .B(n51526), .Z(n51035) );
  XOR U63869 ( .A(n51527), .B(n51035), .Z(n54761) );
  IV U63870 ( .A(n51036), .Z(n51038) );
  NOR U63871 ( .A(n51038), .B(n51037), .Z(n54759) );
  XOR U63872 ( .A(n54761), .B(n54759), .Z(n54764) );
  XOR U63873 ( .A(n54762), .B(n54764), .Z(n51039) );
  NOR U63874 ( .A(n51040), .B(n51039), .Z(n58363) );
  IV U63875 ( .A(n51041), .Z(n51043) );
  NOR U63876 ( .A(n51043), .B(n51042), .Z(n51524) );
  NOR U63877 ( .A(n51524), .B(n54762), .Z(n51044) );
  XOR U63878 ( .A(n54764), .B(n51044), .Z(n51045) );
  NOR U63879 ( .A(n51046), .B(n51045), .Z(n51047) );
  NOR U63880 ( .A(n58363), .B(n51047), .Z(n51048) );
  IV U63881 ( .A(n51048), .Z(n54770) );
  XOR U63882 ( .A(n51521), .B(n54770), .Z(n51519) );
  XOR U63883 ( .A(n51049), .B(n51519), .Z(n51517) );
  XOR U63884 ( .A(n51515), .B(n51517), .Z(n54774) );
  XOR U63885 ( .A(n51512), .B(n54774), .Z(n51050) );
  XOR U63886 ( .A(n51051), .B(n51050), .Z(n54786) );
  IV U63887 ( .A(n51052), .Z(n51054) );
  NOR U63888 ( .A(n51054), .B(n51053), .Z(n54784) );
  IV U63889 ( .A(n51055), .Z(n51057) );
  NOR U63890 ( .A(n51057), .B(n51056), .Z(n51509) );
  NOR U63891 ( .A(n54784), .B(n51509), .Z(n51058) );
  XOR U63892 ( .A(n54786), .B(n51058), .Z(n51505) );
  XOR U63893 ( .A(n51504), .B(n51505), .Z(n51059) );
  NOR U63894 ( .A(n51060), .B(n51059), .Z(n51063) );
  IV U63895 ( .A(n51060), .Z(n51062) );
  XOR U63896 ( .A(n54784), .B(n54786), .Z(n51061) );
  NOR U63897 ( .A(n51062), .B(n51061), .Z(n58355) );
  NOR U63898 ( .A(n51063), .B(n58355), .Z(n54799) );
  XOR U63899 ( .A(n51064), .B(n54799), .Z(n51065) );
  XOR U63900 ( .A(n54800), .B(n51065), .Z(n51501) );
  IV U63901 ( .A(n51066), .Z(n51068) );
  NOR U63902 ( .A(n51068), .B(n51067), .Z(n51072) );
  NOR U63903 ( .A(n51070), .B(n51069), .Z(n51071) );
  NOR U63904 ( .A(n51072), .B(n51071), .Z(n51503) );
  XOR U63905 ( .A(n51501), .B(n51503), .Z(n51494) );
  XOR U63906 ( .A(n51493), .B(n51494), .Z(n51497) );
  XOR U63907 ( .A(n51496), .B(n51497), .Z(n51491) );
  XOR U63908 ( .A(n51490), .B(n51491), .Z(n51482) );
  XOR U63909 ( .A(n51484), .B(n51482), .Z(n51479) );
  XOR U63910 ( .A(n51073), .B(n51479), .Z(n51079) );
  XOR U63911 ( .A(n51074), .B(n51079), .Z(n51082) );
  NOR U63912 ( .A(n51075), .B(n51082), .Z(n51472) );
  IV U63913 ( .A(n51076), .Z(n51077) );
  NOR U63914 ( .A(n51078), .B(n51077), .Z(n51084) );
  IV U63915 ( .A(n51084), .Z(n51081) );
  IV U63916 ( .A(n51079), .Z(n51477) );
  XOR U63917 ( .A(n51475), .B(n51477), .Z(n51080) );
  NOR U63918 ( .A(n51081), .B(n51080), .Z(n54976) );
  IV U63919 ( .A(n51082), .Z(n51083) );
  NOR U63920 ( .A(n51084), .B(n51083), .Z(n51085) );
  NOR U63921 ( .A(n54976), .B(n51085), .Z(n54814) );
  NOR U63922 ( .A(n51086), .B(n54814), .Z(n51087) );
  NOR U63923 ( .A(n51472), .B(n51087), .Z(n51088) );
  IV U63924 ( .A(n51088), .Z(n54819) );
  IV U63925 ( .A(n51089), .Z(n51090) );
  NOR U63926 ( .A(n51091), .B(n51090), .Z(n51469) );
  XOR U63927 ( .A(n54819), .B(n51469), .Z(n51092) );
  XOR U63928 ( .A(n51093), .B(n51092), .Z(n54830) );
  XOR U63929 ( .A(n51094), .B(n54830), .Z(n51460) );
  XOR U63930 ( .A(n51458), .B(n51460), .Z(n51461) );
  XOR U63931 ( .A(n51462), .B(n51461), .Z(n51448) );
  IV U63932 ( .A(n51095), .Z(n51449) );
  NOR U63933 ( .A(n51096), .B(n51449), .Z(n51100) );
  IV U63934 ( .A(n51097), .Z(n51098) );
  NOR U63935 ( .A(n51099), .B(n51098), .Z(n51455) );
  NOR U63936 ( .A(n51100), .B(n51455), .Z(n51101) );
  XOR U63937 ( .A(n51448), .B(n51101), .Z(n51441) );
  NOR U63938 ( .A(n51102), .B(n51440), .Z(n51105) );
  IV U63939 ( .A(n51103), .Z(n51104) );
  NOR U63940 ( .A(n51104), .B(n51111), .Z(n51437) );
  NOR U63941 ( .A(n51105), .B(n51437), .Z(n51106) );
  XOR U63942 ( .A(n51441), .B(n51106), .Z(n51429) );
  IV U63943 ( .A(n51107), .Z(n51109) );
  NOR U63944 ( .A(n51109), .B(n51108), .Z(n51118) );
  IV U63945 ( .A(n51118), .Z(n51431) );
  NOR U63946 ( .A(n51429), .B(n51431), .Z(n51120) );
  IV U63947 ( .A(n51110), .Z(n51112) );
  NOR U63948 ( .A(n51112), .B(n51111), .Z(n51114) );
  IV U63949 ( .A(n51114), .Z(n51113) );
  NOR U63950 ( .A(n51441), .B(n51113), .Z(n58422) );
  NOR U63951 ( .A(n51429), .B(n51114), .Z(n51115) );
  NOR U63952 ( .A(n58422), .B(n51115), .Z(n51116) );
  IV U63953 ( .A(n51116), .Z(n51117) );
  NOR U63954 ( .A(n51118), .B(n51117), .Z(n51119) );
  NOR U63955 ( .A(n51120), .B(n51119), .Z(n51434) );
  NOR U63956 ( .A(n51121), .B(n51434), .Z(n51426) );
  IV U63957 ( .A(n51122), .Z(n51127) );
  IV U63958 ( .A(n51123), .Z(n51124) );
  NOR U63959 ( .A(n51127), .B(n51124), .Z(n51432) );
  XOR U63960 ( .A(n51434), .B(n51432), .Z(n51428) );
  IV U63961 ( .A(n51125), .Z(n51126) );
  NOR U63962 ( .A(n51127), .B(n51126), .Z(n51128) );
  IV U63963 ( .A(n51128), .Z(n51427) );
  XOR U63964 ( .A(n51428), .B(n51427), .Z(n51133) );
  NOR U63965 ( .A(n51129), .B(n51133), .Z(n51130) );
  NOR U63966 ( .A(n51426), .B(n51130), .Z(n51131) );
  NOR U63967 ( .A(n51132), .B(n51131), .Z(n51425) );
  IV U63968 ( .A(n51132), .Z(n51135) );
  IV U63969 ( .A(n51133), .Z(n51134) );
  NOR U63970 ( .A(n51135), .B(n51134), .Z(n58467) );
  NOR U63971 ( .A(n51425), .B(n58467), .Z(n58473) );
  IV U63972 ( .A(n51136), .Z(n51137) );
  NOR U63973 ( .A(n51138), .B(n51137), .Z(n51422) );
  IV U63974 ( .A(n51139), .Z(n51141) );
  NOR U63975 ( .A(n51141), .B(n51140), .Z(n51421) );
  NOR U63976 ( .A(n51422), .B(n51421), .Z(n58474) );
  XOR U63977 ( .A(n58473), .B(n58474), .Z(n51419) );
  XOR U63978 ( .A(n51417), .B(n51419), .Z(n51410) );
  XOR U63979 ( .A(n51142), .B(n51410), .Z(n51404) );
  XOR U63980 ( .A(n51143), .B(n51404), .Z(n51392) );
  XOR U63981 ( .A(n51144), .B(n51392), .Z(n51396) );
  XOR U63982 ( .A(n51395), .B(n51396), .Z(n51391) );
  XOR U63983 ( .A(n51145), .B(n51391), .Z(n51153) );
  IV U63984 ( .A(n51146), .Z(n51148) );
  NOR U63985 ( .A(n51148), .B(n51147), .Z(n51385) );
  IV U63986 ( .A(n51149), .Z(n51151) );
  NOR U63987 ( .A(n51151), .B(n51150), .Z(n51383) );
  NOR U63988 ( .A(n51385), .B(n51383), .Z(n51152) );
  XOR U63989 ( .A(n51153), .B(n51152), .Z(n54843) );
  IV U63990 ( .A(n51154), .Z(n51155) );
  NOR U63991 ( .A(n51155), .B(n51164), .Z(n51161) );
  IV U63992 ( .A(n51161), .Z(n51156) );
  NOR U63993 ( .A(n54843), .B(n51156), .Z(n54953) );
  IV U63994 ( .A(n51157), .Z(n51158) );
  NOR U63995 ( .A(n51159), .B(n51158), .Z(n54841) );
  NOR U63996 ( .A(n54839), .B(n54841), .Z(n51160) );
  XOR U63997 ( .A(n51160), .B(n54843), .Z(n54847) );
  NOR U63998 ( .A(n51161), .B(n54847), .Z(n51162) );
  NOR U63999 ( .A(n54953), .B(n51162), .Z(n51167) );
  IV U64000 ( .A(n51163), .Z(n51165) );
  NOR U64001 ( .A(n51165), .B(n51164), .Z(n51381) );
  NOR U64002 ( .A(n51381), .B(n54846), .Z(n51166) );
  XOR U64003 ( .A(n51167), .B(n51166), .Z(n51380) );
  IV U64004 ( .A(n51168), .Z(n51170) );
  NOR U64005 ( .A(n51170), .B(n51169), .Z(n51171) );
  IV U64006 ( .A(n51171), .Z(n51172) );
  NOR U64007 ( .A(n51173), .B(n51172), .Z(n51376) );
  XOR U64008 ( .A(n51380), .B(n51376), .Z(n51174) );
  XOR U64009 ( .A(n51175), .B(n51174), .Z(n51367) );
  XOR U64010 ( .A(n51368), .B(n51367), .Z(n54855) );
  IV U64011 ( .A(n51176), .Z(n51178) );
  NOR U64012 ( .A(n51178), .B(n51177), .Z(n54854) );
  IV U64013 ( .A(n51179), .Z(n51180) );
  NOR U64014 ( .A(n51181), .B(n51180), .Z(n51370) );
  NOR U64015 ( .A(n54854), .B(n51370), .Z(n51182) );
  XOR U64016 ( .A(n54855), .B(n51182), .Z(n51363) );
  IV U64017 ( .A(n51183), .Z(n51184) );
  NOR U64018 ( .A(n51184), .B(n51186), .Z(n51364) );
  IV U64019 ( .A(n51185), .Z(n51187) );
  NOR U64020 ( .A(n51187), .B(n51186), .Z(n54851) );
  NOR U64021 ( .A(n51364), .B(n54851), .Z(n51188) );
  XOR U64022 ( .A(n51363), .B(n51188), .Z(n51361) );
  IV U64023 ( .A(n51189), .Z(n51192) );
  IV U64024 ( .A(n51190), .Z(n51191) );
  NOR U64025 ( .A(n51192), .B(n51191), .Z(n51358) );
  NOR U64026 ( .A(n51360), .B(n51358), .Z(n51193) );
  XOR U64027 ( .A(n51361), .B(n51193), .Z(n51194) );
  IV U64028 ( .A(n51194), .Z(n51357) );
  IV U64029 ( .A(n51195), .Z(n51198) );
  IV U64030 ( .A(n51196), .Z(n51197) );
  NOR U64031 ( .A(n51198), .B(n51197), .Z(n51355) );
  XOR U64032 ( .A(n51357), .B(n51355), .Z(n54863) );
  XOR U64033 ( .A(n54861), .B(n54863), .Z(n51354) );
  XOR U64034 ( .A(n51352), .B(n51354), .Z(n54870) );
  XOR U64035 ( .A(n54868), .B(n54870), .Z(n54875) );
  XOR U64036 ( .A(n54874), .B(n54875), .Z(n51199) );
  NOR U64037 ( .A(n51200), .B(n51199), .Z(n54877) );
  IV U64038 ( .A(n51201), .Z(n51203) );
  NOR U64039 ( .A(n51203), .B(n51202), .Z(n54871) );
  NOR U64040 ( .A(n54874), .B(n54871), .Z(n51204) );
  XOR U64041 ( .A(n51204), .B(n54875), .Z(n51266) );
  NOR U64042 ( .A(n51205), .B(n51266), .Z(n51206) );
  NOR U64043 ( .A(n54877), .B(n51206), .Z(n51264) );
  NOR U64044 ( .A(n51208), .B(n51207), .Z(n51209) );
  XOR U64045 ( .A(n51210), .B(n51209), .Z(n51211) );
  NOR U64046 ( .A(n51212), .B(n51211), .Z(n51213) );
  NOR U64047 ( .A(n51213), .B(n51251), .Z(n51277) );
  IV U64048 ( .A(n51277), .Z(n51250) );
  XOR U64049 ( .A(n51215), .B(n51214), .Z(n51327) );
  IV U64050 ( .A(n51216), .Z(n51220) );
  NOR U64051 ( .A(n51218), .B(n51217), .Z(n51219) );
  XOR U64052 ( .A(n51220), .B(n51219), .Z(n51247) );
  IV U64053 ( .A(n51221), .Z(n51228) );
  XOR U64054 ( .A(n51223), .B(n51222), .Z(n51233) );
  IV U64055 ( .A(n51224), .Z(n51226) );
  NOR U64056 ( .A(n51226), .B(n51225), .Z(n51235) );
  IV U64057 ( .A(n51235), .Z(n51232) );
  NOR U64058 ( .A(n51233), .B(n51232), .Z(n51304) );
  IV U64059 ( .A(n51304), .Z(n51227) );
  NOR U64060 ( .A(n51228), .B(n51227), .Z(n51306) );
  XOR U64061 ( .A(n51247), .B(n51306), .Z(n51338) );
  NOR U64062 ( .A(n51327), .B(n51338), .Z(n51229) );
  IV U64063 ( .A(n51229), .Z(n51230) );
  NOR U64064 ( .A(n51299), .B(n51230), .Z(n51231) );
  IV U64065 ( .A(n51231), .Z(n51283) );
  XOR U64066 ( .A(n51233), .B(n51232), .Z(n51237) );
  NOR U64067 ( .A(n51235), .B(n51234), .Z(n51236) );
  NOR U64068 ( .A(n51237), .B(n51236), .Z(n51238) );
  NOR U64069 ( .A(n51302), .B(n51238), .Z(n51239) );
  IV U64070 ( .A(n51239), .Z(n51311) );
  IV U64071 ( .A(n51240), .Z(n51242) );
  NOR U64072 ( .A(n51242), .B(n51241), .Z(n51310) );
  IV U64073 ( .A(n51310), .Z(n51243) );
  NOR U64074 ( .A(n51311), .B(n51243), .Z(n51298) );
  IV U64075 ( .A(n51298), .Z(n51244) );
  NOR U64076 ( .A(n51283), .B(n51244), .Z(n51274) );
  IV U64077 ( .A(n51274), .Z(n51245) );
  NOR U64078 ( .A(n51250), .B(n51245), .Z(n51288) );
  IV U64079 ( .A(n51288), .Z(n51259) );
  IV U64080 ( .A(n51306), .Z(n51246) );
  NOR U64081 ( .A(n51247), .B(n51246), .Z(n51331) );
  IV U64082 ( .A(n51331), .Z(n51248) );
  NOR U64083 ( .A(n51327), .B(n51248), .Z(n51275) );
  IV U64084 ( .A(n51275), .Z(n51249) );
  NOR U64085 ( .A(n51250), .B(n51249), .Z(n51260) );
  NOR U64086 ( .A(n51251), .B(n51260), .Z(n51252) );
  XOR U64087 ( .A(n51262), .B(n51252), .Z(n51345) );
  IV U64088 ( .A(n51345), .Z(n51290) );
  NOR U64089 ( .A(n51254), .B(n51253), .Z(n51255) );
  IV U64090 ( .A(n51255), .Z(n51257) );
  XOR U64091 ( .A(n51257), .B(n51256), .Z(n51294) );
  NOR U64092 ( .A(n51290), .B(n51294), .Z(n51258) );
  IV U64093 ( .A(n51258), .Z(n51285) );
  NOR U64094 ( .A(n51259), .B(n51285), .Z(n51271) );
  IV U64095 ( .A(n51271), .Z(n54879) );
  NOR U64096 ( .A(n51264), .B(n54879), .Z(n51273) );
  IV U64097 ( .A(n51260), .Z(n51261) );
  NOR U64098 ( .A(n51262), .B(n51261), .Z(n51292) );
  IV U64099 ( .A(n51292), .Z(n51263) );
  NOR U64100 ( .A(n51263), .B(n51294), .Z(n51265) );
  NOR U64101 ( .A(n51265), .B(n51264), .Z(n51269) );
  IV U64102 ( .A(n51265), .Z(n51268) );
  IV U64103 ( .A(n51266), .Z(n51267) );
  NOR U64104 ( .A(n51268), .B(n51267), .Z(n58578) );
  NOR U64105 ( .A(n51269), .B(n58578), .Z(n51270) );
  IV U64106 ( .A(n51270), .Z(n54880) );
  NOR U64107 ( .A(n51271), .B(n54880), .Z(n51272) );
  NOR U64108 ( .A(n51273), .B(n51272), .Z(n51349) );
  NOR U64109 ( .A(n51275), .B(n51274), .Z(n51276) );
  XOR U64110 ( .A(n51277), .B(n51276), .Z(n51296) );
  IV U64111 ( .A(n51278), .Z(n51280) );
  NOR U64112 ( .A(n51280), .B(n51279), .Z(n51318) );
  IV U64113 ( .A(n51318), .Z(n51281) );
  NOR U64114 ( .A(n51311), .B(n51281), .Z(n51297) );
  IV U64115 ( .A(n51297), .Z(n51282) );
  NOR U64116 ( .A(n51283), .B(n51282), .Z(n51295) );
  IV U64117 ( .A(n51295), .Z(n51284) );
  NOR U64118 ( .A(n51296), .B(n51284), .Z(n51289) );
  IV U64119 ( .A(n51289), .Z(n51286) );
  NOR U64120 ( .A(n51286), .B(n51285), .Z(n51350) );
  IV U64121 ( .A(n51350), .Z(n51287) );
  NOR U64122 ( .A(n51349), .B(n51287), .Z(n54946) );
  NOR U64123 ( .A(n51289), .B(n51288), .Z(n51346) );
  NOR U64124 ( .A(n51346), .B(n51290), .Z(n51291) );
  XOR U64125 ( .A(n51292), .B(n51291), .Z(n51293) );
  XOR U64126 ( .A(n51294), .B(n51293), .Z(n54884) );
  XOR U64127 ( .A(n51296), .B(n51295), .Z(n54886) );
  NOR U64128 ( .A(n51298), .B(n51297), .Z(n51300) );
  NOR U64129 ( .A(n51300), .B(n51299), .Z(n51328) );
  IV U64130 ( .A(n51300), .Z(n51308) );
  XOR U64131 ( .A(n51302), .B(n51301), .Z(n51303) );
  NOR U64132 ( .A(n51304), .B(n51303), .Z(n51305) );
  NOR U64133 ( .A(n51306), .B(n51305), .Z(n51307) );
  NOR U64134 ( .A(n51308), .B(n51307), .Z(n51309) );
  NOR U64135 ( .A(n51328), .B(n51309), .Z(n51334) );
  XOR U64136 ( .A(n51311), .B(n51310), .Z(n51320) );
  IV U64137 ( .A(n51312), .Z(n51314) );
  NOR U64138 ( .A(n51314), .B(n51313), .Z(n51317) );
  IV U64139 ( .A(n51317), .Z(n51315) );
  NOR U64140 ( .A(n51320), .B(n51315), .Z(n51316) );
  IV U64141 ( .A(n51316), .Z(n51335) );
  XOR U64142 ( .A(n51334), .B(n51335), .Z(n54891) );
  NOR U64143 ( .A(n51318), .B(n51317), .Z(n51319) );
  XOR U64144 ( .A(n51320), .B(n51319), .Z(n54927) );
  IV U64145 ( .A(n54927), .Z(n54897) );
  IV U64146 ( .A(n51321), .Z(n51323) );
  NOR U64147 ( .A(n51323), .B(n51322), .Z(n54925) );
  IV U64148 ( .A(n54925), .Z(n51324) );
  NOR U64149 ( .A(n54897), .B(n51324), .Z(n54892) );
  IV U64150 ( .A(n54892), .Z(n51325) );
  NOR U64151 ( .A(n54891), .B(n51325), .Z(n54918) );
  IV U64152 ( .A(n54918), .Z(n51326) );
  XOR U64153 ( .A(n51328), .B(n51338), .Z(n54916) );
  NOR U64154 ( .A(n51326), .B(n54916), .Z(n54901) );
  IV U64155 ( .A(n54901), .Z(n51339) );
  IV U64156 ( .A(n51327), .Z(n51333) );
  IV U64157 ( .A(n51328), .Z(n51329) );
  NOR U64158 ( .A(n51338), .B(n51329), .Z(n51330) );
  NOR U64159 ( .A(n51331), .B(n51330), .Z(n51332) );
  XOR U64160 ( .A(n51333), .B(n51332), .Z(n51343) );
  IV U64161 ( .A(n51334), .Z(n51336) );
  NOR U64162 ( .A(n51336), .B(n51335), .Z(n54921) );
  IV U64163 ( .A(n54921), .Z(n51337) );
  NOR U64164 ( .A(n51338), .B(n51337), .Z(n51341) );
  XOR U64165 ( .A(n51343), .B(n51341), .Z(n54900) );
  NOR U64166 ( .A(n51339), .B(n54900), .Z(n54887) );
  IV U64167 ( .A(n54887), .Z(n51340) );
  NOR U64168 ( .A(n54886), .B(n51340), .Z(n54912) );
  IV U64169 ( .A(n51341), .Z(n51342) );
  NOR U64170 ( .A(n51343), .B(n51342), .Z(n54888) );
  IV U64171 ( .A(n54888), .Z(n51344) );
  NOR U64172 ( .A(n54886), .B(n51344), .Z(n54905) );
  NOR U64173 ( .A(n54912), .B(n54905), .Z(n51347) );
  XOR U64174 ( .A(n51346), .B(n51345), .Z(n54904) );
  NOR U64175 ( .A(n51347), .B(n54904), .Z(n54885) );
  IV U64176 ( .A(n54885), .Z(n51348) );
  NOR U64177 ( .A(n54884), .B(n51348), .Z(n54909) );
  IV U64178 ( .A(n54909), .Z(n51351) );
  XOR U64179 ( .A(n51350), .B(n51349), .Z(n54908) );
  NOR U64180 ( .A(n51351), .B(n54908), .Z(n58601) );
  NOR U64181 ( .A(n54946), .B(n58601), .Z(n54882) );
  IV U64182 ( .A(n51352), .Z(n51353) );
  NOR U64183 ( .A(n51354), .B(n51353), .Z(n54866) );
  IV U64184 ( .A(n54866), .Z(n54860) );
  IV U64185 ( .A(n51355), .Z(n51356) );
  NOR U64186 ( .A(n51357), .B(n51356), .Z(n54865) );
  IV U64187 ( .A(n51358), .Z(n51359) );
  NOR U64188 ( .A(n51359), .B(n51361), .Z(n58565) );
  IV U64189 ( .A(n51360), .Z(n51362) );
  NOR U64190 ( .A(n51362), .B(n51361), .Z(n58535) );
  IV U64191 ( .A(n51363), .Z(n54852) );
  IV U64192 ( .A(n51364), .Z(n51365) );
  NOR U64193 ( .A(n54852), .B(n51365), .Z(n58538) );
  NOR U64194 ( .A(n51366), .B(n51367), .Z(n51373) );
  IV U64195 ( .A(n51367), .Z(n51369) );
  NOR U64196 ( .A(n51369), .B(n51368), .Z(n51371) );
  NOR U64197 ( .A(n51371), .B(n51370), .Z(n51372) );
  NOR U64198 ( .A(n51373), .B(n51372), .Z(n58555) );
  IV U64199 ( .A(n51374), .Z(n51375) );
  NOR U64200 ( .A(n51380), .B(n51375), .Z(n58558) );
  IV U64201 ( .A(n58558), .Z(n58556) );
  IV U64202 ( .A(n51376), .Z(n51377) );
  NOR U64203 ( .A(n51380), .B(n51377), .Z(n58546) );
  IV U64204 ( .A(n51378), .Z(n51379) );
  NOR U64205 ( .A(n51380), .B(n51379), .Z(n58543) );
  IV U64206 ( .A(n51381), .Z(n51382) );
  NOR U64207 ( .A(n54843), .B(n51382), .Z(n58525) );
  IV U64208 ( .A(n58525), .Z(n58524) );
  IV U64209 ( .A(n51383), .Z(n51384) );
  XOR U64210 ( .A(n51390), .B(n51391), .Z(n51386) );
  NOR U64211 ( .A(n51384), .B(n51386), .Z(n58512) );
  IV U64212 ( .A(n58512), .Z(n58516) );
  IV U64213 ( .A(n51385), .Z(n51387) );
  NOR U64214 ( .A(n51387), .B(n51386), .Z(n51388) );
  IV U64215 ( .A(n51388), .Z(n58515) );
  IV U64216 ( .A(n51392), .Z(n51402) );
  IV U64217 ( .A(n51393), .Z(n51394) );
  NOR U64218 ( .A(n51402), .B(n51394), .Z(n51399) );
  IV U64219 ( .A(n51395), .Z(n51397) );
  NOR U64220 ( .A(n51397), .B(n51396), .Z(n51398) );
  NOR U64221 ( .A(n51399), .B(n51398), .Z(n58488) );
  IV U64222 ( .A(n51400), .Z(n51401) );
  NOR U64223 ( .A(n51402), .B(n51401), .Z(n58485) );
  IV U64224 ( .A(n51403), .Z(n51405) );
  NOR U64225 ( .A(n51405), .B(n51404), .Z(n58490) );
  IV U64226 ( .A(n51406), .Z(n51407) );
  NOR U64227 ( .A(n51407), .B(n51410), .Z(n51408) );
  IV U64228 ( .A(n51408), .Z(n58501) );
  IV U64229 ( .A(n51409), .Z(n51413) );
  NOR U64230 ( .A(n51411), .B(n51410), .Z(n51412) );
  IV U64231 ( .A(n51412), .Z(n51415) );
  NOR U64232 ( .A(n51413), .B(n51415), .Z(n58502) );
  IV U64233 ( .A(n58502), .Z(n58500) );
  IV U64234 ( .A(n51414), .Z(n51416) );
  NOR U64235 ( .A(n51416), .B(n51415), .Z(n58458) );
  IV U64236 ( .A(n51417), .Z(n51418) );
  NOR U64237 ( .A(n51419), .B(n51418), .Z(n51420) );
  IV U64238 ( .A(n51420), .Z(n58462) );
  XOR U64239 ( .A(n51422), .B(n51421), .Z(n51423) );
  NOR U64240 ( .A(n58467), .B(n51423), .Z(n51424) );
  NOR U64241 ( .A(n51425), .B(n51424), .Z(n54836) );
  IV U64242 ( .A(n51426), .Z(n58466) );
  NOR U64243 ( .A(n51428), .B(n51427), .Z(n58442) );
  IV U64244 ( .A(n51429), .Z(n51430) );
  NOR U64245 ( .A(n51431), .B(n51430), .Z(n51436) );
  IV U64246 ( .A(n51432), .Z(n51433) );
  NOR U64247 ( .A(n51434), .B(n51433), .Z(n51435) );
  NOR U64248 ( .A(n51436), .B(n51435), .Z(n58440) );
  IV U64249 ( .A(n58440), .Z(n54834) );
  IV U64250 ( .A(n51437), .Z(n51438) );
  NOR U64251 ( .A(n51441), .B(n51438), .Z(n58428) );
  IV U64252 ( .A(n51439), .Z(n51443) );
  NOR U64253 ( .A(n51441), .B(n51440), .Z(n51442) );
  IV U64254 ( .A(n51442), .Z(n51445) );
  NOR U64255 ( .A(n51443), .B(n51445), .Z(n54961) );
  IV U64256 ( .A(n51444), .Z(n51446) );
  NOR U64257 ( .A(n51446), .B(n51445), .Z(n54958) );
  IV U64258 ( .A(n51447), .Z(n51451) );
  IV U64259 ( .A(n51448), .Z(n51457) );
  NOR U64260 ( .A(n51449), .B(n51457), .Z(n51450) );
  IV U64261 ( .A(n51450), .Z(n51453) );
  NOR U64262 ( .A(n51451), .B(n51453), .Z(n58449) );
  IV U64263 ( .A(n51452), .Z(n51454) );
  NOR U64264 ( .A(n51454), .B(n51453), .Z(n55001) );
  IV U64265 ( .A(n51455), .Z(n51456) );
  NOR U64266 ( .A(n51457), .B(n51456), .Z(n54998) );
  IV U64267 ( .A(n51458), .Z(n51459) );
  NOR U64268 ( .A(n51460), .B(n51459), .Z(n51464) );
  NOR U64269 ( .A(n51462), .B(n51461), .Z(n51463) );
  NOR U64270 ( .A(n51464), .B(n51463), .Z(n58447) );
  IV U64271 ( .A(n51465), .Z(n51468) );
  NOR U64272 ( .A(n54830), .B(n51466), .Z(n51467) );
  IV U64273 ( .A(n51467), .Z(n54824) );
  NOR U64274 ( .A(n51468), .B(n54824), .Z(n58425) );
  IV U64275 ( .A(n51469), .Z(n51470) );
  NOR U64276 ( .A(n54819), .B(n51470), .Z(n51471) );
  NOR U64277 ( .A(n51472), .B(n51471), .Z(n54966) );
  IV U64278 ( .A(n51473), .Z(n51474) );
  NOR U64279 ( .A(n51477), .B(n51474), .Z(n54973) );
  IV U64280 ( .A(n51475), .Z(n51476) );
  NOR U64281 ( .A(n51477), .B(n51476), .Z(n54983) );
  IV U64282 ( .A(n51478), .Z(n51480) );
  NOR U64283 ( .A(n51480), .B(n51479), .Z(n54988) );
  IV U64284 ( .A(n51484), .Z(n51481) );
  NOR U64285 ( .A(n51481), .B(n51482), .Z(n51489) );
  IV U64286 ( .A(n51482), .Z(n51483) );
  NOR U64287 ( .A(n51484), .B(n51483), .Z(n51487) );
  IV U64288 ( .A(n51485), .Z(n51486) );
  NOR U64289 ( .A(n51487), .B(n51486), .Z(n51488) );
  NOR U64290 ( .A(n51489), .B(n51488), .Z(n54986) );
  IV U64291 ( .A(n51490), .Z(n51492) );
  NOR U64292 ( .A(n51492), .B(n51491), .Z(n54968) );
  IV U64293 ( .A(n51493), .Z(n51495) );
  NOR U64294 ( .A(n51495), .B(n51494), .Z(n51500) );
  IV U64295 ( .A(n51496), .Z(n51498) );
  NOR U64296 ( .A(n51498), .B(n51497), .Z(n51499) );
  NOR U64297 ( .A(n51500), .B(n51499), .Z(n58389) );
  IV U64298 ( .A(n58389), .Z(n54811) );
  IV U64299 ( .A(n51501), .Z(n51502) );
  NOR U64300 ( .A(n51503), .B(n51502), .Z(n58391) );
  IV U64301 ( .A(n51504), .Z(n51507) );
  IV U64302 ( .A(n51505), .Z(n51506) );
  NOR U64303 ( .A(n51507), .B(n51506), .Z(n51508) );
  IV U64304 ( .A(n51508), .Z(n55019) );
  IV U64305 ( .A(n51509), .Z(n51510) );
  NOR U64306 ( .A(n54786), .B(n51510), .Z(n51511) );
  IV U64307 ( .A(n51511), .Z(n58360) );
  NOR U64308 ( .A(n51512), .B(n54774), .Z(n54792) );
  IV U64309 ( .A(n51513), .Z(n51514) );
  NOR U64310 ( .A(n51514), .B(n54774), .Z(n55028) );
  IV U64311 ( .A(n51515), .Z(n51516) );
  NOR U64312 ( .A(n51517), .B(n51516), .Z(n55029) );
  IV U64313 ( .A(n55029), .Z(n54771) );
  IV U64314 ( .A(n51518), .Z(n51520) );
  NOR U64315 ( .A(n51520), .B(n51519), .Z(n58375) );
  IV U64316 ( .A(n51521), .Z(n51522) );
  NOR U64317 ( .A(n51522), .B(n54770), .Z(n58378) );
  NOR U64318 ( .A(n58363), .B(n58378), .Z(n51523) );
  IV U64319 ( .A(n51523), .Z(n54767) );
  IV U64320 ( .A(n51524), .Z(n51525) );
  NOR U64321 ( .A(n51525), .B(n54764), .Z(n58335) );
  IV U64322 ( .A(n51526), .Z(n51528) );
  IV U64323 ( .A(n51527), .Z(n51530) );
  NOR U64324 ( .A(n51528), .B(n51530), .Z(n58371) );
  IV U64325 ( .A(n51529), .Z(n51531) );
  NOR U64326 ( .A(n51531), .B(n51530), .Z(n51532) );
  IV U64327 ( .A(n51532), .Z(n58324) );
  NOR U64328 ( .A(n51534), .B(n51533), .Z(n54757) );
  IV U64329 ( .A(n54757), .Z(n54751) );
  IV U64330 ( .A(n51535), .Z(n51536) );
  NOR U64331 ( .A(n51536), .B(n54744), .Z(n58346) );
  IV U64332 ( .A(n51537), .Z(n51538) );
  NOR U64333 ( .A(n51539), .B(n51538), .Z(n51540) );
  IV U64334 ( .A(n51540), .Z(n51541) );
  NOR U64335 ( .A(n51542), .B(n51541), .Z(n51543) );
  IV U64336 ( .A(n51543), .Z(n55038) );
  IV U64337 ( .A(n51544), .Z(n51545) );
  NOR U64338 ( .A(n51548), .B(n51545), .Z(n58296) );
  IV U64339 ( .A(n51546), .Z(n51547) );
  NOR U64340 ( .A(n51548), .B(n51547), .Z(n55040) );
  NOR U64341 ( .A(n58296), .B(n55040), .Z(n54741) );
  NOR U64342 ( .A(n54731), .B(n51549), .Z(n54738) );
  IV U64343 ( .A(n51550), .Z(n51551) );
  NOR U64344 ( .A(n54731), .B(n51551), .Z(n54735) );
  IV U64345 ( .A(n51552), .Z(n51553) );
  NOR U64346 ( .A(n51554), .B(n51553), .Z(n54706) );
  IV U64347 ( .A(n54706), .Z(n54701) );
  IV U64348 ( .A(n51555), .Z(n51556) );
  NOR U64349 ( .A(n51556), .B(n54681), .Z(n54686) );
  IV U64350 ( .A(n54686), .Z(n54683) );
  IV U64351 ( .A(n51557), .Z(n51559) );
  IV U64352 ( .A(n51558), .Z(n54671) );
  NOR U64353 ( .A(n51559), .B(n54671), .Z(n51560) );
  NOR U64354 ( .A(n51561), .B(n51560), .Z(n58249) );
  IV U64355 ( .A(n51562), .Z(n51563) );
  NOR U64356 ( .A(n51563), .B(n51565), .Z(n58223) );
  IV U64357 ( .A(n51564), .Z(n51566) );
  NOR U64358 ( .A(n51566), .B(n51565), .Z(n58251) );
  IV U64359 ( .A(n51567), .Z(n54666) );
  NOR U64360 ( .A(n51568), .B(n54666), .Z(n58218) );
  NOR U64361 ( .A(n51570), .B(n51569), .Z(n58215) );
  IV U64362 ( .A(n51571), .Z(n55073) );
  IV U64363 ( .A(n58196), .Z(n54665) );
  IV U64364 ( .A(n51575), .Z(n51580) );
  IV U64365 ( .A(n51576), .Z(n51577) );
  NOR U64366 ( .A(n51580), .B(n51577), .Z(n58198) );
  IV U64367 ( .A(n51578), .Z(n51579) );
  NOR U64368 ( .A(n51580), .B(n51579), .Z(n58201) );
  NOR U64369 ( .A(n51582), .B(n51581), .Z(n54662) );
  IV U64370 ( .A(n54662), .Z(n54655) );
  IV U64371 ( .A(n51583), .Z(n51585) );
  NOR U64372 ( .A(n51585), .B(n51584), .Z(n54660) );
  IV U64373 ( .A(n51586), .Z(n51587) );
  NOR U64374 ( .A(n51587), .B(n54649), .Z(n51592) );
  IV U64375 ( .A(n51588), .Z(n51589) );
  NOR U64376 ( .A(n51590), .B(n51589), .Z(n51591) );
  NOR U64377 ( .A(n51592), .B(n51591), .Z(n55080) );
  IV U64378 ( .A(n51593), .Z(n51594) );
  NOR U64379 ( .A(n54633), .B(n51594), .Z(n58170) );
  IV U64380 ( .A(n51595), .Z(n51598) );
  IV U64381 ( .A(n51596), .Z(n51597) );
  NOR U64382 ( .A(n51598), .B(n51597), .Z(n58164) );
  IV U64383 ( .A(n51599), .Z(n51602) );
  IV U64384 ( .A(n51600), .Z(n51601) );
  NOR U64385 ( .A(n51602), .B(n51601), .Z(n58152) );
  IV U64386 ( .A(n51603), .Z(n51604) );
  NOR U64387 ( .A(n51604), .B(n51606), .Z(n58147) );
  IV U64388 ( .A(n51605), .Z(n51607) );
  NOR U64389 ( .A(n51607), .B(n51606), .Z(n58144) );
  IV U64390 ( .A(n51608), .Z(n51609) );
  NOR U64391 ( .A(n51612), .B(n51609), .Z(n58133) );
  IV U64392 ( .A(n51610), .Z(n51611) );
  NOR U64393 ( .A(n51612), .B(n51611), .Z(n58134) );
  XOR U64394 ( .A(n58133), .B(n58134), .Z(n51613) );
  NOR U64395 ( .A(n58144), .B(n51613), .Z(n51614) );
  IV U64396 ( .A(n51614), .Z(n54630) );
  IV U64397 ( .A(n51615), .Z(n51616) );
  NOR U64398 ( .A(n51617), .B(n51616), .Z(n55089) );
  NOR U64399 ( .A(n51619), .B(n51618), .Z(n51620) );
  NOR U64400 ( .A(n51621), .B(n51620), .Z(n58137) );
  NOR U64401 ( .A(n51623), .B(n51622), .Z(n51624) );
  IV U64402 ( .A(n51624), .Z(n51625) );
  NOR U64403 ( .A(n51625), .B(n51627), .Z(n58121) );
  IV U64404 ( .A(n51626), .Z(n51628) );
  NOR U64405 ( .A(n51628), .B(n51627), .Z(n58124) );
  NOR U64406 ( .A(n51630), .B(n51629), .Z(n51631) );
  NOR U64407 ( .A(n51632), .B(n51631), .Z(n58113) );
  IV U64408 ( .A(n51633), .Z(n51636) );
  IV U64409 ( .A(n51634), .Z(n51635) );
  NOR U64410 ( .A(n51636), .B(n51635), .Z(n58116) );
  IV U64411 ( .A(n51637), .Z(n51640) );
  IV U64412 ( .A(n51638), .Z(n51639) );
  NOR U64413 ( .A(n51640), .B(n51639), .Z(n55103) );
  IV U64414 ( .A(n51641), .Z(n51644) );
  NOR U64415 ( .A(n51647), .B(n51642), .Z(n51643) );
  IV U64416 ( .A(n51643), .Z(n54617) );
  NOR U64417 ( .A(n51644), .B(n54617), .Z(n55097) );
  IV U64418 ( .A(n55097), .Z(n55095) );
  IV U64419 ( .A(n51645), .Z(n51646) );
  NOR U64420 ( .A(n51647), .B(n51646), .Z(n51648) );
  IV U64421 ( .A(n51648), .Z(n51664) );
  NOR U64422 ( .A(n51650), .B(n51649), .Z(n51651) );
  IV U64423 ( .A(n51651), .Z(n51658) );
  XOR U64424 ( .A(n51653), .B(n51652), .Z(n51654) );
  NOR U64425 ( .A(n51655), .B(n51654), .Z(n51656) );
  IV U64426 ( .A(n51656), .Z(n51657) );
  NOR U64427 ( .A(n51658), .B(n51657), .Z(n51659) );
  IV U64428 ( .A(n51659), .Z(n51661) );
  NOR U64429 ( .A(n51661), .B(n51660), .Z(n51662) );
  IV U64430 ( .A(n51662), .Z(n51663) );
  NOR U64431 ( .A(n51664), .B(n51663), .Z(n58088) );
  IV U64432 ( .A(n51665), .Z(n51666) );
  NOR U64433 ( .A(n51669), .B(n51666), .Z(n58085) );
  IV U64434 ( .A(n51667), .Z(n51668) );
  NOR U64435 ( .A(n51669), .B(n51668), .Z(n58102) );
  NOR U64436 ( .A(n51671), .B(n51670), .Z(n51672) );
  IV U64437 ( .A(n51672), .Z(n51673) );
  NOR U64438 ( .A(n54596), .B(n51673), .Z(n58101) );
  NOR U64439 ( .A(n58102), .B(n58101), .Z(n51674) );
  IV U64440 ( .A(n51674), .Z(n54615) );
  IV U64441 ( .A(n51675), .Z(n51677) );
  NOR U64442 ( .A(n51677), .B(n51676), .Z(n54600) );
  NOR U64443 ( .A(n51679), .B(n51678), .Z(n51685) );
  IV U64444 ( .A(n51679), .Z(n51681) );
  NOR U64445 ( .A(n51681), .B(n51680), .Z(n51683) );
  NOR U64446 ( .A(n51683), .B(n51682), .Z(n51684) );
  NOR U64447 ( .A(n51685), .B(n51684), .Z(n55124) );
  IV U64448 ( .A(n51686), .Z(n51687) );
  NOR U64449 ( .A(n51690), .B(n51687), .Z(n55128) );
  IV U64450 ( .A(n51688), .Z(n51689) );
  NOR U64451 ( .A(n51690), .B(n51689), .Z(n51691) );
  IV U64452 ( .A(n51691), .Z(n55129) );
  IV U64453 ( .A(n51692), .Z(n51693) );
  NOR U64454 ( .A(n51694), .B(n51693), .Z(n58067) );
  IV U64455 ( .A(n51695), .Z(n51696) );
  NOR U64456 ( .A(n51699), .B(n51696), .Z(n58073) );
  IV U64457 ( .A(n51697), .Z(n51698) );
  NOR U64458 ( .A(n51699), .B(n51698), .Z(n58029) );
  IV U64459 ( .A(n51700), .Z(n51702) );
  IV U64460 ( .A(n51701), .Z(n51705) );
  NOR U64461 ( .A(n51702), .B(n51705), .Z(n58032) );
  IV U64462 ( .A(n51703), .Z(n51704) );
  NOR U64463 ( .A(n51705), .B(n51704), .Z(n58070) );
  IV U64464 ( .A(n51706), .Z(n51707) );
  NOR U64465 ( .A(n51708), .B(n51707), .Z(n58045) );
  NOR U64466 ( .A(n51710), .B(n51709), .Z(n58026) );
  NOR U64467 ( .A(n58045), .B(n58026), .Z(n51711) );
  IV U64468 ( .A(n51711), .Z(n54590) );
  IV U64469 ( .A(n51712), .Z(n51713) );
  NOR U64470 ( .A(n51713), .B(n51715), .Z(n58042) );
  IV U64471 ( .A(n51714), .Z(n51716) );
  NOR U64472 ( .A(n51716), .B(n51715), .Z(n58021) );
  IV U64473 ( .A(n51717), .Z(n51718) );
  NOR U64474 ( .A(n51718), .B(n55152), .Z(n58018) );
  IV U64475 ( .A(n51719), .Z(n51720) );
  NOR U64476 ( .A(n51720), .B(n55152), .Z(n54589) );
  NOR U64477 ( .A(n51721), .B(n58056), .Z(n51722) );
  NOR U64478 ( .A(n51722), .B(n58057), .Z(n54587) );
  IV U64479 ( .A(n51723), .Z(n51726) );
  IV U64480 ( .A(n51724), .Z(n51725) );
  NOR U64481 ( .A(n51726), .B(n51725), .Z(n58053) );
  IV U64482 ( .A(n51727), .Z(n51731) );
  XOR U64483 ( .A(n54585), .B(n54586), .Z(n51728) );
  NOR U64484 ( .A(n51729), .B(n51728), .Z(n51730) );
  IV U64485 ( .A(n51730), .Z(n51733) );
  NOR U64486 ( .A(n51731), .B(n51733), .Z(n55147) );
  IV U64487 ( .A(n51732), .Z(n51734) );
  NOR U64488 ( .A(n51734), .B(n51733), .Z(n55141) );
  IV U64489 ( .A(n51735), .Z(n51736) );
  NOR U64490 ( .A(n51737), .B(n51736), .Z(n51738) );
  IV U64491 ( .A(n51738), .Z(n55161) );
  IV U64492 ( .A(n51739), .Z(n51740) );
  NOR U64493 ( .A(n51741), .B(n51740), .Z(n55157) );
  IV U64494 ( .A(n51742), .Z(n51743) );
  NOR U64495 ( .A(n51744), .B(n51743), .Z(n54560) );
  IV U64496 ( .A(n54560), .Z(n57972) );
  IV U64497 ( .A(n51745), .Z(n51746) );
  NOR U64498 ( .A(n51746), .B(n51749), .Z(n51747) );
  IV U64499 ( .A(n51747), .Z(n57975) );
  IV U64500 ( .A(n51748), .Z(n51750) );
  NOR U64501 ( .A(n51750), .B(n51749), .Z(n54547) );
  IV U64502 ( .A(n54547), .Z(n54541) );
  IV U64503 ( .A(n51751), .Z(n54544) );
  IV U64504 ( .A(n51752), .Z(n51753) );
  NOR U64505 ( .A(n54544), .B(n51753), .Z(n57996) );
  IV U64506 ( .A(n51754), .Z(n51757) );
  NOR U64507 ( .A(n51759), .B(n54526), .Z(n51755) );
  IV U64508 ( .A(n51755), .Z(n51756) );
  NOR U64509 ( .A(n51757), .B(n51756), .Z(n54528) );
  IV U64510 ( .A(n51758), .Z(n51762) );
  NOR U64511 ( .A(n51759), .B(n51765), .Z(n51760) );
  IV U64512 ( .A(n51760), .Z(n51761) );
  NOR U64513 ( .A(n51762), .B(n51761), .Z(n51763) );
  IV U64514 ( .A(n51763), .Z(n57941) );
  IV U64515 ( .A(n51764), .Z(n51766) );
  NOR U64516 ( .A(n51766), .B(n51765), .Z(n51767) );
  IV U64517 ( .A(n51767), .Z(n57944) );
  IV U64518 ( .A(n51768), .Z(n51769) );
  NOR U64519 ( .A(n51769), .B(n51772), .Z(n54518) );
  IV U64520 ( .A(n54518), .Z(n54515) );
  IV U64521 ( .A(n51770), .Z(n51771) );
  NOR U64522 ( .A(n51771), .B(n51772), .Z(n57952) );
  NOR U64523 ( .A(n51773), .B(n51772), .Z(n57947) );
  IV U64524 ( .A(n51774), .Z(n51776) );
  NOR U64525 ( .A(n51776), .B(n51775), .Z(n51781) );
  IV U64526 ( .A(n51777), .Z(n51779) );
  NOR U64527 ( .A(n51779), .B(n51778), .Z(n51780) );
  NOR U64528 ( .A(n51781), .B(n51780), .Z(n57950) );
  NOR U64529 ( .A(n51782), .B(n57924), .Z(n54513) );
  IV U64530 ( .A(n51783), .Z(n51785) );
  IV U64531 ( .A(n51784), .Z(n51787) );
  NOR U64532 ( .A(n51785), .B(n51787), .Z(n57915) );
  IV U64533 ( .A(n57915), .Z(n57913) );
  IV U64534 ( .A(n51786), .Z(n51788) );
  NOR U64535 ( .A(n51788), .B(n51787), .Z(n57980) );
  IV U64536 ( .A(n51789), .Z(n51790) );
  NOR U64537 ( .A(n51792), .B(n51790), .Z(n57930) );
  IV U64538 ( .A(n51791), .Z(n51793) );
  NOR U64539 ( .A(n51793), .B(n51792), .Z(n55167) );
  IV U64540 ( .A(n51794), .Z(n51795) );
  NOR U64541 ( .A(n51795), .B(n51797), .Z(n57883) );
  IV U64542 ( .A(n51796), .Z(n51798) );
  NOR U64543 ( .A(n51798), .B(n51797), .Z(n55164) );
  NOR U64544 ( .A(n57883), .B(n55164), .Z(n54506) );
  IV U64545 ( .A(n51799), .Z(n51802) );
  IV U64546 ( .A(n51800), .Z(n51801) );
  NOR U64547 ( .A(n51802), .B(n51801), .Z(n57890) );
  IV U64548 ( .A(n57897), .Z(n51806) );
  NOR U64549 ( .A(n57890), .B(n51806), .Z(n54497) );
  IV U64550 ( .A(n51807), .Z(n51808) );
  NOR U64551 ( .A(n51808), .B(n51812), .Z(n57900) );
  IV U64552 ( .A(n51812), .Z(n51809) );
  NOR U64553 ( .A(n51809), .B(n51810), .Z(n51816) );
  IV U64554 ( .A(n51810), .Z(n51811) );
  NOR U64555 ( .A(n51812), .B(n51811), .Z(n51813) );
  NOR U64556 ( .A(n51814), .B(n51813), .Z(n51815) );
  NOR U64557 ( .A(n51816), .B(n51815), .Z(n57895) );
  IV U64558 ( .A(n57895), .Z(n57899) );
  IV U64559 ( .A(n51817), .Z(n51818) );
  NOR U64560 ( .A(n51819), .B(n51818), .Z(n57853) );
  NOR U64561 ( .A(n51822), .B(n51820), .Z(n57856) );
  IV U64562 ( .A(n51821), .Z(n51823) );
  NOR U64563 ( .A(n51823), .B(n51822), .Z(n57861) );
  IV U64564 ( .A(n51824), .Z(n51825) );
  NOR U64565 ( .A(n51825), .B(n51831), .Z(n57864) );
  IV U64566 ( .A(n51826), .Z(n51828) );
  NOR U64567 ( .A(n51828), .B(n51827), .Z(n51829) );
  IV U64568 ( .A(n51829), .Z(n57869) );
  IV U64569 ( .A(n51830), .Z(n51832) );
  NOR U64570 ( .A(n51832), .B(n51831), .Z(n54493) );
  IV U64571 ( .A(n54493), .Z(n54486) );
  IV U64572 ( .A(n51833), .Z(n51835) );
  NOR U64573 ( .A(n51835), .B(n51834), .Z(n54491) );
  IV U64574 ( .A(n51836), .Z(n51837) );
  NOR U64575 ( .A(n51838), .B(n51837), .Z(n55176) );
  IV U64576 ( .A(n51839), .Z(n51841) );
  NOR U64577 ( .A(n51841), .B(n51840), .Z(n55182) );
  NOR U64578 ( .A(n55176), .B(n55182), .Z(n54484) );
  IV U64579 ( .A(n51842), .Z(n51843) );
  NOR U64580 ( .A(n51844), .B(n51843), .Z(n55177) );
  IV U64581 ( .A(n51845), .Z(n51846) );
  NOR U64582 ( .A(n51850), .B(n51846), .Z(n51847) );
  IV U64583 ( .A(n51847), .Z(n55186) );
  IV U64584 ( .A(n51848), .Z(n51849) );
  NOR U64585 ( .A(n51850), .B(n51849), .Z(n55196) );
  IV U64586 ( .A(n55196), .Z(n55189) );
  IV U64587 ( .A(n51851), .Z(n51852) );
  NOR U64588 ( .A(n51853), .B(n51852), .Z(n51856) );
  NOR U64589 ( .A(n51854), .B(n54479), .Z(n51855) );
  NOR U64590 ( .A(n51856), .B(n51855), .Z(n57815) );
  IV U64591 ( .A(n51857), .Z(n51858) );
  NOR U64592 ( .A(n51859), .B(n51858), .Z(n57817) );
  IV U64593 ( .A(n51862), .Z(n51861) );
  NOR U64594 ( .A(n51861), .B(n51860), .Z(n51868) );
  NOR U64595 ( .A(n51863), .B(n51862), .Z(n51866) );
  IV U64596 ( .A(n51864), .Z(n51865) );
  NOR U64597 ( .A(n51866), .B(n51865), .Z(n51867) );
  NOR U64598 ( .A(n51868), .B(n51867), .Z(n57837) );
  IV U64599 ( .A(n51869), .Z(n51870) );
  NOR U64600 ( .A(n51870), .B(n51873), .Z(n57839) );
  IV U64601 ( .A(n51871), .Z(n51872) );
  NOR U64602 ( .A(n51873), .B(n51872), .Z(n51874) );
  IV U64603 ( .A(n51874), .Z(n57836) );
  IV U64604 ( .A(n51875), .Z(n51878) );
  NOR U64605 ( .A(n51876), .B(n51880), .Z(n51877) );
  IV U64606 ( .A(n51877), .Z(n54465) );
  NOR U64607 ( .A(n51878), .B(n54465), .Z(n54467) );
  IV U64608 ( .A(n51879), .Z(n51881) );
  NOR U64609 ( .A(n51881), .B(n51880), .Z(n51882) );
  IV U64610 ( .A(n51882), .Z(n57827) );
  IV U64611 ( .A(n51883), .Z(n51884) );
  NOR U64612 ( .A(n54431), .B(n51884), .Z(n57774) );
  IV U64613 ( .A(n51885), .Z(n51887) );
  NOR U64614 ( .A(n51887), .B(n51886), .Z(n57753) );
  IV U64615 ( .A(n51888), .Z(n51889) );
  NOR U64616 ( .A(n51892), .B(n51889), .Z(n57739) );
  IV U64617 ( .A(n51890), .Z(n51891) );
  NOR U64618 ( .A(n51892), .B(n51891), .Z(n57742) );
  NOR U64619 ( .A(n51893), .B(n51898), .Z(n51894) );
  IV U64620 ( .A(n51894), .Z(n51896) );
  NOR U64621 ( .A(n51896), .B(n51895), .Z(n57734) );
  IV U64622 ( .A(n57734), .Z(n57738) );
  IV U64623 ( .A(n51897), .Z(n51901) );
  NOR U64624 ( .A(n51907), .B(n51898), .Z(n51899) );
  IV U64625 ( .A(n51899), .Z(n51900) );
  NOR U64626 ( .A(n51901), .B(n51900), .Z(n51902) );
  IV U64627 ( .A(n51902), .Z(n57737) );
  IV U64628 ( .A(n51903), .Z(n51904) );
  NOR U64629 ( .A(n51907), .B(n51904), .Z(n57759) );
  IV U64630 ( .A(n51908), .Z(n51905) );
  NOR U64631 ( .A(n51907), .B(n51905), .Z(n51912) );
  IV U64632 ( .A(n51906), .Z(n51910) );
  XOR U64633 ( .A(n51908), .B(n51907), .Z(n51909) );
  NOR U64634 ( .A(n51910), .B(n51909), .Z(n51911) );
  NOR U64635 ( .A(n51912), .B(n51911), .Z(n57783) );
  IV U64636 ( .A(n51913), .Z(n51914) );
  NOR U64637 ( .A(n51914), .B(n54415), .Z(n57780) );
  IV U64638 ( .A(n57780), .Z(n57785) );
  IV U64639 ( .A(n51915), .Z(n51916) );
  NOR U64640 ( .A(n51916), .B(n54415), .Z(n54410) );
  IV U64641 ( .A(n51917), .Z(n51918) );
  NOR U64642 ( .A(n51921), .B(n51918), .Z(n54402) );
  IV U64643 ( .A(n54402), .Z(n54399) );
  IV U64644 ( .A(n51919), .Z(n51920) );
  NOR U64645 ( .A(n51921), .B(n51920), .Z(n55227) );
  IV U64646 ( .A(n51922), .Z(n51924) );
  IV U64647 ( .A(n51923), .Z(n51926) );
  NOR U64648 ( .A(n51924), .B(n51926), .Z(n55224) );
  IV U64649 ( .A(n51925), .Z(n51927) );
  NOR U64650 ( .A(n51927), .B(n51926), .Z(n55216) );
  IV U64651 ( .A(n51928), .Z(n51929) );
  NOR U64652 ( .A(n51931), .B(n51929), .Z(n55219) );
  IV U64653 ( .A(n51930), .Z(n51932) );
  NOR U64654 ( .A(n51932), .B(n51931), .Z(n55232) );
  IV U64655 ( .A(n51933), .Z(n51934) );
  NOR U64656 ( .A(n51935), .B(n51934), .Z(n51939) );
  NOR U64657 ( .A(n51937), .B(n51936), .Z(n51938) );
  NOR U64658 ( .A(n51939), .B(n51938), .Z(n55240) );
  IV U64659 ( .A(n51940), .Z(n51943) );
  IV U64660 ( .A(n51941), .Z(n51942) );
  NOR U64661 ( .A(n51943), .B(n51942), .Z(n55264) );
  IV U64662 ( .A(n51944), .Z(n51946) );
  NOR U64663 ( .A(n51946), .B(n51945), .Z(n55267) );
  IV U64664 ( .A(n51947), .Z(n51950) );
  NOR U64665 ( .A(n51948), .B(n51952), .Z(n51949) );
  IV U64666 ( .A(n51949), .Z(n54370) );
  NOR U64667 ( .A(n51950), .B(n54370), .Z(n55256) );
  IV U64668 ( .A(n51951), .Z(n51953) );
  NOR U64669 ( .A(n51953), .B(n51952), .Z(n54372) );
  IV U64670 ( .A(n51954), .Z(n51955) );
  NOR U64671 ( .A(n51956), .B(n51955), .Z(n51957) );
  IV U64672 ( .A(n51957), .Z(n57699) );
  IV U64673 ( .A(n51958), .Z(n51959) );
  NOR U64674 ( .A(n51959), .B(n54354), .Z(n57700) );
  IV U64675 ( .A(n57700), .Z(n57704) );
  IV U64676 ( .A(n51960), .Z(n51965) );
  IV U64677 ( .A(n51961), .Z(n51962) );
  NOR U64678 ( .A(n51965), .B(n51962), .Z(n57672) );
  IV U64679 ( .A(n51963), .Z(n51964) );
  NOR U64680 ( .A(n51965), .B(n51964), .Z(n57669) );
  IV U64681 ( .A(n51966), .Z(n51967) );
  NOR U64682 ( .A(n51976), .B(n51967), .Z(n57680) );
  IV U64683 ( .A(n51968), .Z(n51969) );
  NOR U64684 ( .A(n51976), .B(n51969), .Z(n57677) );
  IV U64685 ( .A(n51970), .Z(n51973) );
  IV U64686 ( .A(n51971), .Z(n51972) );
  NOR U64687 ( .A(n51973), .B(n51972), .Z(n55279) );
  IV U64688 ( .A(n51974), .Z(n51975) );
  NOR U64689 ( .A(n51976), .B(n51975), .Z(n55280) );
  NOR U64690 ( .A(n55279), .B(n55280), .Z(n51977) );
  IV U64691 ( .A(n51977), .Z(n54352) );
  IV U64692 ( .A(n51978), .Z(n51983) );
  IV U64693 ( .A(n51979), .Z(n51980) );
  NOR U64694 ( .A(n51981), .B(n51980), .Z(n51982) );
  IV U64695 ( .A(n51982), .Z(n54347) );
  NOR U64696 ( .A(n51983), .B(n54347), .Z(n55284) );
  IV U64697 ( .A(n51984), .Z(n51988) );
  NOR U64698 ( .A(n51986), .B(n51985), .Z(n51987) );
  IV U64699 ( .A(n51987), .Z(n54343) );
  NOR U64700 ( .A(n51988), .B(n54343), .Z(n51989) );
  NOR U64701 ( .A(n51990), .B(n51989), .Z(n55291) );
  IV U64702 ( .A(n55291), .Z(n54341) );
  IV U64703 ( .A(n51991), .Z(n51992) );
  NOR U64704 ( .A(n51993), .B(n51992), .Z(n51994) );
  NOR U64705 ( .A(n51995), .B(n51994), .Z(n55290) );
  NOR U64706 ( .A(n51997), .B(n51996), .Z(n55301) );
  IV U64707 ( .A(n51998), .Z(n52000) );
  IV U64708 ( .A(n51999), .Z(n54326) );
  NOR U64709 ( .A(n52000), .B(n54326), .Z(n55320) );
  IV U64710 ( .A(n52001), .Z(n52002) );
  NOR U64711 ( .A(n52002), .B(n54322), .Z(n52003) );
  IV U64712 ( .A(n52003), .Z(n55319) );
  IV U64713 ( .A(n52004), .Z(n52005) );
  NOR U64714 ( .A(n52005), .B(n52011), .Z(n52006) );
  IV U64715 ( .A(n52006), .Z(n57638) );
  IV U64716 ( .A(n52007), .Z(n52009) );
  NOR U64717 ( .A(n52009), .B(n52008), .Z(n52014) );
  IV U64718 ( .A(n52010), .Z(n52012) );
  NOR U64719 ( .A(n52012), .B(n52011), .Z(n52013) );
  NOR U64720 ( .A(n52014), .B(n52013), .Z(n57635) );
  IV U64721 ( .A(n57635), .Z(n54316) );
  NOR U64722 ( .A(n52016), .B(n52015), .Z(n54310) );
  IV U64723 ( .A(n54310), .Z(n54303) );
  IV U64724 ( .A(n52017), .Z(n52018) );
  NOR U64725 ( .A(n54292), .B(n52018), .Z(n55345) );
  NOR U64726 ( .A(n52020), .B(n52019), .Z(n57611) );
  IV U64727 ( .A(n52021), .Z(n52022) );
  NOR U64728 ( .A(n52022), .B(n54280), .Z(n57608) );
  IV U64729 ( .A(n52026), .Z(n52023) );
  NOR U64730 ( .A(n52023), .B(n52024), .Z(n52030) );
  IV U64731 ( .A(n52024), .Z(n52025) );
  NOR U64732 ( .A(n52026), .B(n52025), .Z(n52027) );
  NOR U64733 ( .A(n52028), .B(n52027), .Z(n52029) );
  NOR U64734 ( .A(n52030), .B(n52029), .Z(n55353) );
  IV U64735 ( .A(n52031), .Z(n52032) );
  NOR U64736 ( .A(n52033), .B(n52032), .Z(n55350) );
  IV U64737 ( .A(n52034), .Z(n52035) );
  NOR U64738 ( .A(n52035), .B(n54263), .Z(n55375) );
  IV U64739 ( .A(n52036), .Z(n52037) );
  NOR U64740 ( .A(n52038), .B(n52037), .Z(n57618) );
  IV U64741 ( .A(n52039), .Z(n52043) );
  IV U64742 ( .A(n52040), .Z(n52041) );
  NOR U64743 ( .A(n52043), .B(n52041), .Z(n55369) );
  NOR U64744 ( .A(n57618), .B(n55369), .Z(n54257) );
  IV U64745 ( .A(n52042), .Z(n52046) );
  NOR U64746 ( .A(n52044), .B(n52043), .Z(n52045) );
  IV U64747 ( .A(n52045), .Z(n52048) );
  NOR U64748 ( .A(n52046), .B(n52048), .Z(n55366) );
  IV U64749 ( .A(n52047), .Z(n52049) );
  NOR U64750 ( .A(n52049), .B(n52048), .Z(n55399) );
  IV U64751 ( .A(n52050), .Z(n52051) );
  NOR U64752 ( .A(n52060), .B(n52051), .Z(n52057) );
  IV U64753 ( .A(n52052), .Z(n52055) );
  IV U64754 ( .A(n52053), .Z(n52054) );
  NOR U64755 ( .A(n52055), .B(n52054), .Z(n52056) );
  NOR U64756 ( .A(n52057), .B(n52056), .Z(n55385) );
  IV U64757 ( .A(n52058), .Z(n52059) );
  NOR U64758 ( .A(n52060), .B(n52059), .Z(n55386) );
  IV U64759 ( .A(n52061), .Z(n52064) );
  IV U64760 ( .A(n52062), .Z(n52063) );
  NOR U64761 ( .A(n52064), .B(n52063), .Z(n55394) );
  NOR U64762 ( .A(n55386), .B(n55394), .Z(n54255) );
  IV U64763 ( .A(n52065), .Z(n52066) );
  NOR U64764 ( .A(n54245), .B(n52066), .Z(n55411) );
  IV U64765 ( .A(n52067), .Z(n52069) );
  NOR U64766 ( .A(n52069), .B(n52068), .Z(n55417) );
  IV U64767 ( .A(n52070), .Z(n52071) );
  NOR U64768 ( .A(n52072), .B(n52071), .Z(n57586) );
  IV U64769 ( .A(n52073), .Z(n52075) );
  NOR U64770 ( .A(n52075), .B(n52074), .Z(n55425) );
  NOR U64771 ( .A(n57586), .B(n55425), .Z(n52076) );
  IV U64772 ( .A(n52076), .Z(n54244) );
  IV U64773 ( .A(n52077), .Z(n52079) );
  IV U64774 ( .A(n52078), .Z(n52081) );
  NOR U64775 ( .A(n52079), .B(n52081), .Z(n57587) );
  IV U64776 ( .A(n52080), .Z(n52082) );
  NOR U64777 ( .A(n52082), .B(n52081), .Z(n55414) );
  IV U64778 ( .A(n52083), .Z(n52084) );
  NOR U64779 ( .A(n52084), .B(n52086), .Z(n57570) );
  IV U64780 ( .A(n52085), .Z(n52087) );
  NOR U64781 ( .A(n52087), .B(n52086), .Z(n57564) );
  NOR U64782 ( .A(n52089), .B(n52088), .Z(n52094) );
  IV U64783 ( .A(n52090), .Z(n54231) );
  IV U64784 ( .A(n52091), .Z(n52092) );
  NOR U64785 ( .A(n54231), .B(n52092), .Z(n52093) );
  NOR U64786 ( .A(n52094), .B(n52093), .Z(n57563) );
  IV U64787 ( .A(n52095), .Z(n52096) );
  NOR U64788 ( .A(n52096), .B(n54234), .Z(n55434) );
  IV U64789 ( .A(n52097), .Z(n52098) );
  NOR U64790 ( .A(n52099), .B(n52098), .Z(n55456) );
  IV U64791 ( .A(n52100), .Z(n52102) );
  NOR U64792 ( .A(n52102), .B(n52101), .Z(n55444) );
  NOR U64793 ( .A(n55456), .B(n55444), .Z(n54222) );
  IV U64794 ( .A(n52103), .Z(n52105) );
  IV U64795 ( .A(n52104), .Z(n52115) );
  NOR U64796 ( .A(n52105), .B(n52115), .Z(n52110) );
  IV U64797 ( .A(n52106), .Z(n52108) );
  NOR U64798 ( .A(n52108), .B(n52107), .Z(n52109) );
  NOR U64799 ( .A(n52110), .B(n52109), .Z(n55463) );
  IV U64800 ( .A(n52111), .Z(n52112) );
  NOR U64801 ( .A(n52113), .B(n52112), .Z(n55457) );
  IV U64802 ( .A(n52114), .Z(n52116) );
  NOR U64803 ( .A(n52116), .B(n52115), .Z(n52117) );
  IV U64804 ( .A(n52117), .Z(n55449) );
  NOR U64805 ( .A(n52119), .B(n52118), .Z(n55482) );
  NOR U64806 ( .A(n55482), .B(n55451), .Z(n52120) );
  IV U64807 ( .A(n52120), .Z(n54220) );
  IV U64808 ( .A(n52121), .Z(n54214) );
  IV U64809 ( .A(n52122), .Z(n52123) );
  NOR U64810 ( .A(n54214), .B(n52123), .Z(n52124) );
  IV U64811 ( .A(n52124), .Z(n55472) );
  IV U64812 ( .A(n52128), .Z(n52125) );
  NOR U64813 ( .A(n52126), .B(n52125), .Z(n52133) );
  IV U64814 ( .A(n52127), .Z(n52131) );
  NOR U64815 ( .A(n52129), .B(n52128), .Z(n52130) );
  NOR U64816 ( .A(n52131), .B(n52130), .Z(n52132) );
  NOR U64817 ( .A(n52133), .B(n52132), .Z(n55475) );
  IV U64818 ( .A(n52137), .Z(n52134) );
  NOR U64819 ( .A(n52136), .B(n52134), .Z(n52145) );
  IV U64820 ( .A(n52135), .Z(n52143) );
  IV U64821 ( .A(n52136), .Z(n52138) );
  NOR U64822 ( .A(n52138), .B(n52137), .Z(n52140) );
  NOR U64823 ( .A(n52140), .B(n52139), .Z(n52141) );
  IV U64824 ( .A(n52141), .Z(n52142) );
  NOR U64825 ( .A(n52143), .B(n52142), .Z(n52144) );
  NOR U64826 ( .A(n52145), .B(n52144), .Z(n57513) );
  IV U64827 ( .A(n52146), .Z(n52148) );
  XOR U64828 ( .A(n52154), .B(n52155), .Z(n52147) );
  NOR U64829 ( .A(n52148), .B(n52147), .Z(n54140) );
  IV U64830 ( .A(n52149), .Z(n52150) );
  NOR U64831 ( .A(n52150), .B(n52155), .Z(n54142) );
  IV U64832 ( .A(n54142), .Z(n54134) );
  XOR U64833 ( .A(n54140), .B(n54134), .Z(n54133) );
  IV U64834 ( .A(n52151), .Z(n52153) );
  NOR U64835 ( .A(n52153), .B(n52152), .Z(n52158) );
  IV U64836 ( .A(n52154), .Z(n52156) );
  NOR U64837 ( .A(n52156), .B(n52155), .Z(n52157) );
  NOR U64838 ( .A(n52158), .B(n52157), .Z(n57483) );
  IV U64839 ( .A(n52159), .Z(n52160) );
  NOR U64840 ( .A(n52161), .B(n52160), .Z(n52166) );
  IV U64841 ( .A(n52162), .Z(n52164) );
  NOR U64842 ( .A(n52164), .B(n52163), .Z(n52165) );
  NOR U64843 ( .A(n52166), .B(n52165), .Z(n57485) );
  IV U64844 ( .A(n57485), .Z(n54131) );
  IV U64845 ( .A(n52167), .Z(n52168) );
  NOR U64846 ( .A(n52171), .B(n52168), .Z(n57492) );
  IV U64847 ( .A(n52169), .Z(n52170) );
  NOR U64848 ( .A(n52171), .B(n52170), .Z(n57489) );
  IV U64849 ( .A(n52172), .Z(n52174) );
  IV U64850 ( .A(n52173), .Z(n52178) );
  NOR U64851 ( .A(n52174), .B(n52178), .Z(n55499) );
  IV U64852 ( .A(n52175), .Z(n52176) );
  NOR U64853 ( .A(n52176), .B(n52178), .Z(n55496) );
  IV U64854 ( .A(n52177), .Z(n52179) );
  NOR U64855 ( .A(n52179), .B(n52178), .Z(n52180) );
  NOR U64856 ( .A(n52181), .B(n52180), .Z(n55505) );
  IV U64857 ( .A(n52182), .Z(n52183) );
  NOR U64858 ( .A(n52183), .B(n52185), .Z(n55508) );
  IV U64859 ( .A(n52184), .Z(n52186) );
  NOR U64860 ( .A(n52186), .B(n52185), .Z(n55512) );
  IV U64861 ( .A(n52187), .Z(n52188) );
  NOR U64862 ( .A(n52188), .B(n52190), .Z(n57453) );
  IV U64863 ( .A(n57453), .Z(n57459) );
  IV U64864 ( .A(n52189), .Z(n52191) );
  NOR U64865 ( .A(n52191), .B(n52190), .Z(n57468) );
  IV U64866 ( .A(n52192), .Z(n52198) );
  NOR U64867 ( .A(n52193), .B(n52200), .Z(n52194) );
  IV U64868 ( .A(n52194), .Z(n52195) );
  NOR U64869 ( .A(n52196), .B(n52195), .Z(n52197) );
  IV U64870 ( .A(n52197), .Z(n52205) );
  NOR U64871 ( .A(n52198), .B(n52205), .Z(n57465) );
  IV U64872 ( .A(n52199), .Z(n52203) );
  NOR U64873 ( .A(n52201), .B(n52200), .Z(n52202) );
  IV U64874 ( .A(n52202), .Z(n54111) );
  NOR U64875 ( .A(n52203), .B(n54111), .Z(n52208) );
  IV U64876 ( .A(n52204), .Z(n52206) );
  NOR U64877 ( .A(n52206), .B(n52205), .Z(n52207) );
  NOR U64878 ( .A(n52208), .B(n52207), .Z(n55515) );
  IV U64879 ( .A(n52209), .Z(n52210) );
  NOR U64880 ( .A(n52210), .B(n52213), .Z(n57432) );
  IV U64881 ( .A(n52211), .Z(n52212) );
  NOR U64882 ( .A(n52213), .B(n52212), .Z(n57429) );
  IV U64883 ( .A(n52214), .Z(n52216) );
  NOR U64884 ( .A(n52216), .B(n52215), .Z(n52221) );
  IV U64885 ( .A(n52217), .Z(n52219) );
  NOR U64886 ( .A(n52219), .B(n52218), .Z(n52220) );
  NOR U64887 ( .A(n52221), .B(n52220), .Z(n55542) );
  IV U64888 ( .A(n52222), .Z(n52224) );
  NOR U64889 ( .A(n52224), .B(n52223), .Z(n52229) );
  IV U64890 ( .A(n52225), .Z(n52226) );
  NOR U64891 ( .A(n52227), .B(n52226), .Z(n52228) );
  NOR U64892 ( .A(n52229), .B(n52228), .Z(n55544) );
  IV U64893 ( .A(n52230), .Z(n52231) );
  NOR U64894 ( .A(n52231), .B(n52233), .Z(n57440) );
  IV U64895 ( .A(n52232), .Z(n52234) );
  NOR U64896 ( .A(n52234), .B(n52233), .Z(n57437) );
  IV U64897 ( .A(n52235), .Z(n52237) );
  IV U64898 ( .A(n52236), .Z(n52239) );
  NOR U64899 ( .A(n52237), .B(n52239), .Z(n55525) );
  IV U64900 ( .A(n52238), .Z(n52240) );
  NOR U64901 ( .A(n52240), .B(n52239), .Z(n55522) );
  IV U64902 ( .A(n52241), .Z(n52242) );
  NOR U64903 ( .A(n52243), .B(n52242), .Z(n55534) );
  NOR U64904 ( .A(n52245), .B(n52244), .Z(n55548) );
  NOR U64905 ( .A(n55534), .B(n55548), .Z(n52246) );
  IV U64906 ( .A(n52246), .Z(n54109) );
  IV U64907 ( .A(n52247), .Z(n52252) );
  IV U64908 ( .A(n52248), .Z(n52249) );
  NOR U64909 ( .A(n52252), .B(n52249), .Z(n55536) );
  IV U64910 ( .A(n52250), .Z(n52251) );
  NOR U64911 ( .A(n52252), .B(n52251), .Z(n55535) );
  IV U64912 ( .A(n52253), .Z(n52254) );
  NOR U64913 ( .A(n52255), .B(n52254), .Z(n57407) );
  IV U64914 ( .A(n52256), .Z(n52257) );
  NOR U64915 ( .A(n54104), .B(n52257), .Z(n57397) );
  NOR U64916 ( .A(n52258), .B(n52261), .Z(n52259) );
  IV U64917 ( .A(n52259), .Z(n57404) );
  IV U64918 ( .A(n52260), .Z(n52262) );
  NOR U64919 ( .A(n52262), .B(n52261), .Z(n57376) );
  IV U64920 ( .A(n57376), .Z(n57375) );
  IV U64921 ( .A(n52263), .Z(n52264) );
  NOR U64922 ( .A(n54098), .B(n52264), .Z(n57370) );
  IV U64923 ( .A(n52265), .Z(n52266) );
  NOR U64924 ( .A(n52266), .B(n52271), .Z(n57385) );
  IV U64925 ( .A(n57385), .Z(n57384) );
  IV U64926 ( .A(n52267), .Z(n52268) );
  NOR U64927 ( .A(n52269), .B(n52268), .Z(n52274) );
  IV U64928 ( .A(n52270), .Z(n52272) );
  NOR U64929 ( .A(n52272), .B(n52271), .Z(n52273) );
  NOR U64930 ( .A(n52274), .B(n52273), .Z(n57361) );
  IV U64931 ( .A(n52275), .Z(n52276) );
  NOR U64932 ( .A(n52276), .B(n52282), .Z(n57338) );
  IV U64933 ( .A(n52277), .Z(n52278) );
  NOR U64934 ( .A(n52279), .B(n52278), .Z(n57349) );
  IV U64935 ( .A(n52280), .Z(n52281) );
  NOR U64936 ( .A(n52282), .B(n52281), .Z(n57341) );
  NOR U64937 ( .A(n57349), .B(n57341), .Z(n52283) );
  IV U64938 ( .A(n52283), .Z(n54080) );
  IV U64939 ( .A(n52284), .Z(n52286) );
  IV U64940 ( .A(n52285), .Z(n52289) );
  NOR U64941 ( .A(n52286), .B(n52289), .Z(n57346) );
  IV U64942 ( .A(n52287), .Z(n52288) );
  NOR U64943 ( .A(n52289), .B(n52288), .Z(n57329) );
  NOR U64944 ( .A(n52291), .B(n52290), .Z(n55567) );
  IV U64945 ( .A(n55567), .Z(n55565) );
  NOR U64946 ( .A(n52292), .B(n52294), .Z(n55553) );
  IV U64947 ( .A(n52293), .Z(n52295) );
  NOR U64948 ( .A(n52295), .B(n52294), .Z(n55559) );
  IV U64949 ( .A(n52296), .Z(n52297) );
  NOR U64950 ( .A(n52298), .B(n52297), .Z(n52303) );
  IV U64951 ( .A(n52299), .Z(n52301) );
  NOR U64952 ( .A(n52301), .B(n52300), .Z(n52302) );
  NOR U64953 ( .A(n52303), .B(n52302), .Z(n55551) );
  IV U64954 ( .A(n55551), .Z(n54073) );
  IV U64955 ( .A(n52304), .Z(n52305) );
  NOR U64956 ( .A(n52306), .B(n52305), .Z(n55578) );
  IV U64957 ( .A(n52307), .Z(n52308) );
  NOR U64958 ( .A(n52312), .B(n52308), .Z(n55577) );
  NOR U64959 ( .A(n52310), .B(n52309), .Z(n52311) );
  NOR U64960 ( .A(n52312), .B(n52311), .Z(n55576) );
  IV U64961 ( .A(n52313), .Z(n52315) );
  XOR U64962 ( .A(n52323), .B(n52325), .Z(n52314) );
  NOR U64963 ( .A(n52315), .B(n52314), .Z(n55583) );
  IV U64964 ( .A(n52316), .Z(n52317) );
  NOR U64965 ( .A(n52325), .B(n52317), .Z(n55586) );
  IV U64966 ( .A(n52318), .Z(n52319) );
  NOR U64967 ( .A(n52319), .B(n52325), .Z(n55591) );
  IV U64968 ( .A(n52320), .Z(n52321) );
  NOR U64969 ( .A(n52322), .B(n52321), .Z(n52327) );
  IV U64970 ( .A(n52323), .Z(n52324) );
  NOR U64971 ( .A(n52325), .B(n52324), .Z(n52326) );
  NOR U64972 ( .A(n52327), .B(n52326), .Z(n55595) );
  IV U64973 ( .A(n52328), .Z(n52329) );
  NOR U64974 ( .A(n52330), .B(n52329), .Z(n55607) );
  IV U64975 ( .A(n52331), .Z(n52332) );
  NOR U64976 ( .A(n52333), .B(n52332), .Z(n55597) );
  NOR U64977 ( .A(n55607), .B(n55597), .Z(n54070) );
  NOR U64978 ( .A(n52335), .B(n52334), .Z(n52340) );
  IV U64979 ( .A(n52336), .Z(n52337) );
  NOR U64980 ( .A(n52338), .B(n52337), .Z(n52339) );
  NOR U64981 ( .A(n52340), .B(n52339), .Z(n55605) );
  IV U64982 ( .A(n52341), .Z(n52342) );
  NOR U64983 ( .A(n52343), .B(n52342), .Z(n52344) );
  IV U64984 ( .A(n52344), .Z(n57297) );
  NOR U64985 ( .A(n52345), .B(n52352), .Z(n57298) );
  IV U64986 ( .A(n52346), .Z(n52347) );
  NOR U64987 ( .A(n52347), .B(n52352), .Z(n57264) );
  IV U64988 ( .A(n52348), .Z(n52349) );
  NOR U64989 ( .A(n52349), .B(n52356), .Z(n52354) );
  IV U64990 ( .A(n52350), .Z(n52351) );
  NOR U64991 ( .A(n52352), .B(n52351), .Z(n52353) );
  NOR U64992 ( .A(n52354), .B(n52353), .Z(n57262) );
  IV U64993 ( .A(n57262), .Z(n54069) );
  IV U64994 ( .A(n52355), .Z(n52362) );
  NOR U64995 ( .A(n52357), .B(n52356), .Z(n52358) );
  IV U64996 ( .A(n52358), .Z(n52359) );
  NOR U64997 ( .A(n52360), .B(n52359), .Z(n52361) );
  IV U64998 ( .A(n52361), .Z(n52364) );
  NOR U64999 ( .A(n52362), .B(n52364), .Z(n57303) );
  IV U65000 ( .A(n52363), .Z(n52365) );
  NOR U65001 ( .A(n52365), .B(n52364), .Z(n57306) );
  NOR U65002 ( .A(n52368), .B(n52366), .Z(n57269) );
  IV U65003 ( .A(n52367), .Z(n52369) );
  NOR U65004 ( .A(n52369), .B(n52368), .Z(n57275) );
  IV U65005 ( .A(n52370), .Z(n52371) );
  NOR U65006 ( .A(n52371), .B(n52377), .Z(n57272) );
  IV U65007 ( .A(n52372), .Z(n52374) );
  NOR U65008 ( .A(n52374), .B(n52373), .Z(n52379) );
  IV U65009 ( .A(n52375), .Z(n52376) );
  NOR U65010 ( .A(n52377), .B(n52376), .Z(n52378) );
  NOR U65011 ( .A(n52379), .B(n52378), .Z(n57281) );
  IV U65012 ( .A(n52380), .Z(n52381) );
  NOR U65013 ( .A(n52382), .B(n52381), .Z(n55612) );
  IV U65014 ( .A(n52383), .Z(n52385) );
  NOR U65015 ( .A(n52385), .B(n52384), .Z(n57283) );
  NOR U65016 ( .A(n55612), .B(n57283), .Z(n54068) );
  IV U65017 ( .A(n52386), .Z(n52387) );
  NOR U65018 ( .A(n52387), .B(n54055), .Z(n52388) );
  IV U65019 ( .A(n52388), .Z(n57248) );
  IV U65020 ( .A(n52389), .Z(n52391) );
  IV U65021 ( .A(n52390), .Z(n54051) );
  NOR U65022 ( .A(n52391), .B(n54051), .Z(n55623) );
  IV U65023 ( .A(n52392), .Z(n52394) );
  NOR U65024 ( .A(n52394), .B(n52393), .Z(n54031) );
  IV U65025 ( .A(n52395), .Z(n52397) );
  NOR U65026 ( .A(n52397), .B(n52396), .Z(n52398) );
  NOR U65027 ( .A(n54031), .B(n52398), .Z(n55644) );
  IV U65028 ( .A(n52399), .Z(n52401) );
  NOR U65029 ( .A(n52401), .B(n52400), .Z(n52407) );
  IV U65030 ( .A(n52402), .Z(n52405) );
  NOR U65031 ( .A(n52403), .B(n52412), .Z(n52404) );
  IV U65032 ( .A(n52404), .Z(n54002) );
  NOR U65033 ( .A(n52405), .B(n54002), .Z(n52406) );
  NOR U65034 ( .A(n52407), .B(n52406), .Z(n55660) );
  IV U65035 ( .A(n52408), .Z(n52409) );
  NOR U65036 ( .A(n52410), .B(n52409), .Z(n52415) );
  IV U65037 ( .A(n52411), .Z(n52413) );
  NOR U65038 ( .A(n52413), .B(n52412), .Z(n52414) );
  NOR U65039 ( .A(n52415), .B(n52414), .Z(n57211) );
  NOR U65040 ( .A(n52417), .B(n52416), .Z(n57213) );
  IV U65041 ( .A(n52418), .Z(n52420) );
  NOR U65042 ( .A(n52420), .B(n52419), .Z(n55679) );
  IV U65043 ( .A(n52421), .Z(n52423) );
  NOR U65044 ( .A(n52423), .B(n52422), .Z(n55670) );
  NOR U65045 ( .A(n55679), .B(n55670), .Z(n53997) );
  IV U65046 ( .A(n52424), .Z(n52425) );
  NOR U65047 ( .A(n53995), .B(n52425), .Z(n52426) );
  IV U65048 ( .A(n52426), .Z(n53990) );
  IV U65049 ( .A(n52427), .Z(n52428) );
  NOR U65050 ( .A(n52428), .B(n53987), .Z(n53981) );
  IV U65051 ( .A(n52429), .Z(n52430) );
  NOR U65052 ( .A(n52430), .B(n52437), .Z(n52435) );
  IV U65053 ( .A(n52431), .Z(n52433) );
  NOR U65054 ( .A(n52433), .B(n52432), .Z(n52434) );
  NOR U65055 ( .A(n52435), .B(n52434), .Z(n55686) );
  IV U65056 ( .A(n55686), .Z(n53975) );
  IV U65057 ( .A(n52436), .Z(n52438) );
  NOR U65058 ( .A(n52438), .B(n52437), .Z(n55688) );
  IV U65059 ( .A(n52439), .Z(n52440) );
  NOR U65060 ( .A(n52441), .B(n52440), .Z(n52445) );
  NOR U65061 ( .A(n52443), .B(n52442), .Z(n52444) );
  NOR U65062 ( .A(n52445), .B(n52444), .Z(n55685) );
  IV U65063 ( .A(n55685), .Z(n53974) );
  NOR U65064 ( .A(n52450), .B(n52446), .Z(n57187) );
  IV U65065 ( .A(n52447), .Z(n52448) );
  NOR U65066 ( .A(n52448), .B(n52450), .Z(n57190) );
  IV U65067 ( .A(n52449), .Z(n52451) );
  NOR U65068 ( .A(n52451), .B(n52450), .Z(n55699) );
  IV U65069 ( .A(n52452), .Z(n52453) );
  NOR U65070 ( .A(n52454), .B(n52453), .Z(n52459) );
  IV U65071 ( .A(n52455), .Z(n52457) );
  IV U65072 ( .A(n52456), .Z(n52463) );
  NOR U65073 ( .A(n52457), .B(n52463), .Z(n52458) );
  NOR U65074 ( .A(n52459), .B(n52458), .Z(n55698) );
  NOR U65075 ( .A(n52461), .B(n52460), .Z(n55717) );
  IV U65076 ( .A(n52462), .Z(n52464) );
  NOR U65077 ( .A(n52464), .B(n52463), .Z(n55693) );
  NOR U65078 ( .A(n55717), .B(n55693), .Z(n53972) );
  IV U65079 ( .A(n52465), .Z(n52466) );
  XOR U65080 ( .A(n52467), .B(n53965), .Z(n53969) );
  NOR U65081 ( .A(n52466), .B(n53969), .Z(n55718) );
  IV U65082 ( .A(n52467), .Z(n52468) );
  NOR U65083 ( .A(n52468), .B(n53965), .Z(n52469) );
  IV U65084 ( .A(n52469), .Z(n55712) );
  IV U65085 ( .A(n52470), .Z(n52471) );
  NOR U65086 ( .A(n52472), .B(n52471), .Z(n57162) );
  IV U65087 ( .A(n52473), .Z(n52475) );
  NOR U65088 ( .A(n52475), .B(n52474), .Z(n55705) );
  NOR U65089 ( .A(n57162), .B(n55705), .Z(n53963) );
  IV U65090 ( .A(n52476), .Z(n52477) );
  NOR U65091 ( .A(n53960), .B(n52477), .Z(n53955) );
  IV U65092 ( .A(n52478), .Z(n52479) );
  NOR U65093 ( .A(n52480), .B(n52479), .Z(n53952) );
  IV U65094 ( .A(n53952), .Z(n53946) );
  IV U65095 ( .A(n52481), .Z(n52483) );
  IV U65096 ( .A(n52482), .Z(n52485) );
  NOR U65097 ( .A(n52483), .B(n52485), .Z(n53951) );
  IV U65098 ( .A(n52484), .Z(n52486) );
  NOR U65099 ( .A(n52486), .B(n52485), .Z(n53942) );
  IV U65100 ( .A(n53942), .Z(n53937) );
  IV U65101 ( .A(n52487), .Z(n52488) );
  NOR U65102 ( .A(n52489), .B(n52488), .Z(n57133) );
  NOR U65103 ( .A(n53934), .B(n52490), .Z(n57130) );
  IV U65104 ( .A(n52491), .Z(n57148) );
  IV U65105 ( .A(n55741), .Z(n55734) );
  IV U65106 ( .A(n52492), .Z(n52493) );
  NOR U65107 ( .A(n52493), .B(n53926), .Z(n55729) );
  IV U65108 ( .A(n52494), .Z(n52498) );
  NOR U65109 ( .A(n52496), .B(n52495), .Z(n52497) );
  IV U65110 ( .A(n52497), .Z(n53921) );
  NOR U65111 ( .A(n52498), .B(n53921), .Z(n52499) );
  IV U65112 ( .A(n52499), .Z(n55761) );
  IV U65113 ( .A(n52500), .Z(n52501) );
  NOR U65114 ( .A(n52501), .B(n53903), .Z(n55750) );
  IV U65115 ( .A(n52502), .Z(n52503) );
  NOR U65116 ( .A(n52503), .B(n53903), .Z(n52504) );
  IV U65117 ( .A(n52504), .Z(n55749) );
  IV U65118 ( .A(n52505), .Z(n52507) );
  NOR U65119 ( .A(n52507), .B(n52506), .Z(n52514) );
  IV U65120 ( .A(n52508), .Z(n52512) );
  NOR U65121 ( .A(n52510), .B(n52509), .Z(n52511) );
  IV U65122 ( .A(n52511), .Z(n53895) );
  NOR U65123 ( .A(n52512), .B(n53895), .Z(n52513) );
  NOR U65124 ( .A(n52514), .B(n52513), .Z(n57111) );
  IV U65125 ( .A(n52515), .Z(n52517) );
  NOR U65126 ( .A(n52517), .B(n52516), .Z(n57101) );
  IV U65127 ( .A(n52518), .Z(n52519) );
  NOR U65128 ( .A(n52520), .B(n52519), .Z(n57103) );
  NOR U65129 ( .A(n57101), .B(n57103), .Z(n53893) );
  IV U65130 ( .A(n52521), .Z(n52522) );
  NOR U65131 ( .A(n52523), .B(n52522), .Z(n57084) );
  IV U65132 ( .A(n52524), .Z(n52525) );
  NOR U65133 ( .A(n52526), .B(n52525), .Z(n57106) );
  NOR U65134 ( .A(n57084), .B(n57106), .Z(n53892) );
  NOR U65135 ( .A(n52529), .B(n52527), .Z(n57081) );
  IV U65136 ( .A(n52528), .Z(n52530) );
  NOR U65137 ( .A(n52530), .B(n52529), .Z(n55775) );
  IV U65138 ( .A(n52531), .Z(n53878) );
  IV U65139 ( .A(n52532), .Z(n52533) );
  NOR U65140 ( .A(n53878), .B(n52533), .Z(n55772) );
  IV U65141 ( .A(n52534), .Z(n52539) );
  NOR U65142 ( .A(n52536), .B(n52535), .Z(n52537) );
  IV U65143 ( .A(n52537), .Z(n52538) );
  NOR U65144 ( .A(n52539), .B(n52538), .Z(n57042) );
  IV U65145 ( .A(n52540), .Z(n52542) );
  NOR U65146 ( .A(n52542), .B(n52541), .Z(n57069) );
  IV U65147 ( .A(n52543), .Z(n53844) );
  IV U65148 ( .A(n52546), .Z(n52544) );
  NOR U65149 ( .A(n53844), .B(n52544), .Z(n52550) );
  IV U65150 ( .A(n52545), .Z(n52548) );
  XOR U65151 ( .A(n52546), .B(n53844), .Z(n52547) );
  NOR U65152 ( .A(n52548), .B(n52547), .Z(n52549) );
  NOR U65153 ( .A(n52550), .B(n52549), .Z(n57050) );
  IV U65154 ( .A(n52551), .Z(n52552) );
  NOR U65155 ( .A(n52552), .B(n52554), .Z(n55780) );
  IV U65156 ( .A(n52553), .Z(n52555) );
  NOR U65157 ( .A(n52555), .B(n52554), .Z(n55783) );
  IV U65158 ( .A(n52556), .Z(n52557) );
  NOR U65159 ( .A(n52558), .B(n52557), .Z(n52563) );
  IV U65160 ( .A(n52559), .Z(n52561) );
  IV U65161 ( .A(n52560), .Z(n52565) );
  NOR U65162 ( .A(n52561), .B(n52565), .Z(n52562) );
  NOR U65163 ( .A(n52563), .B(n52562), .Z(n57012) );
  IV U65164 ( .A(n52564), .Z(n52566) );
  NOR U65165 ( .A(n52566), .B(n52565), .Z(n57014) );
  IV U65166 ( .A(n52567), .Z(n52569) );
  NOR U65167 ( .A(n52569), .B(n52568), .Z(n53821) );
  IV U65168 ( .A(n53821), .Z(n53812) );
  IV U65169 ( .A(n52570), .Z(n52571) );
  NOR U65170 ( .A(n52572), .B(n52571), .Z(n57003) );
  IV U65171 ( .A(n52573), .Z(n52575) );
  NOR U65172 ( .A(n52575), .B(n52574), .Z(n55801) );
  NOR U65173 ( .A(n57003), .B(n55801), .Z(n53810) );
  IV U65174 ( .A(n52579), .Z(n52576) );
  NOR U65175 ( .A(n52576), .B(n52577), .Z(n52584) );
  IV U65176 ( .A(n52577), .Z(n52578) );
  NOR U65177 ( .A(n52579), .B(n52578), .Z(n52582) );
  IV U65178 ( .A(n52580), .Z(n52581) );
  NOR U65179 ( .A(n52582), .B(n52581), .Z(n52583) );
  NOR U65180 ( .A(n52584), .B(n52583), .Z(n55799) );
  IV U65181 ( .A(n52585), .Z(n52587) );
  NOR U65182 ( .A(n52587), .B(n52586), .Z(n52598) );
  IV U65183 ( .A(n52588), .Z(n52590) );
  NOR U65184 ( .A(n52590), .B(n52589), .Z(n52595) );
  IV U65185 ( .A(n52591), .Z(n52592) );
  NOR U65186 ( .A(n52593), .B(n52592), .Z(n52594) );
  NOR U65187 ( .A(n52595), .B(n52594), .Z(n52596) );
  IV U65188 ( .A(n52596), .Z(n52597) );
  NOR U65189 ( .A(n52598), .B(n52597), .Z(n57022) );
  NOR U65190 ( .A(n52599), .B(n52603), .Z(n52601) );
  NOR U65191 ( .A(n52601), .B(n52600), .Z(n57020) );
  IV U65192 ( .A(n52602), .Z(n52604) );
  NOR U65193 ( .A(n52604), .B(n52603), .Z(n53808) );
  IV U65194 ( .A(n53808), .Z(n53801) );
  IV U65195 ( .A(n52605), .Z(n52608) );
  NOR U65196 ( .A(n52606), .B(n52612), .Z(n52607) );
  IV U65197 ( .A(n52607), .Z(n53791) );
  NOR U65198 ( .A(n52608), .B(n53791), .Z(n52609) );
  IV U65199 ( .A(n52609), .Z(n56987) );
  IV U65200 ( .A(n52610), .Z(n52611) );
  NOR U65201 ( .A(n52612), .B(n52611), .Z(n52617) );
  IV U65202 ( .A(n52613), .Z(n52614) );
  NOR U65203 ( .A(n52615), .B(n52614), .Z(n52616) );
  NOR U65204 ( .A(n52617), .B(n52616), .Z(n56984) );
  IV U65205 ( .A(n52618), .Z(n52621) );
  NOR U65206 ( .A(n52619), .B(n52623), .Z(n52620) );
  IV U65207 ( .A(n52620), .Z(n53774) );
  NOR U65208 ( .A(n52621), .B(n53774), .Z(n55823) );
  IV U65209 ( .A(n52622), .Z(n52624) );
  NOR U65210 ( .A(n52624), .B(n52623), .Z(n55835) );
  IV U65211 ( .A(n52625), .Z(n52630) );
  IV U65212 ( .A(n52626), .Z(n52627) );
  NOR U65213 ( .A(n52630), .B(n52627), .Z(n55837) );
  IV U65214 ( .A(n52628), .Z(n52629) );
  NOR U65215 ( .A(n52630), .B(n52629), .Z(n55836) );
  IV U65216 ( .A(n52631), .Z(n52632) );
  NOR U65217 ( .A(n53761), .B(n52632), .Z(n56957) );
  IV U65218 ( .A(n52634), .Z(n53757) );
  NOR U65219 ( .A(n52637), .B(n52636), .Z(n56942) );
  IV U65220 ( .A(n52638), .Z(n52640) );
  IV U65221 ( .A(n52639), .Z(n52644) );
  NOR U65222 ( .A(n52640), .B(n52644), .Z(n56939) );
  IV U65223 ( .A(n52641), .Z(n52642) );
  NOR U65224 ( .A(n52642), .B(n52644), .Z(n56916) );
  IV U65225 ( .A(n52643), .Z(n52645) );
  NOR U65226 ( .A(n52645), .B(n52644), .Z(n56922) );
  IV U65227 ( .A(n52646), .Z(n52647) );
  NOR U65228 ( .A(n52647), .B(n52652), .Z(n56901) );
  IV U65229 ( .A(n52648), .Z(n52649) );
  NOR U65230 ( .A(n52650), .B(n52649), .Z(n52655) );
  IV U65231 ( .A(n52651), .Z(n52653) );
  NOR U65232 ( .A(n52653), .B(n52652), .Z(n52654) );
  NOR U65233 ( .A(n52655), .B(n52654), .Z(n56899) );
  IV U65234 ( .A(n56899), .Z(n53750) );
  NOR U65235 ( .A(n53742), .B(n52656), .Z(n56906) );
  IV U65236 ( .A(n52657), .Z(n52658) );
  NOR U65237 ( .A(n53742), .B(n52658), .Z(n56909) );
  IV U65238 ( .A(n52659), .Z(n52660) );
  NOR U65239 ( .A(n52660), .B(n53732), .Z(n53736) );
  IV U65240 ( .A(n53736), .Z(n53723) );
  NOR U65241 ( .A(n52662), .B(n52661), .Z(n56877) );
  IV U65242 ( .A(n52663), .Z(n52665) );
  NOR U65243 ( .A(n52665), .B(n52664), .Z(n52670) );
  IV U65244 ( .A(n52666), .Z(n52667) );
  NOR U65245 ( .A(n52668), .B(n52667), .Z(n52669) );
  NOR U65246 ( .A(n52670), .B(n52669), .Z(n56875) );
  IV U65247 ( .A(n52671), .Z(n52672) );
  NOR U65248 ( .A(n53719), .B(n52672), .Z(n55850) );
  IV U65249 ( .A(n52673), .Z(n52674) );
  NOR U65250 ( .A(n52674), .B(n52677), .Z(n55845) );
  IV U65251 ( .A(n55845), .Z(n55849) );
  IV U65252 ( .A(n52675), .Z(n52676) );
  NOR U65253 ( .A(n52677), .B(n52676), .Z(n55853) );
  NOR U65254 ( .A(n52679), .B(n52678), .Z(n56853) );
  NOR U65255 ( .A(n56853), .B(n52680), .Z(n52681) );
  IV U65256 ( .A(n52681), .Z(n53716) );
  IV U65257 ( .A(n52685), .Z(n52683) );
  NOR U65258 ( .A(n52683), .B(n52682), .Z(n52690) );
  NOR U65259 ( .A(n52685), .B(n52684), .Z(n52688) );
  IV U65260 ( .A(n52686), .Z(n52687) );
  NOR U65261 ( .A(n52688), .B(n52687), .Z(n52689) );
  NOR U65262 ( .A(n52690), .B(n52689), .Z(n55881) );
  IV U65263 ( .A(n52691), .Z(n52692) );
  NOR U65264 ( .A(n52693), .B(n52692), .Z(n55875) );
  IV U65265 ( .A(n52694), .Z(n52695) );
  NOR U65266 ( .A(n52698), .B(n52695), .Z(n55872) );
  IV U65267 ( .A(n52696), .Z(n52700) );
  NOR U65268 ( .A(n52698), .B(n52697), .Z(n52699) );
  IV U65269 ( .A(n52699), .Z(n52702) );
  NOR U65270 ( .A(n52700), .B(n52702), .Z(n56813) );
  IV U65271 ( .A(n52701), .Z(n52703) );
  NOR U65272 ( .A(n52703), .B(n52702), .Z(n56816) );
  IV U65273 ( .A(n52704), .Z(n52706) );
  IV U65274 ( .A(n52705), .Z(n52708) );
  NOR U65275 ( .A(n52706), .B(n52708), .Z(n56808) );
  IV U65276 ( .A(n52707), .Z(n52709) );
  NOR U65277 ( .A(n52709), .B(n52708), .Z(n56805) );
  IV U65278 ( .A(n52710), .Z(n52711) );
  NOR U65279 ( .A(n53683), .B(n52711), .Z(n55885) );
  IV U65280 ( .A(n52712), .Z(n52713) );
  NOR U65281 ( .A(n52714), .B(n52713), .Z(n55882) );
  IV U65282 ( .A(n52715), .Z(n52717) );
  IV U65283 ( .A(n52718), .Z(n53670) );
  NOR U65284 ( .A(n52717), .B(n53670), .Z(n52724) );
  IV U65285 ( .A(n52716), .Z(n52722) );
  XOR U65286 ( .A(n53669), .B(n52718), .Z(n52720) );
  NOR U65287 ( .A(n52718), .B(n52717), .Z(n52719) );
  NOR U65288 ( .A(n52720), .B(n52719), .Z(n52721) );
  NOR U65289 ( .A(n52722), .B(n52721), .Z(n52723) );
  NOR U65290 ( .A(n52724), .B(n52723), .Z(n56791) );
  NOR U65291 ( .A(n52726), .B(n52725), .Z(n53677) );
  IV U65292 ( .A(n53677), .Z(n53668) );
  IV U65293 ( .A(n52727), .Z(n52728) );
  NOR U65294 ( .A(n52729), .B(n52728), .Z(n55914) );
  NOR U65295 ( .A(n55909), .B(n55914), .Z(n53654) );
  IV U65296 ( .A(n52730), .Z(n52731) );
  NOR U65297 ( .A(n52731), .B(n52733), .Z(n52738) );
  IV U65298 ( .A(n52732), .Z(n52736) );
  NOR U65299 ( .A(n52734), .B(n52733), .Z(n52735) );
  IV U65300 ( .A(n52735), .Z(n53644) );
  NOR U65301 ( .A(n52736), .B(n53644), .Z(n52737) );
  NOR U65302 ( .A(n52738), .B(n52737), .Z(n55920) );
  IV U65303 ( .A(n52739), .Z(n52740) );
  NOR U65304 ( .A(n53641), .B(n52740), .Z(n53636) );
  IV U65305 ( .A(n52741), .Z(n52744) );
  IV U65306 ( .A(n52742), .Z(n52743) );
  NOR U65307 ( .A(n52744), .B(n52743), .Z(n55929) );
  IV U65308 ( .A(n52745), .Z(n52747) );
  XOR U65309 ( .A(n52753), .B(n52754), .Z(n52746) );
  NOR U65310 ( .A(n52747), .B(n52746), .Z(n55932) );
  IV U65311 ( .A(n52748), .Z(n52749) );
  NOR U65312 ( .A(n52749), .B(n52754), .Z(n55938) );
  IV U65313 ( .A(n52750), .Z(n52752) );
  NOR U65314 ( .A(n52752), .B(n52751), .Z(n52757) );
  IV U65315 ( .A(n52753), .Z(n52755) );
  NOR U65316 ( .A(n52755), .B(n52754), .Z(n52756) );
  NOR U65317 ( .A(n52757), .B(n52756), .Z(n55961) );
  IV U65318 ( .A(n52758), .Z(n52760) );
  NOR U65319 ( .A(n52760), .B(n52759), .Z(n55953) );
  IV U65320 ( .A(n52761), .Z(n52763) );
  NOR U65321 ( .A(n52763), .B(n52762), .Z(n55965) );
  NOR U65322 ( .A(n55953), .B(n55965), .Z(n53627) );
  IV U65323 ( .A(n52764), .Z(n52766) );
  NOR U65324 ( .A(n52766), .B(n52765), .Z(n52771) );
  IV U65325 ( .A(n52767), .Z(n52769) );
  NOR U65326 ( .A(n52769), .B(n52768), .Z(n52770) );
  NOR U65327 ( .A(n52771), .B(n52770), .Z(n55968) );
  IV U65328 ( .A(n52772), .Z(n52774) );
  NOR U65329 ( .A(n52774), .B(n52773), .Z(n52775) );
  IV U65330 ( .A(n52775), .Z(n55957) );
  IV U65331 ( .A(n52776), .Z(n52777) );
  NOR U65332 ( .A(n52777), .B(n52780), .Z(n52778) );
  IV U65333 ( .A(n52778), .Z(n56753) );
  IV U65334 ( .A(n52779), .Z(n52781) );
  NOR U65335 ( .A(n52781), .B(n52780), .Z(n53625) );
  IV U65336 ( .A(n53625), .Z(n53613) );
  IV U65337 ( .A(n52782), .Z(n52783) );
  NOR U65338 ( .A(n52784), .B(n52783), .Z(n53622) );
  IV U65339 ( .A(n52785), .Z(n52786) );
  NOR U65340 ( .A(n52787), .B(n52786), .Z(n52792) );
  IV U65341 ( .A(n52788), .Z(n52794) );
  IV U65342 ( .A(n52789), .Z(n52790) );
  NOR U65343 ( .A(n52794), .B(n52790), .Z(n52791) );
  NOR U65344 ( .A(n52792), .B(n52791), .Z(n55974) );
  IV U65345 ( .A(n52793), .Z(n52795) );
  NOR U65346 ( .A(n52795), .B(n52794), .Z(n56728) );
  IV U65347 ( .A(n52796), .Z(n52797) );
  NOR U65348 ( .A(n52798), .B(n52797), .Z(n55987) );
  IV U65349 ( .A(n52799), .Z(n52801) );
  NOR U65350 ( .A(n52801), .B(n52800), .Z(n55981) );
  NOR U65351 ( .A(n55987), .B(n55981), .Z(n53573) );
  IV U65352 ( .A(n52802), .Z(n52805) );
  IV U65353 ( .A(n52803), .Z(n52804) );
  NOR U65354 ( .A(n52805), .B(n52804), .Z(n56010) );
  IV U65355 ( .A(n52806), .Z(n52808) );
  NOR U65356 ( .A(n52808), .B(n52807), .Z(n56007) );
  IV U65357 ( .A(n52809), .Z(n52812) );
  NOR U65358 ( .A(n52810), .B(n52818), .Z(n52811) );
  IV U65359 ( .A(n52811), .Z(n52814) );
  NOR U65360 ( .A(n52812), .B(n52814), .Z(n55996) );
  IV U65361 ( .A(n52813), .Z(n52815) );
  NOR U65362 ( .A(n52815), .B(n52814), .Z(n55999) );
  IV U65363 ( .A(n52816), .Z(n52817) );
  NOR U65364 ( .A(n52818), .B(n52817), .Z(n56004) );
  IV U65365 ( .A(n52819), .Z(n52822) );
  IV U65366 ( .A(n52820), .Z(n52821) );
  NOR U65367 ( .A(n52822), .B(n52821), .Z(n56682) );
  IV U65368 ( .A(n52823), .Z(n52826) );
  IV U65369 ( .A(n52824), .Z(n52825) );
  NOR U65370 ( .A(n52826), .B(n52825), .Z(n56679) );
  IV U65371 ( .A(n52827), .Z(n52831) );
  XOR U65372 ( .A(n52839), .B(n52840), .Z(n52828) );
  NOR U65373 ( .A(n52829), .B(n52828), .Z(n52830) );
  IV U65374 ( .A(n52830), .Z(n52835) );
  NOR U65375 ( .A(n52831), .B(n52835), .Z(n56702) );
  IV U65376 ( .A(n52832), .Z(n52833) );
  NOR U65377 ( .A(n52833), .B(n52840), .Z(n52838) );
  IV U65378 ( .A(n52834), .Z(n52836) );
  NOR U65379 ( .A(n52836), .B(n52835), .Z(n52837) );
  NOR U65380 ( .A(n52838), .B(n52837), .Z(n56652) );
  IV U65381 ( .A(n52839), .Z(n52841) );
  NOR U65382 ( .A(n52841), .B(n52840), .Z(n52842) );
  IV U65383 ( .A(n52842), .Z(n56656) );
  IV U65384 ( .A(n52843), .Z(n52845) );
  NOR U65385 ( .A(n52845), .B(n52844), .Z(n53565) );
  IV U65386 ( .A(n52846), .Z(n52850) );
  NOR U65387 ( .A(n52848), .B(n52847), .Z(n52849) );
  IV U65388 ( .A(n52849), .Z(n53546) );
  NOR U65389 ( .A(n52850), .B(n53546), .Z(n56662) );
  IV U65390 ( .A(n52851), .Z(n52852) );
  NOR U65391 ( .A(n52852), .B(n53541), .Z(n52857) );
  XOR U65392 ( .A(n53540), .B(n53541), .Z(n52865) );
  XOR U65393 ( .A(n52864), .B(n52865), .Z(n52855) );
  IV U65394 ( .A(n52853), .Z(n52854) );
  NOR U65395 ( .A(n52855), .B(n52854), .Z(n52856) );
  NOR U65396 ( .A(n52857), .B(n52856), .Z(n56015) );
  IV U65397 ( .A(n56015), .Z(n52862) );
  IV U65398 ( .A(n52858), .Z(n52861) );
  IV U65399 ( .A(n52859), .Z(n52860) );
  NOR U65400 ( .A(n52861), .B(n52860), .Z(n56659) );
  NOR U65401 ( .A(n52862), .B(n56659), .Z(n52863) );
  IV U65402 ( .A(n52863), .Z(n53544) );
  IV U65403 ( .A(n52864), .Z(n52866) );
  NOR U65404 ( .A(n52866), .B(n52865), .Z(n56629) );
  IV U65405 ( .A(n52867), .Z(n52868) );
  NOR U65406 ( .A(n52868), .B(n53535), .Z(n56641) );
  IV U65407 ( .A(n56641), .Z(n56639) );
  IV U65408 ( .A(n52869), .Z(n52871) );
  XOR U65409 ( .A(n53530), .B(n53531), .Z(n52870) );
  NOR U65410 ( .A(n52871), .B(n52870), .Z(n56621) );
  IV U65411 ( .A(n52872), .Z(n52873) );
  NOR U65412 ( .A(n52873), .B(n53531), .Z(n56016) );
  IV U65413 ( .A(n52874), .Z(n52876) );
  NOR U65414 ( .A(n52876), .B(n52875), .Z(n56624) );
  NOR U65415 ( .A(n56016), .B(n56624), .Z(n52877) );
  IV U65416 ( .A(n52877), .Z(n53533) );
  IV U65417 ( .A(n52878), .Z(n52881) );
  IV U65418 ( .A(n52879), .Z(n52880) );
  NOR U65419 ( .A(n52881), .B(n52880), .Z(n53519) );
  IV U65420 ( .A(n52882), .Z(n52883) );
  NOR U65421 ( .A(n52883), .B(n52892), .Z(n52887) );
  NOR U65422 ( .A(n52885), .B(n52884), .Z(n52886) );
  NOR U65423 ( .A(n52887), .B(n52886), .Z(n56603) );
  IV U65424 ( .A(n52888), .Z(n52889) );
  NOR U65425 ( .A(n52890), .B(n52889), .Z(n52895) );
  IV U65426 ( .A(n52891), .Z(n52893) );
  NOR U65427 ( .A(n52893), .B(n52892), .Z(n52894) );
  NOR U65428 ( .A(n52895), .B(n52894), .Z(n56599) );
  IV U65429 ( .A(n52896), .Z(n52897) );
  NOR U65430 ( .A(n52898), .B(n52897), .Z(n53506) );
  IV U65431 ( .A(n52899), .Z(n52900) );
  NOR U65432 ( .A(n52903), .B(n52900), .Z(n56036) );
  IV U65433 ( .A(n52901), .Z(n52902) );
  NOR U65434 ( .A(n52903), .B(n52902), .Z(n56031) );
  IV U65435 ( .A(n52904), .Z(n52907) );
  IV U65436 ( .A(n52905), .Z(n52906) );
  NOR U65437 ( .A(n52907), .B(n52906), .Z(n56028) );
  IV U65438 ( .A(n52908), .Z(n52911) );
  IV U65439 ( .A(n52909), .Z(n52910) );
  NOR U65440 ( .A(n52911), .B(n52910), .Z(n56054) );
  IV U65441 ( .A(n52912), .Z(n52913) );
  NOR U65442 ( .A(n52914), .B(n52913), .Z(n56053) );
  IV U65443 ( .A(n52915), .Z(n52916) );
  NOR U65444 ( .A(n52917), .B(n52916), .Z(n56063) );
  IV U65445 ( .A(n52918), .Z(n52921) );
  IV U65446 ( .A(n52919), .Z(n52920) );
  NOR U65447 ( .A(n52921), .B(n52920), .Z(n52922) );
  NOR U65448 ( .A(n52923), .B(n52922), .Z(n56061) );
  IV U65449 ( .A(n52924), .Z(n52925) );
  NOR U65450 ( .A(n52925), .B(n53471), .Z(n53476) );
  IV U65451 ( .A(n52926), .Z(n52927) );
  NOR U65452 ( .A(n52928), .B(n52927), .Z(n56575) );
  IV U65453 ( .A(n52929), .Z(n52933) );
  IV U65454 ( .A(n52930), .Z(n52931) );
  NOR U65455 ( .A(n52933), .B(n52931), .Z(n56089) );
  IV U65456 ( .A(n52932), .Z(n52934) );
  NOR U65457 ( .A(n52934), .B(n52933), .Z(n56562) );
  IV U65458 ( .A(n52935), .Z(n52936) );
  NOR U65459 ( .A(n52936), .B(n53426), .Z(n52941) );
  IV U65460 ( .A(n52937), .Z(n53422) );
  IV U65461 ( .A(n52938), .Z(n52939) );
  NOR U65462 ( .A(n53422), .B(n52939), .Z(n52940) );
  NOR U65463 ( .A(n52941), .B(n52940), .Z(n56086) );
  IV U65464 ( .A(n52942), .Z(n52944) );
  NOR U65465 ( .A(n52944), .B(n52943), .Z(n53419) );
  IV U65466 ( .A(n53419), .Z(n53416) );
  IV U65467 ( .A(n52948), .Z(n52945) );
  NOR U65468 ( .A(n52945), .B(n52946), .Z(n52952) );
  IV U65469 ( .A(n52946), .Z(n52947) );
  NOR U65470 ( .A(n52948), .B(n52947), .Z(n52949) );
  NOR U65471 ( .A(n52950), .B(n52949), .Z(n52951) );
  NOR U65472 ( .A(n52952), .B(n52951), .Z(n56527) );
  IV U65473 ( .A(n52953), .Z(n52954) );
  NOR U65474 ( .A(n52954), .B(n52967), .Z(n52955) );
  IV U65475 ( .A(n52955), .Z(n52956) );
  NOR U65476 ( .A(n52958), .B(n52956), .Z(n56534) );
  IV U65477 ( .A(n56534), .Z(n56532) );
  IV U65478 ( .A(n52957), .Z(n52959) );
  NOR U65479 ( .A(n52959), .B(n52958), .Z(n52960) );
  NOR U65480 ( .A(n52961), .B(n52960), .Z(n52962) );
  NOR U65481 ( .A(n52962), .B(n52967), .Z(n56513) );
  IV U65482 ( .A(n52963), .Z(n52964) );
  NOR U65483 ( .A(n52965), .B(n52964), .Z(n56095) );
  IV U65484 ( .A(n52966), .Z(n52968) );
  NOR U65485 ( .A(n52968), .B(n52967), .Z(n56510) );
  NOR U65486 ( .A(n56095), .B(n56510), .Z(n53403) );
  IV U65487 ( .A(n52969), .Z(n52970) );
  NOR U65488 ( .A(n53391), .B(n52970), .Z(n56105) );
  NOR U65489 ( .A(n52971), .B(n52976), .Z(n52972) );
  IV U65490 ( .A(n52972), .Z(n56118) );
  IV U65491 ( .A(n52973), .Z(n52974) );
  NOR U65492 ( .A(n52974), .B(n52976), .Z(n56114) );
  IV U65493 ( .A(n52975), .Z(n52977) );
  NOR U65494 ( .A(n52977), .B(n52976), .Z(n56111) );
  IV U65495 ( .A(n52978), .Z(n52979) );
  NOR U65496 ( .A(n52980), .B(n52979), .Z(n52985) );
  IV U65497 ( .A(n52981), .Z(n52983) );
  NOR U65498 ( .A(n52983), .B(n52982), .Z(n52984) );
  NOR U65499 ( .A(n52985), .B(n52984), .Z(n56487) );
  IV U65500 ( .A(n56487), .Z(n53388) );
  IV U65501 ( .A(n52986), .Z(n52988) );
  NOR U65502 ( .A(n52988), .B(n52987), .Z(n56489) );
  IV U65503 ( .A(n52991), .Z(n52999) );
  NOR U65504 ( .A(n52989), .B(n52999), .Z(n52995) );
  IV U65505 ( .A(n52989), .Z(n52990) );
  NOR U65506 ( .A(n52991), .B(n52990), .Z(n52992) );
  NOR U65507 ( .A(n52993), .B(n52992), .Z(n52994) );
  NOR U65508 ( .A(n52995), .B(n52994), .Z(n52996) );
  IV U65509 ( .A(n52996), .Z(n56138) );
  NOR U65510 ( .A(n52997), .B(n53003), .Z(n52998) );
  IV U65511 ( .A(n52998), .Z(n53000) );
  NOR U65512 ( .A(n53000), .B(n52999), .Z(n56139) );
  IV U65513 ( .A(n53001), .Z(n53002) );
  NOR U65514 ( .A(n53003), .B(n53002), .Z(n53004) );
  IV U65515 ( .A(n53004), .Z(n53005) );
  NOR U65516 ( .A(n53007), .B(n53005), .Z(n56144) );
  IV U65517 ( .A(n56144), .Z(n56140) );
  IV U65518 ( .A(n53006), .Z(n53008) );
  NOR U65519 ( .A(n53008), .B(n53007), .Z(n56121) );
  IV U65520 ( .A(n53009), .Z(n53011) );
  NOR U65521 ( .A(n53011), .B(n53010), .Z(n56130) );
  IV U65522 ( .A(n53012), .Z(n53014) );
  NOR U65523 ( .A(n53014), .B(n53013), .Z(n56124) );
  NOR U65524 ( .A(n56130), .B(n56124), .Z(n53371) );
  IV U65525 ( .A(n53021), .Z(n53015) );
  NOR U65526 ( .A(n53016), .B(n53015), .Z(n53019) );
  IV U65527 ( .A(n53017), .Z(n53018) );
  NOR U65528 ( .A(n53019), .B(n53018), .Z(n53022) );
  NOR U65529 ( .A(n53021), .B(n53020), .Z(n56163) );
  NOR U65530 ( .A(n53022), .B(n56163), .Z(n53366) );
  IV U65531 ( .A(n53023), .Z(n53025) );
  IV U65532 ( .A(n53024), .Z(n53032) );
  NOR U65533 ( .A(n53025), .B(n53032), .Z(n56155) );
  IV U65534 ( .A(n53026), .Z(n53028) );
  NOR U65535 ( .A(n53028), .B(n53027), .Z(n56158) );
  NOR U65536 ( .A(n53030), .B(n53029), .Z(n56154) );
  NOR U65537 ( .A(n56158), .B(n56154), .Z(n53360) );
  IV U65538 ( .A(n53031), .Z(n53033) );
  NOR U65539 ( .A(n53033), .B(n53032), .Z(n53355) );
  IV U65540 ( .A(n53034), .Z(n53035) );
  NOR U65541 ( .A(n53035), .B(n53040), .Z(n53331) );
  IV U65542 ( .A(n53036), .Z(n53038) );
  NOR U65543 ( .A(n53038), .B(n53037), .Z(n56456) );
  IV U65544 ( .A(n53039), .Z(n53041) );
  NOR U65545 ( .A(n53041), .B(n53040), .Z(n56457) );
  IV U65546 ( .A(n56457), .Z(n53326) );
  IV U65547 ( .A(n53042), .Z(n53044) );
  NOR U65548 ( .A(n53044), .B(n53043), .Z(n53049) );
  IV U65549 ( .A(n53045), .Z(n53046) );
  NOR U65550 ( .A(n53047), .B(n53046), .Z(n53048) );
  NOR U65551 ( .A(n53049), .B(n53048), .Z(n56168) );
  IV U65552 ( .A(n53050), .Z(n53052) );
  IV U65553 ( .A(n53051), .Z(n53315) );
  NOR U65554 ( .A(n53052), .B(n53315), .Z(n56169) );
  IV U65555 ( .A(n53053), .Z(n53055) );
  IV U65556 ( .A(n53054), .Z(n53298) );
  NOR U65557 ( .A(n53055), .B(n53298), .Z(n53305) );
  IV U65558 ( .A(n53056), .Z(n53057) );
  NOR U65559 ( .A(n53058), .B(n53057), .Z(n53059) );
  IV U65560 ( .A(n53059), .Z(n53060) );
  NOR U65561 ( .A(n53063), .B(n53060), .Z(n56176) );
  IV U65562 ( .A(n53061), .Z(n53062) );
  NOR U65563 ( .A(n53063), .B(n53062), .Z(n56192) );
  IV U65564 ( .A(n53064), .Z(n53067) );
  IV U65565 ( .A(n53065), .Z(n53066) );
  NOR U65566 ( .A(n53067), .B(n53066), .Z(n56428) );
  NOR U65567 ( .A(n56192), .B(n56428), .Z(n53068) );
  IV U65568 ( .A(n53068), .Z(n53296) );
  IV U65569 ( .A(n53069), .Z(n53071) );
  IV U65570 ( .A(n53070), .Z(n53074) );
  NOR U65571 ( .A(n53071), .B(n53074), .Z(n56187) );
  IV U65572 ( .A(n53072), .Z(n53073) );
  NOR U65573 ( .A(n53074), .B(n53073), .Z(n56185) );
  IV U65574 ( .A(n53075), .Z(n53076) );
  NOR U65575 ( .A(n53077), .B(n53076), .Z(n56198) );
  IV U65576 ( .A(n53078), .Z(n53081) );
  IV U65577 ( .A(n53079), .Z(n53080) );
  NOR U65578 ( .A(n53081), .B(n53080), .Z(n56394) );
  IV U65579 ( .A(n53082), .Z(n53083) );
  NOR U65580 ( .A(n53083), .B(n53085), .Z(n56397) );
  IV U65581 ( .A(n56397), .Z(n56401) );
  IV U65582 ( .A(n53084), .Z(n53086) );
  NOR U65583 ( .A(n53086), .B(n53085), .Z(n53087) );
  IV U65584 ( .A(n53087), .Z(n56400) );
  IV U65585 ( .A(n53088), .Z(n53089) );
  NOR U65586 ( .A(n53273), .B(n53089), .Z(n53094) );
  IV U65587 ( .A(n53090), .Z(n53091) );
  NOR U65588 ( .A(n53092), .B(n53091), .Z(n53093) );
  NOR U65589 ( .A(n53094), .B(n53093), .Z(n56207) );
  IV U65590 ( .A(n53095), .Z(n53103) );
  XOR U65591 ( .A(n53101), .B(n53103), .Z(n53098) );
  IV U65592 ( .A(n53096), .Z(n53097) );
  NOR U65593 ( .A(n53098), .B(n53097), .Z(n56209) );
  IV U65594 ( .A(n53099), .Z(n53100) );
  NOR U65595 ( .A(n53103), .B(n53100), .Z(n56220) );
  IV U65596 ( .A(n53101), .Z(n53102) );
  NOR U65597 ( .A(n53103), .B(n53102), .Z(n53108) );
  IV U65598 ( .A(n53104), .Z(n53105) );
  NOR U65599 ( .A(n53106), .B(n53105), .Z(n53107) );
  NOR U65600 ( .A(n53108), .B(n53107), .Z(n56218) );
  IV U65601 ( .A(n53112), .Z(n53110) );
  NOR U65602 ( .A(n53110), .B(n53109), .Z(n53117) );
  NOR U65603 ( .A(n53112), .B(n53111), .Z(n53115) );
  IV U65604 ( .A(n53113), .Z(n53114) );
  NOR U65605 ( .A(n53115), .B(n53114), .Z(n53116) );
  NOR U65606 ( .A(n53117), .B(n53116), .Z(n56370) );
  IV U65607 ( .A(n53118), .Z(n53119) );
  NOR U65608 ( .A(n53119), .B(n53122), .Z(n56372) );
  IV U65609 ( .A(n53120), .Z(n53121) );
  NOR U65610 ( .A(n53122), .B(n53121), .Z(n56377) );
  IV U65611 ( .A(n53123), .Z(n53124) );
  NOR U65612 ( .A(n53263), .B(n53124), .Z(n53125) );
  IV U65613 ( .A(n53125), .Z(n56226) );
  IV U65614 ( .A(n53126), .Z(n53131) );
  IV U65615 ( .A(n53127), .Z(n53128) );
  NOR U65616 ( .A(n53131), .B(n53128), .Z(n56227) );
  IV U65617 ( .A(n53129), .Z(n53130) );
  NOR U65618 ( .A(n53131), .B(n53130), .Z(n56358) );
  IV U65619 ( .A(n53132), .Z(n53135) );
  NOR U65620 ( .A(n53133), .B(n53244), .Z(n53134) );
  IV U65621 ( .A(n53134), .Z(n53256) );
  NOR U65622 ( .A(n53135), .B(n53256), .Z(n56303) );
  IV U65623 ( .A(n53136), .Z(n53137) );
  NOR U65624 ( .A(n53138), .B(n53137), .Z(n56314) );
  NOR U65625 ( .A(n53140), .B(n53139), .Z(n53222) );
  IV U65626 ( .A(n53222), .Z(n53217) );
  IV U65627 ( .A(n53141), .Z(n53143) );
  NOR U65628 ( .A(n53143), .B(n53142), .Z(n56321) );
  IV U65629 ( .A(n53144), .Z(n53145) );
  NOR U65630 ( .A(n53146), .B(n53145), .Z(n53152) );
  IV U65631 ( .A(n53147), .Z(n53150) );
  NOR U65632 ( .A(n53148), .B(n53157), .Z(n53149) );
  IV U65633 ( .A(n53149), .Z(n53154) );
  NOR U65634 ( .A(n53150), .B(n53154), .Z(n53151) );
  NOR U65635 ( .A(n53152), .B(n53151), .Z(n56279) );
  IV U65636 ( .A(n53153), .Z(n53155) );
  NOR U65637 ( .A(n53155), .B(n53154), .Z(n56281) );
  IV U65638 ( .A(n53156), .Z(n53158) );
  NOR U65639 ( .A(n53158), .B(n53157), .Z(n56339) );
  NOR U65640 ( .A(n56281), .B(n56339), .Z(n53215) );
  IV U65641 ( .A(n53159), .Z(n53160) );
  NOR U65642 ( .A(n53161), .B(n53160), .Z(n56270) );
  IV U65643 ( .A(n53162), .Z(n53164) );
  NOR U65644 ( .A(n53164), .B(n53163), .Z(n56342) );
  NOR U65645 ( .A(n56270), .B(n56342), .Z(n53214) );
  IV U65646 ( .A(n53165), .Z(n53167) );
  NOR U65647 ( .A(n53167), .B(n53166), .Z(n53209) );
  IV U65648 ( .A(n53209), .Z(n53203) );
  IV U65649 ( .A(n53168), .Z(n53171) );
  IV U65650 ( .A(n53169), .Z(n53170) );
  NOR U65651 ( .A(n53171), .B(n53170), .Z(n56232) );
  NOR U65652 ( .A(n53202), .B(n53172), .Z(n56288) );
  IV U65653 ( .A(n53173), .Z(n53174) );
  NOR U65654 ( .A(n53198), .B(n53174), .Z(n56242) );
  IV U65655 ( .A(n53175), .Z(n53176) );
  NOR U65656 ( .A(n53177), .B(n53176), .Z(n56255) );
  IV U65657 ( .A(n53178), .Z(n53179) );
  NOR U65658 ( .A(n53180), .B(n53179), .Z(n56250) );
  NOR U65659 ( .A(n56255), .B(n56250), .Z(n53181) );
  IV U65660 ( .A(n53181), .Z(n53196) );
  NOR U65661 ( .A(n53183), .B(n53182), .Z(n53185) );
  NOR U65662 ( .A(n53185), .B(n53184), .Z(n56240) );
  NOR U65663 ( .A(n53187), .B(n53186), .Z(n53188) );
  NOR U65664 ( .A(n53189), .B(n53188), .Z(n56239) );
  XOR U65665 ( .A(n56240), .B(n56239), .Z(n56259) );
  IV U65666 ( .A(n53190), .Z(n53191) );
  NOR U65667 ( .A(n53191), .B(n53193), .Z(n56260) );
  IV U65668 ( .A(n53192), .Z(n53194) );
  NOR U65669 ( .A(n53194), .B(n53193), .Z(n56254) );
  XOR U65670 ( .A(n56260), .B(n56254), .Z(n53195) );
  XOR U65671 ( .A(n56259), .B(n53195), .Z(n56251) );
  XOR U65672 ( .A(n53196), .B(n56251), .Z(n56243) );
  XOR U65673 ( .A(n56242), .B(n56243), .Z(n56247) );
  IV U65674 ( .A(n53197), .Z(n53199) );
  NOR U65675 ( .A(n53199), .B(n53198), .Z(n56245) );
  XOR U65676 ( .A(n56247), .B(n56245), .Z(n56289) );
  XOR U65677 ( .A(n56288), .B(n56289), .Z(n56287) );
  IV U65678 ( .A(n53200), .Z(n53201) );
  NOR U65679 ( .A(n53202), .B(n53201), .Z(n56285) );
  XOR U65680 ( .A(n56287), .B(n56285), .Z(n56233) );
  XOR U65681 ( .A(n56232), .B(n56233), .Z(n56235) );
  NOR U65682 ( .A(n53203), .B(n56235), .Z(n56273) );
  IV U65683 ( .A(n53204), .Z(n53205) );
  NOR U65684 ( .A(n53206), .B(n53205), .Z(n53207) );
  IV U65685 ( .A(n53207), .Z(n56236) );
  XOR U65686 ( .A(n56236), .B(n56235), .Z(n53208) );
  NOR U65687 ( .A(n53209), .B(n53208), .Z(n56272) );
  IV U65688 ( .A(n53210), .Z(n53211) );
  NOR U65689 ( .A(n53212), .B(n53211), .Z(n56271) );
  XOR U65690 ( .A(n56272), .B(n56271), .Z(n53213) );
  NOR U65691 ( .A(n56273), .B(n53213), .Z(n56343) );
  XOR U65692 ( .A(n53214), .B(n56343), .Z(n56340) );
  XOR U65693 ( .A(n53215), .B(n56340), .Z(n56278) );
  XOR U65694 ( .A(n56279), .B(n56278), .Z(n56323) );
  XOR U65695 ( .A(n56321), .B(n56323), .Z(n53216) );
  NOR U65696 ( .A(n53217), .B(n53216), .Z(n56300) );
  IV U65697 ( .A(n53218), .Z(n53220) );
  NOR U65698 ( .A(n53220), .B(n53219), .Z(n56297) );
  NOR U65699 ( .A(n56321), .B(n56297), .Z(n53221) );
  XOR U65700 ( .A(n56323), .B(n53221), .Z(n53227) );
  NOR U65701 ( .A(n53222), .B(n53227), .Z(n53223) );
  NOR U65702 ( .A(n56300), .B(n53223), .Z(n56310) );
  IV U65703 ( .A(n53224), .Z(n53229) );
  IV U65704 ( .A(n53225), .Z(n53226) );
  NOR U65705 ( .A(n53229), .B(n53226), .Z(n53237) );
  IV U65706 ( .A(n53237), .Z(n56311) );
  NOR U65707 ( .A(n56310), .B(n56311), .Z(n53239) );
  IV U65708 ( .A(n53227), .Z(n53232) );
  IV U65709 ( .A(n53228), .Z(n53230) );
  NOR U65710 ( .A(n53230), .B(n53229), .Z(n53233) );
  IV U65711 ( .A(n53233), .Z(n53231) );
  NOR U65712 ( .A(n53232), .B(n53231), .Z(n56325) );
  NOR U65713 ( .A(n56310), .B(n53233), .Z(n53234) );
  NOR U65714 ( .A(n56325), .B(n53234), .Z(n53235) );
  IV U65715 ( .A(n53235), .Z(n53236) );
  NOR U65716 ( .A(n53237), .B(n53236), .Z(n53238) );
  NOR U65717 ( .A(n53239), .B(n53238), .Z(n56315) );
  XOR U65718 ( .A(n56314), .B(n56315), .Z(n56306) );
  IV U65719 ( .A(n56306), .Z(n53247) );
  IV U65720 ( .A(n53240), .Z(n53242) );
  NOR U65721 ( .A(n53242), .B(n53241), .Z(n53252) );
  IV U65722 ( .A(n53252), .Z(n56307) );
  NOR U65723 ( .A(n53247), .B(n56307), .Z(n53254) );
  IV U65724 ( .A(n53243), .Z(n53245) );
  NOR U65725 ( .A(n53245), .B(n53244), .Z(n56313) );
  IV U65726 ( .A(n56313), .Z(n53246) );
  NOR U65727 ( .A(n53246), .B(n56315), .Z(n53249) );
  NOR U65728 ( .A(n53247), .B(n56313), .Z(n53248) );
  NOR U65729 ( .A(n53249), .B(n53248), .Z(n53250) );
  IV U65730 ( .A(n53250), .Z(n53251) );
  NOR U65731 ( .A(n53252), .B(n53251), .Z(n53253) );
  NOR U65732 ( .A(n53254), .B(n53253), .Z(n56304) );
  XOR U65733 ( .A(n56303), .B(n56304), .Z(n56354) );
  IV U65734 ( .A(n53255), .Z(n53257) );
  NOR U65735 ( .A(n53257), .B(n53256), .Z(n56352) );
  XOR U65736 ( .A(n56354), .B(n56352), .Z(n56357) );
  IV U65737 ( .A(n53258), .Z(n53260) );
  NOR U65738 ( .A(n53260), .B(n53259), .Z(n56355) );
  XOR U65739 ( .A(n56357), .B(n56355), .Z(n56359) );
  XOR U65740 ( .A(n56358), .B(n56359), .Z(n56228) );
  XOR U65741 ( .A(n56227), .B(n56228), .Z(n56225) );
  XOR U65742 ( .A(n56226), .B(n56225), .Z(n56333) );
  IV U65743 ( .A(n53261), .Z(n53262) );
  NOR U65744 ( .A(n53263), .B(n53262), .Z(n56334) );
  XOR U65745 ( .A(n56333), .B(n56334), .Z(n56381) );
  IV U65746 ( .A(n53264), .Z(n53265) );
  NOR U65747 ( .A(n53266), .B(n53265), .Z(n56330) );
  IV U65748 ( .A(n53267), .Z(n53269) );
  NOR U65749 ( .A(n53269), .B(n53268), .Z(n56380) );
  NOR U65750 ( .A(n56330), .B(n56380), .Z(n53270) );
  XOR U65751 ( .A(n56381), .B(n53270), .Z(n56378) );
  XOR U65752 ( .A(n56377), .B(n56378), .Z(n56373) );
  XOR U65753 ( .A(n56372), .B(n56373), .Z(n56371) );
  XOR U65754 ( .A(n56370), .B(n56371), .Z(n56217) );
  XOR U65755 ( .A(n56218), .B(n56217), .Z(n56221) );
  XOR U65756 ( .A(n56220), .B(n56221), .Z(n56211) );
  XOR U65757 ( .A(n56209), .B(n56211), .Z(n56208) );
  XOR U65758 ( .A(n56207), .B(n56208), .Z(n53271) );
  IV U65759 ( .A(n53271), .Z(n56215) );
  IV U65760 ( .A(n53272), .Z(n53274) );
  NOR U65761 ( .A(n53274), .B(n53273), .Z(n56214) );
  XOR U65762 ( .A(n56215), .B(n56214), .Z(n56398) );
  XOR U65763 ( .A(n56400), .B(n56398), .Z(n53275) );
  XOR U65764 ( .A(n56401), .B(n53275), .Z(n56395) );
  XOR U65765 ( .A(n56394), .B(n56395), .Z(n56196) );
  XOR U65766 ( .A(n56198), .B(n56196), .Z(n56413) );
  IV U65767 ( .A(n53278), .Z(n53276) );
  NOR U65768 ( .A(n53277), .B(n53276), .Z(n56195) );
  IV U65769 ( .A(n53277), .Z(n53279) );
  NOR U65770 ( .A(n53279), .B(n53278), .Z(n53281) );
  IV U65771 ( .A(n53280), .Z(n56414) );
  NOR U65772 ( .A(n53281), .B(n56414), .Z(n53282) );
  NOR U65773 ( .A(n56195), .B(n53282), .Z(n53283) );
  XOR U65774 ( .A(n56413), .B(n53283), .Z(n56203) );
  IV U65775 ( .A(n53286), .Z(n53284) );
  NOR U65776 ( .A(n53285), .B(n53284), .Z(n53290) );
  IV U65777 ( .A(n53285), .Z(n53287) );
  NOR U65778 ( .A(n53287), .B(n53286), .Z(n56204) );
  NOR U65779 ( .A(n53288), .B(n56204), .Z(n53289) );
  NOR U65780 ( .A(n53290), .B(n53289), .Z(n53291) );
  XOR U65781 ( .A(n56203), .B(n53291), .Z(n56426) );
  IV U65782 ( .A(n53292), .Z(n53293) );
  NOR U65783 ( .A(n53293), .B(n56425), .Z(n53294) );
  XOR U65784 ( .A(n56426), .B(n53294), .Z(n53295) );
  IV U65785 ( .A(n53295), .Z(n56429) );
  XOR U65786 ( .A(n56185), .B(n56429), .Z(n56189) );
  XOR U65787 ( .A(n56187), .B(n56189), .Z(n56193) );
  XOR U65788 ( .A(n53296), .B(n56193), .Z(n56177) );
  XOR U65789 ( .A(n56176), .B(n56177), .Z(n56179) );
  IV U65790 ( .A(n53297), .Z(n53299) );
  NOR U65791 ( .A(n53299), .B(n53298), .Z(n53300) );
  IV U65792 ( .A(n53300), .Z(n56180) );
  XOR U65793 ( .A(n56179), .B(n56180), .Z(n53301) );
  NOR U65794 ( .A(n53305), .B(n53301), .Z(n53307) );
  IV U65795 ( .A(n53302), .Z(n53303) );
  NOR U65796 ( .A(n53313), .B(n53303), .Z(n53309) );
  IV U65797 ( .A(n53309), .Z(n53304) );
  NOR U65798 ( .A(n53307), .B(n53304), .Z(n56183) );
  IV U65799 ( .A(n53305), .Z(n53306) );
  NOR U65800 ( .A(n56179), .B(n53306), .Z(n56184) );
  NOR U65801 ( .A(n56184), .B(n53307), .Z(n53308) );
  NOR U65802 ( .A(n53309), .B(n53308), .Z(n53310) );
  NOR U65803 ( .A(n56183), .B(n53310), .Z(n56438) );
  IV U65804 ( .A(n53311), .Z(n53312) );
  NOR U65805 ( .A(n53313), .B(n53312), .Z(n56441) );
  XOR U65806 ( .A(n56438), .B(n56441), .Z(n53318) );
  IV U65807 ( .A(n53314), .Z(n53316) );
  NOR U65808 ( .A(n53316), .B(n53315), .Z(n53317) );
  IV U65809 ( .A(n53317), .Z(n56443) );
  XOR U65810 ( .A(n53318), .B(n56443), .Z(n56171) );
  XOR U65811 ( .A(n56169), .B(n56171), .Z(n56175) );
  IV U65812 ( .A(n53319), .Z(n53320) );
  NOR U65813 ( .A(n53321), .B(n53320), .Z(n56170) );
  IV U65814 ( .A(n53322), .Z(n53324) );
  NOR U65815 ( .A(n53324), .B(n53323), .Z(n56173) );
  NOR U65816 ( .A(n56170), .B(n56173), .Z(n53325) );
  XOR U65817 ( .A(n56175), .B(n53325), .Z(n56166) );
  XOR U65818 ( .A(n56168), .B(n56166), .Z(n56459) );
  XOR U65819 ( .A(n53326), .B(n56459), .Z(n53327) );
  NOR U65820 ( .A(n56456), .B(n53327), .Z(n53333) );
  IV U65821 ( .A(n56456), .Z(n53328) );
  NOR U65822 ( .A(n53328), .B(n56459), .Z(n53329) );
  NOR U65823 ( .A(n53333), .B(n53329), .Z(n53330) );
  NOR U65824 ( .A(n53331), .B(n53330), .Z(n53334) );
  IV U65825 ( .A(n53331), .Z(n53332) );
  NOR U65826 ( .A(n53333), .B(n53332), .Z(n56461) );
  NOR U65827 ( .A(n53334), .B(n56461), .Z(n53335) );
  IV U65828 ( .A(n53335), .Z(n56464) );
  NOR U65829 ( .A(n53337), .B(n53336), .Z(n56463) );
  XOR U65830 ( .A(n56464), .B(n56463), .Z(n56468) );
  IV U65831 ( .A(n56468), .Z(n53341) );
  IV U65832 ( .A(n53338), .Z(n53339) );
  NOR U65833 ( .A(n53339), .B(n56472), .Z(n53352) );
  IV U65834 ( .A(n53352), .Z(n53340) );
  NOR U65835 ( .A(n53341), .B(n53340), .Z(n53342) );
  NOR U65836 ( .A(n53355), .B(n53342), .Z(n53343) );
  IV U65837 ( .A(n53343), .Z(n53354) );
  IV U65838 ( .A(n53347), .Z(n53344) );
  NOR U65839 ( .A(n53345), .B(n53344), .Z(n56462) );
  NOR U65840 ( .A(n53346), .B(n56462), .Z(n53350) );
  NOR U65841 ( .A(n53348), .B(n53347), .Z(n53349) );
  NOR U65842 ( .A(n53350), .B(n53349), .Z(n53351) );
  XOR U65843 ( .A(n53351), .B(n56468), .Z(n53356) );
  NOR U65844 ( .A(n53352), .B(n53356), .Z(n53353) );
  NOR U65845 ( .A(n53354), .B(n53353), .Z(n53358) );
  IV U65846 ( .A(n53355), .Z(n53357) );
  NOR U65847 ( .A(n53357), .B(n53356), .Z(n56153) );
  NOR U65848 ( .A(n53358), .B(n56153), .Z(n53359) );
  IV U65849 ( .A(n53359), .Z(n56159) );
  XOR U65850 ( .A(n53360), .B(n56159), .Z(n53361) );
  NOR U65851 ( .A(n56155), .B(n53361), .Z(n53364) );
  IV U65852 ( .A(n56155), .Z(n56151) );
  XOR U65853 ( .A(n56154), .B(n56159), .Z(n53362) );
  NOR U65854 ( .A(n56151), .B(n53362), .Z(n53363) );
  NOR U65855 ( .A(n53364), .B(n53363), .Z(n53365) );
  IV U65856 ( .A(n53365), .Z(n56164) );
  XOR U65857 ( .A(n53366), .B(n56164), .Z(n56134) );
  IV U65858 ( .A(n53367), .Z(n53369) );
  IV U65859 ( .A(n53368), .Z(n56131) );
  NOR U65860 ( .A(n53369), .B(n56131), .Z(n53370) );
  XOR U65861 ( .A(n56134), .B(n53370), .Z(n56125) );
  XOR U65862 ( .A(n53371), .B(n56125), .Z(n56122) );
  XOR U65863 ( .A(n56121), .B(n56122), .Z(n56145) );
  XOR U65864 ( .A(n56140), .B(n56145), .Z(n53372) );
  XOR U65865 ( .A(n56139), .B(n53372), .Z(n53373) );
  XOR U65866 ( .A(n56138), .B(n53373), .Z(n56498) );
  IV U65867 ( .A(n53374), .Z(n53378) );
  NOR U65868 ( .A(n53376), .B(n53375), .Z(n53377) );
  IV U65869 ( .A(n53377), .Z(n53384) );
  NOR U65870 ( .A(n53378), .B(n53384), .Z(n53379) );
  IV U65871 ( .A(n53379), .Z(n56497) );
  XOR U65872 ( .A(n56498), .B(n56497), .Z(n56494) );
  IV U65873 ( .A(n53380), .Z(n53381) );
  NOR U65874 ( .A(n53382), .B(n53381), .Z(n53387) );
  IV U65875 ( .A(n53383), .Z(n53385) );
  NOR U65876 ( .A(n53385), .B(n53384), .Z(n53386) );
  NOR U65877 ( .A(n53387), .B(n53386), .Z(n56495) );
  XOR U65878 ( .A(n56494), .B(n56495), .Z(n56490) );
  XOR U65879 ( .A(n56489), .B(n56490), .Z(n56488) );
  XOR U65880 ( .A(n53388), .B(n56488), .Z(n56113) );
  XOR U65881 ( .A(n56111), .B(n56113), .Z(n56115) );
  XOR U65882 ( .A(n56114), .B(n56115), .Z(n56117) );
  XOR U65883 ( .A(n56118), .B(n56117), .Z(n56104) );
  XOR U65884 ( .A(n56105), .B(n56104), .Z(n53395) );
  IV U65885 ( .A(n53389), .Z(n53393) );
  NOR U65886 ( .A(n53391), .B(n53390), .Z(n53392) );
  IV U65887 ( .A(n53392), .Z(n53400) );
  NOR U65888 ( .A(n53393), .B(n53400), .Z(n53394) );
  IV U65889 ( .A(n53394), .Z(n56101) );
  XOR U65890 ( .A(n53395), .B(n56101), .Z(n56096) );
  IV U65891 ( .A(n53396), .Z(n53397) );
  NOR U65892 ( .A(n53398), .B(n53397), .Z(n56106) );
  IV U65893 ( .A(n53399), .Z(n53401) );
  NOR U65894 ( .A(n53401), .B(n53400), .Z(n56092) );
  NOR U65895 ( .A(n56106), .B(n56092), .Z(n53402) );
  XOR U65896 ( .A(n56096), .B(n53402), .Z(n56509) );
  XOR U65897 ( .A(n53403), .B(n56509), .Z(n56515) );
  XOR U65898 ( .A(n56513), .B(n56515), .Z(n56535) );
  XOR U65899 ( .A(n56532), .B(n56535), .Z(n53407) );
  IV U65900 ( .A(n53404), .Z(n53405) );
  NOR U65901 ( .A(n53406), .B(n53405), .Z(n56533) );
  XOR U65902 ( .A(n53407), .B(n56533), .Z(n56524) );
  IV U65903 ( .A(n53408), .Z(n53410) );
  NOR U65904 ( .A(n53410), .B(n53409), .Z(n53415) );
  IV U65905 ( .A(n53411), .Z(n53412) );
  NOR U65906 ( .A(n53413), .B(n53412), .Z(n53414) );
  NOR U65907 ( .A(n53415), .B(n53414), .Z(n56525) );
  XOR U65908 ( .A(n56524), .B(n56525), .Z(n56529) );
  XOR U65909 ( .A(n56527), .B(n56529), .Z(n53417) );
  NOR U65910 ( .A(n53416), .B(n53417), .Z(n56546) );
  IV U65911 ( .A(n53417), .Z(n53418) );
  NOR U65912 ( .A(n53419), .B(n53418), .Z(n56543) );
  IV U65913 ( .A(n53420), .Z(n53421) );
  NOR U65914 ( .A(n53422), .B(n53421), .Z(n56542) );
  XOR U65915 ( .A(n56543), .B(n56542), .Z(n53423) );
  NOR U65916 ( .A(n56546), .B(n53423), .Z(n53424) );
  IV U65917 ( .A(n53424), .Z(n56085) );
  XOR U65918 ( .A(n56086), .B(n56085), .Z(n56565) );
  IV U65919 ( .A(n53433), .Z(n56567) );
  NOR U65920 ( .A(n56565), .B(n56567), .Z(n53435) );
  IV U65921 ( .A(n53425), .Z(n53427) );
  NOR U65922 ( .A(n53427), .B(n53426), .Z(n53429) );
  IV U65923 ( .A(n53429), .Z(n53428) );
  NOR U65924 ( .A(n53428), .B(n56085), .Z(n56087) );
  NOR U65925 ( .A(n56565), .B(n53429), .Z(n53430) );
  NOR U65926 ( .A(n56087), .B(n53430), .Z(n53431) );
  IV U65927 ( .A(n53431), .Z(n53432) );
  NOR U65928 ( .A(n53433), .B(n53432), .Z(n53434) );
  NOR U65929 ( .A(n53435), .B(n53434), .Z(n56563) );
  XOR U65930 ( .A(n56562), .B(n56563), .Z(n56091) );
  XOR U65931 ( .A(n56089), .B(n56091), .Z(n56576) );
  XOR U65932 ( .A(n56575), .B(n56576), .Z(n56072) );
  IV U65933 ( .A(n56072), .Z(n53442) );
  IV U65934 ( .A(n53436), .Z(n53438) );
  NOR U65935 ( .A(n53438), .B(n53437), .Z(n53447) );
  IV U65936 ( .A(n53447), .Z(n56071) );
  NOR U65937 ( .A(n53442), .B(n56071), .Z(n53449) );
  IV U65938 ( .A(n53439), .Z(n53440) );
  NOR U65939 ( .A(n53440), .B(n53451), .Z(n56574) );
  IV U65940 ( .A(n56574), .Z(n53441) );
  NOR U65941 ( .A(n53441), .B(n56576), .Z(n53444) );
  NOR U65942 ( .A(n53442), .B(n56574), .Z(n53443) );
  NOR U65943 ( .A(n53444), .B(n53443), .Z(n53445) );
  IV U65944 ( .A(n53445), .Z(n53446) );
  NOR U65945 ( .A(n53447), .B(n53446), .Z(n53448) );
  NOR U65946 ( .A(n53449), .B(n53448), .Z(n56556) );
  IV U65947 ( .A(n53450), .Z(n53454) );
  NOR U65948 ( .A(n53452), .B(n53451), .Z(n53453) );
  IV U65949 ( .A(n53453), .Z(n53463) );
  NOR U65950 ( .A(n53454), .B(n53463), .Z(n53455) );
  IV U65951 ( .A(n53455), .Z(n56555) );
  XOR U65952 ( .A(n56556), .B(n56555), .Z(n56080) );
  IV U65953 ( .A(n53456), .Z(n53457) );
  NOR U65954 ( .A(n53458), .B(n53457), .Z(n56076) );
  IV U65955 ( .A(n53459), .Z(n53461) );
  NOR U65956 ( .A(n53461), .B(n53460), .Z(n56082) );
  IV U65957 ( .A(n53462), .Z(n53464) );
  NOR U65958 ( .A(n53464), .B(n53463), .Z(n56557) );
  XOR U65959 ( .A(n56082), .B(n56557), .Z(n53465) );
  NOR U65960 ( .A(n56076), .B(n53465), .Z(n53466) );
  XOR U65961 ( .A(n56080), .B(n53466), .Z(n56070) );
  IV U65962 ( .A(n53467), .Z(n53468) );
  NOR U65963 ( .A(n53469), .B(n53468), .Z(n56079) );
  IV U65964 ( .A(n53470), .Z(n53472) );
  NOR U65965 ( .A(n53472), .B(n53471), .Z(n56068) );
  NOR U65966 ( .A(n56079), .B(n56068), .Z(n53473) );
  XOR U65967 ( .A(n56070), .B(n53473), .Z(n53477) );
  NOR U65968 ( .A(n53476), .B(n53477), .Z(n53474) );
  IV U65969 ( .A(n53474), .Z(n53475) );
  NOR U65970 ( .A(n53475), .B(n53480), .Z(n53486) );
  IV U65971 ( .A(n53476), .Z(n53481) );
  XOR U65972 ( .A(n53480), .B(n53481), .Z(n53479) );
  IV U65973 ( .A(n53477), .Z(n53478) );
  NOR U65974 ( .A(n53479), .B(n53478), .Z(n53484) );
  IV U65975 ( .A(n53480), .Z(n53482) );
  NOR U65976 ( .A(n53482), .B(n53481), .Z(n53483) );
  NOR U65977 ( .A(n53484), .B(n53483), .Z(n53485) );
  IV U65978 ( .A(n53485), .Z(n56585) );
  NOR U65979 ( .A(n53486), .B(n56585), .Z(n56060) );
  XOR U65980 ( .A(n56061), .B(n56060), .Z(n56064) );
  XOR U65981 ( .A(n56063), .B(n56064), .Z(n56050) );
  XOR U65982 ( .A(n56053), .B(n56050), .Z(n53487) );
  XOR U65983 ( .A(n56055), .B(n53487), .Z(n53488) );
  XOR U65984 ( .A(n56054), .B(n53488), .Z(n56029) );
  XOR U65985 ( .A(n56028), .B(n56029), .Z(n56032) );
  XOR U65986 ( .A(n56031), .B(n56032), .Z(n56040) );
  XOR U65987 ( .A(n56036), .B(n56040), .Z(n56045) );
  IV U65988 ( .A(n56045), .Z(n53492) );
  IV U65989 ( .A(n53489), .Z(n53490) );
  NOR U65990 ( .A(n53490), .B(n56044), .Z(n53503) );
  IV U65991 ( .A(n53503), .Z(n53491) );
  NOR U65992 ( .A(n53492), .B(n53491), .Z(n53493) );
  NOR U65993 ( .A(n53506), .B(n53493), .Z(n53494) );
  IV U65994 ( .A(n53494), .Z(n53505) );
  IV U65995 ( .A(n53498), .Z(n53495) );
  NOR U65996 ( .A(n53496), .B(n53495), .Z(n56039) );
  NOR U65997 ( .A(n53497), .B(n56039), .Z(n53501) );
  NOR U65998 ( .A(n53499), .B(n53498), .Z(n53500) );
  NOR U65999 ( .A(n53501), .B(n53500), .Z(n53502) );
  XOR U66000 ( .A(n53502), .B(n56045), .Z(n53507) );
  NOR U66001 ( .A(n53503), .B(n53507), .Z(n53504) );
  NOR U66002 ( .A(n53505), .B(n53504), .Z(n53509) );
  IV U66003 ( .A(n53506), .Z(n53508) );
  NOR U66004 ( .A(n53508), .B(n53507), .Z(n56601) );
  NOR U66005 ( .A(n53509), .B(n56601), .Z(n56598) );
  XOR U66006 ( .A(n56599), .B(n56598), .Z(n56604) );
  XOR U66007 ( .A(n56603), .B(n56604), .Z(n56606) );
  NOR U66008 ( .A(n53511), .B(n53510), .Z(n53512) );
  NOR U66009 ( .A(n53513), .B(n53512), .Z(n56605) );
  XOR U66010 ( .A(n56606), .B(n56605), .Z(n53520) );
  NOR U66011 ( .A(n53519), .B(n53520), .Z(n53514) );
  IV U66012 ( .A(n53514), .Z(n53518) );
  IV U66013 ( .A(n53515), .Z(n53516) );
  NOR U66014 ( .A(n53517), .B(n53516), .Z(n53523) );
  NOR U66015 ( .A(n53518), .B(n53523), .Z(n53529) );
  IV U66016 ( .A(n53519), .Z(n53524) );
  XOR U66017 ( .A(n53523), .B(n53524), .Z(n53522) );
  IV U66018 ( .A(n53520), .Z(n53521) );
  NOR U66019 ( .A(n53522), .B(n53521), .Z(n53527) );
  IV U66020 ( .A(n53523), .Z(n53525) );
  NOR U66021 ( .A(n53525), .B(n53524), .Z(n53526) );
  NOR U66022 ( .A(n53527), .B(n53526), .Z(n53528) );
  IV U66023 ( .A(n53528), .Z(n56616) );
  NOR U66024 ( .A(n53529), .B(n56616), .Z(n56020) );
  IV U66025 ( .A(n53530), .Z(n53532) );
  NOR U66026 ( .A(n53532), .B(n53531), .Z(n56019) );
  IV U66027 ( .A(n56019), .Z(n56017) );
  XOR U66028 ( .A(n56020), .B(n56017), .Z(n56625) );
  XOR U66029 ( .A(n53533), .B(n56625), .Z(n56622) );
  XOR U66030 ( .A(n56621), .B(n56622), .Z(n56026) );
  IV U66031 ( .A(n53534), .Z(n53536) );
  NOR U66032 ( .A(n53536), .B(n53535), .Z(n56025) );
  XOR U66033 ( .A(n56026), .B(n56025), .Z(n56643) );
  XOR U66034 ( .A(n56639), .B(n56643), .Z(n56633) );
  IV U66035 ( .A(n53537), .Z(n53539) );
  NOR U66036 ( .A(n53539), .B(n53538), .Z(n56638) );
  IV U66037 ( .A(n53540), .Z(n53542) );
  NOR U66038 ( .A(n53542), .B(n53541), .Z(n56632) );
  NOR U66039 ( .A(n56638), .B(n56632), .Z(n53543) );
  XOR U66040 ( .A(n56633), .B(n53543), .Z(n56630) );
  XOR U66041 ( .A(n56629), .B(n56630), .Z(n56661) );
  XOR U66042 ( .A(n53544), .B(n56661), .Z(n56663) );
  XOR U66043 ( .A(n56662), .B(n56663), .Z(n56666) );
  IV U66044 ( .A(n53545), .Z(n53547) );
  NOR U66045 ( .A(n53547), .B(n53546), .Z(n56665) );
  XOR U66046 ( .A(n56666), .B(n56665), .Z(n56688) );
  IV U66047 ( .A(n53550), .Z(n53548) );
  NOR U66048 ( .A(n53549), .B(n53548), .Z(n53555) );
  NOR U66049 ( .A(n53551), .B(n53550), .Z(n53552) );
  NOR U66050 ( .A(n53553), .B(n53552), .Z(n53554) );
  NOR U66051 ( .A(n53555), .B(n53554), .Z(n53556) );
  IV U66052 ( .A(n53556), .Z(n56687) );
  XOR U66053 ( .A(n56688), .B(n56687), .Z(n53564) );
  NOR U66054 ( .A(n53565), .B(n53564), .Z(n53563) );
  IV U66055 ( .A(n53563), .Z(n53560) );
  IV U66056 ( .A(n53557), .Z(n53558) );
  NOR U66057 ( .A(n53559), .B(n53558), .Z(n53561) );
  NOR U66058 ( .A(n53560), .B(n53561), .Z(n53570) );
  IV U66059 ( .A(n53561), .Z(n53562) );
  NOR U66060 ( .A(n53563), .B(n53562), .Z(n56692) );
  IV U66061 ( .A(n53564), .Z(n53567) );
  IV U66062 ( .A(n53565), .Z(n53566) );
  NOR U66063 ( .A(n53567), .B(n53566), .Z(n53568) );
  NOR U66064 ( .A(n56692), .B(n53568), .Z(n56689) );
  IV U66065 ( .A(n56689), .Z(n53569) );
  NOR U66066 ( .A(n53570), .B(n53569), .Z(n56654) );
  XOR U66067 ( .A(n56656), .B(n56654), .Z(n56653) );
  XOR U66068 ( .A(n56652), .B(n56653), .Z(n53571) );
  IV U66069 ( .A(n53571), .Z(n56704) );
  XOR U66070 ( .A(n56702), .B(n56704), .Z(n53572) );
  XOR U66071 ( .A(n56699), .B(n53572), .Z(n56680) );
  XOR U66072 ( .A(n56679), .B(n56680), .Z(n56683) );
  XOR U66073 ( .A(n56682), .B(n56683), .Z(n56006) );
  XOR U66074 ( .A(n56004), .B(n56006), .Z(n56001) );
  XOR U66075 ( .A(n55999), .B(n56001), .Z(n55998) );
  XOR U66076 ( .A(n55996), .B(n55998), .Z(n55995) );
  XOR U66077 ( .A(n55993), .B(n55995), .Z(n56009) );
  XOR U66078 ( .A(n56007), .B(n56009), .Z(n56011) );
  XOR U66079 ( .A(n56010), .B(n56011), .Z(n55989) );
  XOR U66080 ( .A(n53573), .B(n55989), .Z(n53579) );
  IV U66081 ( .A(n53574), .Z(n53576) );
  NOR U66082 ( .A(n53576), .B(n53575), .Z(n55983) );
  NOR U66083 ( .A(n53581), .B(n53577), .Z(n55990) );
  NOR U66084 ( .A(n55983), .B(n55990), .Z(n53578) );
  XOR U66085 ( .A(n53579), .B(n53578), .Z(n56726) );
  IV U66086 ( .A(n53580), .Z(n53582) );
  NOR U66087 ( .A(n53582), .B(n53581), .Z(n56725) );
  XOR U66088 ( .A(n56726), .B(n56725), .Z(n56729) );
  XOR U66089 ( .A(n56728), .B(n56729), .Z(n55973) );
  XOR U66090 ( .A(n55974), .B(n55973), .Z(n53590) );
  IV U66091 ( .A(n53583), .Z(n53584) );
  NOR U66092 ( .A(n53585), .B(n53584), .Z(n55975) );
  IV U66093 ( .A(n53586), .Z(n53587) );
  NOR U66094 ( .A(n53588), .B(n53587), .Z(n55976) );
  NOR U66095 ( .A(n55975), .B(n55976), .Z(n53589) );
  XOR U66096 ( .A(n53590), .B(n53589), .Z(n53598) );
  IV U66097 ( .A(n53591), .Z(n53592) );
  NOR U66098 ( .A(n53593), .B(n53592), .Z(n53597) );
  IV U66099 ( .A(n53594), .Z(n53595) );
  NOR U66100 ( .A(n53595), .B(n53603), .Z(n53596) );
  NOR U66101 ( .A(n53597), .B(n53596), .Z(n53599) );
  NOR U66102 ( .A(n53598), .B(n53599), .Z(n56742) );
  IV U66103 ( .A(n53598), .Z(n53601) );
  IV U66104 ( .A(n53599), .Z(n53600) );
  NOR U66105 ( .A(n53601), .B(n53600), .Z(n56735) );
  IV U66106 ( .A(n53602), .Z(n53604) );
  NOR U66107 ( .A(n53604), .B(n53603), .Z(n56734) );
  XOR U66108 ( .A(n56735), .B(n56734), .Z(n53605) );
  NOR U66109 ( .A(n56742), .B(n53605), .Z(n53611) );
  IV U66110 ( .A(n53606), .Z(n53607) );
  NOR U66111 ( .A(n53608), .B(n53607), .Z(n53609) );
  NOR U66112 ( .A(n53610), .B(n53609), .Z(n56736) );
  XOR U66113 ( .A(n53611), .B(n56736), .Z(n56745) );
  XOR U66114 ( .A(n53622), .B(n56745), .Z(n53612) );
  NOR U66115 ( .A(n53613), .B(n53612), .Z(n56755) );
  IV U66116 ( .A(n53614), .Z(n53616) );
  NOR U66117 ( .A(n53616), .B(n53615), .Z(n53617) );
  IV U66118 ( .A(n53617), .Z(n56744) );
  IV U66119 ( .A(n53618), .Z(n53620) );
  NOR U66120 ( .A(n53620), .B(n53619), .Z(n53621) );
  NOR U66121 ( .A(n53622), .B(n53621), .Z(n56746) );
  IV U66122 ( .A(n56746), .Z(n53623) );
  XOR U66123 ( .A(n53623), .B(n56745), .Z(n56743) );
  XOR U66124 ( .A(n56744), .B(n56743), .Z(n53624) );
  NOR U66125 ( .A(n53625), .B(n53624), .Z(n53626) );
  NOR U66126 ( .A(n56755), .B(n53626), .Z(n56751) );
  XOR U66127 ( .A(n56753), .B(n56751), .Z(n55956) );
  XOR U66128 ( .A(n55957), .B(n55956), .Z(n55966) );
  XOR U66129 ( .A(n55968), .B(n55966), .Z(n55954) );
  XOR U66130 ( .A(n53627), .B(n55954), .Z(n55960) );
  XOR U66131 ( .A(n55961), .B(n55960), .Z(n55939) );
  XOR U66132 ( .A(n55938), .B(n55939), .Z(n55934) );
  XOR U66133 ( .A(n55932), .B(n55934), .Z(n55931) );
  XOR U66134 ( .A(n55929), .B(n55931), .Z(n55947) );
  IV U66135 ( .A(n53628), .Z(n53629) );
  NOR U66136 ( .A(n53630), .B(n53629), .Z(n53637) );
  IV U66137 ( .A(n53631), .Z(n53632) );
  NOR U66138 ( .A(n53633), .B(n53632), .Z(n53634) );
  NOR U66139 ( .A(n53637), .B(n53634), .Z(n55948) );
  XOR U66140 ( .A(n55947), .B(n55948), .Z(n53635) );
  NOR U66141 ( .A(n53636), .B(n53635), .Z(n55944) );
  IV U66142 ( .A(n53636), .Z(n53639) );
  XOR U66143 ( .A(n53637), .B(n55947), .Z(n53638) );
  NOR U66144 ( .A(n53639), .B(n53638), .Z(n55945) );
  NOR U66145 ( .A(n55944), .B(n55945), .Z(n53648) );
  IV U66146 ( .A(n53640), .Z(n53642) );
  NOR U66147 ( .A(n53642), .B(n53641), .Z(n53647) );
  IV U66148 ( .A(n53643), .Z(n53645) );
  NOR U66149 ( .A(n53645), .B(n53644), .Z(n53646) );
  NOR U66150 ( .A(n53647), .B(n53646), .Z(n55943) );
  XOR U66151 ( .A(n53648), .B(n55943), .Z(n55919) );
  XOR U66152 ( .A(n55920), .B(n55919), .Z(n55921) );
  IV U66153 ( .A(n53649), .Z(n53650) );
  NOR U66154 ( .A(n53651), .B(n53650), .Z(n53652) );
  NOR U66155 ( .A(n53653), .B(n53652), .Z(n55922) );
  XOR U66156 ( .A(n55921), .B(n55922), .Z(n55925) );
  XOR U66157 ( .A(n55924), .B(n55925), .Z(n55915) );
  XOR U66158 ( .A(n53654), .B(n55915), .Z(n53655) );
  IV U66159 ( .A(n53655), .Z(n56783) );
  IV U66160 ( .A(n53658), .Z(n53656) );
  NOR U66161 ( .A(n53657), .B(n53656), .Z(n53664) );
  NOR U66162 ( .A(n53658), .B(n55898), .Z(n56780) );
  NOR U66163 ( .A(n53659), .B(n56780), .Z(n53660) );
  IV U66164 ( .A(n53660), .Z(n53661) );
  NOR U66165 ( .A(n53662), .B(n53661), .Z(n53663) );
  NOR U66166 ( .A(n53664), .B(n53663), .Z(n56778) );
  XOR U66167 ( .A(n56783), .B(n56778), .Z(n55892) );
  IV U66168 ( .A(n53665), .Z(n53667) );
  NOR U66169 ( .A(n53667), .B(n53666), .Z(n55890) );
  XOR U66170 ( .A(n55892), .B(n55890), .Z(n55893) );
  NOR U66171 ( .A(n53668), .B(n55893), .Z(n56796) );
  IV U66172 ( .A(n53669), .Z(n53671) );
  NOR U66173 ( .A(n53671), .B(n53670), .Z(n56793) );
  IV U66174 ( .A(n53672), .Z(n53674) );
  NOR U66175 ( .A(n53674), .B(n53673), .Z(n53675) );
  IV U66176 ( .A(n53675), .Z(n55894) );
  XOR U66177 ( .A(n55894), .B(n55893), .Z(n53676) );
  NOR U66178 ( .A(n53677), .B(n53676), .Z(n56794) );
  XOR U66179 ( .A(n56793), .B(n56794), .Z(n53678) );
  NOR U66180 ( .A(n56796), .B(n53678), .Z(n56790) );
  XOR U66181 ( .A(n56791), .B(n56790), .Z(n55906) );
  IV U66182 ( .A(n53679), .Z(n53680) );
  NOR U66183 ( .A(n53686), .B(n53680), .Z(n53681) );
  IV U66184 ( .A(n53681), .Z(n55905) );
  XOR U66185 ( .A(n55906), .B(n55905), .Z(n55902) );
  IV U66186 ( .A(n53682), .Z(n53684) );
  NOR U66187 ( .A(n53684), .B(n53683), .Z(n53689) );
  IV U66188 ( .A(n53685), .Z(n53687) );
  NOR U66189 ( .A(n53687), .B(n53686), .Z(n53688) );
  NOR U66190 ( .A(n53689), .B(n53688), .Z(n55903) );
  XOR U66191 ( .A(n55902), .B(n55903), .Z(n55884) );
  XOR U66192 ( .A(n55882), .B(n55884), .Z(n55886) );
  XOR U66193 ( .A(n55885), .B(n55886), .Z(n56807) );
  XOR U66194 ( .A(n56805), .B(n56807), .Z(n56809) );
  XOR U66195 ( .A(n56808), .B(n56809), .Z(n56818) );
  XOR U66196 ( .A(n56816), .B(n56818), .Z(n56815) );
  XOR U66197 ( .A(n56813), .B(n56815), .Z(n55874) );
  XOR U66198 ( .A(n55872), .B(n55874), .Z(n55876) );
  XOR U66199 ( .A(n55875), .B(n55876), .Z(n55880) );
  XOR U66200 ( .A(n55881), .B(n55880), .Z(n56833) );
  IV U66201 ( .A(n56833), .Z(n56830) );
  IV U66202 ( .A(n53690), .Z(n53692) );
  NOR U66203 ( .A(n53692), .B(n53691), .Z(n56831) );
  XOR U66204 ( .A(n56830), .B(n56831), .Z(n56846) );
  IV U66205 ( .A(n53693), .Z(n53694) );
  NOR U66206 ( .A(n53695), .B(n53694), .Z(n56829) );
  IV U66207 ( .A(n53696), .Z(n53697) );
  NOR U66208 ( .A(n53697), .B(n53700), .Z(n56845) );
  NOR U66209 ( .A(n56829), .B(n56845), .Z(n53698) );
  XOR U66210 ( .A(n56846), .B(n53698), .Z(n53704) );
  IV U66211 ( .A(n53704), .Z(n53703) );
  IV U66212 ( .A(n53699), .Z(n53701) );
  NOR U66213 ( .A(n53701), .B(n53700), .Z(n53705) );
  IV U66214 ( .A(n53705), .Z(n53702) );
  NOR U66215 ( .A(n53703), .B(n53702), .Z(n56849) );
  NOR U66216 ( .A(n53705), .B(n53704), .Z(n56843) );
  IV U66217 ( .A(n53706), .Z(n53708) );
  NOR U66218 ( .A(n53708), .B(n53707), .Z(n56842) );
  XOR U66219 ( .A(n56843), .B(n56842), .Z(n53709) );
  NOR U66220 ( .A(n56849), .B(n53709), .Z(n55870) );
  IV U66221 ( .A(n53710), .Z(n53711) );
  NOR U66222 ( .A(n53712), .B(n53711), .Z(n56856) );
  NOR U66223 ( .A(n55869), .B(n56856), .Z(n53713) );
  XOR U66224 ( .A(n55870), .B(n53713), .Z(n56855) );
  XOR U66225 ( .A(n53714), .B(n56855), .Z(n53715) );
  XOR U66226 ( .A(n53716), .B(n53715), .Z(n55854) );
  XOR U66227 ( .A(n55853), .B(n55854), .Z(n55848) );
  XOR U66228 ( .A(n55849), .B(n55848), .Z(n53721) );
  IV U66229 ( .A(n53717), .Z(n53718) );
  NOR U66230 ( .A(n53719), .B(n53718), .Z(n53720) );
  IV U66231 ( .A(n53720), .Z(n55846) );
  XOR U66232 ( .A(n53721), .B(n55846), .Z(n55851) );
  XOR U66233 ( .A(n55850), .B(n55851), .Z(n56876) );
  XOR U66234 ( .A(n56875), .B(n56876), .Z(n53722) );
  IV U66235 ( .A(n53722), .Z(n56878) );
  XOR U66236 ( .A(n56877), .B(n56878), .Z(n56873) );
  XOR U66237 ( .A(n56872), .B(n56873), .Z(n53728) );
  NOR U66238 ( .A(n53723), .B(n53728), .Z(n56896) );
  IV U66239 ( .A(n53724), .Z(n53725) );
  NOR U66240 ( .A(n53726), .B(n53725), .Z(n53730) );
  IV U66241 ( .A(n53730), .Z(n53727) );
  NOR U66242 ( .A(n53727), .B(n56878), .Z(n56937) );
  IV U66243 ( .A(n53728), .Z(n53729) );
  NOR U66244 ( .A(n53730), .B(n53729), .Z(n56935) );
  IV U66245 ( .A(n53731), .Z(n53733) );
  NOR U66246 ( .A(n53733), .B(n53732), .Z(n56934) );
  XOR U66247 ( .A(n56935), .B(n56934), .Z(n53734) );
  NOR U66248 ( .A(n56937), .B(n53734), .Z(n53735) );
  NOR U66249 ( .A(n53736), .B(n53735), .Z(n53737) );
  NOR U66250 ( .A(n56896), .B(n53737), .Z(n56891) );
  IV U66251 ( .A(n53738), .Z(n53740) );
  IV U66252 ( .A(n53739), .Z(n53745) );
  NOR U66253 ( .A(n53740), .B(n53745), .Z(n56892) );
  XOR U66254 ( .A(n56891), .B(n56892), .Z(n55842) );
  IV U66255 ( .A(n53741), .Z(n53743) );
  NOR U66256 ( .A(n53743), .B(n53742), .Z(n53748) );
  IV U66257 ( .A(n53744), .Z(n53746) );
  NOR U66258 ( .A(n53746), .B(n53745), .Z(n53747) );
  NOR U66259 ( .A(n53748), .B(n53747), .Z(n55844) );
  XOR U66260 ( .A(n55842), .B(n55844), .Z(n56911) );
  XOR U66261 ( .A(n56909), .B(n56911), .Z(n53749) );
  XOR U66262 ( .A(n56906), .B(n53749), .Z(n56900) );
  XOR U66263 ( .A(n53750), .B(n56900), .Z(n56902) );
  XOR U66264 ( .A(n56901), .B(n56902), .Z(n56921) );
  NOR U66265 ( .A(n53752), .B(n53751), .Z(n53753) );
  NOR U66266 ( .A(n53754), .B(n53753), .Z(n56919) );
  XOR U66267 ( .A(n56921), .B(n56919), .Z(n56923) );
  XOR U66268 ( .A(n56922), .B(n56923), .Z(n56917) );
  XOR U66269 ( .A(n56916), .B(n56917), .Z(n56940) );
  XOR U66270 ( .A(n56939), .B(n56940), .Z(n56943) );
  XOR U66271 ( .A(n56942), .B(n56943), .Z(n56953) );
  IV U66272 ( .A(n53755), .Z(n53756) );
  NOR U66273 ( .A(n53757), .B(n53756), .Z(n56951) );
  XOR U66274 ( .A(n56953), .B(n56951), .Z(n53758) );
  XOR U66275 ( .A(n56952), .B(n53758), .Z(n56959) );
  XOR U66276 ( .A(n56957), .B(n56959), .Z(n53763) );
  IV U66277 ( .A(n53759), .Z(n53760) );
  NOR U66278 ( .A(n53761), .B(n53760), .Z(n53764) );
  IV U66279 ( .A(n53764), .Z(n53762) );
  NOR U66280 ( .A(n53763), .B(n53762), .Z(n56966) );
  IV U66281 ( .A(n53763), .Z(n53765) );
  NOR U66282 ( .A(n53765), .B(n53764), .Z(n56963) );
  IV U66283 ( .A(n53766), .Z(n53768) );
  NOR U66284 ( .A(n53768), .B(n53767), .Z(n56962) );
  XOR U66285 ( .A(n56963), .B(n56962), .Z(n53769) );
  NOR U66286 ( .A(n56966), .B(n53769), .Z(n55831) );
  XOR U66287 ( .A(n55836), .B(n55831), .Z(n53770) );
  XOR U66288 ( .A(n55837), .B(n53770), .Z(n53771) );
  XOR U66289 ( .A(n55835), .B(n53771), .Z(n53772) );
  IV U66290 ( .A(n53772), .Z(n55819) );
  IV U66291 ( .A(n53773), .Z(n53775) );
  NOR U66292 ( .A(n53775), .B(n53774), .Z(n55817) );
  XOR U66293 ( .A(n55819), .B(n55817), .Z(n55824) );
  XOR U66294 ( .A(n55823), .B(n55824), .Z(n55816) );
  IV U66295 ( .A(n53776), .Z(n53779) );
  NOR U66296 ( .A(n53787), .B(n53783), .Z(n53777) );
  IV U66297 ( .A(n53777), .Z(n53778) );
  NOR U66298 ( .A(n53779), .B(n53778), .Z(n55814) );
  XOR U66299 ( .A(n55816), .B(n55814), .Z(n55829) );
  IV U66300 ( .A(n53780), .Z(n53781) );
  NOR U66301 ( .A(n53782), .B(n53781), .Z(n53789) );
  NOR U66302 ( .A(n53784), .B(n53783), .Z(n53785) );
  IV U66303 ( .A(n53785), .Z(n53786) );
  NOR U66304 ( .A(n53787), .B(n53786), .Z(n53788) );
  NOR U66305 ( .A(n53789), .B(n53788), .Z(n55828) );
  XOR U66306 ( .A(n55829), .B(n55828), .Z(n56983) );
  XOR U66307 ( .A(n56984), .B(n56983), .Z(n56986) );
  XOR U66308 ( .A(n56987), .B(n56986), .Z(n55808) );
  IV U66309 ( .A(n53790), .Z(n53792) );
  NOR U66310 ( .A(n53792), .B(n53791), .Z(n55805) );
  XOR U66311 ( .A(n55808), .B(n55805), .Z(n56978) );
  IV U66312 ( .A(n53793), .Z(n53794) );
  NOR U66313 ( .A(n53795), .B(n53794), .Z(n56977) );
  IV U66314 ( .A(n53796), .Z(n53797) );
  NOR U66315 ( .A(n53798), .B(n53797), .Z(n55809) );
  NOR U66316 ( .A(n56977), .B(n55809), .Z(n53799) );
  XOR U66317 ( .A(n56978), .B(n53799), .Z(n56997) );
  XOR U66318 ( .A(n56975), .B(n56997), .Z(n53800) );
  NOR U66319 ( .A(n53801), .B(n53800), .Z(n57000) );
  IV U66320 ( .A(n53802), .Z(n53805) );
  IV U66321 ( .A(n53803), .Z(n53804) );
  NOR U66322 ( .A(n53805), .B(n53804), .Z(n56996) );
  NOR U66323 ( .A(n56996), .B(n56975), .Z(n53806) );
  XOR U66324 ( .A(n56997), .B(n53806), .Z(n53807) );
  NOR U66325 ( .A(n53808), .B(n53807), .Z(n53809) );
  NOR U66326 ( .A(n57000), .B(n53809), .Z(n57019) );
  XOR U66327 ( .A(n57020), .B(n57019), .Z(n57023) );
  XOR U66328 ( .A(n57022), .B(n57023), .Z(n55798) );
  XOR U66329 ( .A(n55799), .B(n55798), .Z(n57005) );
  XOR U66330 ( .A(n53810), .B(n57005), .Z(n53818) );
  IV U66331 ( .A(n53818), .Z(n53811) );
  NOR U66332 ( .A(n53812), .B(n53811), .Z(n55789) );
  IV U66333 ( .A(n53813), .Z(n53815) );
  NOR U66334 ( .A(n53815), .B(n53814), .Z(n53819) );
  IV U66335 ( .A(n53819), .Z(n53817) );
  XOR U66336 ( .A(n55801), .B(n57005), .Z(n53816) );
  NOR U66337 ( .A(n53817), .B(n53816), .Z(n57007) );
  NOR U66338 ( .A(n53819), .B(n53818), .Z(n53820) );
  NOR U66339 ( .A(n57007), .B(n53820), .Z(n53826) );
  NOR U66340 ( .A(n53821), .B(n53826), .Z(n53822) );
  NOR U66341 ( .A(n55789), .B(n53822), .Z(n55793) );
  IV U66342 ( .A(n53823), .Z(n53824) );
  NOR U66343 ( .A(n53824), .B(n53837), .Z(n53833) );
  IV U66344 ( .A(n53833), .Z(n55795) );
  NOR U66345 ( .A(n55793), .B(n55795), .Z(n53835) );
  IV U66346 ( .A(n53838), .Z(n53825) );
  NOR U66347 ( .A(n53825), .B(n53837), .Z(n53829) );
  IV U66348 ( .A(n53829), .Z(n53828) );
  IV U66349 ( .A(n53826), .Z(n53827) );
  NOR U66350 ( .A(n53828), .B(n53827), .Z(n55788) );
  NOR U66351 ( .A(n55793), .B(n53829), .Z(n53830) );
  NOR U66352 ( .A(n55788), .B(n53830), .Z(n53831) );
  IV U66353 ( .A(n53831), .Z(n53832) );
  NOR U66354 ( .A(n53833), .B(n53832), .Z(n53834) );
  NOR U66355 ( .A(n53835), .B(n53834), .Z(n55792) );
  IV U66356 ( .A(n53836), .Z(n53840) );
  XOR U66357 ( .A(n53838), .B(n53837), .Z(n53839) );
  NOR U66358 ( .A(n53840), .B(n53839), .Z(n55790) );
  XOR U66359 ( .A(n55792), .B(n55790), .Z(n57016) );
  XOR U66360 ( .A(n57014), .B(n57016), .Z(n57013) );
  XOR U66361 ( .A(n57012), .B(n57013), .Z(n53841) );
  IV U66362 ( .A(n53841), .Z(n55784) );
  XOR U66363 ( .A(n55783), .B(n55784), .Z(n55782) );
  XOR U66364 ( .A(n55780), .B(n55782), .Z(n57051) );
  XOR U66365 ( .A(n57050), .B(n57051), .Z(n53860) );
  IV U66366 ( .A(n53842), .Z(n53843) );
  NOR U66367 ( .A(n53844), .B(n53843), .Z(n57052) );
  IV U66368 ( .A(n53845), .Z(n53846) );
  NOR U66369 ( .A(n53847), .B(n53846), .Z(n57034) );
  NOR U66370 ( .A(n57052), .B(n57034), .Z(n53848) );
  XOR U66371 ( .A(n53860), .B(n53848), .Z(n53863) );
  IV U66372 ( .A(n53849), .Z(n53852) );
  NOR U66373 ( .A(n53850), .B(n53859), .Z(n53851) );
  IV U66374 ( .A(n53851), .Z(n53855) );
  NOR U66375 ( .A(n53852), .B(n53855), .Z(n53868) );
  IV U66376 ( .A(n53868), .Z(n53853) );
  NOR U66377 ( .A(n53863), .B(n53853), .Z(n57066) );
  IV U66378 ( .A(n53854), .Z(n53856) );
  NOR U66379 ( .A(n53856), .B(n53855), .Z(n57061) );
  IV U66380 ( .A(n53857), .Z(n53858) );
  NOR U66381 ( .A(n53859), .B(n53858), .Z(n53865) );
  IV U66382 ( .A(n53865), .Z(n53862) );
  IV U66383 ( .A(n53860), .Z(n57053) );
  XOR U66384 ( .A(n57052), .B(n57053), .Z(n53861) );
  NOR U66385 ( .A(n53862), .B(n53861), .Z(n57037) );
  IV U66386 ( .A(n53863), .Z(n53864) );
  NOR U66387 ( .A(n53865), .B(n53864), .Z(n53866) );
  NOR U66388 ( .A(n57037), .B(n53866), .Z(n57062) );
  XOR U66389 ( .A(n57061), .B(n57062), .Z(n53867) );
  NOR U66390 ( .A(n53868), .B(n53867), .Z(n53869) );
  NOR U66391 ( .A(n57066), .B(n53869), .Z(n57072) );
  XOR U66392 ( .A(n57069), .B(n57072), .Z(n53876) );
  NOR U66393 ( .A(n53871), .B(n53870), .Z(n53872) );
  IV U66394 ( .A(n53872), .Z(n53874) );
  NOR U66395 ( .A(n53874), .B(n53873), .Z(n53875) );
  IV U66396 ( .A(n53875), .Z(n57074) );
  XOR U66397 ( .A(n53876), .B(n57074), .Z(n57046) );
  XOR U66398 ( .A(n57045), .B(n57046), .Z(n57043) );
  XOR U66399 ( .A(n57042), .B(n57043), .Z(n57093) );
  IV U66400 ( .A(n53877), .Z(n53882) );
  NOR U66401 ( .A(n53879), .B(n53878), .Z(n53880) );
  IV U66402 ( .A(n53880), .Z(n53881) );
  NOR U66403 ( .A(n53882), .B(n53881), .Z(n53883) );
  IV U66404 ( .A(n53883), .Z(n57092) );
  XOR U66405 ( .A(n57093), .B(n57092), .Z(n57089) );
  IV U66406 ( .A(n53884), .Z(n53885) );
  NOR U66407 ( .A(n53886), .B(n53885), .Z(n53891) );
  IV U66408 ( .A(n53887), .Z(n53889) );
  NOR U66409 ( .A(n53889), .B(n53888), .Z(n53890) );
  NOR U66410 ( .A(n53891), .B(n53890), .Z(n57090) );
  XOR U66411 ( .A(n57089), .B(n57090), .Z(n55773) );
  XOR U66412 ( .A(n55772), .B(n55773), .Z(n55776) );
  XOR U66413 ( .A(n55775), .B(n55776), .Z(n57085) );
  XOR U66414 ( .A(n57081), .B(n57085), .Z(n57107) );
  XOR U66415 ( .A(n53892), .B(n57107), .Z(n57100) );
  XOR U66416 ( .A(n53893), .B(n57100), .Z(n57112) );
  XOR U66417 ( .A(n57111), .B(n57112), .Z(n57113) );
  IV U66418 ( .A(n53894), .Z(n53896) );
  NOR U66419 ( .A(n53896), .B(n53895), .Z(n53897) );
  IV U66420 ( .A(n53897), .Z(n57114) );
  XOR U66421 ( .A(n57113), .B(n57114), .Z(n55753) );
  XOR U66422 ( .A(n55749), .B(n55753), .Z(n53898) );
  XOR U66423 ( .A(n55750), .B(n53898), .Z(n53907) );
  IV U66424 ( .A(n53899), .Z(n53900) );
  NOR U66425 ( .A(n53901), .B(n53900), .Z(n53906) );
  IV U66426 ( .A(n53902), .Z(n53904) );
  NOR U66427 ( .A(n53904), .B(n53903), .Z(n53905) );
  NOR U66428 ( .A(n53906), .B(n53905), .Z(n55757) );
  XOR U66429 ( .A(n53907), .B(n55757), .Z(n55765) );
  NOR U66430 ( .A(n53909), .B(n53908), .Z(n55764) );
  IV U66431 ( .A(n53910), .Z(n53911) );
  NOR U66432 ( .A(n53912), .B(n53911), .Z(n53917) );
  IV U66433 ( .A(n53913), .Z(n53914) );
  NOR U66434 ( .A(n53915), .B(n53914), .Z(n53916) );
  NOR U66435 ( .A(n53917), .B(n53916), .Z(n55760) );
  XOR U66436 ( .A(n55764), .B(n55760), .Z(n53918) );
  XOR U66437 ( .A(n55765), .B(n53918), .Z(n53919) );
  XOR U66438 ( .A(n55761), .B(n53919), .Z(n55728) );
  IV U66439 ( .A(n53920), .Z(n53922) );
  NOR U66440 ( .A(n53922), .B(n53921), .Z(n53923) );
  IV U66441 ( .A(n53923), .Z(n55730) );
  XOR U66442 ( .A(n55728), .B(n55730), .Z(n53924) );
  XOR U66443 ( .A(n55729), .B(n53924), .Z(n55739) );
  IV U66444 ( .A(n53925), .Z(n53927) );
  NOR U66445 ( .A(n53927), .B(n53926), .Z(n55735) );
  XOR U66446 ( .A(n55739), .B(n55735), .Z(n53928) );
  XOR U66447 ( .A(n55740), .B(n53928), .Z(n53929) );
  XOR U66448 ( .A(n55734), .B(n53929), .Z(n57143) );
  XOR U66449 ( .A(n57142), .B(n57143), .Z(n57151) );
  XOR U66450 ( .A(n57148), .B(n57151), .Z(n57138) );
  IV U66451 ( .A(n53930), .Z(n53931) );
  NOR U66452 ( .A(n53932), .B(n53931), .Z(n57149) );
  NOR U66453 ( .A(n53934), .B(n53933), .Z(n57139) );
  NOR U66454 ( .A(n57149), .B(n57139), .Z(n53935) );
  XOR U66455 ( .A(n57138), .B(n53935), .Z(n57131) );
  XOR U66456 ( .A(n57130), .B(n57131), .Z(n57134) );
  XOR U66457 ( .A(n57133), .B(n57134), .Z(n53936) );
  NOR U66458 ( .A(n53937), .B(n53936), .Z(n55726) );
  NOR U66459 ( .A(n53939), .B(n53938), .Z(n55723) );
  NOR U66460 ( .A(n57133), .B(n55723), .Z(n53940) );
  XOR U66461 ( .A(n57134), .B(n53940), .Z(n53941) );
  NOR U66462 ( .A(n53942), .B(n53941), .Z(n53943) );
  NOR U66463 ( .A(n55726), .B(n53943), .Z(n53944) );
  IV U66464 ( .A(n53944), .Z(n57170) );
  XOR U66465 ( .A(n53951), .B(n57170), .Z(n53945) );
  NOR U66466 ( .A(n53946), .B(n53945), .Z(n57172) );
  IV U66467 ( .A(n53947), .Z(n53949) );
  NOR U66468 ( .A(n53949), .B(n53948), .Z(n53950) );
  NOR U66469 ( .A(n53951), .B(n53950), .Z(n57169) );
  XOR U66470 ( .A(n57169), .B(n57170), .Z(n53956) );
  NOR U66471 ( .A(n53952), .B(n53956), .Z(n53953) );
  NOR U66472 ( .A(n57172), .B(n53953), .Z(n53954) );
  NOR U66473 ( .A(n53955), .B(n53954), .Z(n57168) );
  IV U66474 ( .A(n53955), .Z(n53958) );
  IV U66475 ( .A(n53956), .Z(n53957) );
  NOR U66476 ( .A(n53958), .B(n53957), .Z(n57166) );
  NOR U66477 ( .A(n57168), .B(n57166), .Z(n53962) );
  IV U66478 ( .A(n53959), .Z(n53961) );
  NOR U66479 ( .A(n53961), .B(n53960), .Z(n57163) );
  XOR U66480 ( .A(n53962), .B(n57163), .Z(n55704) );
  XOR U66481 ( .A(n53963), .B(n55704), .Z(n55711) );
  XOR U66482 ( .A(n55712), .B(n55711), .Z(n55708) );
  IV U66483 ( .A(n53964), .Z(n53966) );
  NOR U66484 ( .A(n53966), .B(n53965), .Z(n53971) );
  IV U66485 ( .A(n53967), .Z(n53968) );
  NOR U66486 ( .A(n53969), .B(n53968), .Z(n53970) );
  NOR U66487 ( .A(n53971), .B(n53970), .Z(n55709) );
  XOR U66488 ( .A(n55708), .B(n55709), .Z(n55716) );
  XOR U66489 ( .A(n55718), .B(n55716), .Z(n55694) );
  XOR U66490 ( .A(n53972), .B(n55694), .Z(n55696) );
  XOR U66491 ( .A(n55698), .B(n55696), .Z(n55700) );
  XOR U66492 ( .A(n55699), .B(n55700), .Z(n57192) );
  XOR U66493 ( .A(n57190), .B(n57192), .Z(n53973) );
  XOR U66494 ( .A(n57187), .B(n53973), .Z(n55684) );
  XOR U66495 ( .A(n53974), .B(n55684), .Z(n55690) );
  XOR U66496 ( .A(n55688), .B(n55690), .Z(n55687) );
  XOR U66497 ( .A(n53975), .B(n55687), .Z(n55682) );
  IV U66498 ( .A(n53976), .Z(n53977) );
  NOR U66499 ( .A(n53978), .B(n53977), .Z(n53979) );
  NOR U66500 ( .A(n53982), .B(n53979), .Z(n55683) );
  XOR U66501 ( .A(n55682), .B(n55683), .Z(n53980) );
  NOR U66502 ( .A(n53981), .B(n53980), .Z(n55676) );
  IV U66503 ( .A(n53981), .Z(n53984) );
  XOR U66504 ( .A(n53982), .B(n55682), .Z(n53983) );
  NOR U66505 ( .A(n53984), .B(n53983), .Z(n55677) );
  NOR U66506 ( .A(n55676), .B(n55677), .Z(n53989) );
  IV U66507 ( .A(n53989), .Z(n53985) );
  NOR U66508 ( .A(n53990), .B(n53985), .Z(n55666) );
  IV U66509 ( .A(n53986), .Z(n53988) );
  NOR U66510 ( .A(n53988), .B(n53987), .Z(n55674) );
  XOR U66511 ( .A(n53989), .B(n55674), .Z(n53992) );
  NOR U66512 ( .A(n55674), .B(n53990), .Z(n53991) );
  NOR U66513 ( .A(n53992), .B(n53991), .Z(n55664) );
  IV U66514 ( .A(n53993), .Z(n53994) );
  NOR U66515 ( .A(n53995), .B(n53994), .Z(n55663) );
  XOR U66516 ( .A(n55664), .B(n55663), .Z(n53996) );
  NOR U66517 ( .A(n55666), .B(n53996), .Z(n55669) );
  XOR U66518 ( .A(n53997), .B(n55669), .Z(n57214) );
  XOR U66519 ( .A(n57213), .B(n57214), .Z(n57212) );
  XOR U66520 ( .A(n57211), .B(n57212), .Z(n55657) );
  IV U66521 ( .A(n55657), .Z(n55655) );
  XOR U66522 ( .A(n55660), .B(n55655), .Z(n57222) );
  IV U66523 ( .A(n53998), .Z(n53999) );
  NOR U66524 ( .A(n54000), .B(n53999), .Z(n57221) );
  IV U66525 ( .A(n54001), .Z(n54003) );
  NOR U66526 ( .A(n54003), .B(n54002), .Z(n55658) );
  NOR U66527 ( .A(n57221), .B(n55658), .Z(n54004) );
  XOR U66528 ( .A(n57222), .B(n54004), .Z(n57219) );
  IV U66529 ( .A(n54005), .Z(n54006) );
  NOR U66530 ( .A(n54007), .B(n54006), .Z(n57218) );
  IV U66531 ( .A(n54008), .Z(n54009) );
  NOR U66532 ( .A(n54010), .B(n54009), .Z(n55639) );
  NOR U66533 ( .A(n57218), .B(n55639), .Z(n54011) );
  XOR U66534 ( .A(n57219), .B(n54011), .Z(n55645) );
  IV U66535 ( .A(n54012), .Z(n54014) );
  NOR U66536 ( .A(n54014), .B(n54013), .Z(n54024) );
  IV U66537 ( .A(n54024), .Z(n55647) );
  NOR U66538 ( .A(n55645), .B(n55647), .Z(n54026) );
  IV U66539 ( .A(n54015), .Z(n54016) );
  NOR U66540 ( .A(n54017), .B(n54016), .Z(n54020) );
  IV U66541 ( .A(n54020), .Z(n54019) );
  XOR U66542 ( .A(n57218), .B(n57219), .Z(n54018) );
  NOR U66543 ( .A(n54019), .B(n54018), .Z(n55641) );
  NOR U66544 ( .A(n55645), .B(n54020), .Z(n54021) );
  NOR U66545 ( .A(n55641), .B(n54021), .Z(n54022) );
  IV U66546 ( .A(n54022), .Z(n54023) );
  NOR U66547 ( .A(n54024), .B(n54023), .Z(n54025) );
  NOR U66548 ( .A(n54026), .B(n54025), .Z(n55643) );
  XOR U66549 ( .A(n55644), .B(n55643), .Z(n55650) );
  IV U66550 ( .A(n54027), .Z(n54028) );
  NOR U66551 ( .A(n54028), .B(n54029), .Z(n54038) );
  IV U66552 ( .A(n54038), .Z(n55651) );
  NOR U66553 ( .A(n55650), .B(n55651), .Z(n54040) );
  NOR U66554 ( .A(n54030), .B(n54029), .Z(n54034) );
  IV U66555 ( .A(n54034), .Z(n54033) );
  XOR U66556 ( .A(n54031), .B(n55643), .Z(n54032) );
  NOR U66557 ( .A(n54033), .B(n54032), .Z(n55654) );
  NOR U66558 ( .A(n55650), .B(n54034), .Z(n54035) );
  NOR U66559 ( .A(n55654), .B(n54035), .Z(n54036) );
  IV U66560 ( .A(n54036), .Z(n54037) );
  NOR U66561 ( .A(n54038), .B(n54037), .Z(n54039) );
  NOR U66562 ( .A(n54040), .B(n54039), .Z(n55633) );
  IV U66563 ( .A(n54041), .Z(n54042) );
  NOR U66564 ( .A(n54043), .B(n54042), .Z(n54044) );
  IV U66565 ( .A(n54044), .Z(n55635) );
  XOR U66566 ( .A(n55633), .B(n55635), .Z(n55627) );
  IV U66567 ( .A(n54045), .Z(n54048) );
  IV U66568 ( .A(n54046), .Z(n54047) );
  NOR U66569 ( .A(n54048), .B(n54047), .Z(n55626) );
  NOR U66570 ( .A(n55634), .B(n55626), .Z(n54049) );
  XOR U66571 ( .A(n55627), .B(n54049), .Z(n55624) );
  XOR U66572 ( .A(n55623), .B(n55624), .Z(n57244) );
  IV U66573 ( .A(n54050), .Z(n54052) );
  NOR U66574 ( .A(n54052), .B(n54051), .Z(n55621) );
  IV U66575 ( .A(n54053), .Z(n54054) );
  NOR U66576 ( .A(n54055), .B(n54054), .Z(n57243) );
  NOR U66577 ( .A(n55621), .B(n57243), .Z(n54056) );
  XOR U66578 ( .A(n57244), .B(n54056), .Z(n57246) );
  XOR U66579 ( .A(n57248), .B(n57246), .Z(n57249) );
  IV U66580 ( .A(n54057), .Z(n54059) );
  NOR U66581 ( .A(n54059), .B(n54058), .Z(n54060) );
  IV U66582 ( .A(n54060), .Z(n57250) );
  XOR U66583 ( .A(n57249), .B(n57250), .Z(n55614) );
  IV U66584 ( .A(n54061), .Z(n54062) );
  NOR U66585 ( .A(n54063), .B(n54062), .Z(n55610) );
  IV U66586 ( .A(n54064), .Z(n54065) );
  NOR U66587 ( .A(n54066), .B(n54065), .Z(n55618) );
  NOR U66588 ( .A(n55610), .B(n55618), .Z(n54067) );
  XOR U66589 ( .A(n55614), .B(n54067), .Z(n57284) );
  XOR U66590 ( .A(n54068), .B(n57284), .Z(n57280) );
  XOR U66591 ( .A(n57281), .B(n57280), .Z(n57274) );
  XOR U66592 ( .A(n57272), .B(n57274), .Z(n57276) );
  XOR U66593 ( .A(n57275), .B(n57276), .Z(n57271) );
  XOR U66594 ( .A(n57269), .B(n57271), .Z(n57307) );
  XOR U66595 ( .A(n57306), .B(n57307), .Z(n57305) );
  XOR U66596 ( .A(n57303), .B(n57305), .Z(n57263) );
  XOR U66597 ( .A(n54069), .B(n57263), .Z(n57265) );
  XOR U66598 ( .A(n57264), .B(n57265), .Z(n57299) );
  XOR U66599 ( .A(n57298), .B(n57299), .Z(n57296) );
  XOR U66600 ( .A(n57297), .B(n57296), .Z(n55603) );
  XOR U66601 ( .A(n55605), .B(n55603), .Z(n55598) );
  XOR U66602 ( .A(n54070), .B(n55598), .Z(n55594) );
  XOR U66603 ( .A(n55595), .B(n55594), .Z(n55593) );
  XOR U66604 ( .A(n55591), .B(n55593), .Z(n55587) );
  XOR U66605 ( .A(n55586), .B(n55587), .Z(n55585) );
  XOR U66606 ( .A(n55583), .B(n55585), .Z(n55573) );
  XOR U66607 ( .A(n55576), .B(n55573), .Z(n54071) );
  XOR U66608 ( .A(n55577), .B(n54071), .Z(n54072) );
  XOR U66609 ( .A(n55578), .B(n54072), .Z(n55552) );
  XOR U66610 ( .A(n54073), .B(n55552), .Z(n55560) );
  XOR U66611 ( .A(n55559), .B(n55560), .Z(n55554) );
  XOR U66612 ( .A(n55553), .B(n55554), .Z(n55568) );
  XOR U66613 ( .A(n55565), .B(n55568), .Z(n57333) );
  IV U66614 ( .A(n54074), .Z(n54075) );
  NOR U66615 ( .A(n54076), .B(n54075), .Z(n55564) );
  NOR U66616 ( .A(n54078), .B(n54077), .Z(n57332) );
  NOR U66617 ( .A(n55564), .B(n57332), .Z(n54079) );
  XOR U66618 ( .A(n57333), .B(n54079), .Z(n57330) );
  XOR U66619 ( .A(n57329), .B(n57330), .Z(n57351) );
  XOR U66620 ( .A(n57346), .B(n57351), .Z(n57342) );
  XOR U66621 ( .A(n54080), .B(n57342), .Z(n57339) );
  XOR U66622 ( .A(n57338), .B(n57339), .Z(n57364) );
  IV U66623 ( .A(n54081), .Z(n54083) );
  NOR U66624 ( .A(n54083), .B(n54082), .Z(n54088) );
  IV U66625 ( .A(n54084), .Z(n54086) );
  NOR U66626 ( .A(n54086), .B(n54085), .Z(n54087) );
  NOR U66627 ( .A(n54088), .B(n54087), .Z(n57363) );
  XOR U66628 ( .A(n57364), .B(n57363), .Z(n57360) );
  XOR U66629 ( .A(n57361), .B(n57360), .Z(n57386) );
  XOR U66630 ( .A(n57384), .B(n57386), .Z(n54092) );
  IV U66631 ( .A(n54089), .Z(n54090) );
  NOR U66632 ( .A(n54090), .B(n54095), .Z(n54091) );
  IV U66633 ( .A(n54091), .Z(n57388) );
  XOR U66634 ( .A(n54092), .B(n57388), .Z(n57369) );
  IV U66635 ( .A(n54093), .Z(n54094) );
  NOR U66636 ( .A(n54095), .B(n54094), .Z(n57367) );
  XOR U66637 ( .A(n57369), .B(n57367), .Z(n57371) );
  XOR U66638 ( .A(n57370), .B(n57371), .Z(n57377) );
  IV U66639 ( .A(n54096), .Z(n54097) );
  NOR U66640 ( .A(n54098), .B(n54097), .Z(n54099) );
  IV U66641 ( .A(n54099), .Z(n57379) );
  XOR U66642 ( .A(n57377), .B(n57379), .Z(n54100) );
  XOR U66643 ( .A(n57375), .B(n54100), .Z(n57403) );
  XOR U66644 ( .A(n57404), .B(n57403), .Z(n57401) );
  IV U66645 ( .A(n54101), .Z(n54102) );
  NOR U66646 ( .A(n54104), .B(n54102), .Z(n57410) );
  IV U66647 ( .A(n54103), .Z(n54106) );
  IV U66648 ( .A(n54104), .Z(n54105) );
  NOR U66649 ( .A(n54106), .B(n54105), .Z(n57400) );
  NOR U66650 ( .A(n57410), .B(n57400), .Z(n54107) );
  XOR U66651 ( .A(n57401), .B(n54107), .Z(n57399) );
  XOR U66652 ( .A(n57397), .B(n57399), .Z(n57409) );
  XOR U66653 ( .A(n57407), .B(n57409), .Z(n55531) );
  XOR U66654 ( .A(n55535), .B(n55531), .Z(n54108) );
  XOR U66655 ( .A(n55536), .B(n54108), .Z(n55549) );
  XOR U66656 ( .A(n54109), .B(n55549), .Z(n55523) );
  XOR U66657 ( .A(n55522), .B(n55523), .Z(n55526) );
  XOR U66658 ( .A(n55525), .B(n55526), .Z(n57438) );
  XOR U66659 ( .A(n57437), .B(n57438), .Z(n57441) );
  XOR U66660 ( .A(n57440), .B(n57441), .Z(n55545) );
  XOR U66661 ( .A(n55544), .B(n55545), .Z(n55541) );
  XOR U66662 ( .A(n55542), .B(n55541), .Z(n57430) );
  XOR U66663 ( .A(n57429), .B(n57430), .Z(n57433) );
  XOR U66664 ( .A(n57432), .B(n57433), .Z(n55518) );
  IV U66665 ( .A(n54110), .Z(n54112) );
  NOR U66666 ( .A(n54112), .B(n54111), .Z(n55517) );
  XOR U66667 ( .A(n55518), .B(n55517), .Z(n55516) );
  XOR U66668 ( .A(n55515), .B(n55516), .Z(n54113) );
  IV U66669 ( .A(n54113), .Z(n57467) );
  XOR U66670 ( .A(n57465), .B(n57467), .Z(n57469) );
  XOR U66671 ( .A(n57468), .B(n57469), .Z(n57455) );
  NOR U66672 ( .A(n57459), .B(n57455), .Z(n54120) );
  IV U66673 ( .A(n57455), .Z(n54114) );
  NOR U66674 ( .A(n57453), .B(n54114), .Z(n54118) );
  IV U66675 ( .A(n54115), .Z(n54123) );
  IV U66676 ( .A(n54116), .Z(n54117) );
  NOR U66677 ( .A(n54123), .B(n54117), .Z(n57451) );
  XOR U66678 ( .A(n54118), .B(n57451), .Z(n54119) );
  NOR U66679 ( .A(n54120), .B(n54119), .Z(n55506) );
  XOR U66680 ( .A(n55512), .B(n55506), .Z(n54124) );
  IV U66681 ( .A(n54121), .Z(n54122) );
  NOR U66682 ( .A(n54123), .B(n54122), .Z(n57452) );
  IV U66683 ( .A(n57452), .Z(n57457) );
  XOR U66684 ( .A(n54124), .B(n57457), .Z(n54125) );
  NOR U66685 ( .A(n55508), .B(n54125), .Z(n54129) );
  IV U66686 ( .A(n55508), .Z(n55509) );
  NOR U66687 ( .A(n55512), .B(n55506), .Z(n54126) );
  IV U66688 ( .A(n54126), .Z(n54127) );
  NOR U66689 ( .A(n55509), .B(n54127), .Z(n54128) );
  NOR U66690 ( .A(n54129), .B(n54128), .Z(n55504) );
  XOR U66691 ( .A(n55505), .B(n55504), .Z(n54130) );
  IV U66692 ( .A(n54130), .Z(n55498) );
  XOR U66693 ( .A(n55496), .B(n55498), .Z(n55500) );
  XOR U66694 ( .A(n55499), .B(n55500), .Z(n57491) );
  XOR U66695 ( .A(n57489), .B(n57491), .Z(n57493) );
  XOR U66696 ( .A(n57492), .B(n57493), .Z(n57486) );
  XOR U66697 ( .A(n54131), .B(n57486), .Z(n57484) );
  XOR U66698 ( .A(n57483), .B(n57484), .Z(n54139) );
  IV U66699 ( .A(n54139), .Z(n54132) );
  NOR U66700 ( .A(n54133), .B(n54132), .Z(n54137) );
  IV U66701 ( .A(n54140), .Z(n54135) );
  NOR U66702 ( .A(n54135), .B(n54134), .Z(n54136) );
  NOR U66703 ( .A(n54137), .B(n54136), .Z(n54138) );
  IV U66704 ( .A(n54138), .Z(n57515) );
  NOR U66705 ( .A(n54140), .B(n54139), .Z(n54141) );
  IV U66706 ( .A(n54141), .Z(n54143) );
  NOR U66707 ( .A(n54143), .B(n54142), .Z(n54144) );
  NOR U66708 ( .A(n57515), .B(n54144), .Z(n57511) );
  IV U66709 ( .A(n54145), .Z(n54147) );
  NOR U66710 ( .A(n54147), .B(n54146), .Z(n54152) );
  IV U66711 ( .A(n54148), .Z(n54149) );
  NOR U66712 ( .A(n54150), .B(n54149), .Z(n54151) );
  NOR U66713 ( .A(n54152), .B(n54151), .Z(n57509) );
  XOR U66714 ( .A(n57511), .B(n57509), .Z(n54153) );
  XOR U66715 ( .A(n57513), .B(n54153), .Z(n54154) );
  IV U66716 ( .A(n54154), .Z(n57503) );
  IV U66717 ( .A(n54155), .Z(n54156) );
  NOR U66718 ( .A(n54165), .B(n54156), .Z(n54157) );
  IV U66719 ( .A(n54157), .Z(n54158) );
  NOR U66720 ( .A(n54159), .B(n54158), .Z(n57501) );
  XOR U66721 ( .A(n57503), .B(n57501), .Z(n57533) );
  IV U66722 ( .A(n57533), .Z(n54167) );
  IV U66723 ( .A(n54160), .Z(n54161) );
  NOR U66724 ( .A(n54162), .B(n54161), .Z(n57532) );
  IV U66725 ( .A(n54163), .Z(n54164) );
  NOR U66726 ( .A(n54165), .B(n54164), .Z(n57504) );
  NOR U66727 ( .A(n57532), .B(n57504), .Z(n54166) );
  XOR U66728 ( .A(n54167), .B(n54166), .Z(n57531) );
  XOR U66729 ( .A(n57531), .B(n57530), .Z(n54171) );
  NOR U66730 ( .A(n54173), .B(n54171), .Z(n54175) );
  IV U66731 ( .A(n54176), .Z(n54172) );
  NOR U66732 ( .A(n54175), .B(n54172), .Z(n55487) );
  IV U66733 ( .A(n54173), .Z(n54174) );
  NOR U66734 ( .A(n57531), .B(n54174), .Z(n55488) );
  NOR U66735 ( .A(n55488), .B(n54175), .Z(n54184) );
  NOR U66736 ( .A(n54176), .B(n54184), .Z(n54177) );
  NOR U66737 ( .A(n55487), .B(n54177), .Z(n55489) );
  IV U66738 ( .A(n54178), .Z(n54179) );
  NOR U66739 ( .A(n54179), .B(n54194), .Z(n55490) );
  IV U66740 ( .A(n55490), .Z(n54180) );
  NOR U66741 ( .A(n55489), .B(n54180), .Z(n54192) );
  IV U66742 ( .A(n54181), .Z(n54182) );
  NOR U66743 ( .A(n54183), .B(n54182), .Z(n54187) );
  IV U66744 ( .A(n54187), .Z(n54186) );
  IV U66745 ( .A(n54184), .Z(n54185) );
  NOR U66746 ( .A(n54186), .B(n54185), .Z(n55495) );
  NOR U66747 ( .A(n55489), .B(n54187), .Z(n54188) );
  NOR U66748 ( .A(n55495), .B(n54188), .Z(n54189) );
  IV U66749 ( .A(n54189), .Z(n54190) );
  NOR U66750 ( .A(n55490), .B(n54190), .Z(n54191) );
  NOR U66751 ( .A(n54192), .B(n54191), .Z(n57526) );
  IV U66752 ( .A(n54193), .Z(n54195) );
  NOR U66753 ( .A(n54195), .B(n54194), .Z(n55491) );
  IV U66754 ( .A(n54196), .Z(n54198) );
  NOR U66755 ( .A(n54198), .B(n54197), .Z(n54199) );
  IV U66756 ( .A(n54199), .Z(n54200) );
  NOR U66757 ( .A(n54204), .B(n54200), .Z(n57525) );
  NOR U66758 ( .A(n55491), .B(n57525), .Z(n54201) );
  XOR U66759 ( .A(n57526), .B(n54201), .Z(n54202) );
  IV U66760 ( .A(n54202), .Z(n57523) );
  NOR U66761 ( .A(n54204), .B(n54203), .Z(n54205) );
  IV U66762 ( .A(n54205), .Z(n54206) );
  NOR U66763 ( .A(n54207), .B(n54206), .Z(n57522) );
  XOR U66764 ( .A(n57523), .B(n57522), .Z(n55476) );
  XOR U66765 ( .A(n55475), .B(n55476), .Z(n54208) );
  IV U66766 ( .A(n54208), .Z(n55470) );
  IV U66767 ( .A(n54209), .Z(n54211) );
  NOR U66768 ( .A(n54211), .B(n54210), .Z(n55468) );
  XOR U66769 ( .A(n55470), .B(n55468), .Z(n55471) );
  XOR U66770 ( .A(n55472), .B(n55471), .Z(n55480) );
  IV U66771 ( .A(n54212), .Z(n54213) );
  NOR U66772 ( .A(n54214), .B(n54213), .Z(n55479) );
  IV U66773 ( .A(n54215), .Z(n54217) );
  NOR U66774 ( .A(n54217), .B(n54216), .Z(n55481) );
  NOR U66775 ( .A(n55479), .B(n55481), .Z(n54218) );
  XOR U66776 ( .A(n55480), .B(n54218), .Z(n54219) );
  XOR U66777 ( .A(n54220), .B(n54219), .Z(n55450) );
  XOR U66778 ( .A(n55449), .B(n55450), .Z(n55461) );
  XOR U66779 ( .A(n55457), .B(n55461), .Z(n54221) );
  XOR U66780 ( .A(n55463), .B(n54221), .Z(n55445) );
  XOR U66781 ( .A(n54222), .B(n55445), .Z(n55432) );
  IV U66782 ( .A(n54223), .Z(n54224) );
  NOR U66783 ( .A(n54225), .B(n54224), .Z(n55441) );
  IV U66784 ( .A(n54226), .Z(n54227) );
  NOR U66785 ( .A(n54227), .B(n54234), .Z(n55431) );
  NOR U66786 ( .A(n55441), .B(n55431), .Z(n54228) );
  XOR U66787 ( .A(n55432), .B(n54228), .Z(n55439) );
  XOR U66788 ( .A(n55434), .B(n55439), .Z(n55429) );
  IV U66789 ( .A(n54229), .Z(n54230) );
  NOR U66790 ( .A(n54231), .B(n54230), .Z(n55428) );
  IV U66791 ( .A(n54232), .Z(n54233) );
  NOR U66792 ( .A(n54234), .B(n54233), .Z(n55438) );
  NOR U66793 ( .A(n55428), .B(n55438), .Z(n54235) );
  XOR U66794 ( .A(n55429), .B(n54235), .Z(n57561) );
  XOR U66795 ( .A(n57563), .B(n57561), .Z(n57565) );
  XOR U66796 ( .A(n57564), .B(n57565), .Z(n57571) );
  XOR U66797 ( .A(n57570), .B(n57571), .Z(n57575) );
  IV U66798 ( .A(n54239), .Z(n54237) );
  NOR U66799 ( .A(n54237), .B(n54236), .Z(n57569) );
  NOR U66800 ( .A(n54239), .B(n54238), .Z(n54240) );
  NOR U66801 ( .A(n54240), .B(n57576), .Z(n54241) );
  NOR U66802 ( .A(n57569), .B(n54241), .Z(n54242) );
  XOR U66803 ( .A(n57575), .B(n54242), .Z(n54243) );
  IV U66804 ( .A(n54243), .Z(n55416) );
  XOR U66805 ( .A(n55414), .B(n55416), .Z(n57588) );
  XOR U66806 ( .A(n57587), .B(n57588), .Z(n55427) );
  XOR U66807 ( .A(n54244), .B(n55427), .Z(n55418) );
  XOR U66808 ( .A(n55417), .B(n55418), .Z(n55422) );
  NOR U66809 ( .A(n54246), .B(n54245), .Z(n55420) );
  XOR U66810 ( .A(n55422), .B(n55420), .Z(n55412) );
  XOR U66811 ( .A(n55411), .B(n55412), .Z(n55408) );
  IV U66812 ( .A(n54247), .Z(n54249) );
  IV U66813 ( .A(n54248), .Z(n54253) );
  NOR U66814 ( .A(n54249), .B(n54253), .Z(n55407) );
  NOR U66815 ( .A(n55410), .B(n55407), .Z(n54250) );
  XOR U66816 ( .A(n55408), .B(n54250), .Z(n54251) );
  IV U66817 ( .A(n54251), .Z(n55396) );
  IV U66818 ( .A(n54252), .Z(n54254) );
  NOR U66819 ( .A(n54254), .B(n54253), .Z(n55393) );
  XOR U66820 ( .A(n55396), .B(n55393), .Z(n55387) );
  XOR U66821 ( .A(n54255), .B(n55387), .Z(n55383) );
  XOR U66822 ( .A(n55385), .B(n55383), .Z(n55403) );
  XOR U66823 ( .A(n55402), .B(n55403), .Z(n54256) );
  XOR U66824 ( .A(n55399), .B(n54256), .Z(n55367) );
  XOR U66825 ( .A(n55366), .B(n55367), .Z(n57619) );
  XOR U66826 ( .A(n54257), .B(n57619), .Z(n55373) );
  IV U66827 ( .A(n54258), .Z(n54260) );
  NOR U66828 ( .A(n54260), .B(n54259), .Z(n54261) );
  IV U66829 ( .A(n54261), .Z(n57617) );
  IV U66830 ( .A(n54262), .Z(n54264) );
  NOR U66831 ( .A(n54264), .B(n54263), .Z(n55378) );
  XOR U66832 ( .A(n57617), .B(n55378), .Z(n54265) );
  XOR U66833 ( .A(n55373), .B(n54265), .Z(n54266) );
  NOR U66834 ( .A(n55375), .B(n54266), .Z(n54270) );
  IV U66835 ( .A(n55375), .Z(n55376) );
  NOR U66836 ( .A(n55378), .B(n55376), .Z(n54267) );
  IV U66837 ( .A(n54267), .Z(n54268) );
  NOR U66838 ( .A(n55373), .B(n54268), .Z(n54269) );
  NOR U66839 ( .A(n54270), .B(n54269), .Z(n55351) );
  XOR U66840 ( .A(n55350), .B(n55351), .Z(n55355) );
  XOR U66841 ( .A(n55353), .B(n55355), .Z(n55359) );
  IV U66842 ( .A(n55359), .Z(n55361) );
  IV U66843 ( .A(n54271), .Z(n54273) );
  NOR U66844 ( .A(n54273), .B(n54272), .Z(n55360) );
  IV U66845 ( .A(n54274), .Z(n54275) );
  NOR U66846 ( .A(n54276), .B(n54275), .Z(n54282) );
  NOR U66847 ( .A(n54278), .B(n54277), .Z(n54279) );
  NOR U66848 ( .A(n54280), .B(n54279), .Z(n54281) );
  NOR U66849 ( .A(n54282), .B(n54281), .Z(n55363) );
  XOR U66850 ( .A(n55360), .B(n55363), .Z(n54283) );
  XOR U66851 ( .A(n55361), .B(n54283), .Z(n57609) );
  XOR U66852 ( .A(n57608), .B(n57609), .Z(n57612) );
  XOR U66853 ( .A(n57611), .B(n57612), .Z(n55344) );
  IV U66854 ( .A(n54284), .Z(n54285) );
  NOR U66855 ( .A(n54292), .B(n54285), .Z(n54286) );
  IV U66856 ( .A(n54286), .Z(n55346) );
  XOR U66857 ( .A(n55344), .B(n55346), .Z(n54287) );
  XOR U66858 ( .A(n55345), .B(n54287), .Z(n54299) );
  NOR U66859 ( .A(n54289), .B(n54288), .Z(n54294) );
  IV U66860 ( .A(n54290), .Z(n54291) );
  NOR U66861 ( .A(n54292), .B(n54291), .Z(n54293) );
  NOR U66862 ( .A(n54294), .B(n54293), .Z(n55340) );
  IV U66863 ( .A(n55340), .Z(n54295) );
  NOR U66864 ( .A(n54299), .B(n54295), .Z(n54298) );
  IV U66865 ( .A(n54296), .Z(n54297) );
  NOR U66866 ( .A(n54298), .B(n54297), .Z(n55341) );
  IV U66867 ( .A(n54299), .Z(n55339) );
  XOR U66868 ( .A(n55340), .B(n55339), .Z(n54305) );
  NOR U66869 ( .A(n54305), .B(n54300), .Z(n54301) );
  NOR U66870 ( .A(n55341), .B(n54301), .Z(n54302) );
  IV U66871 ( .A(n54302), .Z(n54308) );
  NOR U66872 ( .A(n54303), .B(n54308), .Z(n55337) );
  IV U66873 ( .A(n54304), .Z(n54307) );
  IV U66874 ( .A(n54305), .Z(n54306) );
  NOR U66875 ( .A(n54307), .B(n54306), .Z(n55338) );
  NOR U66876 ( .A(n55338), .B(n54308), .Z(n54309) );
  NOR U66877 ( .A(n54310), .B(n54309), .Z(n54311) );
  NOR U66878 ( .A(n55337), .B(n54311), .Z(n57642) );
  NOR U66879 ( .A(n54313), .B(n54312), .Z(n54314) );
  IV U66880 ( .A(n54314), .Z(n57643) );
  XOR U66881 ( .A(n57642), .B(n57643), .Z(n54315) );
  XOR U66882 ( .A(n57644), .B(n54315), .Z(n57636) );
  XOR U66883 ( .A(n54316), .B(n57636), .Z(n57637) );
  XOR U66884 ( .A(n57638), .B(n57637), .Z(n55332) );
  NOR U66885 ( .A(n55333), .B(n54317), .Z(n55313) );
  XOR U66886 ( .A(n55332), .B(n55313), .Z(n55311) );
  IV U66887 ( .A(n54318), .Z(n54320) );
  NOR U66888 ( .A(n54320), .B(n54319), .Z(n55334) );
  IV U66889 ( .A(n54321), .Z(n54323) );
  NOR U66890 ( .A(n54323), .B(n54322), .Z(n55310) );
  NOR U66891 ( .A(n55334), .B(n55310), .Z(n54324) );
  XOR U66892 ( .A(n55311), .B(n54324), .Z(n55317) );
  XOR U66893 ( .A(n55319), .B(n55317), .Z(n55321) );
  XOR U66894 ( .A(n55320), .B(n55321), .Z(n55327) );
  IV U66895 ( .A(n54325), .Z(n54327) );
  NOR U66896 ( .A(n54327), .B(n54326), .Z(n55326) );
  IV U66897 ( .A(n55326), .Z(n55325) );
  XOR U66898 ( .A(n55327), .B(n55325), .Z(n54333) );
  IV U66899 ( .A(n54328), .Z(n54329) );
  NOR U66900 ( .A(n54329), .B(n54335), .Z(n54330) );
  IV U66901 ( .A(n54330), .Z(n54331) );
  NOR U66902 ( .A(n54336), .B(n54331), .Z(n54332) );
  IV U66903 ( .A(n54332), .Z(n55328) );
  XOR U66904 ( .A(n54333), .B(n55328), .Z(n55300) );
  IV U66905 ( .A(n54334), .Z(n54339) );
  NOR U66906 ( .A(n54336), .B(n54335), .Z(n54337) );
  IV U66907 ( .A(n54337), .Z(n54338) );
  NOR U66908 ( .A(n54339), .B(n54338), .Z(n55298) );
  XOR U66909 ( .A(n55300), .B(n55298), .Z(n55302) );
  XOR U66910 ( .A(n55301), .B(n55302), .Z(n55289) );
  XOR U66911 ( .A(n55290), .B(n55289), .Z(n54340) );
  IV U66912 ( .A(n54340), .Z(n55294) );
  XOR U66913 ( .A(n55293), .B(n55294), .Z(n55292) );
  XOR U66914 ( .A(n54341), .B(n55292), .Z(n55276) );
  IV U66915 ( .A(n54342), .Z(n54344) );
  NOR U66916 ( .A(n54344), .B(n54343), .Z(n54345) );
  IV U66917 ( .A(n54345), .Z(n55275) );
  XOR U66918 ( .A(n55276), .B(n55275), .Z(n55272) );
  IV U66919 ( .A(n54346), .Z(n54348) );
  NOR U66920 ( .A(n54348), .B(n54347), .Z(n54349) );
  NOR U66921 ( .A(n54350), .B(n54349), .Z(n55273) );
  XOR U66922 ( .A(n55272), .B(n55273), .Z(n55286) );
  XOR U66923 ( .A(n55284), .B(n55286), .Z(n54351) );
  XOR U66924 ( .A(n54352), .B(n54351), .Z(n57678) );
  XOR U66925 ( .A(n57677), .B(n57678), .Z(n57681) );
  XOR U66926 ( .A(n57680), .B(n57681), .Z(n57670) );
  XOR U66927 ( .A(n57669), .B(n57670), .Z(n57673) );
  XOR U66928 ( .A(n57672), .B(n57673), .Z(n57690) );
  IV U66929 ( .A(n54353), .Z(n54357) );
  NOR U66930 ( .A(n54355), .B(n54354), .Z(n54356) );
  IV U66931 ( .A(n54356), .Z(n54359) );
  NOR U66932 ( .A(n54357), .B(n54359), .Z(n57691) );
  IV U66933 ( .A(n57691), .Z(n57689) );
  XOR U66934 ( .A(n57690), .B(n57689), .Z(n54362) );
  IV U66935 ( .A(n54358), .Z(n54360) );
  NOR U66936 ( .A(n54360), .B(n54359), .Z(n54361) );
  IV U66937 ( .A(n54361), .Z(n57693) );
  XOR U66938 ( .A(n54362), .B(n57693), .Z(n57703) );
  XOR U66939 ( .A(n57704), .B(n57703), .Z(n54367) );
  IV U66940 ( .A(n54363), .Z(n54365) );
  NOR U66941 ( .A(n54365), .B(n54364), .Z(n54366) );
  IV U66942 ( .A(n54366), .Z(n57701) );
  XOR U66943 ( .A(n54367), .B(n57701), .Z(n57698) );
  XOR U66944 ( .A(n57699), .B(n57698), .Z(n54368) );
  NOR U66945 ( .A(n54372), .B(n54368), .Z(n54376) );
  IV U66946 ( .A(n54369), .Z(n54371) );
  NOR U66947 ( .A(n54371), .B(n54370), .Z(n54377) );
  IV U66948 ( .A(n54372), .Z(n54373) );
  NOR U66949 ( .A(n57698), .B(n54373), .Z(n54374) );
  NOR U66950 ( .A(n54377), .B(n54374), .Z(n54375) );
  NOR U66951 ( .A(n54376), .B(n54375), .Z(n55261) );
  IV U66952 ( .A(n54376), .Z(n54378) );
  NOR U66953 ( .A(n54378), .B(n54377), .Z(n54379) );
  NOR U66954 ( .A(n55261), .B(n54379), .Z(n55257) );
  XOR U66955 ( .A(n55256), .B(n55257), .Z(n54382) );
  NOR U66956 ( .A(n54381), .B(n54380), .Z(n55259) );
  XOR U66957 ( .A(n54382), .B(n55259), .Z(n55269) );
  XOR U66958 ( .A(n55267), .B(n55269), .Z(n55266) );
  XOR U66959 ( .A(n55264), .B(n55266), .Z(n55239) );
  XOR U66960 ( .A(n55240), .B(n55239), .Z(n55242) );
  IV U66961 ( .A(n54383), .Z(n54385) );
  IV U66962 ( .A(n54384), .Z(n54387) );
  NOR U66963 ( .A(n54385), .B(n54387), .Z(n55241) );
  XOR U66964 ( .A(n55242), .B(n55241), .Z(n54389) );
  IV U66965 ( .A(n54386), .Z(n54388) );
  NOR U66966 ( .A(n54388), .B(n54387), .Z(n55245) );
  XOR U66967 ( .A(n54389), .B(n55245), .Z(n55236) );
  IV U66968 ( .A(n54390), .Z(n54391) );
  NOR U66969 ( .A(n54392), .B(n54391), .Z(n55246) );
  IV U66970 ( .A(n54393), .Z(n54395) );
  NOR U66971 ( .A(n54395), .B(n54394), .Z(n55235) );
  NOR U66972 ( .A(n55246), .B(n55235), .Z(n54396) );
  XOR U66973 ( .A(n55236), .B(n54396), .Z(n55233) );
  XOR U66974 ( .A(n55232), .B(n55233), .Z(n55220) );
  XOR U66975 ( .A(n55219), .B(n55220), .Z(n54397) );
  XOR U66976 ( .A(n55216), .B(n54397), .Z(n55228) );
  XOR U66977 ( .A(n55224), .B(n55228), .Z(n54398) );
  XOR U66978 ( .A(n55227), .B(n54398), .Z(n54400) );
  NOR U66979 ( .A(n54399), .B(n54400), .Z(n55214) );
  IV U66980 ( .A(n54400), .Z(n54401) );
  NOR U66981 ( .A(n54402), .B(n54401), .Z(n55213) );
  XOR U66982 ( .A(n55213), .B(n55211), .Z(n54403) );
  NOR U66983 ( .A(n55214), .B(n54403), .Z(n54404) );
  IV U66984 ( .A(n54404), .Z(n57730) );
  IV U66985 ( .A(n54405), .Z(n54406) );
  NOR U66986 ( .A(n54407), .B(n54406), .Z(n54408) );
  NOR U66987 ( .A(n54411), .B(n54408), .Z(n57731) );
  XOR U66988 ( .A(n57730), .B(n57731), .Z(n54409) );
  NOR U66989 ( .A(n54410), .B(n54409), .Z(n55208) );
  IV U66990 ( .A(n54410), .Z(n54413) );
  XOR U66991 ( .A(n54411), .B(n57730), .Z(n54412) );
  NOR U66992 ( .A(n54413), .B(n54412), .Z(n55209) );
  NOR U66993 ( .A(n55208), .B(n55209), .Z(n54418) );
  IV U66994 ( .A(n54414), .Z(n54416) );
  NOR U66995 ( .A(n54416), .B(n54415), .Z(n54417) );
  IV U66996 ( .A(n54417), .Z(n55207) );
  XOR U66997 ( .A(n54418), .B(n55207), .Z(n57787) );
  NOR U66998 ( .A(n57785), .B(n57787), .Z(n54425) );
  IV U66999 ( .A(n57787), .Z(n57781) );
  NOR U67000 ( .A(n57780), .B(n57781), .Z(n54423) );
  IV U67001 ( .A(n54419), .Z(n54422) );
  IV U67002 ( .A(n54420), .Z(n54421) );
  NOR U67003 ( .A(n54422), .B(n54421), .Z(n57779) );
  XOR U67004 ( .A(n54423), .B(n57779), .Z(n54424) );
  NOR U67005 ( .A(n54425), .B(n54424), .Z(n54426) );
  XOR U67006 ( .A(n57783), .B(n54426), .Z(n57760) );
  XOR U67007 ( .A(n57759), .B(n57760), .Z(n57735) );
  XOR U67008 ( .A(n57737), .B(n57735), .Z(n54427) );
  XOR U67009 ( .A(n57738), .B(n54427), .Z(n57743) );
  XOR U67010 ( .A(n57742), .B(n57743), .Z(n57740) );
  XOR U67011 ( .A(n57739), .B(n57740), .Z(n57754) );
  XOR U67012 ( .A(n57753), .B(n57754), .Z(n57758) );
  NOR U67013 ( .A(n54429), .B(n54428), .Z(n54435) );
  IV U67014 ( .A(n54429), .Z(n54430) );
  NOR U67015 ( .A(n54431), .B(n54430), .Z(n54432) );
  NOR U67016 ( .A(n54433), .B(n54432), .Z(n54434) );
  NOR U67017 ( .A(n54435), .B(n54434), .Z(n57756) );
  XOR U67018 ( .A(n57758), .B(n57756), .Z(n57775) );
  XOR U67019 ( .A(n57774), .B(n57775), .Z(n57798) );
  IV U67020 ( .A(n54436), .Z(n54437) );
  NOR U67021 ( .A(n54438), .B(n54437), .Z(n57771) );
  NOR U67022 ( .A(n54440), .B(n54439), .Z(n57797) );
  NOR U67023 ( .A(n57771), .B(n57797), .Z(n54441) );
  XOR U67024 ( .A(n57798), .B(n54441), .Z(n57800) );
  IV U67025 ( .A(n54442), .Z(n54443) );
  NOR U67026 ( .A(n54444), .B(n54443), .Z(n54449) );
  IV U67027 ( .A(n54445), .Z(n54446) );
  NOR U67028 ( .A(n54447), .B(n54446), .Z(n54448) );
  NOR U67029 ( .A(n54449), .B(n54448), .Z(n57801) );
  XOR U67030 ( .A(n57800), .B(n57801), .Z(n57804) );
  NOR U67031 ( .A(n54451), .B(n54450), .Z(n57803) );
  IV U67032 ( .A(n54452), .Z(n54453) );
  NOR U67033 ( .A(n54454), .B(n54453), .Z(n55204) );
  NOR U67034 ( .A(n57803), .B(n55204), .Z(n54455) );
  XOR U67035 ( .A(n57804), .B(n54455), .Z(n57823) );
  IV U67036 ( .A(n54456), .Z(n54457) );
  NOR U67037 ( .A(n54458), .B(n54457), .Z(n55203) );
  IV U67038 ( .A(n54459), .Z(n54460) );
  NOR U67039 ( .A(n54461), .B(n54460), .Z(n57822) );
  NOR U67040 ( .A(n55203), .B(n57822), .Z(n54462) );
  XOR U67041 ( .A(n57823), .B(n54462), .Z(n57826) );
  XOR U67042 ( .A(n57827), .B(n57826), .Z(n54463) );
  NOR U67043 ( .A(n54467), .B(n54463), .Z(n54471) );
  IV U67044 ( .A(n54464), .Z(n54466) );
  NOR U67045 ( .A(n54466), .B(n54465), .Z(n54473) );
  IV U67046 ( .A(n54467), .Z(n54468) );
  NOR U67047 ( .A(n57826), .B(n54468), .Z(n54469) );
  NOR U67048 ( .A(n54473), .B(n54469), .Z(n54470) );
  NOR U67049 ( .A(n54471), .B(n54470), .Z(n57850) );
  IV U67050 ( .A(n54471), .Z(n54472) );
  NOR U67051 ( .A(n54473), .B(n54472), .Z(n54474) );
  NOR U67052 ( .A(n57850), .B(n54474), .Z(n57834) );
  XOR U67053 ( .A(n57836), .B(n57834), .Z(n57841) );
  XOR U67054 ( .A(n57839), .B(n57841), .Z(n57838) );
  XOR U67055 ( .A(n57837), .B(n57838), .Z(n54475) );
  IV U67056 ( .A(n54475), .Z(n57819) );
  XOR U67057 ( .A(n57817), .B(n57819), .Z(n57816) );
  XOR U67058 ( .A(n57815), .B(n57816), .Z(n55195) );
  IV U67059 ( .A(n54476), .Z(n54477) );
  NOR U67060 ( .A(n54477), .B(n54479), .Z(n55194) );
  XOR U67061 ( .A(n55195), .B(n55194), .Z(n54481) );
  IV U67062 ( .A(n54478), .Z(n54480) );
  NOR U67063 ( .A(n54480), .B(n54479), .Z(n55190) );
  XOR U67064 ( .A(n54481), .B(n55190), .Z(n54482) );
  XOR U67065 ( .A(n55189), .B(n54482), .Z(n55185) );
  XOR U67066 ( .A(n55186), .B(n55185), .Z(n55178) );
  XOR U67067 ( .A(n55177), .B(n55178), .Z(n54483) );
  XOR U67068 ( .A(n54484), .B(n54483), .Z(n55173) );
  XOR U67069 ( .A(n54491), .B(n55173), .Z(n54485) );
  NOR U67070 ( .A(n54486), .B(n54485), .Z(n55175) );
  IV U67071 ( .A(n54487), .Z(n54489) );
  NOR U67072 ( .A(n54489), .B(n54488), .Z(n54490) );
  NOR U67073 ( .A(n54491), .B(n54490), .Z(n55172) );
  XOR U67074 ( .A(n55173), .B(n55172), .Z(n54492) );
  NOR U67075 ( .A(n54493), .B(n54492), .Z(n54494) );
  NOR U67076 ( .A(n55175), .B(n54494), .Z(n57867) );
  XOR U67077 ( .A(n57869), .B(n57867), .Z(n57865) );
  XOR U67078 ( .A(n57864), .B(n57865), .Z(n57862) );
  XOR U67079 ( .A(n57861), .B(n57862), .Z(n57857) );
  XOR U67080 ( .A(n57856), .B(n57857), .Z(n57854) );
  XOR U67081 ( .A(n57853), .B(n57854), .Z(n57898) );
  XOR U67082 ( .A(n57899), .B(n57898), .Z(n54495) );
  XOR U67083 ( .A(n57900), .B(n54495), .Z(n54496) );
  XOR U67084 ( .A(n54497), .B(n54496), .Z(n57888) );
  IV U67085 ( .A(n57888), .Z(n57889) );
  IV U67086 ( .A(n54498), .Z(n54499) );
  NOR U67087 ( .A(n54500), .B(n54499), .Z(n54505) );
  IV U67088 ( .A(n54501), .Z(n54502) );
  NOR U67089 ( .A(n54503), .B(n54502), .Z(n54504) );
  NOR U67090 ( .A(n54505), .B(n54504), .Z(n57884) );
  XOR U67091 ( .A(n57889), .B(n57884), .Z(n55165) );
  XOR U67092 ( .A(n54506), .B(n55165), .Z(n54507) );
  IV U67093 ( .A(n54507), .Z(n55168) );
  XOR U67094 ( .A(n55167), .B(n55168), .Z(n57935) );
  XOR U67095 ( .A(n57930), .B(n57935), .Z(n57979) );
  IV U67096 ( .A(n54508), .Z(n54509) );
  NOR U67097 ( .A(n54510), .B(n54509), .Z(n57933) );
  NOR U67098 ( .A(n57933), .B(n54511), .Z(n54512) );
  XOR U67099 ( .A(n57979), .B(n54512), .Z(n57981) );
  XOR U67100 ( .A(n57980), .B(n57981), .Z(n57914) );
  XOR U67101 ( .A(n57913), .B(n57914), .Z(n57920) );
  XOR U67102 ( .A(n54513), .B(n57920), .Z(n57951) );
  XOR U67103 ( .A(n57950), .B(n57951), .Z(n54514) );
  IV U67104 ( .A(n54514), .Z(n57948) );
  XOR U67105 ( .A(n57947), .B(n57948), .Z(n57953) );
  XOR U67106 ( .A(n57952), .B(n57953), .Z(n54516) );
  NOR U67107 ( .A(n54515), .B(n54516), .Z(n57966) );
  IV U67108 ( .A(n54516), .Z(n54517) );
  NOR U67109 ( .A(n54518), .B(n54517), .Z(n57963) );
  IV U67110 ( .A(n54519), .Z(n54520) );
  NOR U67111 ( .A(n54521), .B(n54520), .Z(n57962) );
  XOR U67112 ( .A(n57963), .B(n57962), .Z(n54522) );
  NOR U67113 ( .A(n57966), .B(n54522), .Z(n57942) );
  XOR U67114 ( .A(n57944), .B(n57942), .Z(n57940) );
  XOR U67115 ( .A(n57941), .B(n57940), .Z(n54529) );
  NOR U67116 ( .A(n54528), .B(n54529), .Z(n54523) );
  IV U67117 ( .A(n54523), .Z(n54527) );
  IV U67118 ( .A(n54524), .Z(n54525) );
  NOR U67119 ( .A(n54526), .B(n54525), .Z(n54532) );
  NOR U67120 ( .A(n54527), .B(n54532), .Z(n54538) );
  IV U67121 ( .A(n54528), .Z(n54533) );
  XOR U67122 ( .A(n54532), .B(n54533), .Z(n54531) );
  IV U67123 ( .A(n54529), .Z(n54530) );
  NOR U67124 ( .A(n54531), .B(n54530), .Z(n54536) );
  IV U67125 ( .A(n54532), .Z(n54534) );
  NOR U67126 ( .A(n54534), .B(n54533), .Z(n54535) );
  NOR U67127 ( .A(n54536), .B(n54535), .Z(n54537) );
  IV U67128 ( .A(n54537), .Z(n57999) );
  NOR U67129 ( .A(n54538), .B(n57999), .Z(n54539) );
  IV U67130 ( .A(n54539), .Z(n57998) );
  XOR U67131 ( .A(n57996), .B(n57998), .Z(n54540) );
  NOR U67132 ( .A(n54541), .B(n54540), .Z(n57993) );
  IV U67133 ( .A(n54542), .Z(n54543) );
  NOR U67134 ( .A(n54544), .B(n54543), .Z(n57990) );
  NOR U67135 ( .A(n57996), .B(n57990), .Z(n54545) );
  XOR U67136 ( .A(n57998), .B(n54545), .Z(n54546) );
  NOR U67137 ( .A(n54547), .B(n54546), .Z(n54548) );
  NOR U67138 ( .A(n57993), .B(n54548), .Z(n57973) );
  XOR U67139 ( .A(n57975), .B(n57973), .Z(n57971) );
  XOR U67140 ( .A(n57972), .B(n57971), .Z(n54556) );
  IV U67141 ( .A(n54549), .Z(n54550) );
  NOR U67142 ( .A(n54568), .B(n54550), .Z(n54557) );
  IV U67143 ( .A(n54551), .Z(n54553) );
  NOR U67144 ( .A(n54553), .B(n54552), .Z(n54559) );
  NOR U67145 ( .A(n54557), .B(n54559), .Z(n54554) );
  IV U67146 ( .A(n54554), .Z(n54555) );
  NOR U67147 ( .A(n54556), .B(n54555), .Z(n54566) );
  IV U67148 ( .A(n54557), .Z(n54558) );
  NOR U67149 ( .A(n54558), .B(n57971), .Z(n54564) );
  IV U67150 ( .A(n54559), .Z(n54562) );
  XOR U67151 ( .A(n57971), .B(n54560), .Z(n54561) );
  NOR U67152 ( .A(n54562), .B(n54561), .Z(n54563) );
  NOR U67153 ( .A(n54564), .B(n54563), .Z(n54565) );
  IV U67154 ( .A(n54565), .Z(n58013) );
  NOR U67155 ( .A(n54566), .B(n58013), .Z(n54573) );
  IV U67156 ( .A(n54573), .Z(n54571) );
  IV U67157 ( .A(n54567), .Z(n54569) );
  NOR U67158 ( .A(n54569), .B(n54568), .Z(n54572) );
  IV U67159 ( .A(n54572), .Z(n54570) );
  NOR U67160 ( .A(n54571), .B(n54570), .Z(n58004) );
  NOR U67161 ( .A(n54573), .B(n54572), .Z(n58007) );
  NOR U67162 ( .A(n58004), .B(n58007), .Z(n54583) );
  IV U67163 ( .A(n54578), .Z(n54574) );
  NOR U67164 ( .A(n54574), .B(n54576), .Z(n54582) );
  IV U67165 ( .A(n54575), .Z(n54580) );
  IV U67166 ( .A(n54576), .Z(n54577) );
  NOR U67167 ( .A(n54578), .B(n54577), .Z(n54579) );
  NOR U67168 ( .A(n54580), .B(n54579), .Z(n54581) );
  NOR U67169 ( .A(n54582), .B(n54581), .Z(n58003) );
  XOR U67170 ( .A(n54583), .B(n58003), .Z(n55158) );
  XOR U67171 ( .A(n55157), .B(n55158), .Z(n55160) );
  XOR U67172 ( .A(n55161), .B(n55160), .Z(n55138) );
  XOR U67173 ( .A(n55138), .B(n55139), .Z(n55142) );
  XOR U67174 ( .A(n55141), .B(n55142), .Z(n55148) );
  XOR U67175 ( .A(n55147), .B(n55148), .Z(n58054) );
  XOR U67176 ( .A(n58053), .B(n58054), .Z(n55153) );
  XOR U67177 ( .A(n54587), .B(n55153), .Z(n54588) );
  XOR U67178 ( .A(n54589), .B(n54588), .Z(n58020) );
  XOR U67179 ( .A(n58018), .B(n58020), .Z(n58022) );
  XOR U67180 ( .A(n58021), .B(n58022), .Z(n58047) );
  XOR U67181 ( .A(n58042), .B(n58047), .Z(n58027) );
  XOR U67182 ( .A(n54590), .B(n58027), .Z(n58071) );
  XOR U67183 ( .A(n58070), .B(n58071), .Z(n58033) );
  XOR U67184 ( .A(n58032), .B(n58033), .Z(n58030) );
  XOR U67185 ( .A(n58029), .B(n58030), .Z(n58074) );
  XOR U67186 ( .A(n58073), .B(n58074), .Z(n58068) );
  XOR U67187 ( .A(n58067), .B(n58068), .Z(n55132) );
  XOR U67188 ( .A(n55129), .B(n55132), .Z(n54591) );
  XOR U67189 ( .A(n55128), .B(n54591), .Z(n54592) );
  XOR U67190 ( .A(n55124), .B(n54592), .Z(n54601) );
  NOR U67191 ( .A(n54600), .B(n54601), .Z(n54593) );
  IV U67192 ( .A(n54593), .Z(n54599) );
  IV U67193 ( .A(n54594), .Z(n54598) );
  NOR U67194 ( .A(n54596), .B(n54595), .Z(n54597) );
  IV U67195 ( .A(n54597), .Z(n54612) );
  NOR U67196 ( .A(n54598), .B(n54612), .Z(n54604) );
  NOR U67197 ( .A(n54599), .B(n54604), .Z(n54610) );
  IV U67198 ( .A(n54600), .Z(n54605) );
  XOR U67199 ( .A(n54604), .B(n54605), .Z(n54603) );
  IV U67200 ( .A(n54601), .Z(n54602) );
  NOR U67201 ( .A(n54603), .B(n54602), .Z(n54608) );
  IV U67202 ( .A(n54604), .Z(n54606) );
  NOR U67203 ( .A(n54606), .B(n54605), .Z(n54607) );
  NOR U67204 ( .A(n54608), .B(n54607), .Z(n58094) );
  IV U67205 ( .A(n58094), .Z(n54609) );
  NOR U67206 ( .A(n54610), .B(n54609), .Z(n58098) );
  IV U67207 ( .A(n54611), .Z(n54613) );
  NOR U67208 ( .A(n54613), .B(n54612), .Z(n58097) );
  IV U67209 ( .A(n58097), .Z(n58099) );
  XOR U67210 ( .A(n58098), .B(n58099), .Z(n54614) );
  XOR U67211 ( .A(n54615), .B(n54614), .Z(n58086) );
  XOR U67212 ( .A(n58085), .B(n58086), .Z(n58089) );
  XOR U67213 ( .A(n58088), .B(n58089), .Z(n55096) );
  XOR U67214 ( .A(n55095), .B(n55096), .Z(n54619) );
  IV U67215 ( .A(n54616), .Z(n54618) );
  NOR U67216 ( .A(n54618), .B(n54617), .Z(n55098) );
  XOR U67217 ( .A(n54619), .B(n55098), .Z(n55117) );
  IV U67218 ( .A(n54620), .Z(n54621) );
  NOR U67219 ( .A(n54622), .B(n54621), .Z(n54629) );
  NOR U67220 ( .A(n54624), .B(n54623), .Z(n54625) );
  IV U67221 ( .A(n54625), .Z(n54627) );
  NOR U67222 ( .A(n54627), .B(n54626), .Z(n54628) );
  NOR U67223 ( .A(n54629), .B(n54628), .Z(n55119) );
  XOR U67224 ( .A(n55117), .B(n55119), .Z(n55107) );
  XOR U67225 ( .A(n55106), .B(n55107), .Z(n55113) );
  XOR U67226 ( .A(n55112), .B(n55113), .Z(n55104) );
  XOR U67227 ( .A(n55103), .B(n55104), .Z(n58117) );
  XOR U67228 ( .A(n58116), .B(n58117), .Z(n58115) );
  XOR U67229 ( .A(n58113), .B(n58115), .Z(n58126) );
  XOR U67230 ( .A(n58124), .B(n58126), .Z(n58123) );
  XOR U67231 ( .A(n58121), .B(n58123), .Z(n58139) );
  XOR U67232 ( .A(n58137), .B(n58139), .Z(n55091) );
  XOR U67233 ( .A(n55089), .B(n55091), .Z(n58145) );
  XOR U67234 ( .A(n54630), .B(n58145), .Z(n58148) );
  XOR U67235 ( .A(n58147), .B(n58148), .Z(n58156) );
  XOR U67236 ( .A(n58155), .B(n58156), .Z(n58153) );
  XOR U67237 ( .A(n58152), .B(n58153), .Z(n58165) );
  XOR U67238 ( .A(n58164), .B(n58165), .Z(n58177) );
  XOR U67239 ( .A(n58170), .B(n58177), .Z(n58184) );
  IV U67240 ( .A(n54631), .Z(n54632) );
  NOR U67241 ( .A(n54633), .B(n54632), .Z(n58182) );
  IV U67242 ( .A(n54634), .Z(n58178) );
  NOR U67243 ( .A(n54635), .B(n58178), .Z(n54636) );
  NOR U67244 ( .A(n58182), .B(n54636), .Z(n54637) );
  XOR U67245 ( .A(n58184), .B(n54637), .Z(n54647) );
  IV U67246 ( .A(n54647), .Z(n54644) );
  IV U67247 ( .A(n54638), .Z(n54640) );
  NOR U67248 ( .A(n54640), .B(n54639), .Z(n54643) );
  IV U67249 ( .A(n54650), .Z(n54641) );
  NOR U67250 ( .A(n54649), .B(n54641), .Z(n54642) );
  NOR U67251 ( .A(n54643), .B(n54642), .Z(n54645) );
  NOR U67252 ( .A(n54644), .B(n54645), .Z(n58193) );
  IV U67253 ( .A(n54645), .Z(n54646) );
  NOR U67254 ( .A(n54647), .B(n54646), .Z(n58190) );
  IV U67255 ( .A(n54648), .Z(n54652) );
  XOR U67256 ( .A(n54650), .B(n54649), .Z(n54651) );
  NOR U67257 ( .A(n54652), .B(n54651), .Z(n58189) );
  XOR U67258 ( .A(n58190), .B(n58189), .Z(n54653) );
  NOR U67259 ( .A(n58193), .B(n54653), .Z(n55079) );
  XOR U67260 ( .A(n55080), .B(n55079), .Z(n55082) );
  XOR U67261 ( .A(n54660), .B(n55082), .Z(n54654) );
  NOR U67262 ( .A(n54655), .B(n54654), .Z(n55085) );
  IV U67263 ( .A(n54656), .Z(n54657) );
  NOR U67264 ( .A(n54658), .B(n54657), .Z(n54659) );
  NOR U67265 ( .A(n54660), .B(n54659), .Z(n55083) );
  XOR U67266 ( .A(n55082), .B(n55083), .Z(n54661) );
  NOR U67267 ( .A(n54662), .B(n54661), .Z(n54663) );
  NOR U67268 ( .A(n55085), .B(n54663), .Z(n54664) );
  IV U67269 ( .A(n54664), .Z(n58202) );
  XOR U67270 ( .A(n58201), .B(n58202), .Z(n58200) );
  XOR U67271 ( .A(n58198), .B(n58200), .Z(n58197) );
  XOR U67272 ( .A(n54665), .B(n58197), .Z(n55075) );
  XOR U67273 ( .A(n55073), .B(n55075), .Z(n55069) );
  NOR U67274 ( .A(n54667), .B(n54666), .Z(n55068) );
  NOR U67275 ( .A(n55074), .B(n55068), .Z(n54668) );
  XOR U67276 ( .A(n55069), .B(n54668), .Z(n58216) );
  XOR U67277 ( .A(n58215), .B(n58216), .Z(n58220) );
  XOR U67278 ( .A(n58218), .B(n58220), .Z(n58252) );
  XOR U67279 ( .A(n58251), .B(n58252), .Z(n58228) );
  XOR U67280 ( .A(n58223), .B(n58228), .Z(n54669) );
  XOR U67281 ( .A(n58226), .B(n54669), .Z(n58250) );
  XOR U67282 ( .A(n58249), .B(n58250), .Z(n55061) );
  IV U67283 ( .A(n55061), .Z(n55060) );
  IV U67284 ( .A(n54670), .Z(n54672) );
  NOR U67285 ( .A(n54672), .B(n54671), .Z(n55063) );
  XOR U67286 ( .A(n55060), .B(n55063), .Z(n55056) );
  IV U67287 ( .A(n55056), .Z(n54679) );
  IV U67288 ( .A(n54673), .Z(n54674) );
  NOR U67289 ( .A(n54675), .B(n54674), .Z(n55059) );
  IV U67290 ( .A(n54676), .Z(n54677) );
  NOR U67291 ( .A(n54677), .B(n54681), .Z(n55054) );
  NOR U67292 ( .A(n55059), .B(n55054), .Z(n54678) );
  XOR U67293 ( .A(n54679), .B(n54678), .Z(n55052) );
  IV U67294 ( .A(n54680), .Z(n54682) );
  NOR U67295 ( .A(n54682), .B(n54681), .Z(n55051) );
  XOR U67296 ( .A(n55052), .B(n55051), .Z(n54684) );
  NOR U67297 ( .A(n54683), .B(n54684), .Z(n55050) );
  IV U67298 ( .A(n54684), .Z(n54685) );
  NOR U67299 ( .A(n54686), .B(n54685), .Z(n55048) );
  IV U67300 ( .A(n54687), .Z(n54688) );
  NOR U67301 ( .A(n54689), .B(n54688), .Z(n55046) );
  XOR U67302 ( .A(n55048), .B(n55046), .Z(n54690) );
  NOR U67303 ( .A(n55050), .B(n54690), .Z(n58244) );
  NOR U67304 ( .A(n54692), .B(n54691), .Z(n55045) );
  IV U67305 ( .A(n54693), .Z(n54695) );
  IV U67306 ( .A(n54694), .Z(n54698) );
  NOR U67307 ( .A(n54695), .B(n54698), .Z(n58243) );
  NOR U67308 ( .A(n55045), .B(n58243), .Z(n54696) );
  XOR U67309 ( .A(n58244), .B(n54696), .Z(n58261) );
  IV U67310 ( .A(n54697), .Z(n54699) );
  NOR U67311 ( .A(n54699), .B(n54698), .Z(n58241) );
  XOR U67312 ( .A(n58261), .B(n58241), .Z(n54700) );
  NOR U67313 ( .A(n54701), .B(n54700), .Z(n58264) );
  IV U67314 ( .A(n54702), .Z(n54703) );
  NOR U67315 ( .A(n54704), .B(n54703), .Z(n58260) );
  NOR U67316 ( .A(n58260), .B(n58241), .Z(n54705) );
  XOR U67317 ( .A(n58261), .B(n54705), .Z(n58278) );
  NOR U67318 ( .A(n54706), .B(n58278), .Z(n54707) );
  NOR U67319 ( .A(n58264), .B(n54707), .Z(n58274) );
  NOR U67320 ( .A(n54709), .B(n54708), .Z(n58277) );
  IV U67321 ( .A(n54710), .Z(n54713) );
  IV U67322 ( .A(n54711), .Z(n54712) );
  NOR U67323 ( .A(n54713), .B(n54712), .Z(n58273) );
  NOR U67324 ( .A(n58277), .B(n58273), .Z(n54714) );
  XOR U67325 ( .A(n58274), .B(n54714), .Z(n58272) );
  XOR U67326 ( .A(n58270), .B(n58272), .Z(n58314) );
  IV U67327 ( .A(n54715), .Z(n54717) );
  NOR U67328 ( .A(n54717), .B(n54716), .Z(n58269) );
  NOR U67329 ( .A(n58269), .B(n58313), .Z(n54718) );
  XOR U67330 ( .A(n58314), .B(n54718), .Z(n58288) );
  IV U67331 ( .A(n54719), .Z(n54721) );
  NOR U67332 ( .A(n54721), .B(n54720), .Z(n58287) );
  NOR U67333 ( .A(n58310), .B(n58287), .Z(n54722) );
  XOR U67334 ( .A(n58288), .B(n54722), .Z(n58292) );
  IV U67335 ( .A(n54723), .Z(n54725) );
  NOR U67336 ( .A(n54725), .B(n54724), .Z(n58290) );
  XOR U67337 ( .A(n58292), .B(n58290), .Z(n58307) );
  IV U67338 ( .A(n54726), .Z(n54728) );
  NOR U67339 ( .A(n54728), .B(n54727), .Z(n58305) );
  XOR U67340 ( .A(n58307), .B(n58305), .Z(n58304) );
  IV U67341 ( .A(n54729), .Z(n54730) );
  NOR U67342 ( .A(n54731), .B(n54730), .Z(n54732) );
  IV U67343 ( .A(n54732), .Z(n58303) );
  XOR U67344 ( .A(n58304), .B(n58303), .Z(n54733) );
  NOR U67345 ( .A(n54735), .B(n54733), .Z(n54740) );
  IV U67346 ( .A(n54740), .Z(n54734) );
  NOR U67347 ( .A(n54738), .B(n54734), .Z(n58298) );
  IV U67348 ( .A(n54735), .Z(n54736) );
  NOR U67349 ( .A(n58304), .B(n54736), .Z(n54737) );
  NOR U67350 ( .A(n54738), .B(n54737), .Z(n54739) );
  NOR U67351 ( .A(n54740), .B(n54739), .Z(n58295) );
  NOR U67352 ( .A(n58298), .B(n58295), .Z(n55039) );
  XOR U67353 ( .A(n54741), .B(n55039), .Z(n55037) );
  XOR U67354 ( .A(n55038), .B(n55037), .Z(n58343) );
  IV U67355 ( .A(n54745), .Z(n54742) );
  NOR U67356 ( .A(n54742), .B(n54744), .Z(n54749) );
  IV U67357 ( .A(n54743), .Z(n54747) );
  XOR U67358 ( .A(n54745), .B(n54744), .Z(n54746) );
  NOR U67359 ( .A(n54747), .B(n54746), .Z(n54748) );
  NOR U67360 ( .A(n54749), .B(n54748), .Z(n58344) );
  XOR U67361 ( .A(n58343), .B(n58344), .Z(n58347) );
  XOR U67362 ( .A(n58346), .B(n58347), .Z(n54750) );
  NOR U67363 ( .A(n54751), .B(n54750), .Z(n58327) );
  IV U67364 ( .A(n54752), .Z(n54753) );
  NOR U67365 ( .A(n54754), .B(n54753), .Z(n58322) );
  NOR U67366 ( .A(n58346), .B(n58322), .Z(n54755) );
  XOR U67367 ( .A(n58347), .B(n54755), .Z(n54756) );
  NOR U67368 ( .A(n54757), .B(n54756), .Z(n58325) );
  NOR U67369 ( .A(n58327), .B(n58325), .Z(n54758) );
  XOR U67370 ( .A(n58324), .B(n54758), .Z(n58373) );
  XOR U67371 ( .A(n58371), .B(n58373), .Z(n58339) );
  IV U67372 ( .A(n54759), .Z(n54760) );
  NOR U67373 ( .A(n54761), .B(n54760), .Z(n58372) );
  IV U67374 ( .A(n54762), .Z(n54763) );
  NOR U67375 ( .A(n54764), .B(n54763), .Z(n58338) );
  NOR U67376 ( .A(n58372), .B(n58338), .Z(n54765) );
  XOR U67377 ( .A(n58339), .B(n54765), .Z(n54766) );
  IV U67378 ( .A(n54766), .Z(n58336) );
  XOR U67379 ( .A(n58335), .B(n58336), .Z(n58379) );
  XOR U67380 ( .A(n54767), .B(n58379), .Z(n58376) );
  XOR U67381 ( .A(n58375), .B(n58376), .Z(n55026) );
  IV U67382 ( .A(n54768), .Z(n54769) );
  NOR U67383 ( .A(n54770), .B(n54769), .Z(n55025) );
  XOR U67384 ( .A(n55026), .B(n55025), .Z(n55030) );
  XOR U67385 ( .A(n54771), .B(n55030), .Z(n54772) );
  NOR U67386 ( .A(n55028), .B(n54772), .Z(n54779) );
  IV U67387 ( .A(n54773), .Z(n54775) );
  NOR U67388 ( .A(n54775), .B(n54774), .Z(n54781) );
  IV U67389 ( .A(n54781), .Z(n54776) );
  NOR U67390 ( .A(n54779), .B(n54776), .Z(n55033) );
  IV U67391 ( .A(n55028), .Z(n54777) );
  NOR U67392 ( .A(n54777), .B(n55030), .Z(n54778) );
  NOR U67393 ( .A(n54779), .B(n54778), .Z(n54780) );
  NOR U67394 ( .A(n54781), .B(n54780), .Z(n54782) );
  NOR U67395 ( .A(n55033), .B(n54782), .Z(n54789) );
  NOR U67396 ( .A(n54792), .B(n54789), .Z(n54783) );
  IV U67397 ( .A(n54783), .Z(n54787) );
  IV U67398 ( .A(n54784), .Z(n54785) );
  NOR U67399 ( .A(n54786), .B(n54785), .Z(n54788) );
  NOR U67400 ( .A(n54787), .B(n54788), .Z(n54798) );
  IV U67401 ( .A(n54788), .Z(n54793) );
  XOR U67402 ( .A(n54792), .B(n54793), .Z(n54791) );
  IV U67403 ( .A(n54789), .Z(n54790) );
  NOR U67404 ( .A(n54791), .B(n54790), .Z(n54796) );
  IV U67405 ( .A(n54792), .Z(n54794) );
  NOR U67406 ( .A(n54794), .B(n54793), .Z(n54795) );
  NOR U67407 ( .A(n54796), .B(n54795), .Z(n54797) );
  IV U67408 ( .A(n54797), .Z(n58365) );
  NOR U67409 ( .A(n54798), .B(n58365), .Z(n58358) );
  XOR U67410 ( .A(n58360), .B(n58358), .Z(n58356) );
  XOR U67411 ( .A(n58355), .B(n58356), .Z(n55021) );
  XOR U67412 ( .A(n55019), .B(n55021), .Z(n58399) );
  IV U67413 ( .A(n54799), .Z(n54803) );
  IV U67414 ( .A(n54800), .Z(n54801) );
  NOR U67415 ( .A(n54803), .B(n54801), .Z(n55020) );
  IV U67416 ( .A(n54802), .Z(n54806) );
  NOR U67417 ( .A(n54804), .B(n54803), .Z(n54805) );
  IV U67418 ( .A(n54805), .Z(n54809) );
  NOR U67419 ( .A(n54806), .B(n54809), .Z(n58400) );
  NOR U67420 ( .A(n55020), .B(n58400), .Z(n54807) );
  XOR U67421 ( .A(n58399), .B(n54807), .Z(n58397) );
  IV U67422 ( .A(n54808), .Z(n54810) );
  NOR U67423 ( .A(n54810), .B(n54809), .Z(n58396) );
  XOR U67424 ( .A(n58397), .B(n58396), .Z(n58392) );
  XOR U67425 ( .A(n58391), .B(n58392), .Z(n58390) );
  XOR U67426 ( .A(n54811), .B(n58390), .Z(n54969) );
  XOR U67427 ( .A(n54968), .B(n54969), .Z(n54987) );
  XOR U67428 ( .A(n54986), .B(n54987), .Z(n54812) );
  IV U67429 ( .A(n54812), .Z(n54989) );
  XOR U67430 ( .A(n54988), .B(n54989), .Z(n54984) );
  XOR U67431 ( .A(n54983), .B(n54984), .Z(n54978) );
  XOR U67432 ( .A(n54973), .B(n54978), .Z(n54813) );
  XOR U67433 ( .A(n54976), .B(n54813), .Z(n54967) );
  XOR U67434 ( .A(n54966), .B(n54967), .Z(n55006) );
  IV U67435 ( .A(n54814), .Z(n54817) );
  IV U67436 ( .A(n54815), .Z(n54816) );
  NOR U67437 ( .A(n54817), .B(n54816), .Z(n55009) );
  XOR U67438 ( .A(n55006), .B(n55009), .Z(n54822) );
  IV U67439 ( .A(n54818), .Z(n54820) );
  NOR U67440 ( .A(n54820), .B(n54819), .Z(n54821) );
  IV U67441 ( .A(n54821), .Z(n55011) );
  XOR U67442 ( .A(n54822), .B(n55011), .Z(n58426) );
  XOR U67443 ( .A(n58425), .B(n58426), .Z(n58414) );
  IV U67444 ( .A(n54823), .Z(n54825) );
  NOR U67445 ( .A(n54825), .B(n54824), .Z(n58415) );
  IV U67446 ( .A(n58415), .Z(n58413) );
  XOR U67447 ( .A(n58414), .B(n58413), .Z(n54832) );
  NOR U67448 ( .A(n54827), .B(n54826), .Z(n54828) );
  IV U67449 ( .A(n54828), .Z(n54829) );
  NOR U67450 ( .A(n54830), .B(n54829), .Z(n54831) );
  IV U67451 ( .A(n54831), .Z(n58417) );
  XOR U67452 ( .A(n54832), .B(n58417), .Z(n58448) );
  XOR U67453 ( .A(n58447), .B(n58448), .Z(n54833) );
  IV U67454 ( .A(n54833), .Z(n55000) );
  XOR U67455 ( .A(n54998), .B(n55000), .Z(n55002) );
  XOR U67456 ( .A(n55001), .B(n55002), .Z(n58450) );
  XOR U67457 ( .A(n58449), .B(n58450), .Z(n54959) );
  XOR U67458 ( .A(n54958), .B(n54959), .Z(n54962) );
  XOR U67459 ( .A(n54961), .B(n54962), .Z(n58429) );
  XOR U67460 ( .A(n58428), .B(n58429), .Z(n58423) );
  XOR U67461 ( .A(n58422), .B(n58423), .Z(n58441) );
  XOR U67462 ( .A(n54834), .B(n58441), .Z(n58443) );
  XOR U67463 ( .A(n58442), .B(n58443), .Z(n58468) );
  XOR U67464 ( .A(n58466), .B(n58468), .Z(n54835) );
  XOR U67465 ( .A(n54836), .B(n54835), .Z(n58478) );
  XOR U67466 ( .A(n58462), .B(n58478), .Z(n58459) );
  XOR U67467 ( .A(n58458), .B(n58459), .Z(n58504) );
  XOR U67468 ( .A(n58500), .B(n58504), .Z(n54837) );
  XOR U67469 ( .A(n58501), .B(n54837), .Z(n58492) );
  XOR U67470 ( .A(n58490), .B(n58492), .Z(n58486) );
  XOR U67471 ( .A(n58485), .B(n58486), .Z(n58489) );
  XOR U67472 ( .A(n58488), .B(n58489), .Z(n58509) );
  XOR U67473 ( .A(n58510), .B(n58509), .Z(n58513) );
  XOR U67474 ( .A(n58515), .B(n58513), .Z(n54838) );
  XOR U67475 ( .A(n58516), .B(n54838), .Z(n58611) );
  IV U67476 ( .A(n54839), .Z(n54840) );
  NOR U67477 ( .A(n54843), .B(n54840), .Z(n58609) );
  XOR U67478 ( .A(n58611), .B(n58609), .Z(n58526) );
  IV U67479 ( .A(n54841), .Z(n54842) );
  NOR U67480 ( .A(n54843), .B(n54842), .Z(n54844) );
  IV U67481 ( .A(n54844), .Z(n58528) );
  XOR U67482 ( .A(n58526), .B(n58528), .Z(n54845) );
  XOR U67483 ( .A(n58524), .B(n54845), .Z(n54954) );
  XOR U67484 ( .A(n54953), .B(n54954), .Z(n54952) );
  IV U67485 ( .A(n54846), .Z(n54849) );
  IV U67486 ( .A(n54847), .Z(n54848) );
  NOR U67487 ( .A(n54849), .B(n54848), .Z(n54950) );
  XOR U67488 ( .A(n54952), .B(n54950), .Z(n58544) );
  XOR U67489 ( .A(n58543), .B(n58544), .Z(n58547) );
  XOR U67490 ( .A(n58546), .B(n58547), .Z(n58560) );
  XOR U67491 ( .A(n58556), .B(n58560), .Z(n54850) );
  XOR U67492 ( .A(n58555), .B(n54850), .Z(n58606) );
  IV U67493 ( .A(n54851), .Z(n54853) );
  NOR U67494 ( .A(n54853), .B(n54852), .Z(n54858) );
  IV U67495 ( .A(n54854), .Z(n54856) );
  NOR U67496 ( .A(n54856), .B(n54855), .Z(n54857) );
  NOR U67497 ( .A(n54858), .B(n54857), .Z(n58607) );
  XOR U67498 ( .A(n58606), .B(n58607), .Z(n58539) );
  XOR U67499 ( .A(n58538), .B(n58539), .Z(n58537) );
  XOR U67500 ( .A(n58535), .B(n58537), .Z(n58566) );
  XOR U67501 ( .A(n58565), .B(n58566), .Z(n58568) );
  XOR U67502 ( .A(n54865), .B(n58568), .Z(n54859) );
  NOR U67503 ( .A(n54860), .B(n54859), .Z(n58593) );
  IV U67504 ( .A(n54861), .Z(n54862) );
  NOR U67505 ( .A(n54863), .B(n54862), .Z(n54864) );
  NOR U67506 ( .A(n54865), .B(n54864), .Z(n58569) );
  XOR U67507 ( .A(n58569), .B(n58568), .Z(n58589) );
  NOR U67508 ( .A(n54866), .B(n58589), .Z(n54867) );
  NOR U67509 ( .A(n58593), .B(n54867), .Z(n58573) );
  IV U67510 ( .A(n54868), .Z(n54869) );
  NOR U67511 ( .A(n54870), .B(n54869), .Z(n58588) );
  IV U67512 ( .A(n54871), .Z(n54872) );
  NOR U67513 ( .A(n54872), .B(n54875), .Z(n58572) );
  NOR U67514 ( .A(n58588), .B(n58572), .Z(n54873) );
  XOR U67515 ( .A(n58573), .B(n54873), .Z(n58577) );
  IV U67516 ( .A(n54874), .Z(n54876) );
  NOR U67517 ( .A(n54876), .B(n54875), .Z(n54878) );
  NOR U67518 ( .A(n54878), .B(n54877), .Z(n58576) );
  XOR U67519 ( .A(n58577), .B(n58576), .Z(n54944) );
  NOR U67520 ( .A(n54880), .B(n54879), .Z(n54943) );
  NOR U67521 ( .A(n58578), .B(n54943), .Z(n54881) );
  XOR U67522 ( .A(n54944), .B(n54881), .Z(n58602) );
  XOR U67523 ( .A(n54882), .B(n58602), .Z(n54883) );
  IV U67524 ( .A(n54883), .Z(n58600) );
  XOR U67525 ( .A(n54885), .B(n54884), .Z(n54939) );
  IV U67526 ( .A(n54886), .Z(n54890) );
  NOR U67527 ( .A(n54888), .B(n54887), .Z(n54889) );
  XOR U67528 ( .A(n54890), .B(n54889), .Z(n54935) );
  XOR U67529 ( .A(n54892), .B(n54891), .Z(n58627) );
  IV U67530 ( .A(n54893), .Z(n54895) );
  NOR U67531 ( .A(n54895), .B(n54894), .Z(n54924) );
  IV U67532 ( .A(n54924), .Z(n54896) );
  NOR U67533 ( .A(n54897), .B(n54896), .Z(n58626) );
  IV U67534 ( .A(n58626), .Z(n54898) );
  NOR U67535 ( .A(n58627), .B(n54898), .Z(n54917) );
  IV U67536 ( .A(n54917), .Z(n54899) );
  NOR U67537 ( .A(n54916), .B(n54899), .Z(n58632) );
  IV U67538 ( .A(n58632), .Z(n54902) );
  XOR U67539 ( .A(n54901), .B(n54900), .Z(n58633) );
  NOR U67540 ( .A(n54902), .B(n58633), .Z(n54936) );
  IV U67541 ( .A(n54936), .Z(n54903) );
  NOR U67542 ( .A(n54935), .B(n54903), .Z(n54911) );
  IV U67543 ( .A(n54911), .Z(n54906) );
  XOR U67544 ( .A(n54905), .B(n54904), .Z(n54914) );
  NOR U67545 ( .A(n54906), .B(n54914), .Z(n54940) );
  IV U67546 ( .A(n54940), .Z(n54907) );
  NOR U67547 ( .A(n54939), .B(n54907), .Z(n58642) );
  IV U67548 ( .A(n58642), .Z(n54910) );
  XOR U67549 ( .A(n54909), .B(n54908), .Z(n58643) );
  NOR U67550 ( .A(n54910), .B(n58643), .Z(n58598) );
  XOR U67551 ( .A(n58600), .B(n58598), .Z(n58645) );
  NOR U67552 ( .A(n54912), .B(n54911), .Z(n54913) );
  XOR U67553 ( .A(n54914), .B(n54913), .Z(n54915) );
  IV U67554 ( .A(n54915), .Z(n58638) );
  IV U67555 ( .A(n54916), .Z(n54923) );
  NOR U67556 ( .A(n54918), .B(n54917), .Z(n54919) );
  IV U67557 ( .A(n54919), .Z(n54920) );
  NOR U67558 ( .A(n54921), .B(n54920), .Z(n54922) );
  XOR U67559 ( .A(n54923), .B(n54922), .Z(n58630) );
  NOR U67560 ( .A(n54925), .B(n54924), .Z(n54926) );
  XOR U67561 ( .A(n54927), .B(n54926), .Z(n58624) );
  NOR U67562 ( .A(n54929), .B(n54928), .Z(n54930) );
  IV U67563 ( .A(n54930), .Z(n58623) );
  NOR U67564 ( .A(n58624), .B(n58623), .Z(n58625) );
  IV U67565 ( .A(n58625), .Z(n54931) );
  NOR U67566 ( .A(n58627), .B(n54931), .Z(n54932) );
  IV U67567 ( .A(n54932), .Z(n58629) );
  NOR U67568 ( .A(n58630), .B(n58629), .Z(n58631) );
  IV U67569 ( .A(n58631), .Z(n54933) );
  NOR U67570 ( .A(n58633), .B(n54933), .Z(n54934) );
  IV U67571 ( .A(n54934), .Z(n58636) );
  XOR U67572 ( .A(n54936), .B(n54935), .Z(n58635) );
  NOR U67573 ( .A(n58636), .B(n58635), .Z(n54937) );
  IV U67574 ( .A(n54937), .Z(n58637) );
  NOR U67575 ( .A(n58638), .B(n58637), .Z(n54938) );
  IV U67576 ( .A(n54938), .Z(n58640) );
  XOR U67577 ( .A(n54940), .B(n54939), .Z(n58639) );
  NOR U67578 ( .A(n58640), .B(n58639), .Z(n58641) );
  IV U67579 ( .A(n58641), .Z(n54941) );
  NOR U67580 ( .A(n54941), .B(n58643), .Z(n54942) );
  IV U67581 ( .A(n54942), .Z(n58646) );
  NOR U67582 ( .A(n58645), .B(n58646), .Z(n58621) );
  IV U67583 ( .A(n54943), .Z(n54945) );
  IV U67584 ( .A(n54944), .Z(n58579) );
  NOR U67585 ( .A(n54945), .B(n58579), .Z(n54949) );
  IV U67586 ( .A(n54946), .Z(n54947) );
  NOR U67587 ( .A(n54947), .B(n58602), .Z(n54948) );
  NOR U67588 ( .A(n54949), .B(n54948), .Z(n58619) );
  IV U67589 ( .A(n54950), .Z(n54951) );
  NOR U67590 ( .A(n54952), .B(n54951), .Z(n54957) );
  IV U67591 ( .A(n54953), .Z(n54955) );
  NOR U67592 ( .A(n54955), .B(n54954), .Z(n54956) );
  NOR U67593 ( .A(n54957), .B(n54956), .Z(n58534) );
  IV U67594 ( .A(n54958), .Z(n54960) );
  NOR U67595 ( .A(n54960), .B(n54959), .Z(n54965) );
  IV U67596 ( .A(n54961), .Z(n54963) );
  NOR U67597 ( .A(n54963), .B(n54962), .Z(n54964) );
  NOR U67598 ( .A(n54965), .B(n54964), .Z(n58439) );
  NOR U67599 ( .A(n54967), .B(n54966), .Z(n54972) );
  IV U67600 ( .A(n54968), .Z(n54970) );
  NOR U67601 ( .A(n54970), .B(n54969), .Z(n54971) );
  NOR U67602 ( .A(n54972), .B(n54971), .Z(n54982) );
  IV U67603 ( .A(n54976), .Z(n54974) );
  IV U67604 ( .A(n54973), .Z(n54975) );
  NOR U67605 ( .A(n54974), .B(n54975), .Z(n54980) );
  XOR U67606 ( .A(n54976), .B(n54975), .Z(n54977) );
  NOR U67607 ( .A(n54978), .B(n54977), .Z(n54979) );
  NOR U67608 ( .A(n54980), .B(n54979), .Z(n54981) );
  XOR U67609 ( .A(n54982), .B(n54981), .Z(n54997) );
  IV U67610 ( .A(n54983), .Z(n54985) );
  NOR U67611 ( .A(n54985), .B(n54984), .Z(n54995) );
  NOR U67612 ( .A(n54987), .B(n54986), .Z(n54992) );
  IV U67613 ( .A(n54988), .Z(n54990) );
  NOR U67614 ( .A(n54990), .B(n54989), .Z(n54991) );
  NOR U67615 ( .A(n54992), .B(n54991), .Z(n54993) );
  IV U67616 ( .A(n54993), .Z(n54994) );
  NOR U67617 ( .A(n54995), .B(n54994), .Z(n54996) );
  XOR U67618 ( .A(n54997), .B(n54996), .Z(n55017) );
  IV U67619 ( .A(n54998), .Z(n54999) );
  NOR U67620 ( .A(n55000), .B(n54999), .Z(n55005) );
  IV U67621 ( .A(n55001), .Z(n55003) );
  NOR U67622 ( .A(n55003), .B(n55002), .Z(n55004) );
  NOR U67623 ( .A(n55005), .B(n55004), .Z(n55015) );
  IV U67624 ( .A(n55009), .Z(n55007) );
  IV U67625 ( .A(n55006), .Z(n55008) );
  NOR U67626 ( .A(n55007), .B(n55008), .Z(n55013) );
  XOR U67627 ( .A(n55009), .B(n55008), .Z(n55010) );
  NOR U67628 ( .A(n55011), .B(n55010), .Z(n55012) );
  NOR U67629 ( .A(n55013), .B(n55012), .Z(n55014) );
  XOR U67630 ( .A(n55015), .B(n55014), .Z(n55016) );
  XOR U67631 ( .A(n55017), .B(n55016), .Z(n58412) );
  IV U67632 ( .A(n55020), .Z(n55018) );
  NOR U67633 ( .A(n55018), .B(n55019), .Z(n55024) );
  XOR U67634 ( .A(n55020), .B(n55019), .Z(n55022) );
  NOR U67635 ( .A(n55022), .B(n55021), .Z(n55023) );
  NOR U67636 ( .A(n55024), .B(n55023), .Z(n58410) );
  IV U67637 ( .A(n55025), .Z(n55027) );
  NOR U67638 ( .A(n55027), .B(n55026), .Z(n55036) );
  NOR U67639 ( .A(n55029), .B(n55028), .Z(n55031) );
  NOR U67640 ( .A(n55031), .B(n55030), .Z(n55032) );
  NOR U67641 ( .A(n55033), .B(n55032), .Z(n55034) );
  IV U67642 ( .A(n55034), .Z(n55035) );
  NOR U67643 ( .A(n55036), .B(n55035), .Z(n58388) );
  NOR U67644 ( .A(n55038), .B(n55037), .Z(n55044) );
  IV U67645 ( .A(n55039), .Z(n55042) );
  IV U67646 ( .A(n55040), .Z(n55041) );
  NOR U67647 ( .A(n55042), .B(n55041), .Z(n55043) );
  NOR U67648 ( .A(n55044), .B(n55043), .Z(n58334) );
  NOR U67649 ( .A(n55046), .B(n55045), .Z(n55047) );
  NOR U67650 ( .A(n55048), .B(n55047), .Z(n55049) );
  NOR U67651 ( .A(n55050), .B(n55049), .Z(n58268) );
  IV U67652 ( .A(n55051), .Z(n55053) );
  NOR U67653 ( .A(n55053), .B(n55052), .Z(n55058) );
  IV U67654 ( .A(n55054), .Z(n55055) );
  NOR U67655 ( .A(n55056), .B(n55055), .Z(n55057) );
  NOR U67656 ( .A(n55058), .B(n55057), .Z(n58240) );
  IV U67657 ( .A(n55059), .Z(n55062) );
  NOR U67658 ( .A(n55062), .B(n55060), .Z(n55067) );
  XOR U67659 ( .A(n55062), .B(n55061), .Z(n55065) );
  IV U67660 ( .A(n55063), .Z(n55064) );
  NOR U67661 ( .A(n55065), .B(n55064), .Z(n55066) );
  NOR U67662 ( .A(n55067), .B(n55066), .Z(n58238) );
  IV U67663 ( .A(n55068), .Z(n55071) );
  IV U67664 ( .A(n55069), .Z(n55070) );
  NOR U67665 ( .A(n55071), .B(n55070), .Z(n58236) );
  IV U67666 ( .A(n55074), .Z(n55072) );
  NOR U67667 ( .A(n55072), .B(n55073), .Z(n55078) );
  XOR U67668 ( .A(n55074), .B(n55073), .Z(n55076) );
  NOR U67669 ( .A(n55076), .B(n55075), .Z(n55077) );
  NOR U67670 ( .A(n55078), .B(n55077), .Z(n58214) );
  IV U67671 ( .A(n55079), .Z(n55081) );
  NOR U67672 ( .A(n55081), .B(n55080), .Z(n55088) );
  NOR U67673 ( .A(n55083), .B(n55082), .Z(n55084) );
  NOR U67674 ( .A(n55085), .B(n55084), .Z(n55086) );
  IV U67675 ( .A(n55086), .Z(n55087) );
  NOR U67676 ( .A(n55088), .B(n55087), .Z(n58212) );
  IV U67677 ( .A(n55089), .Z(n55090) );
  NOR U67678 ( .A(n55091), .B(n55090), .Z(n55094) );
  IV U67679 ( .A(n58133), .Z(n55092) );
  NOR U67680 ( .A(n55092), .B(n58145), .Z(n55093) );
  NOR U67681 ( .A(n55094), .B(n55093), .Z(n58112) );
  NOR U67682 ( .A(n55095), .B(n55096), .Z(n55102) );
  XOR U67683 ( .A(n55097), .B(n55096), .Z(n55100) );
  IV U67684 ( .A(n55098), .Z(n55099) );
  NOR U67685 ( .A(n55100), .B(n55099), .Z(n55101) );
  NOR U67686 ( .A(n55102), .B(n55101), .Z(n55123) );
  IV U67687 ( .A(n55103), .Z(n55105) );
  NOR U67688 ( .A(n55105), .B(n55104), .Z(n55110) );
  IV U67689 ( .A(n55106), .Z(n55108) );
  NOR U67690 ( .A(n55108), .B(n55107), .Z(n55109) );
  NOR U67691 ( .A(n55110), .B(n55109), .Z(n55111) );
  IV U67692 ( .A(n55111), .Z(n55116) );
  IV U67693 ( .A(n55112), .Z(n55114) );
  NOR U67694 ( .A(n55114), .B(n55113), .Z(n55115) );
  NOR U67695 ( .A(n55116), .B(n55115), .Z(n55121) );
  IV U67696 ( .A(n55117), .Z(n55118) );
  NOR U67697 ( .A(n55119), .B(n55118), .Z(n55120) );
  XOR U67698 ( .A(n55121), .B(n55120), .Z(n55122) );
  XOR U67699 ( .A(n55123), .B(n55122), .Z(n58110) );
  IV U67700 ( .A(n55124), .Z(n55127) );
  IV U67701 ( .A(n55132), .Z(n55125) );
  XOR U67702 ( .A(n55128), .B(n55129), .Z(n55131) );
  XOR U67703 ( .A(n55125), .B(n55131), .Z(n55126) );
  NOR U67704 ( .A(n55127), .B(n55126), .Z(n55137) );
  IV U67705 ( .A(n55128), .Z(n55130) );
  NOR U67706 ( .A(n55130), .B(n55129), .Z(n55134) );
  NOR U67707 ( .A(n55132), .B(n55131), .Z(n55133) );
  NOR U67708 ( .A(n55134), .B(n55133), .Z(n55135) );
  IV U67709 ( .A(n55135), .Z(n55136) );
  NOR U67710 ( .A(n55137), .B(n55136), .Z(n58084) );
  IV U67711 ( .A(n55138), .Z(n55140) );
  NOR U67712 ( .A(n55140), .B(n55139), .Z(n55145) );
  IV U67713 ( .A(n55141), .Z(n55143) );
  NOR U67714 ( .A(n55143), .B(n55142), .Z(n55144) );
  NOR U67715 ( .A(n55145), .B(n55144), .Z(n55146) );
  IV U67716 ( .A(n55146), .Z(n55151) );
  IV U67717 ( .A(n55147), .Z(n55149) );
  NOR U67718 ( .A(n55149), .B(n55148), .Z(n55150) );
  NOR U67719 ( .A(n55151), .B(n55150), .Z(n58017) );
  NOR U67720 ( .A(n55153), .B(n55152), .Z(n55154) );
  IV U67721 ( .A(n55154), .Z(n55155) );
  NOR U67722 ( .A(n55156), .B(n55155), .Z(n58015) );
  IV U67723 ( .A(n55157), .Z(n55159) );
  NOR U67724 ( .A(n55159), .B(n55158), .Z(n55163) );
  NOR U67725 ( .A(n55161), .B(n55160), .Z(n55162) );
  NOR U67726 ( .A(n55163), .B(n55162), .Z(n58011) );
  IV U67727 ( .A(n55164), .Z(n55166) );
  NOR U67728 ( .A(n55166), .B(n55165), .Z(n55171) );
  IV U67729 ( .A(n55167), .Z(n55169) );
  NOR U67730 ( .A(n55169), .B(n55168), .Z(n55170) );
  NOR U67731 ( .A(n55171), .B(n55170), .Z(n57882) );
  NOR U67732 ( .A(n55173), .B(n55172), .Z(n55174) );
  NOR U67733 ( .A(n55175), .B(n55174), .Z(n57880) );
  NOR U67734 ( .A(n55178), .B(n55177), .Z(n55184) );
  NOR U67735 ( .A(n55177), .B(n55176), .Z(n55180) );
  IV U67736 ( .A(n55178), .Z(n55179) );
  NOR U67737 ( .A(n55180), .B(n55179), .Z(n55181) );
  NOR U67738 ( .A(n55182), .B(n55181), .Z(n55183) );
  NOR U67739 ( .A(n55184), .B(n55183), .Z(n55188) );
  NOR U67740 ( .A(n55186), .B(n55185), .Z(n55187) );
  NOR U67741 ( .A(n55188), .B(n55187), .Z(n55202) );
  XOR U67742 ( .A(n55195), .B(n55189), .Z(n55193) );
  XOR U67743 ( .A(n55194), .B(n55193), .Z(n55192) );
  IV U67744 ( .A(n55190), .Z(n55191) );
  NOR U67745 ( .A(n55192), .B(n55191), .Z(n55200) );
  NOR U67746 ( .A(n55194), .B(n55193), .Z(n55198) );
  NOR U67747 ( .A(n55196), .B(n55195), .Z(n55197) );
  NOR U67748 ( .A(n55198), .B(n55197), .Z(n55199) );
  XOR U67749 ( .A(n55200), .B(n55199), .Z(n55201) );
  XOR U67750 ( .A(n55202), .B(n55201), .Z(n57852) );
  NOR U67751 ( .A(n55204), .B(n55203), .Z(n55206) );
  XOR U67752 ( .A(n57803), .B(n57804), .Z(n55205) );
  NOR U67753 ( .A(n55206), .B(n55205), .Z(n57814) );
  NOR U67754 ( .A(n55208), .B(n55207), .Z(n55210) );
  NOR U67755 ( .A(n55210), .B(n55209), .Z(n57729) );
  IV U67756 ( .A(n55211), .Z(n55212) );
  NOR U67757 ( .A(n55213), .B(n55212), .Z(n55215) );
  NOR U67758 ( .A(n55215), .B(n55214), .Z(n57727) );
  IV U67759 ( .A(n55219), .Z(n55217) );
  IV U67760 ( .A(n55216), .Z(n55218) );
  NOR U67761 ( .A(n55217), .B(n55218), .Z(n55223) );
  XOR U67762 ( .A(n55219), .B(n55218), .Z(n55221) );
  NOR U67763 ( .A(n55221), .B(n55220), .Z(n55222) );
  NOR U67764 ( .A(n55223), .B(n55222), .Z(n57725) );
  IV U67765 ( .A(n55227), .Z(n55225) );
  IV U67766 ( .A(n55224), .Z(n55226) );
  NOR U67767 ( .A(n55225), .B(n55226), .Z(n55231) );
  XOR U67768 ( .A(n55227), .B(n55226), .Z(n55229) );
  NOR U67769 ( .A(n55229), .B(n55228), .Z(n55230) );
  NOR U67770 ( .A(n55231), .B(n55230), .Z(n57723) );
  IV U67771 ( .A(n55232), .Z(n55234) );
  NOR U67772 ( .A(n55234), .B(n55233), .Z(n57721) );
  IV U67773 ( .A(n55235), .Z(n55238) );
  IV U67774 ( .A(n55236), .Z(n55237) );
  NOR U67775 ( .A(n55238), .B(n55237), .Z(n57719) );
  NOR U67776 ( .A(n55240), .B(n55239), .Z(n55253) );
  NOR U67777 ( .A(n55241), .B(n55242), .Z(n55251) );
  IV U67778 ( .A(n55241), .Z(n55244) );
  IV U67779 ( .A(n55242), .Z(n55243) );
  NOR U67780 ( .A(n55244), .B(n55243), .Z(n55249) );
  NOR U67781 ( .A(n55246), .B(n55245), .Z(n55247) );
  IV U67782 ( .A(n55247), .Z(n55248) );
  NOR U67783 ( .A(n55249), .B(n55248), .Z(n55250) );
  NOR U67784 ( .A(n55251), .B(n55250), .Z(n55252) );
  NOR U67785 ( .A(n55253), .B(n55252), .Z(n57717) );
  IV U67786 ( .A(n55257), .Z(n55255) );
  IV U67787 ( .A(n55256), .Z(n55254) );
  NOR U67788 ( .A(n55255), .B(n55254), .Z(n55263) );
  NOR U67789 ( .A(n55257), .B(n55256), .Z(n55258) );
  NOR U67790 ( .A(n55259), .B(n55258), .Z(n55260) );
  XOR U67791 ( .A(n55261), .B(n55260), .Z(n55262) );
  NOR U67792 ( .A(n55263), .B(n55262), .Z(n57715) );
  IV U67793 ( .A(n55264), .Z(n55265) );
  NOR U67794 ( .A(n55266), .B(n55265), .Z(n55271) );
  IV U67795 ( .A(n55267), .Z(n55268) );
  NOR U67796 ( .A(n55269), .B(n55268), .Z(n55270) );
  NOR U67797 ( .A(n55271), .B(n55270), .Z(n57713) );
  IV U67798 ( .A(n55272), .Z(n55274) );
  NOR U67799 ( .A(n55274), .B(n55273), .Z(n55278) );
  NOR U67800 ( .A(n55276), .B(n55275), .Z(n55277) );
  NOR U67801 ( .A(n55278), .B(n55277), .Z(n57668) );
  IV U67802 ( .A(n55284), .Z(n55282) );
  XOR U67803 ( .A(n55280), .B(n55279), .Z(n55283) );
  IV U67804 ( .A(n55283), .Z(n55281) );
  NOR U67805 ( .A(n55282), .B(n55281), .Z(n55288) );
  NOR U67806 ( .A(n55284), .B(n55283), .Z(n55285) );
  NOR U67807 ( .A(n55286), .B(n55285), .Z(n55287) );
  NOR U67808 ( .A(n55288), .B(n55287), .Z(n57666) );
  NOR U67809 ( .A(n55290), .B(n55289), .Z(n55309) );
  NOR U67810 ( .A(n55292), .B(n55291), .Z(n55297) );
  IV U67811 ( .A(n55293), .Z(n55295) );
  NOR U67812 ( .A(n55295), .B(n55294), .Z(n55296) );
  NOR U67813 ( .A(n55297), .B(n55296), .Z(n55307) );
  IV U67814 ( .A(n55298), .Z(n55299) );
  NOR U67815 ( .A(n55300), .B(n55299), .Z(n55305) );
  IV U67816 ( .A(n55301), .Z(n55303) );
  NOR U67817 ( .A(n55303), .B(n55302), .Z(n55304) );
  NOR U67818 ( .A(n55305), .B(n55304), .Z(n55306) );
  XOR U67819 ( .A(n55307), .B(n55306), .Z(n55308) );
  XOR U67820 ( .A(n55309), .B(n55308), .Z(n57664) );
  IV U67821 ( .A(n55310), .Z(n55312) );
  NOR U67822 ( .A(n55312), .B(n55311), .Z(n55316) );
  IV U67823 ( .A(n55332), .Z(n55314) );
  NOR U67824 ( .A(n55314), .B(n55313), .Z(n55315) );
  NOR U67825 ( .A(n55316), .B(n55315), .Z(n57662) );
  IV U67826 ( .A(n55317), .Z(n55318) );
  NOR U67827 ( .A(n55319), .B(n55318), .Z(n55324) );
  IV U67828 ( .A(n55320), .Z(n55322) );
  NOR U67829 ( .A(n55322), .B(n55321), .Z(n55323) );
  NOR U67830 ( .A(n55324), .B(n55323), .Z(n57660) );
  NOR U67831 ( .A(n55327), .B(n55325), .Z(n55331) );
  XOR U67832 ( .A(n55327), .B(n55326), .Z(n55329) );
  NOR U67833 ( .A(n55329), .B(n55328), .Z(n55330) );
  NOR U67834 ( .A(n55331), .B(n55330), .Z(n57658) );
  NOR U67835 ( .A(n55333), .B(n55332), .Z(n55336) );
  IV U67836 ( .A(n55334), .Z(n55335) );
  NOR U67837 ( .A(n55336), .B(n55335), .Z(n57656) );
  NOR U67838 ( .A(n55338), .B(n55337), .Z(n57654) );
  NOR U67839 ( .A(n55340), .B(n55339), .Z(n55342) );
  NOR U67840 ( .A(n55342), .B(n55341), .Z(n57634) );
  IV U67841 ( .A(n55345), .Z(n55343) );
  NOR U67842 ( .A(n55343), .B(n55344), .Z(n55349) );
  XOR U67843 ( .A(n55345), .B(n55344), .Z(n55347) );
  NOR U67844 ( .A(n55347), .B(n55346), .Z(n55348) );
  NOR U67845 ( .A(n55349), .B(n55348), .Z(n57632) );
  IV U67846 ( .A(n55350), .Z(n55352) );
  NOR U67847 ( .A(n55352), .B(n55351), .Z(n55357) );
  IV U67848 ( .A(n55353), .Z(n55354) );
  NOR U67849 ( .A(n55355), .B(n55354), .Z(n55356) );
  NOR U67850 ( .A(n55357), .B(n55356), .Z(n57630) );
  IV U67851 ( .A(n55360), .Z(n55358) );
  NOR U67852 ( .A(n55359), .B(n55358), .Z(n55365) );
  NOR U67853 ( .A(n55361), .B(n55360), .Z(n55362) );
  NOR U67854 ( .A(n55363), .B(n55362), .Z(n55364) );
  NOR U67855 ( .A(n55365), .B(n55364), .Z(n57628) );
  IV U67856 ( .A(n55366), .Z(n55368) );
  NOR U67857 ( .A(n55368), .B(n55367), .Z(n55372) );
  IV U67858 ( .A(n55369), .Z(n55370) );
  NOR U67859 ( .A(n57619), .B(n55370), .Z(n55371) );
  NOR U67860 ( .A(n55372), .B(n55371), .Z(n55382) );
  IV U67861 ( .A(n55373), .Z(n57616) );
  XOR U67862 ( .A(n57616), .B(n57617), .Z(n55374) );
  NOR U67863 ( .A(n55375), .B(n55374), .Z(n55380) );
  NOR U67864 ( .A(n57616), .B(n55376), .Z(n55377) );
  NOR U67865 ( .A(n55378), .B(n55377), .Z(n55379) );
  NOR U67866 ( .A(n55380), .B(n55379), .Z(n55381) );
  XOR U67867 ( .A(n55382), .B(n55381), .Z(n57607) );
  IV U67868 ( .A(n55383), .Z(n55384) );
  NOR U67869 ( .A(n55385), .B(n55384), .Z(n55390) );
  IV U67870 ( .A(n55386), .Z(n55388) );
  NOR U67871 ( .A(n55388), .B(n55387), .Z(n55389) );
  NOR U67872 ( .A(n55390), .B(n55389), .Z(n57605) );
  IV U67873 ( .A(n55394), .Z(n55392) );
  IV U67874 ( .A(n55393), .Z(n55391) );
  NOR U67875 ( .A(n55392), .B(n55391), .Z(n55398) );
  NOR U67876 ( .A(n55394), .B(n55393), .Z(n55395) );
  NOR U67877 ( .A(n55396), .B(n55395), .Z(n55397) );
  NOR U67878 ( .A(n55398), .B(n55397), .Z(n57603) );
  IV U67879 ( .A(n55402), .Z(n55400) );
  IV U67880 ( .A(n55399), .Z(n55401) );
  NOR U67881 ( .A(n55400), .B(n55401), .Z(n55406) );
  XOR U67882 ( .A(n55402), .B(n55401), .Z(n55404) );
  NOR U67883 ( .A(n55404), .B(n55403), .Z(n55405) );
  NOR U67884 ( .A(n55406), .B(n55405), .Z(n57601) );
  IV U67885 ( .A(n55407), .Z(n55409) );
  NOR U67886 ( .A(n55409), .B(n55408), .Z(n57599) );
  NOR U67887 ( .A(n55411), .B(n55410), .Z(n55413) );
  NOR U67888 ( .A(n55413), .B(n55412), .Z(n57597) );
  IV U67889 ( .A(n55414), .Z(n55415) );
  NOR U67890 ( .A(n55416), .B(n55415), .Z(n57595) );
  IV U67891 ( .A(n55417), .Z(n55419) );
  NOR U67892 ( .A(n55419), .B(n55418), .Z(n55424) );
  IV U67893 ( .A(n55420), .Z(n55421) );
  NOR U67894 ( .A(n55422), .B(n55421), .Z(n55423) );
  NOR U67895 ( .A(n55424), .B(n55423), .Z(n57593) );
  IV U67896 ( .A(n55425), .Z(n55426) );
  NOR U67897 ( .A(n55427), .B(n55426), .Z(n57585) );
  IV U67898 ( .A(n55428), .Z(n55430) );
  NOR U67899 ( .A(n55430), .B(n55429), .Z(n57560) );
  IV U67900 ( .A(n55431), .Z(n55433) );
  IV U67901 ( .A(n55432), .Z(n55442) );
  NOR U67902 ( .A(n55433), .B(n55442), .Z(n55437) );
  IV U67903 ( .A(n55434), .Z(n55435) );
  NOR U67904 ( .A(n55435), .B(n55439), .Z(n55436) );
  NOR U67905 ( .A(n55437), .B(n55436), .Z(n57558) );
  IV U67906 ( .A(n55438), .Z(n55440) );
  NOR U67907 ( .A(n55440), .B(n55439), .Z(n57556) );
  IV U67908 ( .A(n55441), .Z(n55443) );
  NOR U67909 ( .A(n55443), .B(n55442), .Z(n55448) );
  IV U67910 ( .A(n55444), .Z(n55446) );
  NOR U67911 ( .A(n55446), .B(n55445), .Z(n55447) );
  NOR U67912 ( .A(n55448), .B(n55447), .Z(n57554) );
  NOR U67913 ( .A(n55450), .B(n55449), .Z(n55455) );
  IV U67914 ( .A(n55451), .Z(n55453) );
  IV U67915 ( .A(n55479), .Z(n55477) );
  XOR U67916 ( .A(n55477), .B(n55480), .Z(n55452) );
  NOR U67917 ( .A(n55453), .B(n55452), .Z(n55454) );
  NOR U67918 ( .A(n55455), .B(n55454), .Z(n55467) );
  NOR U67919 ( .A(n55457), .B(n55456), .Z(n55459) );
  IV U67920 ( .A(n55461), .Z(n55458) );
  NOR U67921 ( .A(n55459), .B(n55458), .Z(n55465) );
  IV U67922 ( .A(n55459), .Z(n55460) );
  NOR U67923 ( .A(n55461), .B(n55460), .Z(n55462) );
  NOR U67924 ( .A(n55463), .B(n55462), .Z(n55464) );
  NOR U67925 ( .A(n55465), .B(n55464), .Z(n55466) );
  XOR U67926 ( .A(n55467), .B(n55466), .Z(n57552) );
  IV U67927 ( .A(n55468), .Z(n55469) );
  NOR U67928 ( .A(n55470), .B(n55469), .Z(n55474) );
  NOR U67929 ( .A(n55472), .B(n55471), .Z(n55473) );
  NOR U67930 ( .A(n55474), .B(n55473), .Z(n57550) );
  NOR U67931 ( .A(n55476), .B(n55475), .Z(n57548) );
  IV U67932 ( .A(n55480), .Z(n55478) );
  NOR U67933 ( .A(n55478), .B(n55477), .Z(n55486) );
  NOR U67934 ( .A(n55480), .B(n55479), .Z(n55484) );
  NOR U67935 ( .A(n55482), .B(n55481), .Z(n55483) );
  NOR U67936 ( .A(n55484), .B(n55483), .Z(n55485) );
  NOR U67937 ( .A(n55486), .B(n55485), .Z(n57546) );
  NOR U67938 ( .A(n55488), .B(n55487), .Z(n57544) );
  IV U67939 ( .A(n55489), .Z(n55493) );
  NOR U67940 ( .A(n55491), .B(n55490), .Z(n55492) );
  NOR U67941 ( .A(n55493), .B(n55492), .Z(n55494) );
  NOR U67942 ( .A(n55495), .B(n55494), .Z(n57542) );
  IV U67943 ( .A(n55496), .Z(n55497) );
  NOR U67944 ( .A(n55498), .B(n55497), .Z(n55503) );
  IV U67945 ( .A(n55499), .Z(n55501) );
  NOR U67946 ( .A(n55501), .B(n55500), .Z(n55502) );
  NOR U67947 ( .A(n55503), .B(n55502), .Z(n57482) );
  NOR U67948 ( .A(n55505), .B(n55504), .Z(n57480) );
  IV U67949 ( .A(n55506), .Z(n55510) );
  XOR U67950 ( .A(n55510), .B(n57457), .Z(n55507) );
  NOR U67951 ( .A(n55508), .B(n55507), .Z(n55514) );
  NOR U67952 ( .A(n55510), .B(n55509), .Z(n55511) );
  NOR U67953 ( .A(n55512), .B(n55511), .Z(n55513) );
  NOR U67954 ( .A(n55514), .B(n55513), .Z(n57478) );
  NOR U67955 ( .A(n55516), .B(n55515), .Z(n55521) );
  IV U67956 ( .A(n55517), .Z(n55519) );
  NOR U67957 ( .A(n55519), .B(n55518), .Z(n55520) );
  NOR U67958 ( .A(n55521), .B(n55520), .Z(n57450) );
  IV U67959 ( .A(n55522), .Z(n55524) );
  NOR U67960 ( .A(n55524), .B(n55523), .Z(n55529) );
  IV U67961 ( .A(n55525), .Z(n55527) );
  NOR U67962 ( .A(n55527), .B(n55526), .Z(n55528) );
  NOR U67963 ( .A(n55529), .B(n55528), .Z(n57428) );
  IV U67964 ( .A(n55535), .Z(n55530) );
  XOR U67965 ( .A(n55530), .B(n55536), .Z(n55533) );
  XOR U67966 ( .A(n55534), .B(n55533), .Z(n55532) );
  NOR U67967 ( .A(n55532), .B(n55531), .Z(n55540) );
  NOR U67968 ( .A(n55534), .B(n55533), .Z(n55538) );
  NOR U67969 ( .A(n55536), .B(n55535), .Z(n55537) );
  NOR U67970 ( .A(n55538), .B(n55537), .Z(n55539) );
  XOR U67971 ( .A(n55540), .B(n55539), .Z(n57426) );
  IV U67972 ( .A(n55541), .Z(n55543) );
  NOR U67973 ( .A(n55543), .B(n55542), .Z(n55547) );
  NOR U67974 ( .A(n55545), .B(n55544), .Z(n55546) );
  NOR U67975 ( .A(n55547), .B(n55546), .Z(n57424) );
  IV U67976 ( .A(n55548), .Z(n55550) );
  NOR U67977 ( .A(n55550), .B(n55549), .Z(n57422) );
  NOR U67978 ( .A(n55552), .B(n55551), .Z(n55557) );
  IV U67979 ( .A(n55553), .Z(n55555) );
  NOR U67980 ( .A(n55555), .B(n55554), .Z(n55556) );
  NOR U67981 ( .A(n55557), .B(n55556), .Z(n55558) );
  IV U67982 ( .A(n55558), .Z(n55563) );
  IV U67983 ( .A(n55559), .Z(n55561) );
  NOR U67984 ( .A(n55561), .B(n55560), .Z(n55562) );
  NOR U67985 ( .A(n55563), .B(n55562), .Z(n57328) );
  IV U67986 ( .A(n55564), .Z(n55566) );
  NOR U67987 ( .A(n55565), .B(n55566), .Z(n55571) );
  XOR U67988 ( .A(n55567), .B(n55566), .Z(n55569) );
  NOR U67989 ( .A(n55569), .B(n55568), .Z(n55570) );
  NOR U67990 ( .A(n55571), .B(n55570), .Z(n57326) );
  IV U67991 ( .A(n55577), .Z(n55572) );
  XOR U67992 ( .A(n55572), .B(n55578), .Z(n55575) );
  XOR U67993 ( .A(n55576), .B(n55575), .Z(n55574) );
  NOR U67994 ( .A(n55574), .B(n55573), .Z(n55582) );
  NOR U67995 ( .A(n55576), .B(n55575), .Z(n55580) );
  NOR U67996 ( .A(n55578), .B(n55577), .Z(n55579) );
  NOR U67997 ( .A(n55580), .B(n55579), .Z(n55581) );
  XOR U67998 ( .A(n55582), .B(n55581), .Z(n57324) );
  IV U67999 ( .A(n55583), .Z(n55584) );
  NOR U68000 ( .A(n55585), .B(n55584), .Z(n55590) );
  IV U68001 ( .A(n55586), .Z(n55588) );
  NOR U68002 ( .A(n55588), .B(n55587), .Z(n55589) );
  NOR U68003 ( .A(n55590), .B(n55589), .Z(n57322) );
  IV U68004 ( .A(n55591), .Z(n55592) );
  NOR U68005 ( .A(n55593), .B(n55592), .Z(n57320) );
  IV U68006 ( .A(n55594), .Z(n55596) );
  NOR U68007 ( .A(n55596), .B(n55595), .Z(n55601) );
  IV U68008 ( .A(n55597), .Z(n55599) );
  NOR U68009 ( .A(n55599), .B(n55598), .Z(n55600) );
  NOR U68010 ( .A(n55601), .B(n55600), .Z(n57318) );
  IV U68011 ( .A(n55605), .Z(n55602) );
  NOR U68012 ( .A(n55603), .B(n55602), .Z(n55609) );
  IV U68013 ( .A(n55603), .Z(n55604) );
  NOR U68014 ( .A(n55605), .B(n55604), .Z(n55606) );
  NOR U68015 ( .A(n55607), .B(n55606), .Z(n55608) );
  NOR U68016 ( .A(n55609), .B(n55608), .Z(n57316) );
  IV U68017 ( .A(n55610), .Z(n55613) );
  IV U68018 ( .A(n55614), .Z(n55611) );
  NOR U68019 ( .A(n55613), .B(n55611), .Z(n57261) );
  NOR U68020 ( .A(n55612), .B(n55614), .Z(n55620) );
  IV U68021 ( .A(n55612), .Z(n55616) );
  XOR U68022 ( .A(n55614), .B(n55613), .Z(n55615) );
  NOR U68023 ( .A(n55616), .B(n55615), .Z(n55617) );
  NOR U68024 ( .A(n55618), .B(n55617), .Z(n55619) );
  NOR U68025 ( .A(n55620), .B(n55619), .Z(n57259) );
  IV U68026 ( .A(n55621), .Z(n55622) );
  NOR U68027 ( .A(n57244), .B(n55622), .Z(n57242) );
  IV U68028 ( .A(n55623), .Z(n55625) );
  NOR U68029 ( .A(n55625), .B(n55624), .Z(n55631) );
  IV U68030 ( .A(n55626), .Z(n55629) );
  IV U68031 ( .A(n55627), .Z(n55628) );
  NOR U68032 ( .A(n55629), .B(n55628), .Z(n55630) );
  NOR U68033 ( .A(n55631), .B(n55630), .Z(n57240) );
  IV U68034 ( .A(n55634), .Z(n55632) );
  NOR U68035 ( .A(n55632), .B(n55633), .Z(n55638) );
  XOR U68036 ( .A(n55634), .B(n55633), .Z(n55636) );
  NOR U68037 ( .A(n55636), .B(n55635), .Z(n55637) );
  NOR U68038 ( .A(n55638), .B(n55637), .Z(n57238) );
  IV U68039 ( .A(n55639), .Z(n55640) );
  NOR U68040 ( .A(n57219), .B(n55640), .Z(n55642) );
  NOR U68041 ( .A(n55642), .B(n55641), .Z(n57236) );
  NOR U68042 ( .A(n55644), .B(n55643), .Z(n55649) );
  IV U68043 ( .A(n55645), .Z(n55646) );
  NOR U68044 ( .A(n55647), .B(n55646), .Z(n55648) );
  NOR U68045 ( .A(n55649), .B(n55648), .Z(n57234) );
  IV U68046 ( .A(n55650), .Z(n55652) );
  NOR U68047 ( .A(n55652), .B(n55651), .Z(n55653) );
  NOR U68048 ( .A(n55654), .B(n55653), .Z(n57232) );
  IV U68049 ( .A(n55658), .Z(n55656) );
  NOR U68050 ( .A(n55656), .B(n55655), .Z(n55662) );
  NOR U68051 ( .A(n55658), .B(n55657), .Z(n55659) );
  NOR U68052 ( .A(n55660), .B(n55659), .Z(n55661) );
  NOR U68053 ( .A(n55662), .B(n55661), .Z(n57210) );
  IV U68054 ( .A(n55663), .Z(n55665) );
  NOR U68055 ( .A(n55665), .B(n55664), .Z(n55667) );
  NOR U68056 ( .A(n55667), .B(n55666), .Z(n55668) );
  IV U68057 ( .A(n55668), .Z(n55673) );
  IV U68058 ( .A(n55669), .Z(n55680) );
  IV U68059 ( .A(n55670), .Z(n55671) );
  NOR U68060 ( .A(n55680), .B(n55671), .Z(n55672) );
  NOR U68061 ( .A(n55673), .B(n55672), .Z(n57208) );
  IV U68062 ( .A(n55674), .Z(n55675) );
  NOR U68063 ( .A(n55676), .B(n55675), .Z(n55678) );
  NOR U68064 ( .A(n55678), .B(n55677), .Z(n57206) );
  IV U68065 ( .A(n55679), .Z(n55681) );
  NOR U68066 ( .A(n55681), .B(n55680), .Z(n57204) );
  NOR U68067 ( .A(n55683), .B(n55682), .Z(n57202) );
  NOR U68068 ( .A(n55685), .B(n55684), .Z(n57200) );
  NOR U68069 ( .A(n55687), .B(n55686), .Z(n55692) );
  IV U68070 ( .A(n55688), .Z(n55689) );
  NOR U68071 ( .A(n55690), .B(n55689), .Z(n55691) );
  NOR U68072 ( .A(n55692), .B(n55691), .Z(n57198) );
  IV U68073 ( .A(n55693), .Z(n55695) );
  NOR U68074 ( .A(n55695), .B(n55694), .Z(n57186) );
  IV U68075 ( .A(n55696), .Z(n55697) );
  NOR U68076 ( .A(n55698), .B(n55697), .Z(n55703) );
  IV U68077 ( .A(n55699), .Z(n55701) );
  NOR U68078 ( .A(n55701), .B(n55700), .Z(n55702) );
  NOR U68079 ( .A(n55703), .B(n55702), .Z(n57184) );
  IV U68080 ( .A(n55704), .Z(n55707) );
  IV U68081 ( .A(n55705), .Z(n55706) );
  NOR U68082 ( .A(n55707), .B(n55706), .Z(n57182) );
  IV U68083 ( .A(n55708), .Z(n55710) );
  NOR U68084 ( .A(n55710), .B(n55709), .Z(n55714) );
  NOR U68085 ( .A(n55712), .B(n55711), .Z(n55713) );
  NOR U68086 ( .A(n55714), .B(n55713), .Z(n57180) );
  IV U68087 ( .A(n55717), .Z(n55715) );
  NOR U68088 ( .A(n55715), .B(n55716), .Z(n55722) );
  XOR U68089 ( .A(n55717), .B(n55716), .Z(n55720) );
  IV U68090 ( .A(n55718), .Z(n55719) );
  NOR U68091 ( .A(n55720), .B(n55719), .Z(n55721) );
  NOR U68092 ( .A(n55722), .B(n55721), .Z(n57178) );
  IV U68093 ( .A(n55723), .Z(n55724) );
  NOR U68094 ( .A(n55724), .B(n57134), .Z(n55725) );
  NOR U68095 ( .A(n55726), .B(n55725), .Z(n57161) );
  IV U68096 ( .A(n55729), .Z(n55727) );
  NOR U68097 ( .A(n55727), .B(n55728), .Z(n55733) );
  XOR U68098 ( .A(n55729), .B(n55728), .Z(n55731) );
  NOR U68099 ( .A(n55731), .B(n55730), .Z(n55732) );
  NOR U68100 ( .A(n55733), .B(n55732), .Z(n55747) );
  XOR U68101 ( .A(n55740), .B(n55734), .Z(n55738) );
  XOR U68102 ( .A(n55739), .B(n55738), .Z(n55737) );
  IV U68103 ( .A(n55735), .Z(n55736) );
  NOR U68104 ( .A(n55737), .B(n55736), .Z(n55745) );
  NOR U68105 ( .A(n55739), .B(n55738), .Z(n55743) );
  NOR U68106 ( .A(n55741), .B(n55740), .Z(n55742) );
  NOR U68107 ( .A(n55743), .B(n55742), .Z(n55744) );
  XOR U68108 ( .A(n55745), .B(n55744), .Z(n55746) );
  XOR U68109 ( .A(n55747), .B(n55746), .Z(n57129) );
  IV U68110 ( .A(n55750), .Z(n55748) );
  NOR U68111 ( .A(n55748), .B(n55749), .Z(n55752) );
  XOR U68112 ( .A(n55750), .B(n55749), .Z(n55754) );
  NOR U68113 ( .A(n55754), .B(n55753), .Z(n55751) );
  NOR U68114 ( .A(n55752), .B(n55751), .Z(n55759) );
  IV U68115 ( .A(n55753), .Z(n55755) );
  XOR U68116 ( .A(n55755), .B(n55754), .Z(n55756) );
  NOR U68117 ( .A(n55757), .B(n55756), .Z(n55758) );
  XOR U68118 ( .A(n55759), .B(n55758), .Z(n57127) );
  IV U68119 ( .A(n55760), .Z(n55767) );
  XOR U68120 ( .A(n55765), .B(n55767), .Z(n55763) );
  XOR U68121 ( .A(n55764), .B(n55763), .Z(n55762) );
  NOR U68122 ( .A(n55762), .B(n55761), .Z(n55771) );
  NOR U68123 ( .A(n55764), .B(n55763), .Z(n55769) );
  IV U68124 ( .A(n55765), .Z(n55766) );
  NOR U68125 ( .A(n55767), .B(n55766), .Z(n55768) );
  NOR U68126 ( .A(n55769), .B(n55768), .Z(n55770) );
  XOR U68127 ( .A(n55771), .B(n55770), .Z(n57125) );
  IV U68128 ( .A(n55772), .Z(n55774) );
  NOR U68129 ( .A(n55774), .B(n55773), .Z(n55779) );
  IV U68130 ( .A(n55775), .Z(n55777) );
  NOR U68131 ( .A(n55777), .B(n55776), .Z(n55778) );
  NOR U68132 ( .A(n55779), .B(n55778), .Z(n57080) );
  IV U68133 ( .A(n55780), .Z(n55781) );
  NOR U68134 ( .A(n55782), .B(n55781), .Z(n55787) );
  IV U68135 ( .A(n55783), .Z(n55785) );
  NOR U68136 ( .A(n55785), .B(n55784), .Z(n55786) );
  NOR U68137 ( .A(n55787), .B(n55786), .Z(n57041) );
  NOR U68138 ( .A(n55789), .B(n55788), .Z(n57033) );
  IV U68139 ( .A(n55790), .Z(n55791) );
  NOR U68140 ( .A(n55792), .B(n55791), .Z(n55797) );
  IV U68141 ( .A(n55793), .Z(n55794) );
  NOR U68142 ( .A(n55795), .B(n55794), .Z(n55796) );
  NOR U68143 ( .A(n55797), .B(n55796), .Z(n57031) );
  IV U68144 ( .A(n55798), .Z(n55800) );
  NOR U68145 ( .A(n55800), .B(n55799), .Z(n55804) );
  IV U68146 ( .A(n55801), .Z(n55802) );
  NOR U68147 ( .A(n55802), .B(n57005), .Z(n55803) );
  NOR U68148 ( .A(n55804), .B(n55803), .Z(n57011) );
  IV U68149 ( .A(n55808), .Z(n55806) );
  IV U68150 ( .A(n55805), .Z(n55807) );
  NOR U68151 ( .A(n55806), .B(n55807), .Z(n55813) );
  XOR U68152 ( .A(n55808), .B(n55807), .Z(n55811) );
  IV U68153 ( .A(n55809), .Z(n55810) );
  NOR U68154 ( .A(n55811), .B(n55810), .Z(n55812) );
  NOR U68155 ( .A(n55813), .B(n55812), .Z(n56995) );
  IV U68156 ( .A(n55814), .Z(n55815) );
  NOR U68157 ( .A(n55816), .B(n55815), .Z(n55821) );
  IV U68158 ( .A(n55817), .Z(n55818) );
  NOR U68159 ( .A(n55819), .B(n55818), .Z(n55820) );
  NOR U68160 ( .A(n55821), .B(n55820), .Z(n55822) );
  IV U68161 ( .A(n55822), .Z(n55827) );
  IV U68162 ( .A(n55823), .Z(n55825) );
  NOR U68163 ( .A(n55825), .B(n55824), .Z(n55826) );
  NOR U68164 ( .A(n55827), .B(n55826), .Z(n56974) );
  NOR U68165 ( .A(n55829), .B(n55828), .Z(n56972) );
  XOR U68166 ( .A(n55836), .B(n55837), .Z(n55830) );
  IV U68167 ( .A(n55830), .Z(n55834) );
  XOR U68168 ( .A(n55835), .B(n55834), .Z(n55833) );
  IV U68169 ( .A(n55831), .Z(n55832) );
  NOR U68170 ( .A(n55833), .B(n55832), .Z(n55841) );
  NOR U68171 ( .A(n55835), .B(n55834), .Z(n55839) );
  NOR U68172 ( .A(n55837), .B(n55836), .Z(n55838) );
  NOR U68173 ( .A(n55839), .B(n55838), .Z(n55840) );
  XOR U68174 ( .A(n55841), .B(n55840), .Z(n56970) );
  IV U68175 ( .A(n55842), .Z(n55843) );
  NOR U68176 ( .A(n55844), .B(n55843), .Z(n56890) );
  XOR U68177 ( .A(n55845), .B(n55848), .Z(n55847) );
  NOR U68178 ( .A(n55847), .B(n55846), .Z(n55863) );
  NOR U68179 ( .A(n55849), .B(n55848), .Z(n55860) );
  IV U68180 ( .A(n55850), .Z(n55852) );
  NOR U68181 ( .A(n55852), .B(n55851), .Z(n55857) );
  IV U68182 ( .A(n55853), .Z(n55855) );
  NOR U68183 ( .A(n55855), .B(n55854), .Z(n55856) );
  NOR U68184 ( .A(n55857), .B(n55856), .Z(n55858) );
  IV U68185 ( .A(n55858), .Z(n55859) );
  NOR U68186 ( .A(n55860), .B(n55859), .Z(n55861) );
  IV U68187 ( .A(n55861), .Z(n55862) );
  NOR U68188 ( .A(n55863), .B(n55862), .Z(n56888) );
  NOR U68189 ( .A(n55864), .B(n56855), .Z(n56871) );
  IV U68190 ( .A(n55865), .Z(n55866) );
  NOR U68191 ( .A(n55867), .B(n55866), .Z(n55868) );
  NOR U68192 ( .A(n55869), .B(n55868), .Z(n55871) );
  IV U68193 ( .A(n55870), .Z(n56861) );
  NOR U68194 ( .A(n55871), .B(n56861), .Z(n56869) );
  IV U68195 ( .A(n55872), .Z(n55873) );
  NOR U68196 ( .A(n55874), .B(n55873), .Z(n55879) );
  IV U68197 ( .A(n55875), .Z(n55877) );
  NOR U68198 ( .A(n55877), .B(n55876), .Z(n55878) );
  NOR U68199 ( .A(n55879), .B(n55878), .Z(n56841) );
  NOR U68200 ( .A(n55881), .B(n55880), .Z(n56828) );
  IV U68201 ( .A(n55882), .Z(n55883) );
  NOR U68202 ( .A(n55884), .B(n55883), .Z(n55889) );
  IV U68203 ( .A(n55885), .Z(n55887) );
  NOR U68204 ( .A(n55887), .B(n55886), .Z(n55888) );
  NOR U68205 ( .A(n55889), .B(n55888), .Z(n56826) );
  IV U68206 ( .A(n55890), .Z(n55891) );
  NOR U68207 ( .A(n55892), .B(n55891), .Z(n55896) );
  NOR U68208 ( .A(n55894), .B(n55893), .Z(n55895) );
  NOR U68209 ( .A(n55896), .B(n55895), .Z(n56804) );
  XOR U68210 ( .A(n55909), .B(n55915), .Z(n55897) );
  NOR U68211 ( .A(n55898), .B(n55897), .Z(n55899) );
  IV U68212 ( .A(n55899), .Z(n55912) );
  IV U68213 ( .A(n55900), .Z(n55901) );
  NOR U68214 ( .A(n55912), .B(n55901), .Z(n56789) );
  IV U68215 ( .A(n55902), .Z(n55904) );
  NOR U68216 ( .A(n55904), .B(n55903), .Z(n55908) );
  NOR U68217 ( .A(n55906), .B(n55905), .Z(n55907) );
  NOR U68218 ( .A(n55908), .B(n55907), .Z(n56787) );
  IV U68219 ( .A(n55909), .Z(n55910) );
  NOR U68220 ( .A(n55915), .B(n55910), .Z(n56777) );
  IV U68221 ( .A(n55911), .Z(n55913) );
  NOR U68222 ( .A(n55913), .B(n55912), .Z(n55918) );
  IV U68223 ( .A(n55914), .Z(n55916) );
  NOR U68224 ( .A(n55916), .B(n55915), .Z(n55917) );
  NOR U68225 ( .A(n55918), .B(n55917), .Z(n56775) );
  NOR U68226 ( .A(n55920), .B(n55919), .Z(n56773) );
  IV U68227 ( .A(n55921), .Z(n55923) );
  NOR U68228 ( .A(n55923), .B(n55922), .Z(n55928) );
  IV U68229 ( .A(n55924), .Z(n55926) );
  NOR U68230 ( .A(n55926), .B(n55925), .Z(n55927) );
  NOR U68231 ( .A(n55928), .B(n55927), .Z(n56771) );
  IV U68232 ( .A(n55929), .Z(n55930) );
  NOR U68233 ( .A(n55931), .B(n55930), .Z(n55936) );
  IV U68234 ( .A(n55932), .Z(n55933) );
  NOR U68235 ( .A(n55934), .B(n55933), .Z(n55935) );
  NOR U68236 ( .A(n55936), .B(n55935), .Z(n55937) );
  IV U68237 ( .A(n55937), .Z(n55942) );
  IV U68238 ( .A(n55938), .Z(n55940) );
  NOR U68239 ( .A(n55940), .B(n55939), .Z(n55941) );
  NOR U68240 ( .A(n55942), .B(n55941), .Z(n55952) );
  NOR U68241 ( .A(n55944), .B(n55943), .Z(n55946) );
  NOR U68242 ( .A(n55946), .B(n55945), .Z(n55950) );
  NOR U68243 ( .A(n55948), .B(n55947), .Z(n55949) );
  XOR U68244 ( .A(n55950), .B(n55949), .Z(n55951) );
  XOR U68245 ( .A(n55952), .B(n55951), .Z(n56769) );
  IV U68246 ( .A(n55953), .Z(n55955) );
  NOR U68247 ( .A(n55955), .B(n55954), .Z(n55959) );
  NOR U68248 ( .A(n55957), .B(n55956), .Z(n55958) );
  NOR U68249 ( .A(n55959), .B(n55958), .Z(n56767) );
  IV U68250 ( .A(n55960), .Z(n55962) );
  NOR U68251 ( .A(n55962), .B(n55961), .Z(n56765) );
  IV U68252 ( .A(n55966), .Z(n55964) );
  IV U68253 ( .A(n55965), .Z(n55963) );
  NOR U68254 ( .A(n55964), .B(n55963), .Z(n55970) );
  NOR U68255 ( .A(n55966), .B(n55965), .Z(n55967) );
  NOR U68256 ( .A(n55968), .B(n55967), .Z(n55969) );
  NOR U68257 ( .A(n55970), .B(n55969), .Z(n56763) );
  IV U68258 ( .A(n55973), .Z(n55972) );
  IV U68259 ( .A(n55974), .Z(n55971) );
  NOR U68260 ( .A(n55972), .B(n55971), .Z(n55980) );
  NOR U68261 ( .A(n55974), .B(n55973), .Z(n55978) );
  XOR U68262 ( .A(n55976), .B(n55975), .Z(n55977) );
  NOR U68263 ( .A(n55978), .B(n55977), .Z(n55979) );
  NOR U68264 ( .A(n55980), .B(n55979), .Z(n56724) );
  IV U68265 ( .A(n55981), .Z(n55982) );
  NOR U68266 ( .A(n55982), .B(n55989), .Z(n55986) );
  IV U68267 ( .A(n55983), .Z(n55984) );
  XOR U68268 ( .A(n55987), .B(n55989), .Z(n55991) );
  NOR U68269 ( .A(n55984), .B(n55991), .Z(n55985) );
  NOR U68270 ( .A(n55986), .B(n55985), .Z(n56722) );
  IV U68271 ( .A(n55987), .Z(n55988) );
  NOR U68272 ( .A(n55989), .B(n55988), .Z(n56720) );
  IV U68273 ( .A(n55990), .Z(n55992) );
  NOR U68274 ( .A(n55992), .B(n55991), .Z(n56718) );
  IV U68275 ( .A(n55993), .Z(n55994) );
  NOR U68276 ( .A(n55995), .B(n55994), .Z(n56716) );
  IV U68277 ( .A(n55996), .Z(n55997) );
  NOR U68278 ( .A(n55998), .B(n55997), .Z(n56003) );
  IV U68279 ( .A(n55999), .Z(n56000) );
  NOR U68280 ( .A(n56001), .B(n56000), .Z(n56002) );
  NOR U68281 ( .A(n56003), .B(n56002), .Z(n56714) );
  IV U68282 ( .A(n56004), .Z(n56005) );
  NOR U68283 ( .A(n56006), .B(n56005), .Z(n56712) );
  IV U68284 ( .A(n56007), .Z(n56008) );
  NOR U68285 ( .A(n56009), .B(n56008), .Z(n56014) );
  IV U68286 ( .A(n56010), .Z(n56012) );
  NOR U68287 ( .A(n56012), .B(n56011), .Z(n56013) );
  NOR U68288 ( .A(n56014), .B(n56013), .Z(n56710) );
  NOR U68289 ( .A(n56661), .B(n56015), .Z(n56678) );
  IV U68290 ( .A(n56016), .Z(n56018) );
  NOR U68291 ( .A(n56017), .B(n56018), .Z(n56024) );
  XOR U68292 ( .A(n56019), .B(n56018), .Z(n56022) );
  IV U68293 ( .A(n56020), .Z(n56021) );
  NOR U68294 ( .A(n56022), .B(n56021), .Z(n56023) );
  NOR U68295 ( .A(n56024), .B(n56023), .Z(n56620) );
  IV U68296 ( .A(n56025), .Z(n56027) );
  NOR U68297 ( .A(n56027), .B(n56026), .Z(n56618) );
  IV U68298 ( .A(n56028), .Z(n56030) );
  NOR U68299 ( .A(n56030), .B(n56029), .Z(n56035) );
  IV U68300 ( .A(n56031), .Z(n56033) );
  NOR U68301 ( .A(n56033), .B(n56032), .Z(n56034) );
  NOR U68302 ( .A(n56035), .B(n56034), .Z(n56597) );
  IV U68303 ( .A(n56039), .Z(n56037) );
  IV U68304 ( .A(n56036), .Z(n56038) );
  NOR U68305 ( .A(n56037), .B(n56038), .Z(n56043) );
  XOR U68306 ( .A(n56039), .B(n56038), .Z(n56041) );
  NOR U68307 ( .A(n56041), .B(n56040), .Z(n56042) );
  NOR U68308 ( .A(n56043), .B(n56042), .Z(n56595) );
  NOR U68309 ( .A(n56045), .B(n56044), .Z(n56046) );
  IV U68310 ( .A(n56046), .Z(n56047) );
  NOR U68311 ( .A(n56048), .B(n56047), .Z(n56593) );
  IV U68312 ( .A(n56054), .Z(n56049) );
  XOR U68313 ( .A(n56049), .B(n56055), .Z(n56052) );
  XOR U68314 ( .A(n56053), .B(n56052), .Z(n56051) );
  NOR U68315 ( .A(n56051), .B(n56050), .Z(n56059) );
  NOR U68316 ( .A(n56053), .B(n56052), .Z(n56057) );
  NOR U68317 ( .A(n56055), .B(n56054), .Z(n56056) );
  NOR U68318 ( .A(n56057), .B(n56056), .Z(n56058) );
  XOR U68319 ( .A(n56059), .B(n56058), .Z(n56591) );
  IV U68320 ( .A(n56060), .Z(n56062) );
  NOR U68321 ( .A(n56062), .B(n56061), .Z(n56067) );
  IV U68322 ( .A(n56063), .Z(n56065) );
  NOR U68323 ( .A(n56065), .B(n56064), .Z(n56066) );
  NOR U68324 ( .A(n56067), .B(n56066), .Z(n56589) );
  IV U68325 ( .A(n56068), .Z(n56069) );
  NOR U68326 ( .A(n56070), .B(n56069), .Z(n56587) );
  NOR U68327 ( .A(n56072), .B(n56071), .Z(n56583) );
  IV U68328 ( .A(n56082), .Z(n56074) );
  IV U68329 ( .A(n56080), .Z(n56558) );
  XOR U68330 ( .A(n56557), .B(n56558), .Z(n56073) );
  NOR U68331 ( .A(n56074), .B(n56073), .Z(n56075) );
  NOR U68332 ( .A(n56076), .B(n56075), .Z(n56077) );
  IV U68333 ( .A(n56077), .Z(n56078) );
  NOR U68334 ( .A(n56079), .B(n56078), .Z(n56084) );
  XOR U68335 ( .A(n56557), .B(n56080), .Z(n56081) );
  NOR U68336 ( .A(n56082), .B(n56081), .Z(n56083) );
  NOR U68337 ( .A(n56084), .B(n56083), .Z(n56581) );
  NOR U68338 ( .A(n56086), .B(n56085), .Z(n56088) );
  NOR U68339 ( .A(n56088), .B(n56087), .Z(n56554) );
  IV U68340 ( .A(n56089), .Z(n56090) );
  NOR U68341 ( .A(n56091), .B(n56090), .Z(n56552) );
  IV U68342 ( .A(n56095), .Z(n56093) );
  IV U68343 ( .A(n56092), .Z(n56094) );
  NOR U68344 ( .A(n56093), .B(n56094), .Z(n56099) );
  XOR U68345 ( .A(n56095), .B(n56094), .Z(n56097) );
  NOR U68346 ( .A(n56097), .B(n56096), .Z(n56098) );
  NOR U68347 ( .A(n56099), .B(n56098), .Z(n56523) );
  IV U68348 ( .A(n56105), .Z(n56100) );
  XOR U68349 ( .A(n56100), .B(n56106), .Z(n56103) );
  XOR U68350 ( .A(n56104), .B(n56103), .Z(n56102) );
  NOR U68351 ( .A(n56102), .B(n56101), .Z(n56110) );
  NOR U68352 ( .A(n56104), .B(n56103), .Z(n56108) );
  NOR U68353 ( .A(n56106), .B(n56105), .Z(n56107) );
  NOR U68354 ( .A(n56108), .B(n56107), .Z(n56109) );
  XOR U68355 ( .A(n56110), .B(n56109), .Z(n56521) );
  IV U68356 ( .A(n56111), .Z(n56112) );
  NOR U68357 ( .A(n56113), .B(n56112), .Z(n56508) );
  IV U68358 ( .A(n56114), .Z(n56116) );
  NOR U68359 ( .A(n56116), .B(n56115), .Z(n56120) );
  NOR U68360 ( .A(n56118), .B(n56117), .Z(n56119) );
  NOR U68361 ( .A(n56120), .B(n56119), .Z(n56506) );
  IV U68362 ( .A(n56121), .Z(n56123) );
  NOR U68363 ( .A(n56123), .B(n56122), .Z(n56128) );
  IV U68364 ( .A(n56124), .Z(n56126) );
  IV U68365 ( .A(n56125), .Z(n56129) );
  NOR U68366 ( .A(n56126), .B(n56129), .Z(n56127) );
  NOR U68367 ( .A(n56128), .B(n56127), .Z(n56486) );
  NOR U68368 ( .A(n56130), .B(n56129), .Z(n56136) );
  NOR U68369 ( .A(n56132), .B(n56131), .Z(n56133) );
  NOR U68370 ( .A(n56134), .B(n56133), .Z(n56135) );
  NOR U68371 ( .A(n56136), .B(n56135), .Z(n56150) );
  IV U68372 ( .A(n56139), .Z(n56137) );
  NOR U68373 ( .A(n56137), .B(n56138), .Z(n56142) );
  XOR U68374 ( .A(n56139), .B(n56138), .Z(n56143) );
  NOR U68375 ( .A(n56143), .B(n56140), .Z(n56141) );
  NOR U68376 ( .A(n56142), .B(n56141), .Z(n56148) );
  XOR U68377 ( .A(n56144), .B(n56143), .Z(n56146) );
  NOR U68378 ( .A(n56146), .B(n56145), .Z(n56147) );
  XOR U68379 ( .A(n56148), .B(n56147), .Z(n56149) );
  XOR U68380 ( .A(n56150), .B(n56149), .Z(n56484) );
  NOR U68381 ( .A(n56151), .B(n56159), .Z(n56152) );
  NOR U68382 ( .A(n56153), .B(n56152), .Z(n56482) );
  IV U68383 ( .A(n56154), .Z(n56157) );
  XOR U68384 ( .A(n56155), .B(n56159), .Z(n56156) );
  NOR U68385 ( .A(n56157), .B(n56156), .Z(n56162) );
  IV U68386 ( .A(n56158), .Z(n56160) );
  NOR U68387 ( .A(n56160), .B(n56159), .Z(n56161) );
  NOR U68388 ( .A(n56162), .B(n56161), .Z(n56480) );
  IV U68389 ( .A(n56163), .Z(n56165) );
  NOR U68390 ( .A(n56165), .B(n56164), .Z(n56478) );
  IV U68391 ( .A(n56166), .Z(n56167) );
  NOR U68392 ( .A(n56168), .B(n56167), .Z(n56455) );
  NOR U68393 ( .A(n56170), .B(n56169), .Z(n56172) );
  NOR U68394 ( .A(n56172), .B(n56171), .Z(n56453) );
  IV U68395 ( .A(n56173), .Z(n56174) );
  NOR U68396 ( .A(n56175), .B(n56174), .Z(n56451) );
  IV U68397 ( .A(n56176), .Z(n56178) );
  NOR U68398 ( .A(n56178), .B(n56177), .Z(n56182) );
  NOR U68399 ( .A(n56180), .B(n56179), .Z(n56181) );
  NOR U68400 ( .A(n56182), .B(n56181), .Z(n56449) );
  NOR U68401 ( .A(n56184), .B(n56183), .Z(n56437) );
  IV U68402 ( .A(n56185), .Z(n56186) );
  NOR U68403 ( .A(n56186), .B(n56429), .Z(n56191) );
  IV U68404 ( .A(n56187), .Z(n56188) );
  NOR U68405 ( .A(n56189), .B(n56188), .Z(n56190) );
  NOR U68406 ( .A(n56191), .B(n56190), .Z(n56435) );
  IV U68407 ( .A(n56192), .Z(n56194) );
  NOR U68408 ( .A(n56194), .B(n56193), .Z(n56423) );
  IV U68409 ( .A(n56195), .Z(n56199) );
  XOR U68410 ( .A(n56198), .B(n56199), .Z(n56197) );
  NOR U68411 ( .A(n56197), .B(n56196), .Z(n56202) );
  IV U68412 ( .A(n56198), .Z(n56200) );
  NOR U68413 ( .A(n56200), .B(n56199), .Z(n56201) );
  NOR U68414 ( .A(n56202), .B(n56201), .Z(n56421) );
  IV U68415 ( .A(n56203), .Z(n56206) );
  IV U68416 ( .A(n56204), .Z(n56205) );
  NOR U68417 ( .A(n56206), .B(n56205), .Z(n56412) );
  NOR U68418 ( .A(n56208), .B(n56207), .Z(n56213) );
  IV U68419 ( .A(n56209), .Z(n56210) );
  NOR U68420 ( .A(n56211), .B(n56210), .Z(n56212) );
  NOR U68421 ( .A(n56213), .B(n56212), .Z(n56410) );
  IV U68422 ( .A(n56214), .Z(n56216) );
  NOR U68423 ( .A(n56216), .B(n56215), .Z(n56393) );
  IV U68424 ( .A(n56217), .Z(n56219) );
  NOR U68425 ( .A(n56219), .B(n56218), .Z(n56224) );
  IV U68426 ( .A(n56220), .Z(n56222) );
  NOR U68427 ( .A(n56222), .B(n56221), .Z(n56223) );
  NOR U68428 ( .A(n56224), .B(n56223), .Z(n56391) );
  NOR U68429 ( .A(n56226), .B(n56225), .Z(n56231) );
  IV U68430 ( .A(n56227), .Z(n56229) );
  NOR U68431 ( .A(n56229), .B(n56228), .Z(n56230) );
  NOR U68432 ( .A(n56231), .B(n56230), .Z(n56369) );
  IV U68433 ( .A(n56232), .Z(n56234) );
  NOR U68434 ( .A(n56234), .B(n56233), .Z(n56238) );
  NOR U68435 ( .A(n56236), .B(n56235), .Z(n56237) );
  NOR U68436 ( .A(n56238), .B(n56237), .Z(n56277) );
  IV U68437 ( .A(n56239), .Z(n56241) );
  NOR U68438 ( .A(n56241), .B(n56240), .Z(n56269) );
  IV U68439 ( .A(n56242), .Z(n56244) );
  NOR U68440 ( .A(n56244), .B(n56243), .Z(n56249) );
  IV U68441 ( .A(n56245), .Z(n56246) );
  NOR U68442 ( .A(n56247), .B(n56246), .Z(n56248) );
  NOR U68443 ( .A(n56249), .B(n56248), .Z(n56267) );
  IV U68444 ( .A(n56250), .Z(n56252) );
  NOR U68445 ( .A(n56252), .B(n56251), .Z(n56265) );
  IV U68446 ( .A(n56260), .Z(n56253) );
  NOR U68447 ( .A(n56259), .B(n56253), .Z(n56258) );
  NOR U68448 ( .A(n56255), .B(n56254), .Z(n56256) );
  IV U68449 ( .A(n56256), .Z(n56257) );
  NOR U68450 ( .A(n56258), .B(n56257), .Z(n56263) );
  IV U68451 ( .A(n56259), .Z(n56261) );
  NOR U68452 ( .A(n56261), .B(n56260), .Z(n56262) );
  NOR U68453 ( .A(n56263), .B(n56262), .Z(n56264) );
  NOR U68454 ( .A(n56265), .B(n56264), .Z(n56266) );
  XOR U68455 ( .A(n56267), .B(n56266), .Z(n56268) );
  XOR U68456 ( .A(n56269), .B(n56268), .Z(n56275) );
  XOR U68457 ( .A(n56275), .B(n56274), .Z(n56276) );
  XOR U68458 ( .A(n56277), .B(n56276), .Z(n56296) );
  IV U68459 ( .A(n56278), .Z(n56280) );
  NOR U68460 ( .A(n56280), .B(n56279), .Z(n56284) );
  IV U68461 ( .A(n56281), .Z(n56282) );
  NOR U68462 ( .A(n56282), .B(n56340), .Z(n56283) );
  NOR U68463 ( .A(n56284), .B(n56283), .Z(n56294) );
  IV U68464 ( .A(n56285), .Z(n56286) );
  NOR U68465 ( .A(n56287), .B(n56286), .Z(n56292) );
  IV U68466 ( .A(n56288), .Z(n56290) );
  NOR U68467 ( .A(n56290), .B(n56289), .Z(n56291) );
  NOR U68468 ( .A(n56292), .B(n56291), .Z(n56293) );
  XOR U68469 ( .A(n56294), .B(n56293), .Z(n56295) );
  XOR U68470 ( .A(n56296), .B(n56295), .Z(n56302) );
  IV U68471 ( .A(n56297), .Z(n56298) );
  NOR U68472 ( .A(n56323), .B(n56298), .Z(n56299) );
  NOR U68473 ( .A(n56300), .B(n56299), .Z(n56301) );
  XOR U68474 ( .A(n56302), .B(n56301), .Z(n56329) );
  IV U68475 ( .A(n56303), .Z(n56305) );
  NOR U68476 ( .A(n56305), .B(n56304), .Z(n56309) );
  NOR U68477 ( .A(n56307), .B(n56306), .Z(n56308) );
  NOR U68478 ( .A(n56309), .B(n56308), .Z(n56320) );
  IV U68479 ( .A(n56310), .Z(n56312) );
  NOR U68480 ( .A(n56312), .B(n56311), .Z(n56318) );
  NOR U68481 ( .A(n56314), .B(n56313), .Z(n56316) );
  NOR U68482 ( .A(n56316), .B(n56315), .Z(n56317) );
  NOR U68483 ( .A(n56318), .B(n56317), .Z(n56319) );
  XOR U68484 ( .A(n56320), .B(n56319), .Z(n56327) );
  IV U68485 ( .A(n56321), .Z(n56322) );
  NOR U68486 ( .A(n56323), .B(n56322), .Z(n56324) );
  NOR U68487 ( .A(n56325), .B(n56324), .Z(n56326) );
  XOR U68488 ( .A(n56327), .B(n56326), .Z(n56328) );
  XOR U68489 ( .A(n56329), .B(n56328), .Z(n56351) );
  IV U68490 ( .A(n56333), .Z(n56331) );
  IV U68491 ( .A(n56330), .Z(n56332) );
  NOR U68492 ( .A(n56331), .B(n56332), .Z(n56338) );
  XOR U68493 ( .A(n56333), .B(n56332), .Z(n56336) );
  IV U68494 ( .A(n56334), .Z(n56335) );
  NOR U68495 ( .A(n56336), .B(n56335), .Z(n56337) );
  NOR U68496 ( .A(n56338), .B(n56337), .Z(n56349) );
  IV U68497 ( .A(n56339), .Z(n56341) );
  NOR U68498 ( .A(n56341), .B(n56340), .Z(n56347) );
  IV U68499 ( .A(n56342), .Z(n56345) );
  IV U68500 ( .A(n56343), .Z(n56344) );
  NOR U68501 ( .A(n56345), .B(n56344), .Z(n56346) );
  NOR U68502 ( .A(n56347), .B(n56346), .Z(n56348) );
  XOR U68503 ( .A(n56349), .B(n56348), .Z(n56350) );
  XOR U68504 ( .A(n56351), .B(n56350), .Z(n56367) );
  IV U68505 ( .A(n56352), .Z(n56353) );
  NOR U68506 ( .A(n56354), .B(n56353), .Z(n56365) );
  IV U68507 ( .A(n56355), .Z(n56356) );
  NOR U68508 ( .A(n56357), .B(n56356), .Z(n56362) );
  IV U68509 ( .A(n56358), .Z(n56360) );
  NOR U68510 ( .A(n56360), .B(n56359), .Z(n56361) );
  NOR U68511 ( .A(n56362), .B(n56361), .Z(n56363) );
  IV U68512 ( .A(n56363), .Z(n56364) );
  NOR U68513 ( .A(n56365), .B(n56364), .Z(n56366) );
  XOR U68514 ( .A(n56367), .B(n56366), .Z(n56368) );
  XOR U68515 ( .A(n56369), .B(n56368), .Z(n56389) );
  NOR U68516 ( .A(n56371), .B(n56370), .Z(n56376) );
  IV U68517 ( .A(n56372), .Z(n56374) );
  NOR U68518 ( .A(n56374), .B(n56373), .Z(n56375) );
  NOR U68519 ( .A(n56376), .B(n56375), .Z(n56387) );
  IV U68520 ( .A(n56377), .Z(n56379) );
  NOR U68521 ( .A(n56379), .B(n56378), .Z(n56385) );
  IV U68522 ( .A(n56380), .Z(n56383) );
  IV U68523 ( .A(n56381), .Z(n56382) );
  NOR U68524 ( .A(n56383), .B(n56382), .Z(n56384) );
  NOR U68525 ( .A(n56385), .B(n56384), .Z(n56386) );
  XOR U68526 ( .A(n56387), .B(n56386), .Z(n56388) );
  XOR U68527 ( .A(n56389), .B(n56388), .Z(n56390) );
  XOR U68528 ( .A(n56391), .B(n56390), .Z(n56392) );
  XOR U68529 ( .A(n56393), .B(n56392), .Z(n56408) );
  IV U68530 ( .A(n56394), .Z(n56396) );
  NOR U68531 ( .A(n56396), .B(n56395), .Z(n56406) );
  XOR U68532 ( .A(n56397), .B(n56400), .Z(n56399) );
  NOR U68533 ( .A(n56399), .B(n56398), .Z(n56403) );
  NOR U68534 ( .A(n56401), .B(n56400), .Z(n56402) );
  NOR U68535 ( .A(n56403), .B(n56402), .Z(n56404) );
  IV U68536 ( .A(n56404), .Z(n56405) );
  NOR U68537 ( .A(n56406), .B(n56405), .Z(n56407) );
  XOR U68538 ( .A(n56408), .B(n56407), .Z(n56409) );
  XOR U68539 ( .A(n56410), .B(n56409), .Z(n56411) );
  XOR U68540 ( .A(n56412), .B(n56411), .Z(n56419) );
  NOR U68541 ( .A(n56414), .B(n56413), .Z(n56415) );
  IV U68542 ( .A(n56415), .Z(n56416) );
  NOR U68543 ( .A(n56417), .B(n56416), .Z(n56418) );
  XOR U68544 ( .A(n56419), .B(n56418), .Z(n56420) );
  XOR U68545 ( .A(n56421), .B(n56420), .Z(n56422) );
  XOR U68546 ( .A(n56423), .B(n56422), .Z(n56433) );
  NOR U68547 ( .A(n56425), .B(n56424), .Z(n56427) );
  NOR U68548 ( .A(n56427), .B(n56426), .Z(n56431) );
  NOR U68549 ( .A(n56429), .B(n56428), .Z(n56430) );
  NOR U68550 ( .A(n56431), .B(n56430), .Z(n56432) );
  XOR U68551 ( .A(n56433), .B(n56432), .Z(n56434) );
  XOR U68552 ( .A(n56435), .B(n56434), .Z(n56436) );
  XOR U68553 ( .A(n56437), .B(n56436), .Z(n56447) );
  IV U68554 ( .A(n56441), .Z(n56439) );
  IV U68555 ( .A(n56438), .Z(n56440) );
  NOR U68556 ( .A(n56439), .B(n56440), .Z(n56445) );
  XOR U68557 ( .A(n56441), .B(n56440), .Z(n56442) );
  NOR U68558 ( .A(n56443), .B(n56442), .Z(n56444) );
  NOR U68559 ( .A(n56445), .B(n56444), .Z(n56446) );
  XOR U68560 ( .A(n56447), .B(n56446), .Z(n56448) );
  XOR U68561 ( .A(n56449), .B(n56448), .Z(n56450) );
  XOR U68562 ( .A(n56451), .B(n56450), .Z(n56452) );
  XOR U68563 ( .A(n56453), .B(n56452), .Z(n56454) );
  XOR U68564 ( .A(n56455), .B(n56454), .Z(n56476) );
  NOR U68565 ( .A(n56457), .B(n56456), .Z(n56458) );
  NOR U68566 ( .A(n56459), .B(n56458), .Z(n56460) );
  NOR U68567 ( .A(n56461), .B(n56460), .Z(n56467) );
  NOR U68568 ( .A(n56463), .B(n56462), .Z(n56465) );
  NOR U68569 ( .A(n56465), .B(n56464), .Z(n56466) );
  XOR U68570 ( .A(n56467), .B(n56466), .Z(n56474) );
  NOR U68571 ( .A(n56469), .B(n56468), .Z(n56470) );
  IV U68572 ( .A(n56470), .Z(n56471) );
  NOR U68573 ( .A(n56472), .B(n56471), .Z(n56473) );
  XOR U68574 ( .A(n56474), .B(n56473), .Z(n56475) );
  XOR U68575 ( .A(n56476), .B(n56475), .Z(n56477) );
  XOR U68576 ( .A(n56478), .B(n56477), .Z(n56479) );
  XOR U68577 ( .A(n56480), .B(n56479), .Z(n56481) );
  XOR U68578 ( .A(n56482), .B(n56481), .Z(n56483) );
  XOR U68579 ( .A(n56484), .B(n56483), .Z(n56485) );
  XOR U68580 ( .A(n56486), .B(n56485), .Z(n56504) );
  NOR U68581 ( .A(n56488), .B(n56487), .Z(n56493) );
  IV U68582 ( .A(n56489), .Z(n56491) );
  NOR U68583 ( .A(n56491), .B(n56490), .Z(n56492) );
  NOR U68584 ( .A(n56493), .B(n56492), .Z(n56502) );
  IV U68585 ( .A(n56494), .Z(n56496) );
  NOR U68586 ( .A(n56496), .B(n56495), .Z(n56500) );
  NOR U68587 ( .A(n56498), .B(n56497), .Z(n56499) );
  NOR U68588 ( .A(n56500), .B(n56499), .Z(n56501) );
  XOR U68589 ( .A(n56502), .B(n56501), .Z(n56503) );
  XOR U68590 ( .A(n56504), .B(n56503), .Z(n56505) );
  XOR U68591 ( .A(n56506), .B(n56505), .Z(n56507) );
  XOR U68592 ( .A(n56508), .B(n56507), .Z(n56519) );
  IV U68593 ( .A(n56509), .Z(n56512) );
  IV U68594 ( .A(n56510), .Z(n56511) );
  NOR U68595 ( .A(n56512), .B(n56511), .Z(n56517) );
  IV U68596 ( .A(n56513), .Z(n56514) );
  NOR U68597 ( .A(n56515), .B(n56514), .Z(n56516) );
  XOR U68598 ( .A(n56517), .B(n56516), .Z(n56518) );
  XOR U68599 ( .A(n56519), .B(n56518), .Z(n56520) );
  XOR U68600 ( .A(n56521), .B(n56520), .Z(n56522) );
  XOR U68601 ( .A(n56523), .B(n56522), .Z(n56550) );
  IV U68602 ( .A(n56524), .Z(n56526) );
  NOR U68603 ( .A(n56526), .B(n56525), .Z(n56531) );
  IV U68604 ( .A(n56527), .Z(n56528) );
  NOR U68605 ( .A(n56529), .B(n56528), .Z(n56530) );
  NOR U68606 ( .A(n56531), .B(n56530), .Z(n56541) );
  NOR U68607 ( .A(n56535), .B(n56532), .Z(n56539) );
  IV U68608 ( .A(n56533), .Z(n56537) );
  XOR U68609 ( .A(n56535), .B(n56534), .Z(n56536) );
  NOR U68610 ( .A(n56537), .B(n56536), .Z(n56538) );
  NOR U68611 ( .A(n56539), .B(n56538), .Z(n56540) );
  XOR U68612 ( .A(n56541), .B(n56540), .Z(n56548) );
  IV U68613 ( .A(n56542), .Z(n56544) );
  NOR U68614 ( .A(n56544), .B(n56543), .Z(n56545) );
  NOR U68615 ( .A(n56546), .B(n56545), .Z(n56547) );
  XOR U68616 ( .A(n56548), .B(n56547), .Z(n56549) );
  XOR U68617 ( .A(n56550), .B(n56549), .Z(n56551) );
  XOR U68618 ( .A(n56552), .B(n56551), .Z(n56553) );
  XOR U68619 ( .A(n56554), .B(n56553), .Z(n56573) );
  NOR U68620 ( .A(n56556), .B(n56555), .Z(n56561) );
  IV U68621 ( .A(n56557), .Z(n56559) );
  NOR U68622 ( .A(n56559), .B(n56558), .Z(n56560) );
  NOR U68623 ( .A(n56561), .B(n56560), .Z(n56571) );
  IV U68624 ( .A(n56562), .Z(n56564) );
  NOR U68625 ( .A(n56564), .B(n56563), .Z(n56569) );
  IV U68626 ( .A(n56565), .Z(n56566) );
  NOR U68627 ( .A(n56567), .B(n56566), .Z(n56568) );
  NOR U68628 ( .A(n56569), .B(n56568), .Z(n56570) );
  XOR U68629 ( .A(n56571), .B(n56570), .Z(n56572) );
  XOR U68630 ( .A(n56573), .B(n56572), .Z(n56579) );
  NOR U68631 ( .A(n56575), .B(n56574), .Z(n56577) );
  NOR U68632 ( .A(n56577), .B(n56576), .Z(n56578) );
  XOR U68633 ( .A(n56579), .B(n56578), .Z(n56580) );
  XOR U68634 ( .A(n56581), .B(n56580), .Z(n56582) );
  XOR U68635 ( .A(n56583), .B(n56582), .Z(n56584) );
  XOR U68636 ( .A(n56585), .B(n56584), .Z(n56586) );
  XOR U68637 ( .A(n56587), .B(n56586), .Z(n56588) );
  XOR U68638 ( .A(n56589), .B(n56588), .Z(n56590) );
  XOR U68639 ( .A(n56591), .B(n56590), .Z(n56592) );
  XOR U68640 ( .A(n56593), .B(n56592), .Z(n56594) );
  XOR U68641 ( .A(n56595), .B(n56594), .Z(n56596) );
  XOR U68642 ( .A(n56597), .B(n56596), .Z(n56614) );
  IV U68643 ( .A(n56598), .Z(n56600) );
  NOR U68644 ( .A(n56600), .B(n56599), .Z(n56602) );
  NOR U68645 ( .A(n56602), .B(n56601), .Z(n56612) );
  NOR U68646 ( .A(n56604), .B(n56603), .Z(n56610) );
  IV U68647 ( .A(n56605), .Z(n56608) );
  IV U68648 ( .A(n56606), .Z(n56607) );
  NOR U68649 ( .A(n56608), .B(n56607), .Z(n56609) );
  NOR U68650 ( .A(n56610), .B(n56609), .Z(n56611) );
  XOR U68651 ( .A(n56612), .B(n56611), .Z(n56613) );
  XOR U68652 ( .A(n56614), .B(n56613), .Z(n56615) );
  XOR U68653 ( .A(n56616), .B(n56615), .Z(n56617) );
  XOR U68654 ( .A(n56618), .B(n56617), .Z(n56619) );
  XOR U68655 ( .A(n56620), .B(n56619), .Z(n56651) );
  IV U68656 ( .A(n56621), .Z(n56623) );
  NOR U68657 ( .A(n56623), .B(n56622), .Z(n56628) );
  IV U68658 ( .A(n56624), .Z(n56626) );
  NOR U68659 ( .A(n56626), .B(n56625), .Z(n56627) );
  NOR U68660 ( .A(n56628), .B(n56627), .Z(n56649) );
  IV U68661 ( .A(n56629), .Z(n56631) );
  NOR U68662 ( .A(n56631), .B(n56630), .Z(n56637) );
  IV U68663 ( .A(n56632), .Z(n56635) );
  IV U68664 ( .A(n56633), .Z(n56634) );
  NOR U68665 ( .A(n56635), .B(n56634), .Z(n56636) );
  NOR U68666 ( .A(n56637), .B(n56636), .Z(n56647) );
  IV U68667 ( .A(n56638), .Z(n56640) );
  NOR U68668 ( .A(n56639), .B(n56640), .Z(n56645) );
  XOR U68669 ( .A(n56641), .B(n56640), .Z(n56642) );
  NOR U68670 ( .A(n56643), .B(n56642), .Z(n56644) );
  NOR U68671 ( .A(n56645), .B(n56644), .Z(n56646) );
  XOR U68672 ( .A(n56647), .B(n56646), .Z(n56648) );
  XOR U68673 ( .A(n56649), .B(n56648), .Z(n56650) );
  XOR U68674 ( .A(n56651), .B(n56650), .Z(n56676) );
  NOR U68675 ( .A(n56653), .B(n56652), .Z(n56658) );
  IV U68676 ( .A(n56654), .Z(n56655) );
  NOR U68677 ( .A(n56656), .B(n56655), .Z(n56657) );
  NOR U68678 ( .A(n56658), .B(n56657), .Z(n56674) );
  IV U68679 ( .A(n56659), .Z(n56660) );
  NOR U68680 ( .A(n56661), .B(n56660), .Z(n56672) );
  IV U68681 ( .A(n56662), .Z(n56664) );
  NOR U68682 ( .A(n56664), .B(n56663), .Z(n56669) );
  IV U68683 ( .A(n56665), .Z(n56667) );
  NOR U68684 ( .A(n56667), .B(n56666), .Z(n56668) );
  NOR U68685 ( .A(n56669), .B(n56668), .Z(n56670) );
  IV U68686 ( .A(n56670), .Z(n56671) );
  NOR U68687 ( .A(n56672), .B(n56671), .Z(n56673) );
  XOR U68688 ( .A(n56674), .B(n56673), .Z(n56675) );
  XOR U68689 ( .A(n56676), .B(n56675), .Z(n56677) );
  XOR U68690 ( .A(n56678), .B(n56677), .Z(n56698) );
  IV U68691 ( .A(n56679), .Z(n56681) );
  NOR U68692 ( .A(n56681), .B(n56680), .Z(n56686) );
  IV U68693 ( .A(n56682), .Z(n56684) );
  NOR U68694 ( .A(n56684), .B(n56683), .Z(n56685) );
  NOR U68695 ( .A(n56686), .B(n56685), .Z(n56696) );
  NOR U68696 ( .A(n56688), .B(n56687), .Z(n56690) );
  NOR U68697 ( .A(n56689), .B(n56690), .Z(n56694) );
  IV U68698 ( .A(n56690), .Z(n56691) );
  NOR U68699 ( .A(n56692), .B(n56691), .Z(n56693) );
  NOR U68700 ( .A(n56694), .B(n56693), .Z(n56695) );
  XOR U68701 ( .A(n56696), .B(n56695), .Z(n56697) );
  XOR U68702 ( .A(n56698), .B(n56697), .Z(n56708) );
  IV U68703 ( .A(n56702), .Z(n56700) );
  IV U68704 ( .A(n56699), .Z(n56701) );
  NOR U68705 ( .A(n56700), .B(n56701), .Z(n56706) );
  XOR U68706 ( .A(n56702), .B(n56701), .Z(n56703) );
  NOR U68707 ( .A(n56704), .B(n56703), .Z(n56705) );
  NOR U68708 ( .A(n56706), .B(n56705), .Z(n56707) );
  XOR U68709 ( .A(n56708), .B(n56707), .Z(n56709) );
  XOR U68710 ( .A(n56710), .B(n56709), .Z(n56711) );
  XOR U68711 ( .A(n56712), .B(n56711), .Z(n56713) );
  XOR U68712 ( .A(n56714), .B(n56713), .Z(n56715) );
  XOR U68713 ( .A(n56716), .B(n56715), .Z(n56717) );
  XOR U68714 ( .A(n56718), .B(n56717), .Z(n56719) );
  XOR U68715 ( .A(n56720), .B(n56719), .Z(n56721) );
  XOR U68716 ( .A(n56722), .B(n56721), .Z(n56723) );
  XOR U68717 ( .A(n56724), .B(n56723), .Z(n56761) );
  IV U68718 ( .A(n56725), .Z(n56727) );
  NOR U68719 ( .A(n56727), .B(n56726), .Z(n56732) );
  IV U68720 ( .A(n56728), .Z(n56730) );
  NOR U68721 ( .A(n56730), .B(n56729), .Z(n56731) );
  NOR U68722 ( .A(n56732), .B(n56731), .Z(n56759) );
  NOR U68723 ( .A(n56735), .B(n56736), .Z(n56733) );
  NOR U68724 ( .A(n56734), .B(n56733), .Z(n56740) );
  IV U68725 ( .A(n56735), .Z(n56738) );
  IV U68726 ( .A(n56736), .Z(n56737) );
  NOR U68727 ( .A(n56738), .B(n56737), .Z(n56739) );
  NOR U68728 ( .A(n56740), .B(n56739), .Z(n56741) );
  NOR U68729 ( .A(n56742), .B(n56741), .Z(n56750) );
  NOR U68730 ( .A(n56744), .B(n56743), .Z(n56748) );
  NOR U68731 ( .A(n56746), .B(n56745), .Z(n56747) );
  NOR U68732 ( .A(n56748), .B(n56747), .Z(n56749) );
  XOR U68733 ( .A(n56750), .B(n56749), .Z(n56757) );
  IV U68734 ( .A(n56751), .Z(n56752) );
  NOR U68735 ( .A(n56753), .B(n56752), .Z(n56754) );
  NOR U68736 ( .A(n56755), .B(n56754), .Z(n56756) );
  XOR U68737 ( .A(n56757), .B(n56756), .Z(n56758) );
  XOR U68738 ( .A(n56759), .B(n56758), .Z(n56760) );
  XOR U68739 ( .A(n56761), .B(n56760), .Z(n56762) );
  XOR U68740 ( .A(n56763), .B(n56762), .Z(n56764) );
  XOR U68741 ( .A(n56765), .B(n56764), .Z(n56766) );
  XOR U68742 ( .A(n56767), .B(n56766), .Z(n56768) );
  XOR U68743 ( .A(n56769), .B(n56768), .Z(n56770) );
  XOR U68744 ( .A(n56771), .B(n56770), .Z(n56772) );
  XOR U68745 ( .A(n56773), .B(n56772), .Z(n56774) );
  XOR U68746 ( .A(n56775), .B(n56774), .Z(n56776) );
  XOR U68747 ( .A(n56777), .B(n56776), .Z(n56785) );
  IV U68748 ( .A(n56778), .Z(n56779) );
  NOR U68749 ( .A(n56780), .B(n56779), .Z(n56781) );
  IV U68750 ( .A(n56781), .Z(n56782) );
  NOR U68751 ( .A(n56783), .B(n56782), .Z(n56784) );
  XOR U68752 ( .A(n56785), .B(n56784), .Z(n56786) );
  XOR U68753 ( .A(n56787), .B(n56786), .Z(n56788) );
  XOR U68754 ( .A(n56789), .B(n56788), .Z(n56802) );
  IV U68755 ( .A(n56790), .Z(n56792) );
  NOR U68756 ( .A(n56792), .B(n56791), .Z(n56800) );
  IV U68757 ( .A(n56793), .Z(n56795) );
  NOR U68758 ( .A(n56795), .B(n56794), .Z(n56797) );
  NOR U68759 ( .A(n56797), .B(n56796), .Z(n56798) );
  IV U68760 ( .A(n56798), .Z(n56799) );
  NOR U68761 ( .A(n56800), .B(n56799), .Z(n56801) );
  XOR U68762 ( .A(n56802), .B(n56801), .Z(n56803) );
  XOR U68763 ( .A(n56804), .B(n56803), .Z(n56824) );
  IV U68764 ( .A(n56805), .Z(n56806) );
  NOR U68765 ( .A(n56807), .B(n56806), .Z(n56812) );
  IV U68766 ( .A(n56808), .Z(n56810) );
  NOR U68767 ( .A(n56810), .B(n56809), .Z(n56811) );
  NOR U68768 ( .A(n56812), .B(n56811), .Z(n56822) );
  IV U68769 ( .A(n56813), .Z(n56814) );
  NOR U68770 ( .A(n56815), .B(n56814), .Z(n56820) );
  IV U68771 ( .A(n56816), .Z(n56817) );
  NOR U68772 ( .A(n56818), .B(n56817), .Z(n56819) );
  NOR U68773 ( .A(n56820), .B(n56819), .Z(n56821) );
  XOR U68774 ( .A(n56822), .B(n56821), .Z(n56823) );
  XOR U68775 ( .A(n56824), .B(n56823), .Z(n56825) );
  XOR U68776 ( .A(n56826), .B(n56825), .Z(n56827) );
  XOR U68777 ( .A(n56828), .B(n56827), .Z(n56839) );
  IV U68778 ( .A(n56829), .Z(n56832) );
  NOR U68779 ( .A(n56830), .B(n56832), .Z(n56837) );
  IV U68780 ( .A(n56831), .Z(n56835) );
  XOR U68781 ( .A(n56833), .B(n56832), .Z(n56834) );
  NOR U68782 ( .A(n56835), .B(n56834), .Z(n56836) );
  NOR U68783 ( .A(n56837), .B(n56836), .Z(n56838) );
  XOR U68784 ( .A(n56839), .B(n56838), .Z(n56840) );
  XOR U68785 ( .A(n56841), .B(n56840), .Z(n56867) );
  IV U68786 ( .A(n56842), .Z(n56844) );
  NOR U68787 ( .A(n56844), .B(n56843), .Z(n56852) );
  IV U68788 ( .A(n56845), .Z(n56847) );
  NOR U68789 ( .A(n56847), .B(n56846), .Z(n56848) );
  NOR U68790 ( .A(n56849), .B(n56848), .Z(n56850) );
  IV U68791 ( .A(n56850), .Z(n56851) );
  NOR U68792 ( .A(n56852), .B(n56851), .Z(n56865) );
  IV U68793 ( .A(n56853), .Z(n56854) );
  NOR U68794 ( .A(n56855), .B(n56854), .Z(n56863) );
  IV U68795 ( .A(n56856), .Z(n56858) );
  NOR U68796 ( .A(n56858), .B(n56857), .Z(n56859) );
  IV U68797 ( .A(n56859), .Z(n56860) );
  NOR U68798 ( .A(n56861), .B(n56860), .Z(n56862) );
  NOR U68799 ( .A(n56863), .B(n56862), .Z(n56864) );
  XOR U68800 ( .A(n56865), .B(n56864), .Z(n56866) );
  XOR U68801 ( .A(n56867), .B(n56866), .Z(n56868) );
  XOR U68802 ( .A(n56869), .B(n56868), .Z(n56870) );
  XOR U68803 ( .A(n56871), .B(n56870), .Z(n56886) );
  IV U68804 ( .A(n56872), .Z(n56874) );
  NOR U68805 ( .A(n56874), .B(n56873), .Z(n56884) );
  NOR U68806 ( .A(n56876), .B(n56875), .Z(n56881) );
  IV U68807 ( .A(n56877), .Z(n56879) );
  NOR U68808 ( .A(n56879), .B(n56878), .Z(n56880) );
  NOR U68809 ( .A(n56881), .B(n56880), .Z(n56882) );
  IV U68810 ( .A(n56882), .Z(n56883) );
  NOR U68811 ( .A(n56884), .B(n56883), .Z(n56885) );
  XOR U68812 ( .A(n56886), .B(n56885), .Z(n56887) );
  XOR U68813 ( .A(n56888), .B(n56887), .Z(n56889) );
  XOR U68814 ( .A(n56890), .B(n56889), .Z(n56898) );
  IV U68815 ( .A(n56891), .Z(n56894) );
  IV U68816 ( .A(n56892), .Z(n56893) );
  NOR U68817 ( .A(n56894), .B(n56893), .Z(n56895) );
  NOR U68818 ( .A(n56896), .B(n56895), .Z(n56897) );
  XOR U68819 ( .A(n56898), .B(n56897), .Z(n56933) );
  NOR U68820 ( .A(n56900), .B(n56899), .Z(n56905) );
  IV U68821 ( .A(n56901), .Z(n56903) );
  NOR U68822 ( .A(n56903), .B(n56902), .Z(n56904) );
  NOR U68823 ( .A(n56905), .B(n56904), .Z(n56915) );
  IV U68824 ( .A(n56909), .Z(n56907) );
  IV U68825 ( .A(n56906), .Z(n56908) );
  NOR U68826 ( .A(n56907), .B(n56908), .Z(n56913) );
  XOR U68827 ( .A(n56909), .B(n56908), .Z(n56910) );
  NOR U68828 ( .A(n56911), .B(n56910), .Z(n56912) );
  NOR U68829 ( .A(n56913), .B(n56912), .Z(n56914) );
  XOR U68830 ( .A(n56915), .B(n56914), .Z(n56931) );
  IV U68831 ( .A(n56916), .Z(n56918) );
  NOR U68832 ( .A(n56918), .B(n56917), .Z(n56929) );
  IV U68833 ( .A(n56919), .Z(n56920) );
  NOR U68834 ( .A(n56921), .B(n56920), .Z(n56926) );
  IV U68835 ( .A(n56922), .Z(n56924) );
  NOR U68836 ( .A(n56924), .B(n56923), .Z(n56925) );
  NOR U68837 ( .A(n56926), .B(n56925), .Z(n56927) );
  IV U68838 ( .A(n56927), .Z(n56928) );
  NOR U68839 ( .A(n56929), .B(n56928), .Z(n56930) );
  XOR U68840 ( .A(n56931), .B(n56930), .Z(n56932) );
  XOR U68841 ( .A(n56933), .B(n56932), .Z(n56950) );
  IV U68842 ( .A(n56934), .Z(n56936) );
  NOR U68843 ( .A(n56936), .B(n56935), .Z(n56938) );
  NOR U68844 ( .A(n56938), .B(n56937), .Z(n56948) );
  IV U68845 ( .A(n56939), .Z(n56941) );
  NOR U68846 ( .A(n56941), .B(n56940), .Z(n56946) );
  IV U68847 ( .A(n56942), .Z(n56944) );
  NOR U68848 ( .A(n56944), .B(n56943), .Z(n56945) );
  NOR U68849 ( .A(n56946), .B(n56945), .Z(n56947) );
  XOR U68850 ( .A(n56948), .B(n56947), .Z(n56949) );
  XOR U68851 ( .A(n56950), .B(n56949), .Z(n56956) );
  NOR U68852 ( .A(n56952), .B(n56951), .Z(n56954) );
  NOR U68853 ( .A(n56954), .B(n56953), .Z(n56955) );
  XOR U68854 ( .A(n56956), .B(n56955), .Z(n56961) );
  IV U68855 ( .A(n56957), .Z(n56958) );
  NOR U68856 ( .A(n56959), .B(n56958), .Z(n56960) );
  XOR U68857 ( .A(n56961), .B(n56960), .Z(n56968) );
  IV U68858 ( .A(n56962), .Z(n56964) );
  NOR U68859 ( .A(n56964), .B(n56963), .Z(n56965) );
  NOR U68860 ( .A(n56966), .B(n56965), .Z(n56967) );
  XOR U68861 ( .A(n56968), .B(n56967), .Z(n56969) );
  XOR U68862 ( .A(n56970), .B(n56969), .Z(n56971) );
  XOR U68863 ( .A(n56972), .B(n56971), .Z(n56973) );
  XOR U68864 ( .A(n56974), .B(n56973), .Z(n56993) );
  IV U68865 ( .A(n56975), .Z(n56976) );
  NOR U68866 ( .A(n56976), .B(n56997), .Z(n56982) );
  IV U68867 ( .A(n56977), .Z(n56980) );
  IV U68868 ( .A(n56978), .Z(n56979) );
  NOR U68869 ( .A(n56980), .B(n56979), .Z(n56981) );
  NOR U68870 ( .A(n56982), .B(n56981), .Z(n56991) );
  IV U68871 ( .A(n56983), .Z(n56985) );
  NOR U68872 ( .A(n56985), .B(n56984), .Z(n56989) );
  NOR U68873 ( .A(n56987), .B(n56986), .Z(n56988) );
  NOR U68874 ( .A(n56989), .B(n56988), .Z(n56990) );
  XOR U68875 ( .A(n56991), .B(n56990), .Z(n56992) );
  XOR U68876 ( .A(n56993), .B(n56992), .Z(n56994) );
  XOR U68877 ( .A(n56995), .B(n56994), .Z(n57002) );
  IV U68878 ( .A(n56996), .Z(n56998) );
  NOR U68879 ( .A(n56998), .B(n56997), .Z(n56999) );
  NOR U68880 ( .A(n57000), .B(n56999), .Z(n57001) );
  XOR U68881 ( .A(n57002), .B(n57001), .Z(n57009) );
  IV U68882 ( .A(n57003), .Z(n57004) );
  NOR U68883 ( .A(n57005), .B(n57004), .Z(n57006) );
  NOR U68884 ( .A(n57007), .B(n57006), .Z(n57008) );
  XOR U68885 ( .A(n57009), .B(n57008), .Z(n57010) );
  XOR U68886 ( .A(n57011), .B(n57010), .Z(n57029) );
  NOR U68887 ( .A(n57013), .B(n57012), .Z(n57018) );
  IV U68888 ( .A(n57014), .Z(n57015) );
  NOR U68889 ( .A(n57016), .B(n57015), .Z(n57017) );
  NOR U68890 ( .A(n57018), .B(n57017), .Z(n57027) );
  IV U68891 ( .A(n57019), .Z(n57021) );
  NOR U68892 ( .A(n57021), .B(n57020), .Z(n57025) );
  NOR U68893 ( .A(n57023), .B(n57022), .Z(n57024) );
  NOR U68894 ( .A(n57025), .B(n57024), .Z(n57026) );
  XOR U68895 ( .A(n57027), .B(n57026), .Z(n57028) );
  XOR U68896 ( .A(n57029), .B(n57028), .Z(n57030) );
  XOR U68897 ( .A(n57031), .B(n57030), .Z(n57032) );
  XOR U68898 ( .A(n57033), .B(n57032), .Z(n57039) );
  IV U68899 ( .A(n57034), .Z(n57035) );
  NOR U68900 ( .A(n57053), .B(n57035), .Z(n57036) );
  NOR U68901 ( .A(n57037), .B(n57036), .Z(n57038) );
  XOR U68902 ( .A(n57039), .B(n57038), .Z(n57040) );
  XOR U68903 ( .A(n57041), .B(n57040), .Z(n57060) );
  IV U68904 ( .A(n57042), .Z(n57044) );
  NOR U68905 ( .A(n57044), .B(n57043), .Z(n57049) );
  IV U68906 ( .A(n57045), .Z(n57047) );
  NOR U68907 ( .A(n57047), .B(n57046), .Z(n57048) );
  NOR U68908 ( .A(n57049), .B(n57048), .Z(n57058) );
  NOR U68909 ( .A(n57051), .B(n57050), .Z(n57056) );
  IV U68910 ( .A(n57052), .Z(n57054) );
  NOR U68911 ( .A(n57054), .B(n57053), .Z(n57055) );
  NOR U68912 ( .A(n57056), .B(n57055), .Z(n57057) );
  XOR U68913 ( .A(n57058), .B(n57057), .Z(n57059) );
  XOR U68914 ( .A(n57060), .B(n57059), .Z(n57068) );
  IV U68915 ( .A(n57061), .Z(n57064) );
  IV U68916 ( .A(n57062), .Z(n57063) );
  NOR U68917 ( .A(n57064), .B(n57063), .Z(n57065) );
  NOR U68918 ( .A(n57066), .B(n57065), .Z(n57067) );
  XOR U68919 ( .A(n57068), .B(n57067), .Z(n57078) );
  IV U68920 ( .A(n57072), .Z(n57070) );
  IV U68921 ( .A(n57069), .Z(n57071) );
  NOR U68922 ( .A(n57070), .B(n57071), .Z(n57076) );
  XOR U68923 ( .A(n57072), .B(n57071), .Z(n57073) );
  NOR U68924 ( .A(n57074), .B(n57073), .Z(n57075) );
  NOR U68925 ( .A(n57076), .B(n57075), .Z(n57077) );
  XOR U68926 ( .A(n57078), .B(n57077), .Z(n57079) );
  XOR U68927 ( .A(n57080), .B(n57079), .Z(n57099) );
  IV U68928 ( .A(n57084), .Z(n57082) );
  IV U68929 ( .A(n57081), .Z(n57083) );
  NOR U68930 ( .A(n57082), .B(n57083), .Z(n57088) );
  XOR U68931 ( .A(n57084), .B(n57083), .Z(n57086) );
  NOR U68932 ( .A(n57086), .B(n57085), .Z(n57087) );
  NOR U68933 ( .A(n57088), .B(n57087), .Z(n57097) );
  IV U68934 ( .A(n57089), .Z(n57091) );
  NOR U68935 ( .A(n57091), .B(n57090), .Z(n57095) );
  NOR U68936 ( .A(n57093), .B(n57092), .Z(n57094) );
  NOR U68937 ( .A(n57095), .B(n57094), .Z(n57096) );
  XOR U68938 ( .A(n57097), .B(n57096), .Z(n57098) );
  XOR U68939 ( .A(n57099), .B(n57098), .Z(n57123) );
  IV U68940 ( .A(n57100), .Z(n57104) );
  IV U68941 ( .A(n57101), .Z(n57102) );
  NOR U68942 ( .A(n57104), .B(n57102), .Z(n57121) );
  IV U68943 ( .A(n57103), .Z(n57105) );
  NOR U68944 ( .A(n57105), .B(n57104), .Z(n57110) );
  IV U68945 ( .A(n57106), .Z(n57108) );
  NOR U68946 ( .A(n57108), .B(n57107), .Z(n57109) );
  NOR U68947 ( .A(n57110), .B(n57109), .Z(n57119) );
  NOR U68948 ( .A(n57112), .B(n57111), .Z(n57117) );
  IV U68949 ( .A(n57113), .Z(n57115) );
  NOR U68950 ( .A(n57115), .B(n57114), .Z(n57116) );
  NOR U68951 ( .A(n57117), .B(n57116), .Z(n57118) );
  XOR U68952 ( .A(n57119), .B(n57118), .Z(n57120) );
  XOR U68953 ( .A(n57121), .B(n57120), .Z(n57122) );
  XOR U68954 ( .A(n57123), .B(n57122), .Z(n57124) );
  XOR U68955 ( .A(n57125), .B(n57124), .Z(n57126) );
  XOR U68956 ( .A(n57127), .B(n57126), .Z(n57128) );
  XOR U68957 ( .A(n57129), .B(n57128), .Z(n57159) );
  IV U68958 ( .A(n57130), .Z(n57132) );
  NOR U68959 ( .A(n57132), .B(n57131), .Z(n57137) );
  IV U68960 ( .A(n57133), .Z(n57135) );
  NOR U68961 ( .A(n57135), .B(n57134), .Z(n57136) );
  NOR U68962 ( .A(n57137), .B(n57136), .Z(n57157) );
  IV U68963 ( .A(n57138), .Z(n57141) );
  IV U68964 ( .A(n57139), .Z(n57140) );
  NOR U68965 ( .A(n57141), .B(n57140), .Z(n57146) );
  IV U68966 ( .A(n57142), .Z(n57144) );
  NOR U68967 ( .A(n57144), .B(n57143), .Z(n57145) );
  NOR U68968 ( .A(n57146), .B(n57145), .Z(n57155) );
  IV U68969 ( .A(n57149), .Z(n57147) );
  NOR U68970 ( .A(n57147), .B(n57148), .Z(n57153) );
  XOR U68971 ( .A(n57149), .B(n57148), .Z(n57150) );
  NOR U68972 ( .A(n57151), .B(n57150), .Z(n57152) );
  NOR U68973 ( .A(n57153), .B(n57152), .Z(n57154) );
  XOR U68974 ( .A(n57155), .B(n57154), .Z(n57156) );
  XOR U68975 ( .A(n57157), .B(n57156), .Z(n57158) );
  XOR U68976 ( .A(n57159), .B(n57158), .Z(n57160) );
  XOR U68977 ( .A(n57161), .B(n57160), .Z(n57176) );
  NOR U68978 ( .A(n57163), .B(n57162), .Z(n57164) );
  IV U68979 ( .A(n57164), .Z(n57165) );
  NOR U68980 ( .A(n57166), .B(n57165), .Z(n57167) );
  NOR U68981 ( .A(n57168), .B(n57167), .Z(n57174) );
  NOR U68982 ( .A(n57170), .B(n57169), .Z(n57171) );
  NOR U68983 ( .A(n57172), .B(n57171), .Z(n57173) );
  XOR U68984 ( .A(n57174), .B(n57173), .Z(n57175) );
  XOR U68985 ( .A(n57176), .B(n57175), .Z(n57177) );
  XOR U68986 ( .A(n57178), .B(n57177), .Z(n57179) );
  XOR U68987 ( .A(n57180), .B(n57179), .Z(n57181) );
  XOR U68988 ( .A(n57182), .B(n57181), .Z(n57183) );
  XOR U68989 ( .A(n57184), .B(n57183), .Z(n57185) );
  XOR U68990 ( .A(n57186), .B(n57185), .Z(n57196) );
  IV U68991 ( .A(n57190), .Z(n57188) );
  IV U68992 ( .A(n57187), .Z(n57189) );
  NOR U68993 ( .A(n57188), .B(n57189), .Z(n57194) );
  XOR U68994 ( .A(n57190), .B(n57189), .Z(n57191) );
  NOR U68995 ( .A(n57192), .B(n57191), .Z(n57193) );
  NOR U68996 ( .A(n57194), .B(n57193), .Z(n57195) );
  XOR U68997 ( .A(n57196), .B(n57195), .Z(n57197) );
  XOR U68998 ( .A(n57198), .B(n57197), .Z(n57199) );
  XOR U68999 ( .A(n57200), .B(n57199), .Z(n57201) );
  XOR U69000 ( .A(n57202), .B(n57201), .Z(n57203) );
  XOR U69001 ( .A(n57204), .B(n57203), .Z(n57205) );
  XOR U69002 ( .A(n57206), .B(n57205), .Z(n57207) );
  XOR U69003 ( .A(n57208), .B(n57207), .Z(n57209) );
  XOR U69004 ( .A(n57210), .B(n57209), .Z(n57230) );
  NOR U69005 ( .A(n57212), .B(n57211), .Z(n57217) );
  IV U69006 ( .A(n57213), .Z(n57215) );
  NOR U69007 ( .A(n57215), .B(n57214), .Z(n57216) );
  NOR U69008 ( .A(n57217), .B(n57216), .Z(n57228) );
  IV U69009 ( .A(n57218), .Z(n57220) );
  NOR U69010 ( .A(n57220), .B(n57219), .Z(n57226) );
  IV U69011 ( .A(n57221), .Z(n57224) );
  IV U69012 ( .A(n57222), .Z(n57223) );
  NOR U69013 ( .A(n57224), .B(n57223), .Z(n57225) );
  NOR U69014 ( .A(n57226), .B(n57225), .Z(n57227) );
  XOR U69015 ( .A(n57228), .B(n57227), .Z(n57229) );
  XOR U69016 ( .A(n57230), .B(n57229), .Z(n57231) );
  XOR U69017 ( .A(n57232), .B(n57231), .Z(n57233) );
  XOR U69018 ( .A(n57234), .B(n57233), .Z(n57235) );
  XOR U69019 ( .A(n57236), .B(n57235), .Z(n57237) );
  XOR U69020 ( .A(n57238), .B(n57237), .Z(n57239) );
  XOR U69021 ( .A(n57240), .B(n57239), .Z(n57241) );
  XOR U69022 ( .A(n57242), .B(n57241), .Z(n57257) );
  IV U69023 ( .A(n57243), .Z(n57245) );
  NOR U69024 ( .A(n57245), .B(n57244), .Z(n57255) );
  IV U69025 ( .A(n57246), .Z(n57247) );
  NOR U69026 ( .A(n57248), .B(n57247), .Z(n57252) );
  NOR U69027 ( .A(n57250), .B(n57249), .Z(n57251) );
  NOR U69028 ( .A(n57252), .B(n57251), .Z(n57253) );
  IV U69029 ( .A(n57253), .Z(n57254) );
  NOR U69030 ( .A(n57255), .B(n57254), .Z(n57256) );
  XOR U69031 ( .A(n57257), .B(n57256), .Z(n57258) );
  XOR U69032 ( .A(n57259), .B(n57258), .Z(n57260) );
  XOR U69033 ( .A(n57261), .B(n57260), .Z(n57295) );
  NOR U69034 ( .A(n57263), .B(n57262), .Z(n57268) );
  IV U69035 ( .A(n57264), .Z(n57266) );
  NOR U69036 ( .A(n57266), .B(n57265), .Z(n57267) );
  NOR U69037 ( .A(n57268), .B(n57267), .Z(n57293) );
  IV U69038 ( .A(n57269), .Z(n57270) );
  NOR U69039 ( .A(n57271), .B(n57270), .Z(n57291) );
  IV U69040 ( .A(n57272), .Z(n57273) );
  NOR U69041 ( .A(n57274), .B(n57273), .Z(n57279) );
  IV U69042 ( .A(n57275), .Z(n57277) );
  NOR U69043 ( .A(n57277), .B(n57276), .Z(n57278) );
  NOR U69044 ( .A(n57279), .B(n57278), .Z(n57289) );
  IV U69045 ( .A(n57280), .Z(n57282) );
  NOR U69046 ( .A(n57282), .B(n57281), .Z(n57287) );
  IV U69047 ( .A(n57283), .Z(n57285) );
  NOR U69048 ( .A(n57285), .B(n57284), .Z(n57286) );
  NOR U69049 ( .A(n57287), .B(n57286), .Z(n57288) );
  XOR U69050 ( .A(n57289), .B(n57288), .Z(n57290) );
  XOR U69051 ( .A(n57291), .B(n57290), .Z(n57292) );
  XOR U69052 ( .A(n57293), .B(n57292), .Z(n57294) );
  XOR U69053 ( .A(n57295), .B(n57294), .Z(n57314) );
  NOR U69054 ( .A(n57297), .B(n57296), .Z(n57302) );
  IV U69055 ( .A(n57298), .Z(n57300) );
  NOR U69056 ( .A(n57300), .B(n57299), .Z(n57301) );
  NOR U69057 ( .A(n57302), .B(n57301), .Z(n57312) );
  IV U69058 ( .A(n57303), .Z(n57304) );
  NOR U69059 ( .A(n57305), .B(n57304), .Z(n57310) );
  IV U69060 ( .A(n57306), .Z(n57308) );
  NOR U69061 ( .A(n57308), .B(n57307), .Z(n57309) );
  NOR U69062 ( .A(n57310), .B(n57309), .Z(n57311) );
  XOR U69063 ( .A(n57312), .B(n57311), .Z(n57313) );
  XOR U69064 ( .A(n57314), .B(n57313), .Z(n57315) );
  XOR U69065 ( .A(n57316), .B(n57315), .Z(n57317) );
  XOR U69066 ( .A(n57318), .B(n57317), .Z(n57319) );
  XOR U69067 ( .A(n57320), .B(n57319), .Z(n57321) );
  XOR U69068 ( .A(n57322), .B(n57321), .Z(n57323) );
  XOR U69069 ( .A(n57324), .B(n57323), .Z(n57325) );
  XOR U69070 ( .A(n57326), .B(n57325), .Z(n57327) );
  XOR U69071 ( .A(n57328), .B(n57327), .Z(n57359) );
  IV U69072 ( .A(n57329), .Z(n57331) );
  NOR U69073 ( .A(n57331), .B(n57330), .Z(n57337) );
  IV U69074 ( .A(n57332), .Z(n57335) );
  IV U69075 ( .A(n57333), .Z(n57334) );
  NOR U69076 ( .A(n57335), .B(n57334), .Z(n57336) );
  NOR U69077 ( .A(n57337), .B(n57336), .Z(n57357) );
  IV U69078 ( .A(n57338), .Z(n57340) );
  NOR U69079 ( .A(n57340), .B(n57339), .Z(n57345) );
  IV U69080 ( .A(n57341), .Z(n57343) );
  NOR U69081 ( .A(n57343), .B(n57342), .Z(n57344) );
  NOR U69082 ( .A(n57345), .B(n57344), .Z(n57355) );
  IV U69083 ( .A(n57349), .Z(n57347) );
  IV U69084 ( .A(n57346), .Z(n57348) );
  NOR U69085 ( .A(n57347), .B(n57348), .Z(n57353) );
  XOR U69086 ( .A(n57349), .B(n57348), .Z(n57350) );
  NOR U69087 ( .A(n57351), .B(n57350), .Z(n57352) );
  NOR U69088 ( .A(n57353), .B(n57352), .Z(n57354) );
  XOR U69089 ( .A(n57355), .B(n57354), .Z(n57356) );
  XOR U69090 ( .A(n57357), .B(n57356), .Z(n57358) );
  XOR U69091 ( .A(n57359), .B(n57358), .Z(n57396) );
  IV U69092 ( .A(n57360), .Z(n57362) );
  NOR U69093 ( .A(n57362), .B(n57361), .Z(n57366) );
  NOR U69094 ( .A(n57364), .B(n57363), .Z(n57365) );
  NOR U69095 ( .A(n57366), .B(n57365), .Z(n57394) );
  IV U69096 ( .A(n57367), .Z(n57368) );
  NOR U69097 ( .A(n57369), .B(n57368), .Z(n57374) );
  IV U69098 ( .A(n57370), .Z(n57372) );
  NOR U69099 ( .A(n57372), .B(n57371), .Z(n57373) );
  NOR U69100 ( .A(n57374), .B(n57373), .Z(n57383) );
  NOR U69101 ( .A(n57377), .B(n57375), .Z(n57381) );
  XOR U69102 ( .A(n57377), .B(n57376), .Z(n57378) );
  NOR U69103 ( .A(n57379), .B(n57378), .Z(n57380) );
  NOR U69104 ( .A(n57381), .B(n57380), .Z(n57382) );
  XOR U69105 ( .A(n57383), .B(n57382), .Z(n57392) );
  NOR U69106 ( .A(n57386), .B(n57384), .Z(n57390) );
  XOR U69107 ( .A(n57386), .B(n57385), .Z(n57387) );
  NOR U69108 ( .A(n57388), .B(n57387), .Z(n57389) );
  NOR U69109 ( .A(n57390), .B(n57389), .Z(n57391) );
  XOR U69110 ( .A(n57392), .B(n57391), .Z(n57393) );
  XOR U69111 ( .A(n57394), .B(n57393), .Z(n57395) );
  XOR U69112 ( .A(n57396), .B(n57395), .Z(n57420) );
  IV U69113 ( .A(n57397), .Z(n57398) );
  NOR U69114 ( .A(n57399), .B(n57398), .Z(n57418) );
  IV U69115 ( .A(n57400), .Z(n57402) );
  IV U69116 ( .A(n57401), .Z(n57411) );
  NOR U69117 ( .A(n57402), .B(n57411), .Z(n57406) );
  NOR U69118 ( .A(n57404), .B(n57403), .Z(n57405) );
  NOR U69119 ( .A(n57406), .B(n57405), .Z(n57416) );
  IV U69120 ( .A(n57407), .Z(n57408) );
  NOR U69121 ( .A(n57409), .B(n57408), .Z(n57414) );
  IV U69122 ( .A(n57410), .Z(n57412) );
  NOR U69123 ( .A(n57412), .B(n57411), .Z(n57413) );
  NOR U69124 ( .A(n57414), .B(n57413), .Z(n57415) );
  XOR U69125 ( .A(n57416), .B(n57415), .Z(n57417) );
  XOR U69126 ( .A(n57418), .B(n57417), .Z(n57419) );
  XOR U69127 ( .A(n57420), .B(n57419), .Z(n57421) );
  XOR U69128 ( .A(n57422), .B(n57421), .Z(n57423) );
  XOR U69129 ( .A(n57424), .B(n57423), .Z(n57425) );
  XOR U69130 ( .A(n57426), .B(n57425), .Z(n57427) );
  XOR U69131 ( .A(n57428), .B(n57427), .Z(n57448) );
  IV U69132 ( .A(n57429), .Z(n57431) );
  NOR U69133 ( .A(n57431), .B(n57430), .Z(n57436) );
  IV U69134 ( .A(n57432), .Z(n57434) );
  NOR U69135 ( .A(n57434), .B(n57433), .Z(n57435) );
  NOR U69136 ( .A(n57436), .B(n57435), .Z(n57446) );
  IV U69137 ( .A(n57437), .Z(n57439) );
  NOR U69138 ( .A(n57439), .B(n57438), .Z(n57444) );
  IV U69139 ( .A(n57440), .Z(n57442) );
  NOR U69140 ( .A(n57442), .B(n57441), .Z(n57443) );
  NOR U69141 ( .A(n57444), .B(n57443), .Z(n57445) );
  XOR U69142 ( .A(n57446), .B(n57445), .Z(n57447) );
  XOR U69143 ( .A(n57448), .B(n57447), .Z(n57449) );
  XOR U69144 ( .A(n57450), .B(n57449), .Z(n57476) );
  IV U69145 ( .A(n57451), .Z(n57456) );
  XOR U69146 ( .A(n57452), .B(n57456), .Z(n57458) );
  XOR U69147 ( .A(n57453), .B(n57458), .Z(n57454) );
  NOR U69148 ( .A(n57455), .B(n57454), .Z(n57464) );
  NOR U69149 ( .A(n57457), .B(n57456), .Z(n57461) );
  NOR U69150 ( .A(n57459), .B(n57458), .Z(n57460) );
  NOR U69151 ( .A(n57461), .B(n57460), .Z(n57462) );
  IV U69152 ( .A(n57462), .Z(n57463) );
  NOR U69153 ( .A(n57464), .B(n57463), .Z(n57474) );
  IV U69154 ( .A(n57465), .Z(n57466) );
  NOR U69155 ( .A(n57467), .B(n57466), .Z(n57472) );
  IV U69156 ( .A(n57468), .Z(n57470) );
  NOR U69157 ( .A(n57470), .B(n57469), .Z(n57471) );
  NOR U69158 ( .A(n57472), .B(n57471), .Z(n57473) );
  XOR U69159 ( .A(n57474), .B(n57473), .Z(n57475) );
  XOR U69160 ( .A(n57476), .B(n57475), .Z(n57477) );
  XOR U69161 ( .A(n57478), .B(n57477), .Z(n57479) );
  XOR U69162 ( .A(n57480), .B(n57479), .Z(n57481) );
  XOR U69163 ( .A(n57482), .B(n57481), .Z(n57500) );
  NOR U69164 ( .A(n57484), .B(n57483), .Z(n57488) );
  NOR U69165 ( .A(n57486), .B(n57485), .Z(n57487) );
  NOR U69166 ( .A(n57488), .B(n57487), .Z(n57498) );
  IV U69167 ( .A(n57489), .Z(n57490) );
  NOR U69168 ( .A(n57491), .B(n57490), .Z(n57496) );
  IV U69169 ( .A(n57492), .Z(n57494) );
  NOR U69170 ( .A(n57494), .B(n57493), .Z(n57495) );
  NOR U69171 ( .A(n57496), .B(n57495), .Z(n57497) );
  XOR U69172 ( .A(n57498), .B(n57497), .Z(n57499) );
  XOR U69173 ( .A(n57500), .B(n57499), .Z(n57521) );
  IV U69174 ( .A(n57501), .Z(n57502) );
  NOR U69175 ( .A(n57503), .B(n57502), .Z(n57507) );
  IV U69176 ( .A(n57504), .Z(n57505) );
  NOR U69177 ( .A(n57533), .B(n57505), .Z(n57506) );
  NOR U69178 ( .A(n57507), .B(n57506), .Z(n57519) );
  IV U69179 ( .A(n57511), .Z(n57508) );
  NOR U69180 ( .A(n57509), .B(n57508), .Z(n57517) );
  IV U69181 ( .A(n57509), .Z(n57510) );
  NOR U69182 ( .A(n57511), .B(n57510), .Z(n57512) );
  NOR U69183 ( .A(n57513), .B(n57512), .Z(n57514) );
  XOR U69184 ( .A(n57515), .B(n57514), .Z(n57516) );
  NOR U69185 ( .A(n57517), .B(n57516), .Z(n57518) );
  XOR U69186 ( .A(n57519), .B(n57518), .Z(n57520) );
  XOR U69187 ( .A(n57521), .B(n57520), .Z(n57540) );
  IV U69188 ( .A(n57522), .Z(n57524) );
  NOR U69189 ( .A(n57524), .B(n57523), .Z(n57529) );
  IV U69190 ( .A(n57525), .Z(n57527) );
  NOR U69191 ( .A(n57527), .B(n57526), .Z(n57528) );
  NOR U69192 ( .A(n57529), .B(n57528), .Z(n57538) );
  NOR U69193 ( .A(n57531), .B(n57530), .Z(n57536) );
  IV U69194 ( .A(n57532), .Z(n57534) );
  NOR U69195 ( .A(n57534), .B(n57533), .Z(n57535) );
  NOR U69196 ( .A(n57536), .B(n57535), .Z(n57537) );
  XOR U69197 ( .A(n57538), .B(n57537), .Z(n57539) );
  XOR U69198 ( .A(n57540), .B(n57539), .Z(n57541) );
  XOR U69199 ( .A(n57542), .B(n57541), .Z(n57543) );
  XOR U69200 ( .A(n57544), .B(n57543), .Z(n57545) );
  XOR U69201 ( .A(n57546), .B(n57545), .Z(n57547) );
  XOR U69202 ( .A(n57548), .B(n57547), .Z(n57549) );
  XOR U69203 ( .A(n57550), .B(n57549), .Z(n57551) );
  XOR U69204 ( .A(n57552), .B(n57551), .Z(n57553) );
  XOR U69205 ( .A(n57554), .B(n57553), .Z(n57555) );
  XOR U69206 ( .A(n57556), .B(n57555), .Z(n57557) );
  XOR U69207 ( .A(n57558), .B(n57557), .Z(n57559) );
  XOR U69208 ( .A(n57560), .B(n57559), .Z(n57583) );
  IV U69209 ( .A(n57561), .Z(n57562) );
  NOR U69210 ( .A(n57563), .B(n57562), .Z(n57568) );
  IV U69211 ( .A(n57564), .Z(n57566) );
  NOR U69212 ( .A(n57566), .B(n57565), .Z(n57567) );
  NOR U69213 ( .A(n57568), .B(n57567), .Z(n57574) );
  NOR U69214 ( .A(n57570), .B(n57569), .Z(n57572) );
  NOR U69215 ( .A(n57572), .B(n57571), .Z(n57573) );
  XOR U69216 ( .A(n57574), .B(n57573), .Z(n57581) );
  NOR U69217 ( .A(n57576), .B(n57575), .Z(n57577) );
  IV U69218 ( .A(n57577), .Z(n57578) );
  NOR U69219 ( .A(n57579), .B(n57578), .Z(n57580) );
  XOR U69220 ( .A(n57581), .B(n57580), .Z(n57582) );
  XOR U69221 ( .A(n57583), .B(n57582), .Z(n57584) );
  XOR U69222 ( .A(n57585), .B(n57584), .Z(n57591) );
  NOR U69223 ( .A(n57587), .B(n57586), .Z(n57589) );
  NOR U69224 ( .A(n57589), .B(n57588), .Z(n57590) );
  XOR U69225 ( .A(n57591), .B(n57590), .Z(n57592) );
  XOR U69226 ( .A(n57593), .B(n57592), .Z(n57594) );
  XOR U69227 ( .A(n57595), .B(n57594), .Z(n57596) );
  XOR U69228 ( .A(n57597), .B(n57596), .Z(n57598) );
  XOR U69229 ( .A(n57599), .B(n57598), .Z(n57600) );
  XOR U69230 ( .A(n57601), .B(n57600), .Z(n57602) );
  XOR U69231 ( .A(n57603), .B(n57602), .Z(n57604) );
  XOR U69232 ( .A(n57605), .B(n57604), .Z(n57606) );
  XOR U69233 ( .A(n57607), .B(n57606), .Z(n57626) );
  IV U69234 ( .A(n57608), .Z(n57610) );
  NOR U69235 ( .A(n57610), .B(n57609), .Z(n57615) );
  IV U69236 ( .A(n57611), .Z(n57613) );
  NOR U69237 ( .A(n57613), .B(n57612), .Z(n57614) );
  NOR U69238 ( .A(n57615), .B(n57614), .Z(n57624) );
  NOR U69239 ( .A(n57617), .B(n57616), .Z(n57622) );
  IV U69240 ( .A(n57618), .Z(n57620) );
  NOR U69241 ( .A(n57620), .B(n57619), .Z(n57621) );
  NOR U69242 ( .A(n57622), .B(n57621), .Z(n57623) );
  XOR U69243 ( .A(n57624), .B(n57623), .Z(n57625) );
  XOR U69244 ( .A(n57626), .B(n57625), .Z(n57627) );
  XOR U69245 ( .A(n57628), .B(n57627), .Z(n57629) );
  XOR U69246 ( .A(n57630), .B(n57629), .Z(n57631) );
  XOR U69247 ( .A(n57632), .B(n57631), .Z(n57633) );
  XOR U69248 ( .A(n57634), .B(n57633), .Z(n57652) );
  NOR U69249 ( .A(n57636), .B(n57635), .Z(n57640) );
  NOR U69250 ( .A(n57638), .B(n57637), .Z(n57639) );
  NOR U69251 ( .A(n57640), .B(n57639), .Z(n57650) );
  IV U69252 ( .A(n57644), .Z(n57641) );
  NOR U69253 ( .A(n57641), .B(n57643), .Z(n57648) );
  IV U69254 ( .A(n57642), .Z(n57646) );
  XOR U69255 ( .A(n57644), .B(n57643), .Z(n57645) );
  NOR U69256 ( .A(n57646), .B(n57645), .Z(n57647) );
  NOR U69257 ( .A(n57648), .B(n57647), .Z(n57649) );
  XOR U69258 ( .A(n57650), .B(n57649), .Z(n57651) );
  XOR U69259 ( .A(n57652), .B(n57651), .Z(n57653) );
  XOR U69260 ( .A(n57654), .B(n57653), .Z(n57655) );
  XOR U69261 ( .A(n57656), .B(n57655), .Z(n57657) );
  XOR U69262 ( .A(n57658), .B(n57657), .Z(n57659) );
  XOR U69263 ( .A(n57660), .B(n57659), .Z(n57661) );
  XOR U69264 ( .A(n57662), .B(n57661), .Z(n57663) );
  XOR U69265 ( .A(n57664), .B(n57663), .Z(n57665) );
  XOR U69266 ( .A(n57666), .B(n57665), .Z(n57667) );
  XOR U69267 ( .A(n57668), .B(n57667), .Z(n57688) );
  IV U69268 ( .A(n57669), .Z(n57671) );
  NOR U69269 ( .A(n57671), .B(n57670), .Z(n57676) );
  IV U69270 ( .A(n57672), .Z(n57674) );
  NOR U69271 ( .A(n57674), .B(n57673), .Z(n57675) );
  NOR U69272 ( .A(n57676), .B(n57675), .Z(n57686) );
  IV U69273 ( .A(n57677), .Z(n57679) );
  NOR U69274 ( .A(n57679), .B(n57678), .Z(n57684) );
  IV U69275 ( .A(n57680), .Z(n57682) );
  NOR U69276 ( .A(n57682), .B(n57681), .Z(n57683) );
  NOR U69277 ( .A(n57684), .B(n57683), .Z(n57685) );
  XOR U69278 ( .A(n57686), .B(n57685), .Z(n57687) );
  XOR U69279 ( .A(n57688), .B(n57687), .Z(n57697) );
  NOR U69280 ( .A(n57689), .B(n57690), .Z(n57695) );
  XOR U69281 ( .A(n57691), .B(n57690), .Z(n57692) );
  NOR U69282 ( .A(n57693), .B(n57692), .Z(n57694) );
  NOR U69283 ( .A(n57695), .B(n57694), .Z(n57696) );
  XOR U69284 ( .A(n57697), .B(n57696), .Z(n57711) );
  NOR U69285 ( .A(n57699), .B(n57698), .Z(n57709) );
  XOR U69286 ( .A(n57700), .B(n57703), .Z(n57702) );
  NOR U69287 ( .A(n57702), .B(n57701), .Z(n57706) );
  NOR U69288 ( .A(n57704), .B(n57703), .Z(n57705) );
  NOR U69289 ( .A(n57706), .B(n57705), .Z(n57707) );
  IV U69290 ( .A(n57707), .Z(n57708) );
  NOR U69291 ( .A(n57709), .B(n57708), .Z(n57710) );
  XOR U69292 ( .A(n57711), .B(n57710), .Z(n57712) );
  XOR U69293 ( .A(n57713), .B(n57712), .Z(n57714) );
  XOR U69294 ( .A(n57715), .B(n57714), .Z(n57716) );
  XOR U69295 ( .A(n57717), .B(n57716), .Z(n57718) );
  XOR U69296 ( .A(n57719), .B(n57718), .Z(n57720) );
  XOR U69297 ( .A(n57721), .B(n57720), .Z(n57722) );
  XOR U69298 ( .A(n57723), .B(n57722), .Z(n57724) );
  XOR U69299 ( .A(n57725), .B(n57724), .Z(n57726) );
  XOR U69300 ( .A(n57727), .B(n57726), .Z(n57728) );
  XOR U69301 ( .A(n57729), .B(n57728), .Z(n57733) );
  NOR U69302 ( .A(n57731), .B(n57730), .Z(n57732) );
  XOR U69303 ( .A(n57733), .B(n57732), .Z(n57770) );
  XOR U69304 ( .A(n57734), .B(n57737), .Z(n57736) );
  NOR U69305 ( .A(n57736), .B(n57735), .Z(n57752) );
  NOR U69306 ( .A(n57738), .B(n57737), .Z(n57749) );
  IV U69307 ( .A(n57739), .Z(n57741) );
  NOR U69308 ( .A(n57741), .B(n57740), .Z(n57746) );
  IV U69309 ( .A(n57742), .Z(n57744) );
  NOR U69310 ( .A(n57744), .B(n57743), .Z(n57745) );
  NOR U69311 ( .A(n57746), .B(n57745), .Z(n57747) );
  IV U69312 ( .A(n57747), .Z(n57748) );
  NOR U69313 ( .A(n57749), .B(n57748), .Z(n57750) );
  IV U69314 ( .A(n57750), .Z(n57751) );
  NOR U69315 ( .A(n57752), .B(n57751), .Z(n57768) );
  IV U69316 ( .A(n57753), .Z(n57755) );
  NOR U69317 ( .A(n57755), .B(n57754), .Z(n57766) );
  IV U69318 ( .A(n57756), .Z(n57757) );
  NOR U69319 ( .A(n57758), .B(n57757), .Z(n57763) );
  IV U69320 ( .A(n57759), .Z(n57761) );
  NOR U69321 ( .A(n57761), .B(n57760), .Z(n57762) );
  NOR U69322 ( .A(n57763), .B(n57762), .Z(n57764) );
  IV U69323 ( .A(n57764), .Z(n57765) );
  NOR U69324 ( .A(n57766), .B(n57765), .Z(n57767) );
  XOR U69325 ( .A(n57768), .B(n57767), .Z(n57769) );
  XOR U69326 ( .A(n57770), .B(n57769), .Z(n57796) );
  IV U69327 ( .A(n57774), .Z(n57772) );
  IV U69328 ( .A(n57771), .Z(n57773) );
  NOR U69329 ( .A(n57772), .B(n57773), .Z(n57778) );
  XOR U69330 ( .A(n57774), .B(n57773), .Z(n57776) );
  NOR U69331 ( .A(n57776), .B(n57775), .Z(n57777) );
  NOR U69332 ( .A(n57778), .B(n57777), .Z(n57794) );
  IV U69333 ( .A(n57779), .Z(n57784) );
  XOR U69334 ( .A(n57780), .B(n57784), .Z(n57786) );
  XOR U69335 ( .A(n57781), .B(n57786), .Z(n57782) );
  NOR U69336 ( .A(n57783), .B(n57782), .Z(n57792) );
  NOR U69337 ( .A(n57785), .B(n57784), .Z(n57789) );
  NOR U69338 ( .A(n57787), .B(n57786), .Z(n57788) );
  NOR U69339 ( .A(n57789), .B(n57788), .Z(n57790) );
  IV U69340 ( .A(n57790), .Z(n57791) );
  NOR U69341 ( .A(n57792), .B(n57791), .Z(n57793) );
  XOR U69342 ( .A(n57794), .B(n57793), .Z(n57795) );
  XOR U69343 ( .A(n57796), .B(n57795), .Z(n57812) );
  IV U69344 ( .A(n57797), .Z(n57799) );
  NOR U69345 ( .A(n57799), .B(n57798), .Z(n57810) );
  IV U69346 ( .A(n57800), .Z(n57802) );
  NOR U69347 ( .A(n57802), .B(n57801), .Z(n57807) );
  IV U69348 ( .A(n57803), .Z(n57805) );
  NOR U69349 ( .A(n57805), .B(n57804), .Z(n57806) );
  NOR U69350 ( .A(n57807), .B(n57806), .Z(n57808) );
  IV U69351 ( .A(n57808), .Z(n57809) );
  NOR U69352 ( .A(n57810), .B(n57809), .Z(n57811) );
  XOR U69353 ( .A(n57812), .B(n57811), .Z(n57813) );
  XOR U69354 ( .A(n57814), .B(n57813), .Z(n57833) );
  NOR U69355 ( .A(n57816), .B(n57815), .Z(n57821) );
  IV U69356 ( .A(n57817), .Z(n57818) );
  NOR U69357 ( .A(n57819), .B(n57818), .Z(n57820) );
  NOR U69358 ( .A(n57821), .B(n57820), .Z(n57831) );
  IV U69359 ( .A(n57822), .Z(n57825) );
  IV U69360 ( .A(n57823), .Z(n57824) );
  NOR U69361 ( .A(n57825), .B(n57824), .Z(n57829) );
  NOR U69362 ( .A(n57827), .B(n57826), .Z(n57828) );
  NOR U69363 ( .A(n57829), .B(n57828), .Z(n57830) );
  XOR U69364 ( .A(n57831), .B(n57830), .Z(n57832) );
  XOR U69365 ( .A(n57833), .B(n57832), .Z(n57848) );
  IV U69366 ( .A(n57834), .Z(n57835) );
  NOR U69367 ( .A(n57836), .B(n57835), .Z(n57846) );
  NOR U69368 ( .A(n57838), .B(n57837), .Z(n57843) );
  IV U69369 ( .A(n57839), .Z(n57840) );
  NOR U69370 ( .A(n57841), .B(n57840), .Z(n57842) );
  NOR U69371 ( .A(n57843), .B(n57842), .Z(n57844) );
  IV U69372 ( .A(n57844), .Z(n57845) );
  NOR U69373 ( .A(n57846), .B(n57845), .Z(n57847) );
  XOR U69374 ( .A(n57848), .B(n57847), .Z(n57849) );
  XOR U69375 ( .A(n57850), .B(n57849), .Z(n57851) );
  XOR U69376 ( .A(n57852), .B(n57851), .Z(n57878) );
  IV U69377 ( .A(n57853), .Z(n57855) );
  NOR U69378 ( .A(n57855), .B(n57854), .Z(n57860) );
  IV U69379 ( .A(n57856), .Z(n57858) );
  NOR U69380 ( .A(n57858), .B(n57857), .Z(n57859) );
  NOR U69381 ( .A(n57860), .B(n57859), .Z(n57876) );
  IV U69382 ( .A(n57861), .Z(n57863) );
  NOR U69383 ( .A(n57863), .B(n57862), .Z(n57874) );
  IV U69384 ( .A(n57864), .Z(n57866) );
  NOR U69385 ( .A(n57866), .B(n57865), .Z(n57871) );
  IV U69386 ( .A(n57867), .Z(n57868) );
  NOR U69387 ( .A(n57869), .B(n57868), .Z(n57870) );
  NOR U69388 ( .A(n57871), .B(n57870), .Z(n57872) );
  IV U69389 ( .A(n57872), .Z(n57873) );
  NOR U69390 ( .A(n57874), .B(n57873), .Z(n57875) );
  XOR U69391 ( .A(n57876), .B(n57875), .Z(n57877) );
  XOR U69392 ( .A(n57878), .B(n57877), .Z(n57879) );
  XOR U69393 ( .A(n57880), .B(n57879), .Z(n57881) );
  XOR U69394 ( .A(n57882), .B(n57881), .Z(n57911) );
  IV U69395 ( .A(n57883), .Z(n57886) );
  IV U69396 ( .A(n57884), .Z(n57887) );
  XOR U69397 ( .A(n57888), .B(n57887), .Z(n57885) );
  NOR U69398 ( .A(n57886), .B(n57885), .Z(n57894) );
  NOR U69399 ( .A(n57888), .B(n57887), .Z(n57892) );
  NOR U69400 ( .A(n57890), .B(n57889), .Z(n57891) );
  NOR U69401 ( .A(n57892), .B(n57891), .Z(n57893) );
  NOR U69402 ( .A(n57894), .B(n57893), .Z(n57909) );
  XOR U69403 ( .A(n57895), .B(n57898), .Z(n57901) );
  XOR U69404 ( .A(n57900), .B(n57901), .Z(n57896) );
  NOR U69405 ( .A(n57897), .B(n57896), .Z(n57907) );
  NOR U69406 ( .A(n57899), .B(n57898), .Z(n57904) );
  IV U69407 ( .A(n57900), .Z(n57902) );
  NOR U69408 ( .A(n57902), .B(n57901), .Z(n57903) );
  NOR U69409 ( .A(n57904), .B(n57903), .Z(n57905) );
  IV U69410 ( .A(n57905), .Z(n57906) );
  NOR U69411 ( .A(n57907), .B(n57906), .Z(n57908) );
  XOR U69412 ( .A(n57909), .B(n57908), .Z(n57910) );
  XOR U69413 ( .A(n57911), .B(n57910), .Z(n57929) );
  IV U69414 ( .A(n57914), .Z(n57912) );
  NOR U69415 ( .A(n57913), .B(n57912), .Z(n57927) );
  NOR U69416 ( .A(n57915), .B(n57914), .Z(n57918) );
  IV U69417 ( .A(n57916), .Z(n57917) );
  NOR U69418 ( .A(n57918), .B(n57917), .Z(n57923) );
  IV U69419 ( .A(n57919), .Z(n57921) );
  NOR U69420 ( .A(n57921), .B(n57920), .Z(n57922) );
  NOR U69421 ( .A(n57923), .B(n57922), .Z(n57925) );
  NOR U69422 ( .A(n57925), .B(n57924), .Z(n57926) );
  NOR U69423 ( .A(n57927), .B(n57926), .Z(n57928) );
  XOR U69424 ( .A(n57929), .B(n57928), .Z(n57939) );
  IV U69425 ( .A(n57933), .Z(n57931) );
  IV U69426 ( .A(n57930), .Z(n57932) );
  NOR U69427 ( .A(n57931), .B(n57932), .Z(n57937) );
  XOR U69428 ( .A(n57933), .B(n57932), .Z(n57934) );
  NOR U69429 ( .A(n57935), .B(n57934), .Z(n57936) );
  NOR U69430 ( .A(n57937), .B(n57936), .Z(n57938) );
  XOR U69431 ( .A(n57939), .B(n57938), .Z(n57970) );
  NOR U69432 ( .A(n57941), .B(n57940), .Z(n57946) );
  IV U69433 ( .A(n57942), .Z(n57943) );
  NOR U69434 ( .A(n57944), .B(n57943), .Z(n57945) );
  NOR U69435 ( .A(n57946), .B(n57945), .Z(n57961) );
  IV U69436 ( .A(n57947), .Z(n57949) );
  NOR U69437 ( .A(n57949), .B(n57948), .Z(n57959) );
  NOR U69438 ( .A(n57951), .B(n57950), .Z(n57956) );
  IV U69439 ( .A(n57952), .Z(n57954) );
  NOR U69440 ( .A(n57954), .B(n57953), .Z(n57955) );
  NOR U69441 ( .A(n57956), .B(n57955), .Z(n57957) );
  IV U69442 ( .A(n57957), .Z(n57958) );
  NOR U69443 ( .A(n57959), .B(n57958), .Z(n57960) );
  XOR U69444 ( .A(n57961), .B(n57960), .Z(n57968) );
  IV U69445 ( .A(n57962), .Z(n57964) );
  NOR U69446 ( .A(n57964), .B(n57963), .Z(n57965) );
  NOR U69447 ( .A(n57966), .B(n57965), .Z(n57967) );
  XOR U69448 ( .A(n57968), .B(n57967), .Z(n57969) );
  XOR U69449 ( .A(n57970), .B(n57969), .Z(n57989) );
  NOR U69450 ( .A(n57972), .B(n57971), .Z(n57977) );
  IV U69451 ( .A(n57973), .Z(n57974) );
  NOR U69452 ( .A(n57975), .B(n57974), .Z(n57976) );
  NOR U69453 ( .A(n57977), .B(n57976), .Z(n57987) );
  NOR U69454 ( .A(n57979), .B(n57978), .Z(n57985) );
  IV U69455 ( .A(n57980), .Z(n57983) );
  IV U69456 ( .A(n57981), .Z(n57982) );
  NOR U69457 ( .A(n57983), .B(n57982), .Z(n57984) );
  NOR U69458 ( .A(n57985), .B(n57984), .Z(n57986) );
  XOR U69459 ( .A(n57987), .B(n57986), .Z(n57988) );
  XOR U69460 ( .A(n57989), .B(n57988), .Z(n57995) );
  IV U69461 ( .A(n57990), .Z(n57991) );
  NOR U69462 ( .A(n57998), .B(n57991), .Z(n57992) );
  NOR U69463 ( .A(n57993), .B(n57992), .Z(n57994) );
  XOR U69464 ( .A(n57995), .B(n57994), .Z(n58002) );
  IV U69465 ( .A(n57996), .Z(n57997) );
  NOR U69466 ( .A(n57998), .B(n57997), .Z(n58000) );
  NOR U69467 ( .A(n58000), .B(n57999), .Z(n58001) );
  XOR U69468 ( .A(n58002), .B(n58001), .Z(n58009) );
  IV U69469 ( .A(n58003), .Z(n58005) );
  NOR U69470 ( .A(n58005), .B(n58004), .Z(n58006) );
  NOR U69471 ( .A(n58007), .B(n58006), .Z(n58008) );
  XOR U69472 ( .A(n58009), .B(n58008), .Z(n58010) );
  XOR U69473 ( .A(n58011), .B(n58010), .Z(n58012) );
  XOR U69474 ( .A(n58013), .B(n58012), .Z(n58014) );
  XOR U69475 ( .A(n58015), .B(n58014), .Z(n58016) );
  XOR U69476 ( .A(n58017), .B(n58016), .Z(n58066) );
  IV U69477 ( .A(n58018), .Z(n58019) );
  NOR U69478 ( .A(n58020), .B(n58019), .Z(n58025) );
  IV U69479 ( .A(n58021), .Z(n58023) );
  NOR U69480 ( .A(n58023), .B(n58022), .Z(n58024) );
  NOR U69481 ( .A(n58025), .B(n58024), .Z(n58041) );
  IV U69482 ( .A(n58026), .Z(n58028) );
  NOR U69483 ( .A(n58028), .B(n58027), .Z(n58039) );
  IV U69484 ( .A(n58029), .Z(n58031) );
  NOR U69485 ( .A(n58031), .B(n58030), .Z(n58036) );
  IV U69486 ( .A(n58032), .Z(n58034) );
  NOR U69487 ( .A(n58034), .B(n58033), .Z(n58035) );
  NOR U69488 ( .A(n58036), .B(n58035), .Z(n58037) );
  IV U69489 ( .A(n58037), .Z(n58038) );
  NOR U69490 ( .A(n58039), .B(n58038), .Z(n58040) );
  XOR U69491 ( .A(n58041), .B(n58040), .Z(n58051) );
  IV U69492 ( .A(n58045), .Z(n58043) );
  IV U69493 ( .A(n58042), .Z(n58044) );
  NOR U69494 ( .A(n58043), .B(n58044), .Z(n58049) );
  XOR U69495 ( .A(n58045), .B(n58044), .Z(n58046) );
  NOR U69496 ( .A(n58047), .B(n58046), .Z(n58048) );
  NOR U69497 ( .A(n58049), .B(n58048), .Z(n58050) );
  XOR U69498 ( .A(n58051), .B(n58050), .Z(n58064) );
  IV U69499 ( .A(n58054), .Z(n58052) );
  NOR U69500 ( .A(n58053), .B(n58052), .Z(n58062) );
  IV U69501 ( .A(n58053), .Z(n58055) );
  NOR U69502 ( .A(n58055), .B(n58054), .Z(n58060) );
  IV U69503 ( .A(n58056), .Z(n58058) );
  NOR U69504 ( .A(n58058), .B(n58057), .Z(n58059) );
  NOR U69505 ( .A(n58060), .B(n58059), .Z(n58061) );
  NOR U69506 ( .A(n58062), .B(n58061), .Z(n58063) );
  XOR U69507 ( .A(n58064), .B(n58063), .Z(n58065) );
  XOR U69508 ( .A(n58066), .B(n58065), .Z(n58082) );
  IV U69509 ( .A(n58067), .Z(n58069) );
  NOR U69510 ( .A(n58069), .B(n58068), .Z(n58080) );
  IV U69511 ( .A(n58070), .Z(n58072) );
  NOR U69512 ( .A(n58072), .B(n58071), .Z(n58077) );
  IV U69513 ( .A(n58073), .Z(n58075) );
  NOR U69514 ( .A(n58075), .B(n58074), .Z(n58076) );
  NOR U69515 ( .A(n58077), .B(n58076), .Z(n58078) );
  IV U69516 ( .A(n58078), .Z(n58079) );
  NOR U69517 ( .A(n58080), .B(n58079), .Z(n58081) );
  XOR U69518 ( .A(n58082), .B(n58081), .Z(n58083) );
  XOR U69519 ( .A(n58084), .B(n58083), .Z(n58096) );
  IV U69520 ( .A(n58085), .Z(n58087) );
  NOR U69521 ( .A(n58087), .B(n58086), .Z(n58092) );
  IV U69522 ( .A(n58088), .Z(n58090) );
  NOR U69523 ( .A(n58090), .B(n58089), .Z(n58091) );
  NOR U69524 ( .A(n58092), .B(n58091), .Z(n58093) );
  XOR U69525 ( .A(n58094), .B(n58093), .Z(n58095) );
  XOR U69526 ( .A(n58096), .B(n58095), .Z(n58108) );
  NOR U69527 ( .A(n58098), .B(n58097), .Z(n58106) );
  IV U69528 ( .A(n58098), .Z(n58100) );
  NOR U69529 ( .A(n58100), .B(n58099), .Z(n58104) );
  XOR U69530 ( .A(n58102), .B(n58101), .Z(n58103) );
  NOR U69531 ( .A(n58104), .B(n58103), .Z(n58105) );
  NOR U69532 ( .A(n58106), .B(n58105), .Z(n58107) );
  XOR U69533 ( .A(n58108), .B(n58107), .Z(n58109) );
  XOR U69534 ( .A(n58110), .B(n58109), .Z(n58111) );
  XOR U69535 ( .A(n58112), .B(n58111), .Z(n58132) );
  IV U69536 ( .A(n58113), .Z(n58114) );
  NOR U69537 ( .A(n58115), .B(n58114), .Z(n58120) );
  IV U69538 ( .A(n58116), .Z(n58118) );
  NOR U69539 ( .A(n58118), .B(n58117), .Z(n58119) );
  NOR U69540 ( .A(n58120), .B(n58119), .Z(n58130) );
  IV U69541 ( .A(n58121), .Z(n58122) );
  NOR U69542 ( .A(n58123), .B(n58122), .Z(n58128) );
  IV U69543 ( .A(n58124), .Z(n58125) );
  NOR U69544 ( .A(n58126), .B(n58125), .Z(n58127) );
  NOR U69545 ( .A(n58128), .B(n58127), .Z(n58129) );
  XOR U69546 ( .A(n58130), .B(n58129), .Z(n58131) );
  XOR U69547 ( .A(n58132), .B(n58131), .Z(n58143) );
  XOR U69548 ( .A(n58133), .B(n58145), .Z(n58136) );
  IV U69549 ( .A(n58134), .Z(n58135) );
  NOR U69550 ( .A(n58136), .B(n58135), .Z(n58141) );
  IV U69551 ( .A(n58137), .Z(n58138) );
  NOR U69552 ( .A(n58139), .B(n58138), .Z(n58140) );
  NOR U69553 ( .A(n58141), .B(n58140), .Z(n58142) );
  XOR U69554 ( .A(n58143), .B(n58142), .Z(n58163) );
  IV U69555 ( .A(n58144), .Z(n58146) );
  NOR U69556 ( .A(n58146), .B(n58145), .Z(n58151) );
  IV U69557 ( .A(n58147), .Z(n58149) );
  NOR U69558 ( .A(n58149), .B(n58148), .Z(n58150) );
  NOR U69559 ( .A(n58151), .B(n58150), .Z(n58161) );
  IV U69560 ( .A(n58152), .Z(n58154) );
  NOR U69561 ( .A(n58154), .B(n58153), .Z(n58159) );
  IV U69562 ( .A(n58155), .Z(n58157) );
  NOR U69563 ( .A(n58157), .B(n58156), .Z(n58158) );
  NOR U69564 ( .A(n58159), .B(n58158), .Z(n58160) );
  XOR U69565 ( .A(n58161), .B(n58160), .Z(n58162) );
  XOR U69566 ( .A(n58163), .B(n58162), .Z(n58175) );
  IV U69567 ( .A(n58164), .Z(n58166) );
  NOR U69568 ( .A(n58166), .B(n58165), .Z(n58173) );
  IV U69569 ( .A(n58167), .Z(n58168) );
  NOR U69570 ( .A(n58168), .B(n58178), .Z(n58169) );
  NOR U69571 ( .A(n58170), .B(n58169), .Z(n58171) );
  NOR U69572 ( .A(n58171), .B(n58177), .Z(n58172) );
  NOR U69573 ( .A(n58173), .B(n58172), .Z(n58174) );
  XOR U69574 ( .A(n58175), .B(n58174), .Z(n58188) );
  IV U69575 ( .A(n58176), .Z(n58181) );
  NOR U69576 ( .A(n58178), .B(n58177), .Z(n58179) );
  IV U69577 ( .A(n58179), .Z(n58180) );
  NOR U69578 ( .A(n58181), .B(n58180), .Z(n58186) );
  IV U69579 ( .A(n58182), .Z(n58183) );
  NOR U69580 ( .A(n58184), .B(n58183), .Z(n58185) );
  NOR U69581 ( .A(n58186), .B(n58185), .Z(n58187) );
  XOR U69582 ( .A(n58188), .B(n58187), .Z(n58195) );
  IV U69583 ( .A(n58189), .Z(n58191) );
  NOR U69584 ( .A(n58191), .B(n58190), .Z(n58192) );
  NOR U69585 ( .A(n58193), .B(n58192), .Z(n58194) );
  XOR U69586 ( .A(n58195), .B(n58194), .Z(n58210) );
  NOR U69587 ( .A(n58197), .B(n58196), .Z(n58208) );
  IV U69588 ( .A(n58198), .Z(n58199) );
  NOR U69589 ( .A(n58200), .B(n58199), .Z(n58205) );
  IV U69590 ( .A(n58201), .Z(n58203) );
  NOR U69591 ( .A(n58203), .B(n58202), .Z(n58204) );
  NOR U69592 ( .A(n58205), .B(n58204), .Z(n58206) );
  IV U69593 ( .A(n58206), .Z(n58207) );
  NOR U69594 ( .A(n58208), .B(n58207), .Z(n58209) );
  XOR U69595 ( .A(n58210), .B(n58209), .Z(n58211) );
  XOR U69596 ( .A(n58212), .B(n58211), .Z(n58213) );
  XOR U69597 ( .A(n58214), .B(n58213), .Z(n58234) );
  IV U69598 ( .A(n58215), .Z(n58217) );
  NOR U69599 ( .A(n58217), .B(n58216), .Z(n58222) );
  IV U69600 ( .A(n58218), .Z(n58219) );
  NOR U69601 ( .A(n58220), .B(n58219), .Z(n58221) );
  NOR U69602 ( .A(n58222), .B(n58221), .Z(n58232) );
  IV U69603 ( .A(n58226), .Z(n58224) );
  IV U69604 ( .A(n58223), .Z(n58225) );
  NOR U69605 ( .A(n58224), .B(n58225), .Z(n58230) );
  XOR U69606 ( .A(n58226), .B(n58225), .Z(n58227) );
  NOR U69607 ( .A(n58228), .B(n58227), .Z(n58229) );
  NOR U69608 ( .A(n58230), .B(n58229), .Z(n58231) );
  XOR U69609 ( .A(n58232), .B(n58231), .Z(n58233) );
  XOR U69610 ( .A(n58234), .B(n58233), .Z(n58235) );
  XOR U69611 ( .A(n58236), .B(n58235), .Z(n58237) );
  XOR U69612 ( .A(n58238), .B(n58237), .Z(n58239) );
  XOR U69613 ( .A(n58240), .B(n58239), .Z(n58259) );
  IV U69614 ( .A(n58241), .Z(n58242) );
  NOR U69615 ( .A(n58242), .B(n58261), .Z(n58248) );
  IV U69616 ( .A(n58243), .Z(n58246) );
  IV U69617 ( .A(n58244), .Z(n58245) );
  NOR U69618 ( .A(n58246), .B(n58245), .Z(n58247) );
  NOR U69619 ( .A(n58248), .B(n58247), .Z(n58257) );
  NOR U69620 ( .A(n58250), .B(n58249), .Z(n58255) );
  IV U69621 ( .A(n58251), .Z(n58253) );
  NOR U69622 ( .A(n58253), .B(n58252), .Z(n58254) );
  NOR U69623 ( .A(n58255), .B(n58254), .Z(n58256) );
  XOR U69624 ( .A(n58257), .B(n58256), .Z(n58258) );
  XOR U69625 ( .A(n58259), .B(n58258), .Z(n58266) );
  IV U69626 ( .A(n58260), .Z(n58262) );
  NOR U69627 ( .A(n58262), .B(n58261), .Z(n58263) );
  NOR U69628 ( .A(n58264), .B(n58263), .Z(n58265) );
  XOR U69629 ( .A(n58266), .B(n58265), .Z(n58267) );
  XOR U69630 ( .A(n58268), .B(n58267), .Z(n58286) );
  NOR U69631 ( .A(n58270), .B(n58269), .Z(n58271) );
  NOR U69632 ( .A(n58272), .B(n58271), .Z(n58284) );
  IV U69633 ( .A(n58273), .Z(n58276) );
  IV U69634 ( .A(n58274), .Z(n58275) );
  NOR U69635 ( .A(n58276), .B(n58275), .Z(n58282) );
  IV U69636 ( .A(n58277), .Z(n58280) );
  IV U69637 ( .A(n58278), .Z(n58279) );
  NOR U69638 ( .A(n58280), .B(n58279), .Z(n58281) );
  NOR U69639 ( .A(n58282), .B(n58281), .Z(n58283) );
  XOR U69640 ( .A(n58284), .B(n58283), .Z(n58285) );
  XOR U69641 ( .A(n58286), .B(n58285), .Z(n58302) );
  IV U69642 ( .A(n58287), .Z(n58289) );
  IV U69643 ( .A(n58288), .Z(n58311) );
  NOR U69644 ( .A(n58289), .B(n58311), .Z(n58294) );
  IV U69645 ( .A(n58290), .Z(n58291) );
  NOR U69646 ( .A(n58292), .B(n58291), .Z(n58293) );
  NOR U69647 ( .A(n58294), .B(n58293), .Z(n58300) );
  NOR U69648 ( .A(n58296), .B(n58295), .Z(n58297) );
  NOR U69649 ( .A(n58298), .B(n58297), .Z(n58299) );
  XOR U69650 ( .A(n58300), .B(n58299), .Z(n58301) );
  XOR U69651 ( .A(n58302), .B(n58301), .Z(n58321) );
  NOR U69652 ( .A(n58304), .B(n58303), .Z(n58309) );
  IV U69653 ( .A(n58305), .Z(n58306) );
  NOR U69654 ( .A(n58307), .B(n58306), .Z(n58308) );
  NOR U69655 ( .A(n58309), .B(n58308), .Z(n58319) );
  IV U69656 ( .A(n58310), .Z(n58312) );
  NOR U69657 ( .A(n58312), .B(n58311), .Z(n58317) );
  IV U69658 ( .A(n58313), .Z(n58315) );
  NOR U69659 ( .A(n58315), .B(n58314), .Z(n58316) );
  NOR U69660 ( .A(n58317), .B(n58316), .Z(n58318) );
  XOR U69661 ( .A(n58319), .B(n58318), .Z(n58320) );
  XOR U69662 ( .A(n58321), .B(n58320), .Z(n58332) );
  IV U69663 ( .A(n58322), .Z(n58323) );
  NOR U69664 ( .A(n58323), .B(n58347), .Z(n58330) );
  NOR U69665 ( .A(n58325), .B(n58324), .Z(n58326) );
  NOR U69666 ( .A(n58327), .B(n58326), .Z(n58328) );
  IV U69667 ( .A(n58328), .Z(n58329) );
  NOR U69668 ( .A(n58330), .B(n58329), .Z(n58331) );
  XOR U69669 ( .A(n58332), .B(n58331), .Z(n58333) );
  XOR U69670 ( .A(n58334), .B(n58333), .Z(n58354) );
  IV U69671 ( .A(n58335), .Z(n58337) );
  NOR U69672 ( .A(n58337), .B(n58336), .Z(n58342) );
  IV U69673 ( .A(n58338), .Z(n58340) );
  NOR U69674 ( .A(n58340), .B(n58339), .Z(n58341) );
  NOR U69675 ( .A(n58342), .B(n58341), .Z(n58352) );
  IV U69676 ( .A(n58343), .Z(n58345) );
  NOR U69677 ( .A(n58345), .B(n58344), .Z(n58350) );
  IV U69678 ( .A(n58346), .Z(n58348) );
  NOR U69679 ( .A(n58348), .B(n58347), .Z(n58349) );
  NOR U69680 ( .A(n58350), .B(n58349), .Z(n58351) );
  XOR U69681 ( .A(n58352), .B(n58351), .Z(n58353) );
  XOR U69682 ( .A(n58354), .B(n58353), .Z(n58370) );
  IV U69683 ( .A(n58355), .Z(n58357) );
  NOR U69684 ( .A(n58357), .B(n58356), .Z(n58362) );
  IV U69685 ( .A(n58358), .Z(n58359) );
  NOR U69686 ( .A(n58360), .B(n58359), .Z(n58361) );
  NOR U69687 ( .A(n58362), .B(n58361), .Z(n58368) );
  IV U69688 ( .A(n58363), .Z(n58364) );
  NOR U69689 ( .A(n58364), .B(n58379), .Z(n58366) );
  NOR U69690 ( .A(n58366), .B(n58365), .Z(n58367) );
  XOR U69691 ( .A(n58368), .B(n58367), .Z(n58369) );
  XOR U69692 ( .A(n58370), .B(n58369), .Z(n58386) );
  NOR U69693 ( .A(n58372), .B(n58371), .Z(n58374) );
  NOR U69694 ( .A(n58374), .B(n58373), .Z(n58384) );
  IV U69695 ( .A(n58375), .Z(n58377) );
  NOR U69696 ( .A(n58377), .B(n58376), .Z(n58382) );
  IV U69697 ( .A(n58378), .Z(n58380) );
  NOR U69698 ( .A(n58380), .B(n58379), .Z(n58381) );
  NOR U69699 ( .A(n58382), .B(n58381), .Z(n58383) );
  XOR U69700 ( .A(n58384), .B(n58383), .Z(n58385) );
  XOR U69701 ( .A(n58386), .B(n58385), .Z(n58387) );
  XOR U69702 ( .A(n58388), .B(n58387), .Z(n58408) );
  NOR U69703 ( .A(n58390), .B(n58389), .Z(n58395) );
  IV U69704 ( .A(n58391), .Z(n58393) );
  NOR U69705 ( .A(n58393), .B(n58392), .Z(n58394) );
  NOR U69706 ( .A(n58395), .B(n58394), .Z(n58406) );
  IV U69707 ( .A(n58396), .Z(n58398) );
  NOR U69708 ( .A(n58398), .B(n58397), .Z(n58404) );
  IV U69709 ( .A(n58399), .Z(n58402) );
  IV U69710 ( .A(n58400), .Z(n58401) );
  NOR U69711 ( .A(n58402), .B(n58401), .Z(n58403) );
  NOR U69712 ( .A(n58404), .B(n58403), .Z(n58405) );
  XOR U69713 ( .A(n58406), .B(n58405), .Z(n58407) );
  XOR U69714 ( .A(n58408), .B(n58407), .Z(n58409) );
  XOR U69715 ( .A(n58410), .B(n58409), .Z(n58411) );
  XOR U69716 ( .A(n58412), .B(n58411), .Z(n58421) );
  NOR U69717 ( .A(n58413), .B(n58414), .Z(n58419) );
  XOR U69718 ( .A(n58415), .B(n58414), .Z(n58416) );
  NOR U69719 ( .A(n58417), .B(n58416), .Z(n58418) );
  NOR U69720 ( .A(n58419), .B(n58418), .Z(n58420) );
  XOR U69721 ( .A(n58421), .B(n58420), .Z(n58437) );
  IV U69722 ( .A(n58422), .Z(n58424) );
  NOR U69723 ( .A(n58424), .B(n58423), .Z(n58435) );
  IV U69724 ( .A(n58425), .Z(n58427) );
  NOR U69725 ( .A(n58427), .B(n58426), .Z(n58432) );
  IV U69726 ( .A(n58428), .Z(n58430) );
  NOR U69727 ( .A(n58430), .B(n58429), .Z(n58431) );
  NOR U69728 ( .A(n58432), .B(n58431), .Z(n58433) );
  IV U69729 ( .A(n58433), .Z(n58434) );
  NOR U69730 ( .A(n58435), .B(n58434), .Z(n58436) );
  XOR U69731 ( .A(n58437), .B(n58436), .Z(n58438) );
  XOR U69732 ( .A(n58439), .B(n58438), .Z(n58457) );
  NOR U69733 ( .A(n58441), .B(n58440), .Z(n58446) );
  IV U69734 ( .A(n58442), .Z(n58444) );
  NOR U69735 ( .A(n58444), .B(n58443), .Z(n58445) );
  NOR U69736 ( .A(n58446), .B(n58445), .Z(n58455) );
  NOR U69737 ( .A(n58448), .B(n58447), .Z(n58453) );
  IV U69738 ( .A(n58449), .Z(n58451) );
  NOR U69739 ( .A(n58451), .B(n58450), .Z(n58452) );
  NOR U69740 ( .A(n58453), .B(n58452), .Z(n58454) );
  XOR U69741 ( .A(n58455), .B(n58454), .Z(n58456) );
  XOR U69742 ( .A(n58457), .B(n58456), .Z(n58484) );
  IV U69743 ( .A(n58458), .Z(n58460) );
  NOR U69744 ( .A(n58460), .B(n58459), .Z(n58464) );
  IV U69745 ( .A(n58478), .Z(n58461) );
  NOR U69746 ( .A(n58462), .B(n58461), .Z(n58463) );
  NOR U69747 ( .A(n58464), .B(n58463), .Z(n58482) );
  IV U69748 ( .A(n58467), .Z(n58465) );
  NOR U69749 ( .A(n58465), .B(n58466), .Z(n58471) );
  XOR U69750 ( .A(n58467), .B(n58466), .Z(n58469) );
  NOR U69751 ( .A(n58469), .B(n58468), .Z(n58470) );
  NOR U69752 ( .A(n58471), .B(n58470), .Z(n58472) );
  IV U69753 ( .A(n58472), .Z(n58480) );
  IV U69754 ( .A(n58473), .Z(n58475) );
  NOR U69755 ( .A(n58475), .B(n58474), .Z(n58476) );
  IV U69756 ( .A(n58476), .Z(n58477) );
  NOR U69757 ( .A(n58478), .B(n58477), .Z(n58479) );
  NOR U69758 ( .A(n58480), .B(n58479), .Z(n58481) );
  XOR U69759 ( .A(n58482), .B(n58481), .Z(n58483) );
  XOR U69760 ( .A(n58484), .B(n58483), .Z(n58499) );
  IV U69761 ( .A(n58485), .Z(n58487) );
  NOR U69762 ( .A(n58487), .B(n58486), .Z(n58497) );
  NOR U69763 ( .A(n58489), .B(n58488), .Z(n58494) );
  IV U69764 ( .A(n58490), .Z(n58491) );
  NOR U69765 ( .A(n58492), .B(n58491), .Z(n58493) );
  NOR U69766 ( .A(n58494), .B(n58493), .Z(n58495) );
  IV U69767 ( .A(n58495), .Z(n58496) );
  NOR U69768 ( .A(n58497), .B(n58496), .Z(n58498) );
  XOR U69769 ( .A(n58499), .B(n58498), .Z(n58508) );
  NOR U69770 ( .A(n58500), .B(n58501), .Z(n58506) );
  XOR U69771 ( .A(n58502), .B(n58501), .Z(n58503) );
  NOR U69772 ( .A(n58504), .B(n58503), .Z(n58505) );
  NOR U69773 ( .A(n58506), .B(n58505), .Z(n58507) );
  XOR U69774 ( .A(n58508), .B(n58507), .Z(n58523) );
  IV U69775 ( .A(n58509), .Z(n58511) );
  NOR U69776 ( .A(n58511), .B(n58510), .Z(n58521) );
  XOR U69777 ( .A(n58512), .B(n58515), .Z(n58514) );
  NOR U69778 ( .A(n58514), .B(n58513), .Z(n58518) );
  NOR U69779 ( .A(n58516), .B(n58515), .Z(n58517) );
  NOR U69780 ( .A(n58518), .B(n58517), .Z(n58519) );
  IV U69781 ( .A(n58519), .Z(n58520) );
  NOR U69782 ( .A(n58521), .B(n58520), .Z(n58522) );
  XOR U69783 ( .A(n58523), .B(n58522), .Z(n58532) );
  NOR U69784 ( .A(n58526), .B(n58524), .Z(n58530) );
  XOR U69785 ( .A(n58526), .B(n58525), .Z(n58527) );
  NOR U69786 ( .A(n58528), .B(n58527), .Z(n58529) );
  NOR U69787 ( .A(n58530), .B(n58529), .Z(n58531) );
  XOR U69788 ( .A(n58532), .B(n58531), .Z(n58533) );
  XOR U69789 ( .A(n58534), .B(n58533), .Z(n58554) );
  IV U69790 ( .A(n58535), .Z(n58536) );
  NOR U69791 ( .A(n58537), .B(n58536), .Z(n58542) );
  IV U69792 ( .A(n58538), .Z(n58540) );
  NOR U69793 ( .A(n58540), .B(n58539), .Z(n58541) );
  NOR U69794 ( .A(n58542), .B(n58541), .Z(n58552) );
  IV U69795 ( .A(n58543), .Z(n58545) );
  NOR U69796 ( .A(n58545), .B(n58544), .Z(n58550) );
  IV U69797 ( .A(n58546), .Z(n58548) );
  NOR U69798 ( .A(n58548), .B(n58547), .Z(n58549) );
  NOR U69799 ( .A(n58550), .B(n58549), .Z(n58551) );
  XOR U69800 ( .A(n58552), .B(n58551), .Z(n58553) );
  XOR U69801 ( .A(n58554), .B(n58553), .Z(n58564) );
  IV U69802 ( .A(n58555), .Z(n58557) );
  NOR U69803 ( .A(n58556), .B(n58557), .Z(n58562) );
  XOR U69804 ( .A(n58558), .B(n58557), .Z(n58559) );
  NOR U69805 ( .A(n58560), .B(n58559), .Z(n58561) );
  NOR U69806 ( .A(n58562), .B(n58561), .Z(n58563) );
  XOR U69807 ( .A(n58564), .B(n58563), .Z(n58597) );
  IV U69808 ( .A(n58565), .Z(n58567) );
  NOR U69809 ( .A(n58567), .B(n58566), .Z(n58571) );
  NOR U69810 ( .A(n58569), .B(n58568), .Z(n58570) );
  NOR U69811 ( .A(n58571), .B(n58570), .Z(n58587) );
  IV U69812 ( .A(n58572), .Z(n58575) );
  IV U69813 ( .A(n58573), .Z(n58574) );
  NOR U69814 ( .A(n58575), .B(n58574), .Z(n58585) );
  NOR U69815 ( .A(n58577), .B(n58576), .Z(n58582) );
  IV U69816 ( .A(n58578), .Z(n58580) );
  NOR U69817 ( .A(n58580), .B(n58579), .Z(n58581) );
  NOR U69818 ( .A(n58582), .B(n58581), .Z(n58583) );
  IV U69819 ( .A(n58583), .Z(n58584) );
  NOR U69820 ( .A(n58585), .B(n58584), .Z(n58586) );
  XOR U69821 ( .A(n58587), .B(n58586), .Z(n58595) );
  IV U69822 ( .A(n58588), .Z(n58591) );
  IV U69823 ( .A(n58589), .Z(n58590) );
  NOR U69824 ( .A(n58591), .B(n58590), .Z(n58592) );
  NOR U69825 ( .A(n58593), .B(n58592), .Z(n58594) );
  XOR U69826 ( .A(n58595), .B(n58594), .Z(n58596) );
  XOR U69827 ( .A(n58597), .B(n58596), .Z(n58617) );
  IV U69828 ( .A(n58598), .Z(n58599) );
  NOR U69829 ( .A(n58600), .B(n58599), .Z(n58605) );
  IV U69830 ( .A(n58601), .Z(n58603) );
  NOR U69831 ( .A(n58603), .B(n58602), .Z(n58604) );
  NOR U69832 ( .A(n58605), .B(n58604), .Z(n58615) );
  IV U69833 ( .A(n58606), .Z(n58608) );
  NOR U69834 ( .A(n58608), .B(n58607), .Z(n58613) );
  IV U69835 ( .A(n58609), .Z(n58610) );
  NOR U69836 ( .A(n58611), .B(n58610), .Z(n58612) );
  NOR U69837 ( .A(n58613), .B(n58612), .Z(n58614) );
  XOR U69838 ( .A(n58615), .B(n58614), .Z(n58616) );
  XOR U69839 ( .A(n58617), .B(n58616), .Z(n58618) );
  XOR U69840 ( .A(n58619), .B(n58618), .Z(n58620) );
  XOR U69841 ( .A(n58621), .B(n58620), .Z(n58622) );
  IV U69842 ( .A(n58622), .Z(o[10]) );
  XOR U69843 ( .A(n58624), .B(n58623), .Z(o[1]) );
  NOR U69844 ( .A(n58626), .B(n58625), .Z(n58628) );
  XOR U69845 ( .A(n58628), .B(n58627), .Z(o[2]) );
  XOR U69846 ( .A(n58630), .B(n58629), .Z(o[3]) );
  NOR U69847 ( .A(n58632), .B(n58631), .Z(n58634) );
  XOR U69848 ( .A(n58634), .B(n58633), .Z(o[4]) );
  XOR U69849 ( .A(n58636), .B(n58635), .Z(o[5]) );
  XOR U69850 ( .A(n58638), .B(n58637), .Z(o[6]) );
  XOR U69851 ( .A(n58640), .B(n58639), .Z(o[7]) );
  NOR U69852 ( .A(n58642), .B(n58641), .Z(n58644) );
  XOR U69853 ( .A(n58644), .B(n58643), .Z(o[8]) );
  XOR U69854 ( .A(n58646), .B(n58645), .Z(o[9]) );
endmodule

