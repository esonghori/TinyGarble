
module mult_N128_CC4 ( clk, rst, a, b, c );
  input [127:0] a;
  input [31:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511;
  wire   [255:0] sreg;

  DFF \sreg_reg[223]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[222]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[221]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[220]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[219]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[218]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[217]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[216]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[215]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[214]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[213]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[212]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[211]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[210]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[209]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[208]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[207]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[206]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[205]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[204]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[203]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[202]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[201]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[200]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[199]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[198]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[197]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[196]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[195]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[194]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[193]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[192]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[191]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U35 ( .A(n4931), .B(n4932), .Z(n1) );
  NANDN U36 ( .A(n4930), .B(n4929), .Z(n2) );
  NAND U37 ( .A(n1), .B(n2), .Z(n5116) );
  NAND U38 ( .A(n7562), .B(n7563), .Z(n3) );
  NANDN U39 ( .A(n7565), .B(n7564), .Z(n4) );
  AND U40 ( .A(n3), .B(n4), .Z(n7725) );
  NAND U41 ( .A(n9881), .B(n9882), .Z(n5) );
  NANDN U42 ( .A(n9884), .B(n9883), .Z(n6) );
  AND U43 ( .A(n5), .B(n6), .Z(n10042) );
  XNOR U44 ( .A(n19061), .B(n19062), .Z(n19064) );
  XNOR U45 ( .A(n19067), .B(n19068), .Z(n19070) );
  NAND U46 ( .A(n19167), .B(n19166), .Z(n7) );
  NAND U47 ( .A(n19164), .B(n19165), .Z(n8) );
  NAND U48 ( .A(n7), .B(n8), .Z(n19254) );
  XNOR U49 ( .A(n4233), .B(n4232), .Z(n4234) );
  XNOR U50 ( .A(n5682), .B(n5681), .Z(n5683) );
  XNOR U51 ( .A(n6562), .B(n6561), .Z(n6563) );
  XNOR U52 ( .A(n6992), .B(n6991), .Z(n6993) );
  XNOR U53 ( .A(n7567), .B(n7566), .Z(n7568) );
  XNOR U54 ( .A(n7990), .B(n7989), .Z(n7991) );
  XNOR U55 ( .A(n8439), .B(n8438), .Z(n8440) );
  XNOR U56 ( .A(n9612), .B(n9611), .Z(n9613) );
  XNOR U57 ( .A(n9886), .B(n9885), .Z(n9887) );
  XNOR U58 ( .A(n11212), .B(n11211), .Z(n11213) );
  XNOR U59 ( .A(n11921), .B(n11920), .Z(n11922) );
  XNOR U60 ( .A(n12792), .B(n12791), .Z(n12793) );
  XNOR U61 ( .A(n13078), .B(n13077), .Z(n13079) );
  XNOR U62 ( .A(n13372), .B(n13371), .Z(n13373) );
  XNOR U63 ( .A(n13940), .B(n13939), .Z(n13941) );
  NAND U64 ( .A(n2187), .B(n2186), .Z(n9) );
  NANDN U65 ( .A(n2185), .B(n2184), .Z(n10) );
  NAND U66 ( .A(n9), .B(n10), .Z(n2229) );
  NAND U67 ( .A(n3185), .B(n3186), .Z(n11) );
  NANDN U68 ( .A(n3188), .B(n3187), .Z(n12) );
  AND U69 ( .A(n11), .B(n12), .Z(n3412) );
  NAND U70 ( .A(n4228), .B(n4229), .Z(n13) );
  NANDN U71 ( .A(n4231), .B(n4230), .Z(n14) );
  AND U72 ( .A(n13), .B(n14), .Z(n4385) );
  NAND U73 ( .A(n4928), .B(n4927), .Z(n15) );
  NANDN U74 ( .A(n4926), .B(n4925), .Z(n16) );
  NAND U75 ( .A(n15), .B(n16), .Z(n5117) );
  NAND U76 ( .A(n5398), .B(n5397), .Z(n17) );
  NANDN U77 ( .A(n5396), .B(n5395), .Z(n18) );
  AND U78 ( .A(n17), .B(n18), .Z(n5548) );
  NAND U79 ( .A(n5677), .B(n5678), .Z(n19) );
  NANDN U80 ( .A(n5680), .B(n5679), .Z(n20) );
  AND U81 ( .A(n19), .B(n20), .Z(n5842) );
  NAND U82 ( .A(n6557), .B(n6558), .Z(n21) );
  NANDN U83 ( .A(n6560), .B(n6559), .Z(n22) );
  AND U84 ( .A(n21), .B(n22), .Z(n6722) );
  NAND U85 ( .A(n6712), .B(n6713), .Z(n23) );
  NANDN U86 ( .A(n6715), .B(n6714), .Z(n24) );
  AND U87 ( .A(n23), .B(n24), .Z(n6866) );
  NAND U88 ( .A(n6987), .B(n6988), .Z(n25) );
  NANDN U89 ( .A(n6990), .B(n6989), .Z(n26) );
  AND U90 ( .A(n25), .B(n26), .Z(n7152) );
  NAND U91 ( .A(n7142), .B(n7143), .Z(n27) );
  NANDN U92 ( .A(n7145), .B(n7144), .Z(n28) );
  AND U93 ( .A(n27), .B(n28), .Z(n7295) );
  NAND U94 ( .A(n7438), .B(n7437), .Z(n29) );
  NANDN U95 ( .A(n7436), .B(n7435), .Z(n30) );
  AND U96 ( .A(n29), .B(n30), .Z(n7572) );
  NAND U97 ( .A(n7738), .B(n7737), .Z(n31) );
  NANDN U98 ( .A(n7736), .B(n7735), .Z(n32) );
  NAND U99 ( .A(n31), .B(n32), .Z(n7913) );
  NAND U100 ( .A(n7724), .B(n7723), .Z(n33) );
  NANDN U101 ( .A(n7722), .B(n7721), .Z(n34) );
  AND U102 ( .A(n33), .B(n34), .Z(n7856) );
  NAND U103 ( .A(n7985), .B(n7986), .Z(n35) );
  NANDN U104 ( .A(n7988), .B(n7987), .Z(n36) );
  AND U105 ( .A(n35), .B(n36), .Z(n8150) );
  NAND U106 ( .A(n8434), .B(n8435), .Z(n37) );
  NANDN U107 ( .A(n8437), .B(n8436), .Z(n38) );
  AND U108 ( .A(n37), .B(n38), .Z(n8590) );
  NAND U109 ( .A(n9167), .B(n9166), .Z(n39) );
  NANDN U110 ( .A(n9165), .B(n9164), .Z(n40) );
  AND U111 ( .A(n39), .B(n40), .Z(n9317) );
  NAND U112 ( .A(n9607), .B(n9608), .Z(n41) );
  NANDN U113 ( .A(n9610), .B(n9609), .Z(n42) );
  AND U114 ( .A(n41), .B(n42), .Z(n9760) );
  NAND U115 ( .A(n9759), .B(n9758), .Z(n43) );
  NANDN U116 ( .A(n9757), .B(n9756), .Z(n44) );
  AND U117 ( .A(n43), .B(n44), .Z(n9891) );
  NAND U118 ( .A(n10055), .B(n10054), .Z(n45) );
  NANDN U119 ( .A(n10053), .B(n10052), .Z(n46) );
  NAND U120 ( .A(n45), .B(n46), .Z(n10233) );
  NAND U121 ( .A(n11207), .B(n11208), .Z(n47) );
  NANDN U122 ( .A(n11210), .B(n11209), .Z(n48) );
  AND U123 ( .A(n47), .B(n48), .Z(n11362) );
  NAND U124 ( .A(n11492), .B(n11491), .Z(n49) );
  NANDN U125 ( .A(n11490), .B(n11489), .Z(n50) );
  AND U126 ( .A(n49), .B(n50), .Z(n11640) );
  NAND U127 ( .A(n11916), .B(n11917), .Z(n51) );
  NANDN U128 ( .A(n11919), .B(n11918), .Z(n52) );
  AND U129 ( .A(n51), .B(n52), .Z(n12086) );
  NAND U130 ( .A(n12365), .B(n12364), .Z(n53) );
  NANDN U131 ( .A(n12363), .B(n12362), .Z(n54) );
  AND U132 ( .A(n53), .B(n54), .Z(n12465) );
  XNOR U133 ( .A(n12797), .B(n12798), .Z(n12800) );
  NAND U134 ( .A(n12787), .B(n12788), .Z(n55) );
  NANDN U135 ( .A(n12790), .B(n12789), .Z(n56) );
  AND U136 ( .A(n55), .B(n56), .Z(n12952) );
  NAND U137 ( .A(n12951), .B(n12950), .Z(n57) );
  NANDN U138 ( .A(n12949), .B(n12948), .Z(n58) );
  AND U139 ( .A(n57), .B(n58), .Z(n13083) );
  NAND U140 ( .A(n13073), .B(n13074), .Z(n59) );
  NANDN U141 ( .A(n13076), .B(n13075), .Z(n60) );
  AND U142 ( .A(n59), .B(n60), .Z(n13236) );
  NAND U143 ( .A(n13367), .B(n13368), .Z(n61) );
  NANDN U144 ( .A(n13370), .B(n13369), .Z(n62) );
  AND U145 ( .A(n61), .B(n62), .Z(n13522) );
  NAND U146 ( .A(n13799), .B(n13798), .Z(n63) );
  NANDN U147 ( .A(n13797), .B(n13796), .Z(n64) );
  AND U148 ( .A(n63), .B(n64), .Z(n13945) );
  NAND U149 ( .A(n13935), .B(n13936), .Z(n65) );
  NANDN U150 ( .A(n13938), .B(n13937), .Z(n66) );
  AND U151 ( .A(n65), .B(n66), .Z(n14094) );
  NAND U152 ( .A(n14084), .B(n14085), .Z(n67) );
  NANDN U153 ( .A(n14087), .B(n14086), .Z(n68) );
  AND U154 ( .A(n67), .B(n68), .Z(n14233) );
  NAND U155 ( .A(n14232), .B(n14231), .Z(n69) );
  NANDN U156 ( .A(n14230), .B(n14229), .Z(n70) );
  AND U157 ( .A(n69), .B(n70), .Z(n14318) );
  NAND U158 ( .A(n14419), .B(n14418), .Z(n71) );
  NANDN U159 ( .A(n14417), .B(n14416), .Z(n72) );
  AND U160 ( .A(n71), .B(n72), .Z(n14507) );
  XNOR U161 ( .A(n15086), .B(n15087), .Z(n15089) );
  XNOR U162 ( .A(n16277), .B(n16276), .Z(n16278) );
  XNOR U163 ( .A(n16527), .B(n16526), .Z(n16528) );
  OR U164 ( .A(b[1]), .B(n17139), .Z(n73) );
  NAND U165 ( .A(n17140), .B(n17141), .Z(n74) );
  NAND U166 ( .A(n73), .B(n74), .Z(n17293) );
  NAND U167 ( .A(n7728), .B(n7727), .Z(n75) );
  NANDN U168 ( .A(n7726), .B(n7725), .Z(n76) );
  NAND U169 ( .A(n75), .B(n76), .Z(n7931) );
  NAND U170 ( .A(n10045), .B(n10044), .Z(n77) );
  NANDN U171 ( .A(n10043), .B(n10042), .Z(n78) );
  NAND U172 ( .A(n77), .B(n78), .Z(n10251) );
  NAND U173 ( .A(n16272), .B(n16273), .Z(n79) );
  NANDN U174 ( .A(n16275), .B(n16274), .Z(n80) );
  AND U175 ( .A(n79), .B(n80), .Z(n16427) );
  XOR U176 ( .A(n16768), .B(n16769), .Z(n16770) );
  NAND U177 ( .A(n1137), .B(n1136), .Z(n81) );
  NANDN U178 ( .A(n1135), .B(n1134), .Z(n82) );
  NAND U179 ( .A(n81), .B(n82), .Z(n1173) );
  NAND U180 ( .A(n1407), .B(n1406), .Z(n83) );
  NANDN U181 ( .A(n1405), .B(n1404), .Z(n84) );
  NAND U182 ( .A(n83), .B(n84), .Z(n1559) );
  NAND U183 ( .A(n1595), .B(n1594), .Z(n85) );
  NANDN U184 ( .A(n1597), .B(n1596), .Z(n86) );
  NAND U185 ( .A(n85), .B(n86), .Z(n1664) );
  XNOR U186 ( .A(n19064), .B(n19063), .Z(n19069) );
  NAND U187 ( .A(n16959), .B(n16960), .Z(n87) );
  NANDN U188 ( .A(n16958), .B(n16957), .Z(n88) );
  NAND U189 ( .A(n87), .B(n88), .Z(n17098) );
  XOR U190 ( .A(n18425), .B(n18426), .Z(n89) );
  NANDN U191 ( .A(n18427), .B(n89), .Z(n90) );
  NAND U192 ( .A(n18425), .B(n18426), .Z(n91) );
  AND U193 ( .A(n90), .B(n91), .Z(n18457) );
  NAND U194 ( .A(n18532), .B(n18531), .Z(n92) );
  NANDN U195 ( .A(n18530), .B(n18529), .Z(n93) );
  AND U196 ( .A(n92), .B(n93), .Z(n18626) );
  NAND U197 ( .A(n18785), .B(n18784), .Z(n94) );
  NANDN U198 ( .A(n18783), .B(n18782), .Z(n95) );
  NAND U199 ( .A(n94), .B(n95), .Z(n18814) );
  NAND U200 ( .A(n19335), .B(n19334), .Z(n96) );
  NANDN U201 ( .A(n19333), .B(n19382), .Z(n97) );
  NAND U202 ( .A(n96), .B(n97), .Z(n19366) );
  NANDN U203 ( .A(a[0]), .B(n16990), .Z(n98) );
  NANDN U204 ( .A(b[2]), .B(n17151), .Z(n99) );
  NAND U205 ( .A(n99), .B(n98), .Z(n100) );
  NANDN U206 ( .A(n578), .B(n100), .Z(n631) );
  NAND U207 ( .A(n19163), .B(n19162), .Z(n101) );
  NANDN U208 ( .A(n19161), .B(n19160), .Z(n102) );
  NAND U209 ( .A(n101), .B(n102), .Z(n19257) );
  XOR U210 ( .A(n19204), .B(n19205), .Z(n103) );
  NANDN U211 ( .A(n19206), .B(n103), .Z(n104) );
  NAND U212 ( .A(n19204), .B(n19205), .Z(n105) );
  AND U213 ( .A(n104), .B(n105), .Z(n19262) );
  NAND U214 ( .A(n19460), .B(n19459), .Z(n106) );
  XOR U215 ( .A(n19459), .B(n19460), .Z(n107) );
  NAND U216 ( .A(n107), .B(n19458), .Z(n108) );
  NAND U217 ( .A(n106), .B(n108), .Z(n19492) );
  ANDN U218 ( .B(n19483), .A(n2539), .Z(n2623) );
  NAND U219 ( .A(n2804), .B(n2805), .Z(n109) );
  NANDN U220 ( .A(n2803), .B(n2802), .Z(n110) );
  AND U221 ( .A(n109), .B(n110), .Z(n2900) );
  XNOR U222 ( .A(n3789), .B(n3790), .Z(n3792) );
  XNOR U223 ( .A(n3904), .B(n3905), .Z(n3907) );
  XNOR U224 ( .A(n3898), .B(n3899), .Z(n3901) );
  XNOR U225 ( .A(n4051), .B(n4052), .Z(n4054) );
  XNOR U226 ( .A(n4045), .B(n4046), .Z(n4048) );
  XNOR U227 ( .A(n4518), .B(n4519), .Z(n4521) );
  XOR U228 ( .A(n4636), .B(n4637), .Z(n4638) );
  XOR U229 ( .A(n4630), .B(n4631), .Z(n4632) );
  XNOR U230 ( .A(n4797), .B(n4798), .Z(n4800) );
  XNOR U231 ( .A(n4791), .B(n4792), .Z(n4794) );
  XNOR U232 ( .A(n5234), .B(n5235), .Z(n5237) );
  XNOR U233 ( .A(n5228), .B(n5229), .Z(n5231) );
  XNOR U234 ( .A(n5378), .B(n5377), .Z(n5379) );
  XNOR U235 ( .A(n5536), .B(n5537), .Z(n5539) );
  XNOR U236 ( .A(n5830), .B(n5831), .Z(n5833) );
  XNOR U237 ( .A(n6124), .B(n6125), .Z(n6127) );
  XNOR U238 ( .A(n6408), .B(n6409), .Z(n6411) );
  XNOR U239 ( .A(n6717), .B(n6716), .Z(n6718) );
  XNOR U240 ( .A(n6854), .B(n6855), .Z(n6857) );
  XNOR U241 ( .A(n7147), .B(n7146), .Z(n7148) );
  XNOR U242 ( .A(n7283), .B(n7284), .Z(n7286) );
  XNOR U243 ( .A(n7844), .B(n7845), .Z(n7847) );
  XNOR U244 ( .A(n8273), .B(n8274), .Z(n8276) );
  XNOR U245 ( .A(n8872), .B(n8873), .Z(n8875) );
  XNOR U246 ( .A(n9002), .B(n9003), .Z(n9005) );
  XNOR U247 ( .A(n8996), .B(n8997), .Z(n8999) );
  XNOR U248 ( .A(n9460), .B(n9461), .Z(n9463) );
  XNOR U249 ( .A(n10305), .B(n10306), .Z(n10308) );
  XNOR U250 ( .A(n10603), .B(n10604), .Z(n10606) );
  XOR U251 ( .A(n10735), .B(n10736), .Z(n10737) );
  XOR U252 ( .A(n10729), .B(n10730), .Z(n10731) );
  XNOR U253 ( .A(n10884), .B(n10885), .Z(n10887) );
  XNOR U254 ( .A(n10878), .B(n10879), .Z(n10881) );
  XNOR U255 ( .A(n11350), .B(n11351), .Z(n11353) );
  XNOR U256 ( .A(n11472), .B(n11471), .Z(n11473) );
  XNOR U257 ( .A(n11628), .B(n11629), .Z(n11631) );
  XNOR U258 ( .A(n11761), .B(n11762), .Z(n11764) );
  XNOR U259 ( .A(n11755), .B(n11756), .Z(n11758) );
  XOR U260 ( .A(n12189), .B(n12190), .Z(n12191) );
  XNOR U261 ( .A(n12184), .B(n12183), .Z(n12185) );
  XNOR U262 ( .A(n12345), .B(n12344), .Z(n12346) );
  XOR U263 ( .A(n12622), .B(n12623), .Z(n12624) );
  XNOR U264 ( .A(n12617), .B(n12616), .Z(n12618) );
  XNOR U265 ( .A(n13224), .B(n13225), .Z(n13227) );
  XNOR U266 ( .A(n13643), .B(n13644), .Z(n13646) );
  XNOR U267 ( .A(n13779), .B(n13778), .Z(n13780) );
  XNOR U268 ( .A(n14089), .B(n14088), .Z(n14090) );
  XNOR U269 ( .A(n14399), .B(n14398), .Z(n14400) );
  XNOR U270 ( .A(n14649), .B(n14650), .Z(n14652) );
  XNOR U271 ( .A(n15369), .B(n15370), .Z(n15372) );
  XNOR U272 ( .A(n15827), .B(n15828), .Z(n15830) );
  XNOR U273 ( .A(n16111), .B(n16112), .Z(n16114) );
  NAND U274 ( .A(n2303), .B(n2304), .Z(n111) );
  NANDN U275 ( .A(n2302), .B(n2301), .Z(n112) );
  AND U276 ( .A(n111), .B(n112), .Z(n2378) );
  XOR U277 ( .A(n3213), .B(n3214), .Z(n3215) );
  XNOR U278 ( .A(n3493), .B(n3494), .Z(n3496) );
  XOR U279 ( .A(n3642), .B(n3643), .Z(n3644) );
  XOR U280 ( .A(n3801), .B(n3802), .Z(n3803) );
  XOR U281 ( .A(n4530), .B(n4531), .Z(n4532) );
  NAND U282 ( .A(n4398), .B(n4397), .Z(n113) );
  NANDN U283 ( .A(n4396), .B(n4395), .Z(n114) );
  NAND U284 ( .A(n113), .B(n114), .Z(n4595) );
  XNOR U285 ( .A(n4827), .B(n4828), .Z(n4830) );
  NANDN U286 ( .A(n4922), .B(n4921), .Z(n115) );
  NANDN U287 ( .A(n4924), .B(n4923), .Z(n116) );
  NAND U288 ( .A(n115), .B(n116), .Z(n5118) );
  NAND U289 ( .A(n5561), .B(n5560), .Z(n117) );
  NANDN U290 ( .A(n5559), .B(n5558), .Z(n118) );
  NAND U291 ( .A(n117), .B(n118), .Z(n5752) );
  NAND U292 ( .A(n5855), .B(n5854), .Z(n119) );
  NANDN U293 ( .A(n5853), .B(n5852), .Z(n120) );
  NAND U294 ( .A(n119), .B(n120), .Z(n6054) );
  XNOR U295 ( .A(n6136), .B(n6137), .Z(n6139) );
  XNOR U296 ( .A(n6420), .B(n6421), .Z(n6423) );
  NAND U297 ( .A(n6735), .B(n6734), .Z(n121) );
  NANDN U298 ( .A(n6733), .B(n6732), .Z(n122) );
  NAND U299 ( .A(n121), .B(n122), .Z(n6807) );
  NAND U300 ( .A(n6879), .B(n6878), .Z(n123) );
  NANDN U301 ( .A(n6877), .B(n6876), .Z(n124) );
  NAND U302 ( .A(n123), .B(n124), .Z(n7062) );
  NAND U303 ( .A(n7165), .B(n7164), .Z(n125) );
  NANDN U304 ( .A(n7163), .B(n7162), .Z(n126) );
  NAND U305 ( .A(n125), .B(n126), .Z(n7237) );
  NAND U306 ( .A(n7308), .B(n7307), .Z(n127) );
  NANDN U307 ( .A(n7306), .B(n7305), .Z(n128) );
  NAND U308 ( .A(n127), .B(n128), .Z(n7504) );
  NAND U309 ( .A(n7869), .B(n7868), .Z(n129) );
  NANDN U310 ( .A(n7867), .B(n7866), .Z(n130) );
  NAND U311 ( .A(n129), .B(n130), .Z(n8059) );
  XNOR U312 ( .A(n8285), .B(n8286), .Z(n8288) );
  XOR U313 ( .A(n8735), .B(n8736), .Z(n8737) );
  NAND U314 ( .A(n8603), .B(n8602), .Z(n131) );
  NANDN U315 ( .A(n8601), .B(n8600), .Z(n132) );
  NAND U316 ( .A(n131), .B(n132), .Z(n8801) );
  XOR U317 ( .A(n8884), .B(n8885), .Z(n8886) );
  XOR U318 ( .A(n9472), .B(n9473), .Z(n9474) );
  NAND U319 ( .A(n9773), .B(n9772), .Z(n133) );
  NANDN U320 ( .A(n9771), .B(n9770), .Z(n134) );
  NAND U321 ( .A(n133), .B(n134), .Z(n9948) );
  NAND U322 ( .A(n10041), .B(n10040), .Z(n135) );
  NANDN U323 ( .A(n10039), .B(n10038), .Z(n136) );
  AND U324 ( .A(n135), .B(n136), .Z(n10174) );
  XNOR U325 ( .A(n10317), .B(n10318), .Z(n10320) );
  XNOR U326 ( .A(n10615), .B(n10616), .Z(n10618) );
  XNOR U327 ( .A(n10914), .B(n10915), .Z(n10917) );
  XNOR U328 ( .A(n11217), .B(n11218), .Z(n11220) );
  NAND U329 ( .A(n11653), .B(n11652), .Z(n137) );
  NANDN U330 ( .A(n11651), .B(n11650), .Z(n138) );
  NAND U331 ( .A(n137), .B(n138), .Z(n11858) );
  NAND U332 ( .A(n12099), .B(n12098), .Z(n139) );
  NANDN U333 ( .A(n12097), .B(n12096), .Z(n140) );
  NAND U334 ( .A(n139), .B(n140), .Z(n12178) );
  XNOR U335 ( .A(n12366), .B(n12367), .Z(n12369) );
  NAND U336 ( .A(n12478), .B(n12477), .Z(n141) );
  NANDN U337 ( .A(n12476), .B(n12475), .Z(n142) );
  NAND U338 ( .A(n141), .B(n142), .Z(n12611) );
  NAND U339 ( .A(n12965), .B(n12964), .Z(n143) );
  NANDN U340 ( .A(n12963), .B(n12962), .Z(n144) );
  NAND U341 ( .A(n143), .B(n144), .Z(n13140) );
  NAND U342 ( .A(n13096), .B(n13095), .Z(n145) );
  NANDN U343 ( .A(n13094), .B(n13093), .Z(n146) );
  NAND U344 ( .A(n145), .B(n146), .Z(n13178) );
  XOR U345 ( .A(n13655), .B(n13656), .Z(n13657) );
  NAND U346 ( .A(n13535), .B(n13534), .Z(n147) );
  NANDN U347 ( .A(n13533), .B(n13532), .Z(n148) );
  NAND U348 ( .A(n147), .B(n148), .Z(n13719) );
  NAND U349 ( .A(n13958), .B(n13957), .Z(n149) );
  NANDN U350 ( .A(n13956), .B(n13955), .Z(n150) );
  NAND U351 ( .A(n149), .B(n150), .Z(n14039) );
  NAND U352 ( .A(n14246), .B(n14245), .Z(n151) );
  NANDN U353 ( .A(n14244), .B(n14243), .Z(n152) );
  NAND U354 ( .A(n151), .B(n152), .Z(n14421) );
  XOR U355 ( .A(n14655), .B(n14656), .Z(n14657) );
  NAND U356 ( .A(n14520), .B(n14519), .Z(n153) );
  NANDN U357 ( .A(n14518), .B(n14517), .Z(n154) );
  NAND U358 ( .A(n153), .B(n154), .Z(n14720) );
  NAND U359 ( .A(n14645), .B(n14646), .Z(n155) );
  NANDN U360 ( .A(n14648), .B(n14647), .Z(n156) );
  AND U361 ( .A(n155), .B(n156), .Z(n14802) );
  XOR U362 ( .A(n15246), .B(n15247), .Z(n15248) );
  XOR U363 ( .A(n15381), .B(n15382), .Z(n15383) );
  XNOR U364 ( .A(n15690), .B(n15691), .Z(n15693) );
  XOR U365 ( .A(n15839), .B(n15840), .Z(n15841) );
  XNOR U366 ( .A(n16123), .B(n16124), .Z(n16126) );
  NOR U367 ( .A(b[17]), .B(b[18]), .Z(n157) );
  NAND U368 ( .A(n18834), .B(n2921), .Z(n158) );
  NANDN U369 ( .A(n157), .B(n158), .Z(n159) );
  ANDN U370 ( .B(n159), .A(n581), .Z(n1532) );
  NAND U371 ( .A(n1645), .B(n1646), .Z(n160) );
  NANDN U372 ( .A(n1644), .B(n1643), .Z(n161) );
  AND U373 ( .A(n160), .B(n161), .Z(n1739) );
  NAND U374 ( .A(n1540), .B(n1539), .Z(n162) );
  NANDN U375 ( .A(n1538), .B(n1537), .Z(n163) );
  NAND U376 ( .A(n162), .B(n163), .Z(n1601) );
  NAND U377 ( .A(n2021), .B(n2020), .Z(n164) );
  NANDN U378 ( .A(n2019), .B(n2018), .Z(n165) );
  NAND U379 ( .A(n164), .B(n165), .Z(n2113) );
  NAND U380 ( .A(n3415), .B(n3414), .Z(n166) );
  NANDN U381 ( .A(n3413), .B(n3412), .Z(n167) );
  AND U382 ( .A(n166), .B(n167), .Z(n3571) );
  OR U383 ( .A(n3867), .B(n3868), .Z(n168) );
  NAND U384 ( .A(n3866), .B(n3865), .Z(n169) );
  NAND U385 ( .A(n168), .B(n169), .Z(n4007) );
  XNOR U386 ( .A(n4449), .B(n4450), .Z(n4444) );
  NAND U387 ( .A(n4388), .B(n4387), .Z(n170) );
  NANDN U388 ( .A(n4386), .B(n4385), .Z(n171) );
  NAND U389 ( .A(n170), .B(n171), .Z(n4477) );
  OR U390 ( .A(n5550), .B(n5551), .Z(n172) );
  NAND U391 ( .A(n5549), .B(n5548), .Z(n173) );
  NAND U392 ( .A(n172), .B(n173), .Z(n5757) );
  XNOR U393 ( .A(n5906), .B(n5907), .Z(n5901) );
  NAND U394 ( .A(n5845), .B(n5844), .Z(n174) );
  NANDN U395 ( .A(n5843), .B(n5842), .Z(n175) );
  NAND U396 ( .A(n174), .B(n175), .Z(n5934) );
  XNOR U397 ( .A(n6786), .B(n6787), .Z(n6781) );
  NAND U398 ( .A(n6725), .B(n6724), .Z(n176) );
  NANDN U399 ( .A(n6723), .B(n6722), .Z(n177) );
  NAND U400 ( .A(n176), .B(n177), .Z(n6929) );
  NAND U401 ( .A(n6869), .B(n6868), .Z(n178) );
  NANDN U402 ( .A(n6867), .B(n6866), .Z(n179) );
  NAND U403 ( .A(n178), .B(n179), .Z(n7074) );
  XNOR U404 ( .A(n7216), .B(n7217), .Z(n7211) );
  NAND U405 ( .A(n7155), .B(n7154), .Z(n180) );
  NANDN U406 ( .A(n7153), .B(n7152), .Z(n181) );
  NAND U407 ( .A(n180), .B(n181), .Z(n7359) );
  NAND U408 ( .A(n7298), .B(n7297), .Z(n182) );
  NANDN U409 ( .A(n7296), .B(n7295), .Z(n183) );
  NAND U410 ( .A(n182), .B(n183), .Z(n7388) );
  OR U411 ( .A(n7858), .B(n7859), .Z(n184) );
  NAND U412 ( .A(n7857), .B(n7856), .Z(n185) );
  NAND U413 ( .A(n184), .B(n185), .Z(n8065) );
  XNOR U414 ( .A(n8216), .B(n8217), .Z(n8211) );
  NAND U415 ( .A(n8153), .B(n8152), .Z(n186) );
  NANDN U416 ( .A(n8151), .B(n8150), .Z(n187) );
  NAND U417 ( .A(n186), .B(n187), .Z(n8364) );
  XNOR U418 ( .A(n8654), .B(n8655), .Z(n8649) );
  NAND U419 ( .A(n8593), .B(n8592), .Z(n188) );
  NANDN U420 ( .A(n8591), .B(n8590), .Z(n189) );
  NAND U421 ( .A(n188), .B(n189), .Z(n8682) );
  OR U422 ( .A(n9319), .B(n9320), .Z(n190) );
  NAND U423 ( .A(n9318), .B(n9317), .Z(n191) );
  NAND U424 ( .A(n190), .B(n191), .Z(n9414) );
  XNOR U425 ( .A(n9824), .B(n9825), .Z(n9819) );
  NAND U426 ( .A(n9763), .B(n9762), .Z(n192) );
  NANDN U427 ( .A(n9761), .B(n9760), .Z(n193) );
  NAND U428 ( .A(n192), .B(n193), .Z(n9966) );
  NAND U429 ( .A(n11311), .B(n11310), .Z(n194) );
  NANDN U430 ( .A(n11313), .B(n11312), .Z(n195) );
  NAND U431 ( .A(n194), .B(n195), .Z(n11564) );
  OR U432 ( .A(n11642), .B(n11643), .Z(n196) );
  NAND U433 ( .A(n11641), .B(n11640), .Z(n197) );
  NAND U434 ( .A(n196), .B(n197), .Z(n11733) );
  XNOR U435 ( .A(n12150), .B(n12151), .Z(n12145) );
  NAND U436 ( .A(n12089), .B(n12088), .Z(n198) );
  NANDN U437 ( .A(n12087), .B(n12086), .Z(n199) );
  NAND U438 ( .A(n198), .B(n199), .Z(n12298) );
  OR U439 ( .A(n12467), .B(n12468), .Z(n200) );
  NAND U440 ( .A(n12466), .B(n12465), .Z(n201) );
  NAND U441 ( .A(n200), .B(n201), .Z(n12724) );
  NANDN U442 ( .A(n12609), .B(n12608), .Z(n202) );
  NANDN U443 ( .A(n12607), .B(n12606), .Z(n203) );
  NAND U444 ( .A(n202), .B(n203), .Z(n12873) );
  XNOR U445 ( .A(n13016), .B(n13017), .Z(n13011) );
  NAND U446 ( .A(n12955), .B(n12954), .Z(n204) );
  NANDN U447 ( .A(n12953), .B(n12952), .Z(n205) );
  NAND U448 ( .A(n204), .B(n205), .Z(n13158) );
  OR U449 ( .A(n13085), .B(n13086), .Z(n206) );
  NAND U450 ( .A(n13084), .B(n13083), .Z(n207) );
  NAND U451 ( .A(n206), .B(n207), .Z(n13292) );
  NAND U452 ( .A(n13187), .B(n13186), .Z(n208) );
  NAND U453 ( .A(n13184), .B(n13185), .Z(n209) );
  NAND U454 ( .A(n208), .B(n209), .Z(n13320) );
  XNOR U455 ( .A(n13586), .B(n13587), .Z(n13581) );
  NAND U456 ( .A(n13525), .B(n13524), .Z(n210) );
  NANDN U457 ( .A(n13523), .B(n13522), .Z(n211) );
  NAND U458 ( .A(n210), .B(n211), .Z(n13732) );
  OR U459 ( .A(n13947), .B(n13948), .Z(n212) );
  NAND U460 ( .A(n13946), .B(n13945), .Z(n213) );
  NAND U461 ( .A(n212), .B(n213), .Z(n14150) );
  NAND U462 ( .A(n14047), .B(n14046), .Z(n214) );
  NAND U463 ( .A(n14044), .B(n14045), .Z(n215) );
  NAND U464 ( .A(n214), .B(n215), .Z(n14290) );
  NAND U465 ( .A(n14236), .B(n14235), .Z(n216) );
  NANDN U466 ( .A(n14234), .B(n14233), .Z(n217) );
  NAND U467 ( .A(n216), .B(n217), .Z(n14439) );
  OR U468 ( .A(n14509), .B(n14510), .Z(n218) );
  NAND U469 ( .A(n14508), .B(n14507), .Z(n219) );
  NAND U470 ( .A(n218), .B(n219), .Z(n14599) );
  NAND U471 ( .A(n15150), .B(n15149), .Z(n220) );
  NANDN U472 ( .A(n15148), .B(n15147), .Z(n221) );
  NAND U473 ( .A(n220), .B(n221), .Z(n15187) );
  XNOR U474 ( .A(n16493), .B(n16494), .Z(n16488) );
  NAND U475 ( .A(n16589), .B(n16588), .Z(n222) );
  NANDN U476 ( .A(n16587), .B(n16586), .Z(n223) );
  NAND U477 ( .A(n222), .B(n223), .Z(n16781) );
  NAND U478 ( .A(n17291), .B(n17290), .Z(n224) );
  NANDN U479 ( .A(n17293), .B(n17292), .Z(n225) );
  NAND U480 ( .A(n224), .B(n225), .Z(n17391) );
  NANDN U481 ( .A(n1258), .B(n1257), .Z(n226) );
  NANDN U482 ( .A(n1260), .B(n1259), .Z(n227) );
  NAND U483 ( .A(n226), .B(n227), .Z(n1328) );
  NAND U484 ( .A(n1587), .B(n1586), .Z(n228) );
  NANDN U485 ( .A(n1585), .B(n1584), .Z(n229) );
  NAND U486 ( .A(n228), .B(n229), .Z(n1666) );
  XOR U487 ( .A(n3166), .B(n3165), .Z(n230) );
  NANDN U488 ( .A(n3164), .B(n230), .Z(n231) );
  NAND U489 ( .A(n3166), .B(n3165), .Z(n232) );
  AND U490 ( .A(n231), .B(n232), .Z(n3295) );
  NANDN U491 ( .A(n7782), .B(n7781), .Z(n233) );
  NANDN U492 ( .A(n7784), .B(n7783), .Z(n234) );
  NAND U493 ( .A(n233), .B(n234), .Z(n7802) );
  NANDN U494 ( .A(n7933), .B(n7932), .Z(n235) );
  NANDN U495 ( .A(n7931), .B(n7930), .Z(n236) );
  AND U496 ( .A(n235), .B(n236), .Z(n7943) );
  NANDN U497 ( .A(n10100), .B(n10099), .Z(n237) );
  NANDN U498 ( .A(n10102), .B(n10101), .Z(n238) );
  NAND U499 ( .A(n237), .B(n238), .Z(n10120) );
  NANDN U500 ( .A(n10253), .B(n10252), .Z(n239) );
  NANDN U501 ( .A(n10251), .B(n10250), .Z(n240) );
  AND U502 ( .A(n239), .B(n240), .Z(n10263) );
  NAND U503 ( .A(n14576), .B(n14577), .Z(n241) );
  NANDN U504 ( .A(n14575), .B(n14574), .Z(n242) );
  NAND U505 ( .A(n241), .B(n242), .Z(n14593) );
  NAND U506 ( .A(n16430), .B(n16429), .Z(n243) );
  NANDN U507 ( .A(n16428), .B(n16427), .Z(n244) );
  NAND U508 ( .A(n243), .B(n244), .Z(n16640) );
  NAND U509 ( .A(n16789), .B(n16788), .Z(n245) );
  NANDN U510 ( .A(n16787), .B(n16786), .Z(n246) );
  NAND U511 ( .A(n245), .B(n246), .Z(n16802) );
  XOR U512 ( .A(n16807), .B(n16808), .Z(n16809) );
  XOR U513 ( .A(n17352), .B(n17353), .Z(n17354) );
  NANDN U514 ( .A(n17663), .B(n17662), .Z(n247) );
  NANDN U515 ( .A(n17661), .B(n17660), .Z(n248) );
  NAND U516 ( .A(n247), .B(n248), .Z(n17780) );
  NAND U517 ( .A(n18528), .B(n18527), .Z(n249) );
  NANDN U518 ( .A(n18526), .B(n18525), .Z(n250) );
  NAND U519 ( .A(n249), .B(n250), .Z(n18620) );
  NAND U520 ( .A(n18564), .B(n18563), .Z(n251) );
  NANDN U521 ( .A(n18562), .B(n18561), .Z(n252) );
  NAND U522 ( .A(n251), .B(n252), .Z(n18646) );
  XOR U523 ( .A(n19049), .B(n19050), .Z(n19051) );
  NAND U524 ( .A(n1099), .B(n1098), .Z(n253) );
  NANDN U525 ( .A(n1097), .B(n1096), .Z(n254) );
  NAND U526 ( .A(n253), .B(n254), .Z(n1165) );
  OR U527 ( .A(n1082), .B(n1083), .Z(n255) );
  NAND U528 ( .A(n1080), .B(n1081), .Z(n256) );
  AND U529 ( .A(n255), .B(n256), .Z(n1091) );
  NAND U530 ( .A(n1561), .B(n1560), .Z(n257) );
  NANDN U531 ( .A(n1559), .B(n1558), .Z(n258) );
  NAND U532 ( .A(n257), .B(n258), .Z(n1569) );
  XOR U533 ( .A(n19151), .B(n19152), .Z(n19153) );
  XOR U534 ( .A(n19109), .B(n19110), .Z(n19111) );
  NAND U535 ( .A(n636), .B(n635), .Z(n259) );
  XOR U536 ( .A(n635), .B(n636), .Z(n260) );
  NANDN U537 ( .A(n634), .B(n260), .Z(n261) );
  NAND U538 ( .A(n259), .B(n261), .Z(n661) );
  OR U539 ( .A(n1037), .B(n1038), .Z(n262) );
  NAND U540 ( .A(n1036), .B(n1035), .Z(n263) );
  NAND U541 ( .A(n262), .B(n263), .Z(n1084) );
  NAND U542 ( .A(n2208), .B(n2209), .Z(n264) );
  NANDN U543 ( .A(n2207), .B(n2206), .Z(n265) );
  NAND U544 ( .A(n264), .B(n265), .Z(n2328) );
  NAND U545 ( .A(n3151), .B(n3150), .Z(n266) );
  NANDN U546 ( .A(n3149), .B(n3148), .Z(n267) );
  NAND U547 ( .A(n266), .B(n267), .Z(n3293) );
  NAND U548 ( .A(n4026), .B(n4025), .Z(n268) );
  NAND U549 ( .A(n4023), .B(n4024), .Z(n269) );
  NAND U550 ( .A(n268), .B(n269), .Z(n4173) );
  NAND U551 ( .A(n7662), .B(n7661), .Z(n270) );
  NAND U552 ( .A(n7659), .B(n7660), .Z(n271) );
  NAND U553 ( .A(n270), .B(n271), .Z(n7799) );
  NAND U554 ( .A(n9979), .B(n9978), .Z(n272) );
  NAND U555 ( .A(n9976), .B(n9977), .Z(n273) );
  NAND U556 ( .A(n272), .B(n273), .Z(n10117) );
  NAND U557 ( .A(n11005), .B(n11004), .Z(n274) );
  NAND U558 ( .A(n11002), .B(n11003), .Z(n275) );
  NAND U559 ( .A(n274), .B(n275), .Z(n11152) );
  NAND U560 ( .A(n14452), .B(n14451), .Z(n276) );
  NAND U561 ( .A(n14449), .B(n14450), .Z(n277) );
  NAND U562 ( .A(n276), .B(n277), .Z(n14592) );
  NAND U563 ( .A(n18459), .B(n18458), .Z(n278) );
  NANDN U564 ( .A(n18457), .B(n18456), .Z(n279) );
  NAND U565 ( .A(n278), .B(n279), .Z(n18628) );
  NAND U566 ( .A(n18731), .B(n18730), .Z(n280) );
  NANDN U567 ( .A(n18729), .B(n18728), .Z(n281) );
  NAND U568 ( .A(n280), .B(n281), .Z(n18809) );
  NANDN U569 ( .A(n19320), .B(n19319), .Z(n282) );
  NANDN U570 ( .A(n19322), .B(n19321), .Z(n283) );
  NAND U571 ( .A(n282), .B(n283), .Z(n19353) );
  NAND U572 ( .A(n19332), .B(n19331), .Z(n284) );
  NANDN U573 ( .A(n19330), .B(n19329), .Z(n285) );
  NAND U574 ( .A(n284), .B(n285), .Z(n19359) );
  OR U575 ( .A(n19366), .B(n19367), .Z(n286) );
  NAND U576 ( .A(n19365), .B(n19364), .Z(n287) );
  NAND U577 ( .A(n286), .B(n287), .Z(n19415) );
  NAND U578 ( .A(n17095), .B(n17096), .Z(n288) );
  NANDN U579 ( .A(n17094), .B(n17093), .Z(n289) );
  AND U580 ( .A(n288), .B(n289), .Z(n17231) );
  NAND U581 ( .A(n19262), .B(n19260), .Z(n290) );
  XOR U582 ( .A(n19260), .B(n19262), .Z(n291) );
  NANDN U583 ( .A(n19261), .B(n291), .Z(n292) );
  NAND U584 ( .A(n290), .B(n292), .Z(n19266) );
  NAND U585 ( .A(n19492), .B(n19490), .Z(n293) );
  XOR U586 ( .A(n19490), .B(n19492), .Z(n294) );
  NANDN U587 ( .A(n19491), .B(n294), .Z(n295) );
  NAND U588 ( .A(n293), .B(n295), .Z(n19504) );
  NANDN U589 ( .A(n2921), .B(b[29]), .Z(n296) );
  ANDN U590 ( .B(n296), .A(n585), .Z(n297) );
  XNOR U591 ( .A(b[29]), .B(n2921), .Z(n298) );
  NAND U592 ( .A(n298), .B(b[30]), .Z(n299) );
  NAND U593 ( .A(n297), .B(n299), .Z(n2904) );
  XNOR U594 ( .A(n3328), .B(n3329), .Z(n3331) );
  XNOR U595 ( .A(n3322), .B(n3323), .Z(n3325) );
  XOR U596 ( .A(n3316), .B(n3317), .Z(n3318) );
  XNOR U597 ( .A(n3311), .B(n3310), .Z(n3312) );
  XNOR U598 ( .A(n3481), .B(n3482), .Z(n3484) );
  XNOR U599 ( .A(n3630), .B(n3631), .Z(n3633) );
  XOR U600 ( .A(n3892), .B(n3893), .Z(n3894) );
  XNOR U601 ( .A(n3887), .B(n3886), .Z(n3888) );
  XOR U602 ( .A(n4039), .B(n4040), .Z(n4041) );
  XNOR U603 ( .A(n4034), .B(n4033), .Z(n4035) );
  XNOR U604 ( .A(n4373), .B(n4374), .Z(n4376) );
  XNOR U605 ( .A(n4648), .B(n4649), .Z(n4651) );
  XNOR U606 ( .A(n4642), .B(n4643), .Z(n4645) );
  XOR U607 ( .A(n4785), .B(n4786), .Z(n4787) );
  XNOR U608 ( .A(n4780), .B(n4779), .Z(n4781) );
  XOR U609 ( .A(n4917), .B(n4918), .Z(n4966) );
  XNOR U610 ( .A(n5110), .B(n5111), .Z(n5113) );
  XOR U611 ( .A(n5222), .B(n5223), .Z(n5224) );
  XOR U612 ( .A(n5216), .B(n5217), .Z(n5218) );
  XNOR U613 ( .A(n5957), .B(n5958), .Z(n5960) );
  XNOR U614 ( .A(n5951), .B(n5952), .Z(n5954) );
  XOR U615 ( .A(n5945), .B(n5946), .Z(n5947) );
  XNOR U616 ( .A(n5940), .B(n5939), .Z(n5941) );
  XNOR U617 ( .A(n6243), .B(n6244), .Z(n6246) );
  XNOR U618 ( .A(n6237), .B(n6238), .Z(n6240) );
  XOR U619 ( .A(n6231), .B(n6232), .Z(n6233) );
  XNOR U620 ( .A(n6226), .B(n6225), .Z(n6227) );
  XOR U621 ( .A(n7417), .B(n7418), .Z(n7419) );
  XNOR U622 ( .A(n7704), .B(n7703), .Z(n7705) );
  XNOR U623 ( .A(n8120), .B(n8121), .Z(n8123) );
  XNOR U624 ( .A(n8114), .B(n8115), .Z(n8117) );
  XOR U625 ( .A(n8108), .B(n8109), .Z(n8110) );
  XNOR U626 ( .A(n8103), .B(n8102), .Z(n8104) );
  XNOR U627 ( .A(n8578), .B(n8579), .Z(n8581) );
  XNOR U628 ( .A(n8723), .B(n8724), .Z(n8726) );
  XOR U629 ( .A(n8990), .B(n8991), .Z(n8992) );
  XOR U630 ( .A(n8984), .B(n8985), .Z(n8986) );
  XOR U631 ( .A(n9146), .B(n9147), .Z(n9148) );
  XNOR U632 ( .A(n9305), .B(n9306), .Z(n9308) );
  XNOR U633 ( .A(n9739), .B(n9738), .Z(n9740) );
  XNOR U634 ( .A(n10021), .B(n10020), .Z(n10022) );
  XNOR U635 ( .A(n10144), .B(n10145), .Z(n10147) );
  XNOR U636 ( .A(n10138), .B(n10139), .Z(n10141) );
  XOR U637 ( .A(n10132), .B(n10133), .Z(n10134) );
  XOR U638 ( .A(n10126), .B(n10127), .Z(n10128) );
  XNOR U639 ( .A(n10448), .B(n10449), .Z(n10451) );
  XNOR U640 ( .A(n10442), .B(n10443), .Z(n10445) );
  XOR U641 ( .A(n10436), .B(n10437), .Z(n10438) );
  XNOR U642 ( .A(n10431), .B(n10430), .Z(n10432) );
  XNOR U643 ( .A(n10747), .B(n10748), .Z(n10750) );
  XNOR U644 ( .A(n10741), .B(n10742), .Z(n10744) );
  XOR U645 ( .A(n10872), .B(n10873), .Z(n10874) );
  XNOR U646 ( .A(n10867), .B(n10866), .Z(n10868) );
  XNOR U647 ( .A(n11030), .B(n11031), .Z(n11033) );
  XNOR U648 ( .A(n11024), .B(n11025), .Z(n11027) );
  XOR U649 ( .A(n11018), .B(n11019), .Z(n11020) );
  XOR U650 ( .A(n11012), .B(n11013), .Z(n11014) );
  XOR U651 ( .A(n11749), .B(n11750), .Z(n11751) );
  XNOR U652 ( .A(n11744), .B(n11743), .Z(n11745) );
  XNOR U653 ( .A(n12080), .B(n12081), .Z(n12083) );
  XNOR U654 ( .A(n12201), .B(n12202), .Z(n12204) );
  XNOR U655 ( .A(n12195), .B(n12196), .Z(n12198) );
  XNOR U656 ( .A(n12563), .B(n12564), .Z(n12566) );
  XNOR U657 ( .A(n12634), .B(n12635), .Z(n12637) );
  XNOR U658 ( .A(n12628), .B(n12629), .Z(n12631) );
  XNOR U659 ( .A(n12931), .B(n12930), .Z(n12932) );
  XNOR U660 ( .A(n13510), .B(n13511), .Z(n13513) );
  XNOR U661 ( .A(n14212), .B(n14211), .Z(n14213) );
  XNOR U662 ( .A(n14495), .B(n14496), .Z(n14498) );
  XNOR U663 ( .A(n14652), .B(n14651), .Z(n14664) );
  XNOR U664 ( .A(n14796), .B(n14797), .Z(n14799) );
  XNOR U665 ( .A(n14919), .B(n14920), .Z(n14922) );
  XNOR U666 ( .A(n14913), .B(n14914), .Z(n14916) );
  XOR U667 ( .A(n14907), .B(n14908), .Z(n14909) );
  XNOR U668 ( .A(n14902), .B(n14901), .Z(n14903) );
  XNOR U669 ( .A(n15074), .B(n15075), .Z(n15077) );
  XNOR U670 ( .A(n15234), .B(n15235), .Z(n15237) );
  XNOR U671 ( .A(n15501), .B(n15502), .Z(n15504) );
  XNOR U672 ( .A(n15495), .B(n15496), .Z(n15498) );
  XOR U673 ( .A(n15489), .B(n15490), .Z(n15491) );
  XOR U674 ( .A(n15483), .B(n15484), .Z(n15485) );
  XNOR U675 ( .A(n15678), .B(n15679), .Z(n15681) );
  XNOR U676 ( .A(n15956), .B(n15957), .Z(n15959) );
  XNOR U677 ( .A(n15950), .B(n15951), .Z(n15953) );
  XOR U678 ( .A(n15944), .B(n15945), .Z(n15946) );
  XNOR U679 ( .A(n15939), .B(n15938), .Z(n15940) );
  ANDN U680 ( .B(n2921), .A(n582), .Z(n300) );
  AND U681 ( .A(n19015), .B(n300), .Z(n301) );
  NOR U682 ( .A(n582), .B(b[20]), .Z(n302) );
  NAND U683 ( .A(n302), .B(n581), .Z(n303) );
  NANDN U684 ( .A(n301), .B(n303), .Z(n1719) );
  XNOR U685 ( .A(n2022), .B(n2023), .Z(n2025) );
  NAND U686 ( .A(n2780), .B(n2779), .Z(n304) );
  NANDN U687 ( .A(n2778), .B(n2777), .Z(n305) );
  NAND U688 ( .A(n304), .B(n305), .Z(n2879) );
  NAND U689 ( .A(n3123), .B(n3122), .Z(n306) );
  NANDN U690 ( .A(n3121), .B(n3120), .Z(n307) );
  NAND U691 ( .A(n306), .B(n307), .Z(n3279) );
  NAND U692 ( .A(n3050), .B(n3049), .Z(n308) );
  NANDN U693 ( .A(n3048), .B(n3047), .Z(n309) );
  NAND U694 ( .A(n308), .B(n309), .Z(n3273) );
  NAND U695 ( .A(n3657), .B(n3656), .Z(n310) );
  NANDN U696 ( .A(n3655), .B(n3654), .Z(n311) );
  NAND U697 ( .A(n310), .B(n311), .Z(n3866) );
  XOR U698 ( .A(n3934), .B(n3935), .Z(n3936) );
  NAND U699 ( .A(n3816), .B(n3815), .Z(n312) );
  NANDN U700 ( .A(n3814), .B(n3813), .Z(n313) );
  NAND U701 ( .A(n312), .B(n313), .Z(n4001) );
  XNOR U702 ( .A(n4081), .B(n4082), .Z(n4084) );
  XNOR U703 ( .A(n4238), .B(n4239), .Z(n4241) );
  XOR U704 ( .A(n4678), .B(n4679), .Z(n4680) );
  NAND U705 ( .A(n4545), .B(n4544), .Z(n314) );
  NANDN U706 ( .A(n4543), .B(n4542), .Z(n315) );
  NAND U707 ( .A(n314), .B(n315), .Z(n4745) );
  XNOR U708 ( .A(n4957), .B(n4958), .Z(n4960) );
  XNOR U709 ( .A(n5399), .B(n5400), .Z(n5402) );
  XOR U710 ( .A(n5687), .B(n5688), .Z(n5689) );
  NAND U711 ( .A(n5702), .B(n5701), .Z(n316) );
  NANDN U712 ( .A(n5700), .B(n5699), .Z(n317) );
  NAND U713 ( .A(n316), .B(n317), .Z(n5785) );
  XOR U714 ( .A(n5987), .B(n5988), .Z(n5989) );
  XOR U715 ( .A(n6273), .B(n6274), .Z(n6275) );
  XOR U716 ( .A(n6567), .B(n6568), .Z(n6569) );
  NAND U717 ( .A(n6582), .B(n6581), .Z(n318) );
  NANDN U718 ( .A(n6580), .B(n6579), .Z(n319) );
  NAND U719 ( .A(n318), .B(n319), .Z(n6667) );
  XOR U720 ( .A(n6997), .B(n6998), .Z(n6999) );
  NAND U721 ( .A(n7012), .B(n7011), .Z(n320) );
  NANDN U722 ( .A(n7010), .B(n7009), .Z(n321) );
  NAND U723 ( .A(n320), .B(n321), .Z(n7097) );
  XOR U724 ( .A(n7439), .B(n7440), .Z(n7441) );
  NAND U725 ( .A(n7454), .B(n7453), .Z(n322) );
  NANDN U726 ( .A(n7452), .B(n7451), .Z(n323) );
  NAND U727 ( .A(n322), .B(n323), .Z(n7630) );
  XOR U728 ( .A(n7995), .B(n7996), .Z(n7997) );
  NAND U729 ( .A(n8010), .B(n8009), .Z(n324) );
  NANDN U730 ( .A(n8008), .B(n8007), .Z(n325) );
  NAND U731 ( .A(n324), .B(n325), .Z(n8093) );
  XOR U732 ( .A(n8444), .B(n8445), .Z(n8446) );
  NAND U733 ( .A(n8459), .B(n8458), .Z(n326) );
  NANDN U734 ( .A(n8457), .B(n8456), .Z(n327) );
  NAND U735 ( .A(n326), .B(n327), .Z(n8533) );
  XOR U736 ( .A(n9032), .B(n9033), .Z(n9034) );
  NAND U737 ( .A(n8899), .B(n8898), .Z(n328) );
  NANDN U738 ( .A(n8897), .B(n8896), .Z(n329) );
  NAND U739 ( .A(n328), .B(n329), .Z(n9100) );
  XNOR U740 ( .A(n9168), .B(n9169), .Z(n9171) );
  XOR U741 ( .A(n9617), .B(n9618), .Z(n9619) );
  NAND U742 ( .A(n9487), .B(n9486), .Z(n330) );
  NANDN U743 ( .A(n9485), .B(n9484), .Z(n331) );
  NAND U744 ( .A(n330), .B(n331), .Z(n9682) );
  NAND U745 ( .A(n9632), .B(n9631), .Z(n332) );
  NANDN U746 ( .A(n9630), .B(n9629), .Z(n333) );
  NAND U747 ( .A(n332), .B(n333), .Z(n9705) );
  NAND U748 ( .A(n9904), .B(n9903), .Z(n334) );
  NANDN U749 ( .A(n9902), .B(n9901), .Z(n335) );
  NAND U750 ( .A(n334), .B(n335), .Z(n9986) );
  XOR U751 ( .A(n10478), .B(n10479), .Z(n10480) );
  XOR U752 ( .A(n10777), .B(n10778), .Z(n10779) );
  XNOR U753 ( .A(n11060), .B(n11061), .Z(n11063) );
  XOR U754 ( .A(n11493), .B(n11494), .Z(n11495) );
  NAND U755 ( .A(n11375), .B(n11374), .Z(n336) );
  NANDN U756 ( .A(n11373), .B(n11372), .Z(n337) );
  NAND U757 ( .A(n336), .B(n337), .Z(n11558) );
  NAND U758 ( .A(n11508), .B(n11507), .Z(n338) );
  NANDN U759 ( .A(n11506), .B(n11505), .Z(n339) );
  NAND U760 ( .A(n338), .B(n339), .Z(n11697) );
  XOR U761 ( .A(n11791), .B(n11792), .Z(n11793) );
  XNOR U762 ( .A(n11926), .B(n11927), .Z(n11929) );
  XOR U763 ( .A(n13377), .B(n13378), .Z(n13379) );
  NAND U764 ( .A(n13249), .B(n13248), .Z(n340) );
  NANDN U765 ( .A(n13247), .B(n13246), .Z(n341) );
  NAND U766 ( .A(n340), .B(n341), .Z(n13442) );
  NAND U767 ( .A(n13392), .B(n13391), .Z(n342) );
  NANDN U768 ( .A(n13390), .B(n13389), .Z(n343) );
  NAND U769 ( .A(n342), .B(n343), .Z(n13465) );
  XOR U770 ( .A(n13800), .B(n13801), .Z(n13802) );
  NAND U771 ( .A(n13670), .B(n13669), .Z(n344) );
  NANDN U772 ( .A(n13668), .B(n13667), .Z(n345) );
  NAND U773 ( .A(n344), .B(n345), .Z(n13865) );
  NAND U774 ( .A(n13815), .B(n13814), .Z(n346) );
  NANDN U775 ( .A(n13813), .B(n13812), .Z(n347) );
  NAND U776 ( .A(n346), .B(n347), .Z(n14002) );
  NAND U777 ( .A(n14107), .B(n14106), .Z(n348) );
  NANDN U778 ( .A(n14105), .B(n14104), .Z(n349) );
  NAND U779 ( .A(n348), .B(n349), .Z(n14178) );
  NAND U780 ( .A(n14331), .B(n14330), .Z(n350) );
  NANDN U781 ( .A(n14329), .B(n14328), .Z(n351) );
  NAND U782 ( .A(n350), .B(n351), .Z(n14564) );
  NAND U783 ( .A(n14670), .B(n14669), .Z(n352) );
  NANDN U784 ( .A(n14668), .B(n14667), .Z(n353) );
  NAND U785 ( .A(n352), .B(n353), .Z(n14743) );
  NAND U786 ( .A(n15261), .B(n15260), .Z(n354) );
  NANDN U787 ( .A(n15259), .B(n15258), .Z(n355) );
  NAND U788 ( .A(n354), .B(n355), .Z(n15449) );
  XOR U789 ( .A(n15531), .B(n15532), .Z(n15533) );
  XOR U790 ( .A(n15986), .B(n15987), .Z(n15988) );
  NAND U791 ( .A(n15854), .B(n15853), .Z(n356) );
  NANDN U792 ( .A(n15852), .B(n15851), .Z(n357) );
  NAND U793 ( .A(n356), .B(n357), .Z(n16053) );
  XOR U794 ( .A(n16282), .B(n16283), .Z(n16284) );
  XNOR U795 ( .A(n16908), .B(n16909), .Z(n16911) );
  XNOR U796 ( .A(n17602), .B(n17603), .Z(n17615) );
  XOR U797 ( .A(n18505), .B(n18506), .Z(n18507) );
  NANDN U798 ( .A(a[0]), .B(n18336), .Z(n358) );
  OR U799 ( .A(b[11]), .B(b[12]), .Z(n359) );
  NAND U800 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U801 ( .A(n580), .B(n360), .Z(n1056) );
  NAND U802 ( .A(n1898), .B(n1899), .Z(n361) );
  NANDN U803 ( .A(n1897), .B(n1896), .Z(n362) );
  AND U804 ( .A(n361), .B(n362), .Z(n1980) );
  NAND U805 ( .A(n2231), .B(n2230), .Z(n363) );
  NANDN U806 ( .A(n2229), .B(n2228), .Z(n364) );
  NAND U807 ( .A(n363), .B(n364), .Z(n2426) );
  XOR U808 ( .A(n3422), .B(n3423), .Z(n3424) );
  NAND U809 ( .A(n3309), .B(n3308), .Z(n365) );
  NAND U810 ( .A(n3306), .B(n3307), .Z(n366) );
  NAND U811 ( .A(n365), .B(n366), .Z(n3566) );
  XNOR U812 ( .A(n3720), .B(n3721), .Z(n3715) );
  XNOR U813 ( .A(n3749), .B(n3750), .Z(n3744) );
  XNOR U814 ( .A(n4014), .B(n4015), .Z(n4009) );
  NAND U815 ( .A(n4334), .B(n4333), .Z(n367) );
  NANDN U816 ( .A(n4336), .B(n4335), .Z(n368) );
  NAND U817 ( .A(n367), .B(n368), .Z(n4471) );
  XNOR U818 ( .A(n4626), .B(n4627), .Z(n4621) );
  NAND U819 ( .A(n4891), .B(n4890), .Z(n369) );
  NAND U820 ( .A(n4888), .B(n4889), .Z(n370) );
  NAND U821 ( .A(n369), .B(n370), .Z(n5030) );
  OR U822 ( .A(n5117), .B(n5116), .Z(n371) );
  NANDN U823 ( .A(n5119), .B(n5118), .Z(n372) );
  NAND U824 ( .A(n371), .B(n372), .Z(n5331) );
  NAND U825 ( .A(n5613), .B(n5612), .Z(n373) );
  NANDN U826 ( .A(n5611), .B(n5610), .Z(n374) );
  NAND U827 ( .A(n373), .B(n374), .Z(n5762) );
  NAND U828 ( .A(n5791), .B(n5790), .Z(n375) );
  NANDN U829 ( .A(n5793), .B(n5792), .Z(n376) );
  NAND U830 ( .A(n375), .B(n376), .Z(n5928) );
  XNOR U831 ( .A(n6353), .B(n6354), .Z(n6348) );
  XNOR U832 ( .A(n6645), .B(n6646), .Z(n6640) );
  NAND U833 ( .A(n6673), .B(n6672), .Z(n377) );
  NANDN U834 ( .A(n6675), .B(n6674), .Z(n378) );
  NAND U835 ( .A(n377), .B(n378), .Z(n6923) );
  NAND U836 ( .A(n6816), .B(n6815), .Z(n379) );
  NAND U837 ( .A(n6813), .B(n6814), .Z(n380) );
  NAND U838 ( .A(n379), .B(n380), .Z(n7068) );
  NAND U839 ( .A(n7103), .B(n7102), .Z(n381) );
  NANDN U840 ( .A(n7105), .B(n7104), .Z(n382) );
  NAND U841 ( .A(n381), .B(n382), .Z(n7353) );
  NAND U842 ( .A(n7246), .B(n7245), .Z(n383) );
  NAND U843 ( .A(n7243), .B(n7244), .Z(n384) );
  NAND U844 ( .A(n383), .B(n384), .Z(n7382) );
  OR U845 ( .A(n7574), .B(n7575), .Z(n385) );
  NAND U846 ( .A(n7573), .B(n7572), .Z(n386) );
  NAND U847 ( .A(n385), .B(n386), .Z(n7781) );
  NAND U848 ( .A(n7678), .B(n7677), .Z(n387) );
  NAND U849 ( .A(n7675), .B(n7676), .Z(n388) );
  NAND U850 ( .A(n387), .B(n388), .Z(n7925) );
  NAND U851 ( .A(n8099), .B(n8098), .Z(n389) );
  NANDN U852 ( .A(n8101), .B(n8100), .Z(n390) );
  NAND U853 ( .A(n389), .B(n390), .Z(n8358) );
  XNOR U854 ( .A(n8394), .B(n8395), .Z(n8389) );
  NAND U855 ( .A(n8539), .B(n8538), .Z(n391) );
  NANDN U856 ( .A(n8541), .B(n8540), .Z(n392) );
  NAND U857 ( .A(n391), .B(n392), .Z(n8676) );
  XNOR U858 ( .A(n8832), .B(n8833), .Z(n8827) );
  XNOR U859 ( .A(n8980), .B(n8981), .Z(n8975) );
  XNOR U860 ( .A(n9567), .B(n9568), .Z(n9562) );
  NAND U861 ( .A(n9711), .B(n9710), .Z(n393) );
  NANDN U862 ( .A(n9713), .B(n9712), .Z(n394) );
  NAND U863 ( .A(n393), .B(n394), .Z(n9960) );
  OR U864 ( .A(n9893), .B(n9894), .Z(n395) );
  NAND U865 ( .A(n9892), .B(n9891), .Z(n396) );
  NAND U866 ( .A(n395), .B(n396), .Z(n10099) );
  NAND U867 ( .A(n9995), .B(n9994), .Z(n397) );
  NAND U868 ( .A(n9992), .B(n9993), .Z(n398) );
  NAND U869 ( .A(n397), .B(n398), .Z(n10245) );
  OR U870 ( .A(n10176), .B(n10177), .Z(n399) );
  NAND U871 ( .A(n10175), .B(n10174), .Z(n400) );
  NAND U872 ( .A(n399), .B(n400), .Z(n10389) );
  XNOR U873 ( .A(n10426), .B(n10427), .Z(n10421) );
  XNOR U874 ( .A(n10725), .B(n10726), .Z(n10720) );
  NAND U875 ( .A(n10978), .B(n10977), .Z(n401) );
  NAND U876 ( .A(n10975), .B(n10976), .Z(n402) );
  NAND U877 ( .A(n401), .B(n402), .Z(n11133) );
  XNOR U878 ( .A(n11426), .B(n11427), .Z(n11421) );
  NAND U879 ( .A(n11365), .B(n11364), .Z(n403) );
  NANDN U880 ( .A(n11363), .B(n11362), .Z(n404) );
  NAND U881 ( .A(n403), .B(n404), .Z(n11570) );
  OR U882 ( .A(n11308), .B(n11309), .Z(n405) );
  NAND U883 ( .A(n11307), .B(n11306), .Z(n406) );
  NAND U884 ( .A(n405), .B(n406), .Z(n11563) );
  NAND U885 ( .A(n11705), .B(n11704), .Z(n407) );
  NANDN U886 ( .A(n11703), .B(n11702), .Z(n408) );
  NAND U887 ( .A(n407), .B(n408), .Z(n11738) );
  NAND U888 ( .A(n12034), .B(n12033), .Z(n409) );
  NANDN U889 ( .A(n12036), .B(n12035), .Z(n410) );
  NAND U890 ( .A(n409), .B(n410), .Z(n12292) );
  NAND U891 ( .A(n12429), .B(n12428), .Z(n411) );
  NANDN U892 ( .A(n12427), .B(n12426), .Z(n412) );
  NAND U893 ( .A(n411), .B(n412), .Z(n12580) );
  NAND U894 ( .A(n12578), .B(n12577), .Z(n413) );
  NANDN U895 ( .A(n12576), .B(n12575), .Z(n414) );
  NAND U896 ( .A(n413), .B(n414), .Z(n12729) );
  NAND U897 ( .A(n12860), .B(n12859), .Z(n415) );
  NANDN U898 ( .A(n12858), .B(n12857), .Z(n416) );
  NAND U899 ( .A(n415), .B(n416), .Z(n13009) );
  NAND U900 ( .A(n12903), .B(n12902), .Z(n417) );
  NANDN U901 ( .A(n12905), .B(n12904), .Z(n418) );
  NAND U902 ( .A(n417), .B(n418), .Z(n13152) );
  NAND U903 ( .A(n13239), .B(n13238), .Z(n419) );
  NANDN U904 ( .A(n13237), .B(n13236), .Z(n420) );
  NAND U905 ( .A(n419), .B(n420), .Z(n13326) );
  NAND U906 ( .A(n13471), .B(n13470), .Z(n421) );
  NANDN U907 ( .A(n13473), .B(n13472), .Z(n422) );
  NAND U908 ( .A(n421), .B(n422), .Z(n13726) );
  XNOR U909 ( .A(n13878), .B(n13879), .Z(n13873) );
  NAND U910 ( .A(n14010), .B(n14009), .Z(n423) );
  NANDN U911 ( .A(n14008), .B(n14007), .Z(n424) );
  NAND U912 ( .A(n423), .B(n424), .Z(n14155) );
  NAND U913 ( .A(n14097), .B(n14096), .Z(n425) );
  NANDN U914 ( .A(n14095), .B(n14094), .Z(n426) );
  NAND U915 ( .A(n425), .B(n426), .Z(n14296) );
  NAND U916 ( .A(n14186), .B(n14185), .Z(n427) );
  NAND U917 ( .A(n14183), .B(n14184), .Z(n428) );
  NAND U918 ( .A(n427), .B(n428), .Z(n14433) );
  OR U919 ( .A(n14320), .B(n14321), .Z(n429) );
  NAND U920 ( .A(n14319), .B(n14318), .Z(n430) );
  NAND U921 ( .A(n429), .B(n430), .Z(n14574) );
  NAND U922 ( .A(n14573), .B(n14572), .Z(n431) );
  NANDN U923 ( .A(n14571), .B(n14570), .Z(n432) );
  NAND U924 ( .A(n431), .B(n432), .Z(n14604) );
  XNOR U925 ( .A(n14868), .B(n14869), .Z(n14863) );
  NANDN U926 ( .A(n14803), .B(n14802), .Z(n433) );
  NANDN U927 ( .A(n14805), .B(n14804), .Z(n434) );
  NAND U928 ( .A(n433), .B(n434), .Z(n15016) );
  XNOR U929 ( .A(n15194), .B(n15195), .Z(n15189) );
  XNOR U930 ( .A(n15462), .B(n15463), .Z(n15457) );
  XNOR U931 ( .A(n15611), .B(n15612), .Z(n15606) );
  XNOR U932 ( .A(n15787), .B(n15788), .Z(n15782) );
  XNOR U933 ( .A(n15934), .B(n15935), .Z(n15929) );
  XNOR U934 ( .A(n16232), .B(n16233), .Z(n16227) );
  NAND U935 ( .A(n16297), .B(n16296), .Z(n435) );
  NANDN U936 ( .A(n16295), .B(n16294), .Z(n436) );
  NAND U937 ( .A(n435), .B(n436), .Z(n16369) );
  XNOR U938 ( .A(n16762), .B(n16763), .Z(n16765) );
  XNOR U939 ( .A(n16756), .B(n16757), .Z(n16758) );
  NAND U940 ( .A(n17921), .B(n17920), .Z(n437) );
  NANDN U941 ( .A(n17923), .B(n17922), .Z(n438) );
  NAND U942 ( .A(n437), .B(n438), .Z(n18111) );
  NANDN U943 ( .A(n18402), .B(n18401), .Z(n439) );
  NANDN U944 ( .A(n18404), .B(n18403), .Z(n440) );
  NAND U945 ( .A(n439), .B(n440), .Z(n18460) );
  NANDN U946 ( .A(n2921), .B(b[9]), .Z(n441) );
  AND U947 ( .A(b[11]), .B(n441), .Z(n442) );
  XNOR U948 ( .A(n2921), .B(b[9]), .Z(n443) );
  NAND U949 ( .A(n443), .B(b[10]), .Z(n444) );
  AND U950 ( .A(n442), .B(n444), .Z(n922) );
  NAND U951 ( .A(n1191), .B(n1190), .Z(n445) );
  NANDN U952 ( .A(n1189), .B(n1188), .Z(n446) );
  NAND U953 ( .A(n445), .B(n446), .Z(n1237) );
  NAND U954 ( .A(n1385), .B(n1384), .Z(n447) );
  NANDN U955 ( .A(n1383), .B(n1382), .Z(n448) );
  AND U956 ( .A(n447), .B(n448), .Z(n1398) );
  NAND U957 ( .A(n1601), .B(n1600), .Z(n449) );
  NAND U958 ( .A(n1598), .B(n1599), .Z(n450) );
  NAND U959 ( .A(n449), .B(n450), .Z(n1668) );
  NANDN U960 ( .A(n2438), .B(n2437), .Z(n451) );
  NANDN U961 ( .A(n2436), .B(n2435), .Z(n452) );
  AND U962 ( .A(n451), .B(n452), .Z(n2457) );
  NAND U963 ( .A(n2595), .B(n2594), .Z(n453) );
  NANDN U964 ( .A(n2593), .B(n2592), .Z(n454) );
  NAND U965 ( .A(n453), .B(n454), .Z(n2727) );
  NANDN U966 ( .A(n5758), .B(n5757), .Z(n455) );
  NANDN U967 ( .A(n5760), .B(n5759), .Z(n456) );
  NAND U968 ( .A(n455), .B(n456), .Z(n5778) );
  NANDN U969 ( .A(n8066), .B(n8065), .Z(n457) );
  NANDN U970 ( .A(n8068), .B(n8067), .Z(n458) );
  NAND U971 ( .A(n457), .B(n458), .Z(n8086) );
  NANDN U972 ( .A(n9415), .B(n9414), .Z(n459) );
  NANDN U973 ( .A(n9417), .B(n9416), .Z(n460) );
  NAND U974 ( .A(n459), .B(n460), .Z(n9553) );
  NANDN U975 ( .A(n11734), .B(n11733), .Z(n461) );
  NANDN U976 ( .A(n11736), .B(n11735), .Z(n462) );
  NAND U977 ( .A(n461), .B(n462), .Z(n11874) );
  NAND U978 ( .A(n12726), .B(n12727), .Z(n463) );
  NANDN U979 ( .A(n12725), .B(n12724), .Z(n464) );
  NAND U980 ( .A(n463), .B(n464), .Z(n12745) );
  NANDN U981 ( .A(n13293), .B(n13292), .Z(n465) );
  NANDN U982 ( .A(n13295), .B(n13294), .Z(n466) );
  NAND U983 ( .A(n465), .B(n466), .Z(n13313) );
  NANDN U984 ( .A(n14151), .B(n14150), .Z(n467) );
  NANDN U985 ( .A(n14153), .B(n14152), .Z(n468) );
  NAND U986 ( .A(n467), .B(n468), .Z(n14171) );
  NANDN U987 ( .A(n14600), .B(n14599), .Z(n469) );
  NANDN U988 ( .A(n14602), .B(n14601), .Z(n470) );
  NAND U989 ( .A(n469), .B(n470), .Z(n14736) );
  NAND U990 ( .A(n16376), .B(n16375), .Z(n471) );
  NANDN U991 ( .A(n16378), .B(n16377), .Z(n472) );
  NAND U992 ( .A(n471), .B(n472), .Z(n16634) );
  NAND U993 ( .A(n17667), .B(n17666), .Z(n473) );
  NANDN U994 ( .A(n17665), .B(n17664), .Z(n474) );
  NAND U995 ( .A(n473), .B(n474), .Z(n17867) );
  NAND U996 ( .A(n18035), .B(n18034), .Z(n475) );
  NANDN U997 ( .A(n18033), .B(n18032), .Z(n476) );
  NAND U998 ( .A(n475), .B(n476), .Z(n18229) );
  NAND U999 ( .A(n696), .B(n695), .Z(n477) );
  NANDN U1000 ( .A(n694), .B(n693), .Z(n478) );
  NAND U1001 ( .A(n477), .B(n478), .Z(n738) );
  NANDN U1002 ( .A(n847), .B(n846), .Z(n479) );
  NANDN U1003 ( .A(n849), .B(n848), .Z(n480) );
  AND U1004 ( .A(n479), .B(n480), .Z(n857) );
  NANDN U1005 ( .A(n1326), .B(n1325), .Z(n481) );
  NANDN U1006 ( .A(n1328), .B(n1327), .Z(n482) );
  NAND U1007 ( .A(n481), .B(n482), .Z(n1392) );
  NANDN U1008 ( .A(n1664), .B(n1663), .Z(n483) );
  NANDN U1009 ( .A(n1666), .B(n1665), .Z(n484) );
  NAND U1010 ( .A(n483), .B(n484), .Z(n1756) );
  NAND U1011 ( .A(n16665), .B(n16664), .Z(n485) );
  NANDN U1012 ( .A(n16663), .B(n16662), .Z(n486) );
  NAND U1013 ( .A(n485), .B(n486), .Z(n16932) );
  XNOR U1014 ( .A(n17075), .B(n17076), .Z(n17078) );
  NAND U1015 ( .A(n17351), .B(n17350), .Z(n487) );
  NAND U1016 ( .A(n17348), .B(n17349), .Z(n488) );
  NAND U1017 ( .A(n487), .B(n488), .Z(n17372) );
  NAND U1018 ( .A(n17387), .B(n17386), .Z(n489) );
  NANDN U1019 ( .A(n17385), .B(n17384), .Z(n490) );
  NAND U1020 ( .A(n489), .B(n490), .Z(n17511) );
  NAND U1021 ( .A(n17652), .B(n17653), .Z(n491) );
  NANDN U1022 ( .A(n17651), .B(n17650), .Z(n492) );
  NAND U1023 ( .A(n491), .B(n492), .Z(n17774) );
  NANDN U1024 ( .A(n18648), .B(n18647), .Z(n493) );
  NANDN U1025 ( .A(n18646), .B(n18645), .Z(n494) );
  NAND U1026 ( .A(n493), .B(n494), .Z(n18793) );
  OR U1027 ( .A(n18970), .B(n18971), .Z(n495) );
  NAND U1028 ( .A(n18969), .B(n18968), .Z(n496) );
  NAND U1029 ( .A(n495), .B(n496), .Z(n19033) );
  XNOR U1030 ( .A(n19070), .B(n19069), .Z(n19046) );
  NAND U1031 ( .A(n19270), .B(n19269), .Z(n497) );
  NANDN U1032 ( .A(n19268), .B(n19267), .Z(n498) );
  NAND U1033 ( .A(n497), .B(n498), .Z(n19322) );
  NANDN U1034 ( .A(n1569), .B(n1568), .Z(n499) );
  NANDN U1035 ( .A(n1571), .B(n1570), .Z(n500) );
  NAND U1036 ( .A(n499), .B(n500), .Z(n1657) );
  NAND U1037 ( .A(n3293), .B(n3292), .Z(n501) );
  NANDN U1038 ( .A(n3291), .B(n3290), .Z(n502) );
  NAND U1039 ( .A(n501), .B(n502), .Z(n3436) );
  NAND U1040 ( .A(n4173), .B(n4172), .Z(n503) );
  NAND U1041 ( .A(n4170), .B(n4171), .Z(n504) );
  NAND U1042 ( .A(n503), .B(n504), .Z(n4318) );
  NAND U1043 ( .A(n5049), .B(n5048), .Z(n505) );
  NAND U1044 ( .A(n5046), .B(n5047), .Z(n506) );
  NAND U1045 ( .A(n505), .B(n506), .Z(n5195) );
  NAND U1046 ( .A(n5634), .B(n5633), .Z(n507) );
  NAND U1047 ( .A(n5631), .B(n5632), .Z(n508) );
  NAND U1048 ( .A(n507), .B(n508), .Z(n5775) );
  NAND U1049 ( .A(n6365), .B(n6364), .Z(n509) );
  NAND U1050 ( .A(n6362), .B(n6363), .Z(n510) );
  NAND U1051 ( .A(n509), .B(n510), .Z(n6512) );
  NAND U1052 ( .A(n7942), .B(n7941), .Z(n511) );
  NAND U1053 ( .A(n7939), .B(n7940), .Z(n512) );
  NAND U1054 ( .A(n511), .B(n512), .Z(n8083) );
  NAND U1055 ( .A(n9407), .B(n9406), .Z(n513) );
  NAND U1056 ( .A(n9404), .B(n9405), .Z(n514) );
  NAND U1057 ( .A(n513), .B(n514), .Z(n9550) );
  NAND U1058 ( .A(n10262), .B(n10261), .Z(n515) );
  NAND U1059 ( .A(n10259), .B(n10260), .Z(n516) );
  NAND U1060 ( .A(n515), .B(n516), .Z(n10409) );
  NAND U1061 ( .A(n11152), .B(n11151), .Z(n517) );
  NAND U1062 ( .A(n11149), .B(n11150), .Z(n518) );
  NAND U1063 ( .A(n517), .B(n518), .Z(n11297) );
  NAND U1064 ( .A(n11726), .B(n11725), .Z(n519) );
  NAND U1065 ( .A(n11723), .B(n11724), .Z(n520) );
  NAND U1066 ( .A(n519), .B(n520), .Z(n11871) );
  NAND U1067 ( .A(n12599), .B(n12598), .Z(n521) );
  NAND U1068 ( .A(n12596), .B(n12597), .Z(n522) );
  NAND U1069 ( .A(n521), .B(n522), .Z(n12742) );
  NAND U1070 ( .A(n13171), .B(n13170), .Z(n523) );
  NAND U1071 ( .A(n13168), .B(n13169), .Z(n524) );
  NAND U1072 ( .A(n523), .B(n524), .Z(n13310) );
  NAND U1073 ( .A(n14031), .B(n14030), .Z(n525) );
  NAND U1074 ( .A(n14028), .B(n14029), .Z(n526) );
  NAND U1075 ( .A(n525), .B(n526), .Z(n14168) );
  NAND U1076 ( .A(n14592), .B(n14591), .Z(n527) );
  NAND U1077 ( .A(n14589), .B(n14590), .Z(n528) );
  NAND U1078 ( .A(n527), .B(n528), .Z(n14733) );
  NAND U1079 ( .A(n15623), .B(n15622), .Z(n529) );
  NAND U1080 ( .A(n15620), .B(n15621), .Z(n530) );
  NAND U1081 ( .A(n529), .B(n530), .Z(n15770) );
  NANDN U1082 ( .A(n18713), .B(n18712), .Z(n531) );
  NANDN U1083 ( .A(n18711), .B(n18710), .Z(n532) );
  AND U1084 ( .A(n531), .B(n532), .Z(n18717) );
  NAND U1085 ( .A(n19411), .B(n19412), .Z(n533) );
  NANDN U1086 ( .A(n19410), .B(n19451), .Z(n534) );
  AND U1087 ( .A(n533), .B(n534), .Z(n19430) );
  XOR U1088 ( .A(n632), .B(n631), .Z(n535) );
  NANDN U1089 ( .A(n630), .B(n535), .Z(n536) );
  NAND U1090 ( .A(n632), .B(n631), .Z(n537) );
  AND U1091 ( .A(n536), .B(n537), .Z(n636) );
  NAND U1092 ( .A(n816), .B(n815), .Z(n538) );
  NANDN U1093 ( .A(n814), .B(n813), .Z(n539) );
  NAND U1094 ( .A(n538), .B(n539), .Z(n853) );
  NAND U1095 ( .A(n1163), .B(n1162), .Z(n540) );
  NANDN U1096 ( .A(n1161), .B(n1160), .Z(n541) );
  NAND U1097 ( .A(n540), .B(n541), .Z(n1227) );
  NAND U1098 ( .A(n2330), .B(n2329), .Z(n542) );
  NAND U1099 ( .A(n2327), .B(n2328), .Z(n543) );
  NAND U1100 ( .A(n542), .B(n543), .Z(n2448) );
  NAND U1101 ( .A(n17232), .B(n17230), .Z(n544) );
  XOR U1102 ( .A(n17230), .B(n17232), .Z(n545) );
  NANDN U1103 ( .A(n17231), .B(n545), .Z(n546) );
  NAND U1104 ( .A(n544), .B(n546), .Z(n17369) );
  NAND U1105 ( .A(n18542), .B(n18541), .Z(n547) );
  XOR U1106 ( .A(n18541), .B(n18542), .Z(n548) );
  NAND U1107 ( .A(n548), .B(n18540), .Z(n549) );
  NAND U1108 ( .A(n547), .B(n549), .Z(n18635) );
  NAND U1109 ( .A(n18881), .B(n18880), .Z(n550) );
  XOR U1110 ( .A(n18880), .B(n18881), .Z(n551) );
  NANDN U1111 ( .A(n18882), .B(n551), .Z(n552) );
  NAND U1112 ( .A(n550), .B(n552), .Z(n18958) );
  XNOR U1113 ( .A(n19209), .B(n19210), .Z(n19204) );
  NAND U1114 ( .A(n19266), .B(n19265), .Z(n553) );
  XOR U1115 ( .A(n19265), .B(n19266), .Z(n554) );
  NAND U1116 ( .A(n554), .B(n19264), .Z(n555) );
  NAND U1117 ( .A(n553), .B(n555), .Z(n19315) );
  XOR U1118 ( .A(n19395), .B(n19394), .Z(n556) );
  NANDN U1119 ( .A(n19393), .B(n556), .Z(n557) );
  NAND U1120 ( .A(n19395), .B(n19394), .Z(n558) );
  AND U1121 ( .A(n557), .B(n558), .Z(n19425) );
  XNOR U1122 ( .A(n584), .B(b[31]), .Z(n559) );
  ANDN U1123 ( .B(n559), .A(b[30]), .Z(n560) );
  NOR U1124 ( .A(n560), .B(n19502), .Z(n561) );
  NANDN U1125 ( .A(b[29]), .B(n585), .Z(n562) );
  AND U1126 ( .A(n561), .B(n562), .Z(n563) );
  NANDN U1127 ( .A(n19505), .B(n19503), .Z(n564) );
  XNOR U1128 ( .A(n19505), .B(n19503), .Z(n565) );
  NAND U1129 ( .A(n565), .B(n19504), .Z(n566) );
  NAND U1130 ( .A(n564), .B(n566), .Z(n567) );
  XNOR U1131 ( .A(n563), .B(n567), .Z(n568) );
  OR U1132 ( .A(n19506), .B(n19507), .Z(n569) );
  XNOR U1133 ( .A(n19507), .B(n19508), .Z(n570) );
  NANDN U1134 ( .A(n19509), .B(n570), .Z(n571) );
  AND U1135 ( .A(n569), .B(n571), .Z(n572) );
  ANDN U1136 ( .B(n19511), .A(n19510), .Z(n573) );
  XNOR U1137 ( .A(n568), .B(n572), .Z(n574) );
  XNOR U1138 ( .A(n573), .B(n574), .Z(c[255]) );
  XOR U1139 ( .A(b[27]), .B(b[28]), .Z(n575) );
  IV U1140 ( .A(n575), .Z(n576) );
  IV U1141 ( .A(b[0]), .Z(n577) );
  IV U1142 ( .A(b[3]), .Z(n578) );
  IV U1143 ( .A(b[9]), .Z(n579) );
  IV U1144 ( .A(b[13]), .Z(n580) );
  IV U1145 ( .A(b[19]), .Z(n581) );
  IV U1146 ( .A(b[21]), .Z(n582) );
  IV U1147 ( .A(b[27]), .Z(n583) );
  IV U1148 ( .A(b[29]), .Z(n584) );
  IV U1149 ( .A(b[31]), .Z(n585) );
  NANDN U1150 ( .A(n577), .B(a[0]), .Z(n587) );
  XNOR U1151 ( .A(n587), .B(sreg[96]), .Z(c[96]) );
  IV U1152 ( .A(b[1]), .Z(n17151) );
  ANDN U1153 ( .B(a[0]), .A(n17151), .Z(n586) );
  NANDN U1154 ( .A(n577), .B(a[1]), .Z(n592) );
  XNOR U1155 ( .A(n586), .B(n592), .Z(n595) );
  XNOR U1156 ( .A(sreg[97]), .B(n595), .Z(n597) );
  NANDN U1157 ( .A(n587), .B(sreg[96]), .Z(n596) );
  XOR U1158 ( .A(n597), .B(n596), .Z(c[97]) );
  NANDN U1159 ( .A(n577), .B(a[2]), .Z(n588) );
  XOR U1160 ( .A(n17151), .B(n588), .Z(n590) );
  NANDN U1161 ( .A(b[0]), .B(a[1]), .Z(n589) );
  AND U1162 ( .A(n590), .B(n589), .Z(n600) );
  IV U1163 ( .A(a[0]), .Z(n2921) );
  NANDN U1164 ( .A(n2921), .B(b[2]), .Z(n591) );
  XOR U1165 ( .A(n17151), .B(n591), .Z(n594) );
  OR U1166 ( .A(n592), .B(a[0]), .Z(n593) );
  AND U1167 ( .A(n594), .B(n593), .Z(n601) );
  XOR U1168 ( .A(n600), .B(n601), .Z(n611) );
  NAND U1169 ( .A(sreg[97]), .B(n595), .Z(n599) );
  OR U1170 ( .A(n597), .B(n596), .Z(n598) );
  NAND U1171 ( .A(n599), .B(n598), .Z(n610) );
  XNOR U1172 ( .A(n610), .B(sreg[98]), .Z(n612) );
  XNOR U1173 ( .A(n611), .B(n612), .Z(c[98]) );
  NAND U1174 ( .A(n601), .B(n600), .Z(n632) );
  XNOR U1175 ( .A(n17151), .B(b[2]), .Z(n16990) );
  NANDN U1176 ( .A(n577), .B(a[3]), .Z(n602) );
  XOR U1177 ( .A(n17151), .B(n602), .Z(n604) );
  NANDN U1178 ( .A(b[0]), .B(a[2]), .Z(n603) );
  AND U1179 ( .A(n604), .B(n603), .Z(n620) );
  XNOR U1180 ( .A(n578), .B(a[0]), .Z(n606) );
  XNOR U1181 ( .A(n578), .B(b[1]), .Z(n626) );
  XNOR U1182 ( .A(n578), .B(b[2]), .Z(n625) );
  AND U1183 ( .A(n626), .B(n625), .Z(n605) );
  NAND U1184 ( .A(n606), .B(n605), .Z(n608) );
  XNOR U1185 ( .A(b[3]), .B(a[1]), .Z(n627) );
  NANDN U1186 ( .A(n627), .B(n16990), .Z(n607) );
  AND U1187 ( .A(n608), .B(n607), .Z(n621) );
  XNOR U1188 ( .A(n620), .B(n621), .Z(n630) );
  XNOR U1189 ( .A(n631), .B(n630), .Z(n609) );
  XNOR U1190 ( .A(n632), .B(n609), .Z(n615) );
  XNOR U1191 ( .A(sreg[99]), .B(n615), .Z(n617) );
  NAND U1192 ( .A(n610), .B(sreg[98]), .Z(n614) );
  NANDN U1193 ( .A(n612), .B(n611), .Z(n613) );
  AND U1194 ( .A(n614), .B(n613), .Z(n616) );
  XOR U1195 ( .A(n617), .B(n616), .Z(c[99]) );
  NAND U1196 ( .A(sreg[99]), .B(n615), .Z(n619) );
  OR U1197 ( .A(n617), .B(n616), .Z(n618) );
  NAND U1198 ( .A(n619), .B(n618), .Z(n654) );
  XNOR U1199 ( .A(n654), .B(sreg[100]), .Z(n656) );
  NANDN U1200 ( .A(n621), .B(n620), .Z(n634) );
  NANDN U1201 ( .A(n577), .B(a[4]), .Z(n622) );
  XOR U1202 ( .A(n17151), .B(n622), .Z(n624) );
  NANDN U1203 ( .A(b[0]), .B(a[3]), .Z(n623) );
  AND U1204 ( .A(n624), .B(n623), .Z(n648) );
  NAND U1205 ( .A(n626), .B(n625), .Z(n16988) );
  OR U1206 ( .A(n627), .B(n16988), .Z(n629) );
  XNOR U1207 ( .A(b[3]), .B(a[2]), .Z(n645) );
  NANDN U1208 ( .A(n645), .B(n16990), .Z(n628) );
  AND U1209 ( .A(n629), .B(n628), .Z(n649) );
  XOR U1210 ( .A(n648), .B(n649), .Z(n651) );
  XOR U1211 ( .A(b[3]), .B(b[4]), .Z(n17310) );
  NANDN U1212 ( .A(n2921), .B(n17310), .Z(n650) );
  XOR U1213 ( .A(n651), .B(n650), .Z(n635) );
  XOR U1214 ( .A(n635), .B(n636), .Z(n633) );
  XNOR U1215 ( .A(n634), .B(n633), .Z(n655) );
  XNOR U1216 ( .A(n656), .B(n655), .Z(c[100]) );
  NANDN U1217 ( .A(n577), .B(a[5]), .Z(n637) );
  XOR U1218 ( .A(n17151), .B(n637), .Z(n639) );
  NANDN U1219 ( .A(b[0]), .B(a[4]), .Z(n638) );
  AND U1220 ( .A(n639), .B(n638), .Z(n665) );
  XOR U1221 ( .A(b[5]), .B(a[1]), .Z(n673) );
  AND U1222 ( .A(n17310), .B(n673), .Z(n644) );
  XNOR U1223 ( .A(b[5]), .B(n2921), .Z(n642) );
  XOR U1224 ( .A(b[5]), .B(b[4]), .Z(n641) );
  XNOR U1225 ( .A(b[5]), .B(n578), .Z(n640) );
  AND U1226 ( .A(n641), .B(n640), .Z(n17311) );
  NAND U1227 ( .A(n642), .B(n17311), .Z(n643) );
  NANDN U1228 ( .A(n644), .B(n643), .Z(n666) );
  XNOR U1229 ( .A(n665), .B(n666), .Z(n679) );
  NANDN U1230 ( .A(n578), .B(b[4]), .Z(n17442) );
  AND U1231 ( .A(n17442), .B(b[5]), .Z(n17733) );
  NAND U1232 ( .A(n17733), .B(n650), .Z(n676) );
  XNOR U1233 ( .A(b[3]), .B(a[3]), .Z(n667) );
  NANDN U1234 ( .A(n667), .B(n16990), .Z(n647) );
  OR U1235 ( .A(n645), .B(n16988), .Z(n646) );
  NAND U1236 ( .A(n647), .B(n646), .Z(n677) );
  XNOR U1237 ( .A(n676), .B(n677), .Z(n678) );
  XOR U1238 ( .A(n679), .B(n678), .Z(n660) );
  NANDN U1239 ( .A(n649), .B(n648), .Z(n653) );
  OR U1240 ( .A(n651), .B(n650), .Z(n652) );
  AND U1241 ( .A(n653), .B(n652), .Z(n659) );
  XOR U1242 ( .A(n660), .B(n659), .Z(n662) );
  XOR U1243 ( .A(n661), .B(n662), .Z(n682) );
  XNOR U1244 ( .A(sreg[101]), .B(n682), .Z(n684) );
  NAND U1245 ( .A(n654), .B(sreg[100]), .Z(n658) );
  NANDN U1246 ( .A(n656), .B(n655), .Z(n657) );
  AND U1247 ( .A(n658), .B(n657), .Z(n683) );
  XOR U1248 ( .A(n684), .B(n683), .Z(c[101]) );
  OR U1249 ( .A(n660), .B(n659), .Z(n664) );
  NAND U1250 ( .A(n662), .B(n661), .Z(n663) );
  NAND U1251 ( .A(n664), .B(n663), .Z(n690) );
  AND U1252 ( .A(n666), .B(n665), .Z(n716) );
  OR U1253 ( .A(n667), .B(n16988), .Z(n669) );
  XNOR U1254 ( .A(b[3]), .B(a[4]), .Z(n710) );
  NANDN U1255 ( .A(n710), .B(n16990), .Z(n668) );
  NAND U1256 ( .A(n669), .B(n668), .Z(n696) );
  XOR U1257 ( .A(b[5]), .B(b[6]), .Z(n17555) );
  NANDN U1258 ( .A(n2921), .B(n17555), .Z(n694) );
  NANDN U1259 ( .A(n577), .B(a[6]), .Z(n670) );
  XOR U1260 ( .A(n17151), .B(n670), .Z(n672) );
  NANDN U1261 ( .A(b[0]), .B(a[5]), .Z(n671) );
  AND U1262 ( .A(n672), .B(n671), .Z(n693) );
  XNOR U1263 ( .A(n694), .B(n693), .Z(n695) );
  XNOR U1264 ( .A(n696), .B(n695), .Z(n713) );
  XOR U1265 ( .A(b[5]), .B(a[2]), .Z(n697) );
  NAND U1266 ( .A(n17310), .B(n697), .Z(n675) );
  NAND U1267 ( .A(n17311), .B(n673), .Z(n674) );
  NAND U1268 ( .A(n675), .B(n674), .Z(n714) );
  XNOR U1269 ( .A(n713), .B(n714), .Z(n715) );
  XOR U1270 ( .A(n716), .B(n715), .Z(n687) );
  NANDN U1271 ( .A(n677), .B(n676), .Z(n681) );
  NAND U1272 ( .A(n679), .B(n678), .Z(n680) );
  NAND U1273 ( .A(n681), .B(n680), .Z(n688) );
  XNOR U1274 ( .A(n687), .B(n688), .Z(n689) );
  XNOR U1275 ( .A(n690), .B(n689), .Z(n721) );
  NAND U1276 ( .A(sreg[101]), .B(n682), .Z(n686) );
  OR U1277 ( .A(n684), .B(n683), .Z(n685) );
  NAND U1278 ( .A(n686), .B(n685), .Z(n719) );
  XNOR U1279 ( .A(n719), .B(sreg[102]), .Z(n720) );
  XOR U1280 ( .A(n721), .B(n720), .Z(c[102]) );
  NANDN U1281 ( .A(n688), .B(n687), .Z(n692) );
  NAND U1282 ( .A(n690), .B(n689), .Z(n691) );
  NAND U1283 ( .A(n692), .B(n691), .Z(n732) );
  XOR U1284 ( .A(b[5]), .B(a[3]), .Z(n758) );
  NAND U1285 ( .A(n758), .B(n17310), .Z(n699) );
  NAND U1286 ( .A(n697), .B(n17311), .Z(n698) );
  NAND U1287 ( .A(n699), .B(n698), .Z(n754) );
  XOR U1288 ( .A(b[7]), .B(a[1]), .Z(n747) );
  AND U1289 ( .A(n17555), .B(n747), .Z(n704) );
  XNOR U1290 ( .A(b[7]), .B(n2921), .Z(n702) );
  XOR U1291 ( .A(b[7]), .B(b[5]), .Z(n701) );
  XOR U1292 ( .A(b[7]), .B(b[6]), .Z(n700) );
  AND U1293 ( .A(n701), .B(n700), .Z(n17553) );
  NAND U1294 ( .A(n702), .B(n17553), .Z(n703) );
  NANDN U1295 ( .A(n704), .B(n703), .Z(n753) );
  XNOR U1296 ( .A(n754), .B(n753), .Z(n744) );
  OR U1297 ( .A(b[5]), .B(b[6]), .Z(n705) );
  NANDN U1298 ( .A(n2921), .B(n705), .Z(n706) );
  NAND U1299 ( .A(b[6]), .B(b[5]), .Z(n17711) );
  AND U1300 ( .A(n17711), .B(b[7]), .Z(n17972) );
  NAND U1301 ( .A(n706), .B(n17972), .Z(n741) );
  NANDN U1302 ( .A(n577), .B(a[7]), .Z(n707) );
  XOR U1303 ( .A(n17151), .B(n707), .Z(n709) );
  NANDN U1304 ( .A(b[0]), .B(a[6]), .Z(n708) );
  AND U1305 ( .A(n709), .B(n708), .Z(n742) );
  XNOR U1306 ( .A(n741), .B(n742), .Z(n743) );
  XOR U1307 ( .A(n744), .B(n743), .Z(n735) );
  XNOR U1308 ( .A(b[3]), .B(a[5]), .Z(n750) );
  NANDN U1309 ( .A(n750), .B(n16990), .Z(n712) );
  OR U1310 ( .A(n710), .B(n16988), .Z(n711) );
  AND U1311 ( .A(n712), .B(n711), .Z(n736) );
  XNOR U1312 ( .A(n735), .B(n736), .Z(n737) );
  XNOR U1313 ( .A(n738), .B(n737), .Z(n729) );
  NANDN U1314 ( .A(n714), .B(n713), .Z(n718) );
  NANDN U1315 ( .A(n716), .B(n715), .Z(n717) );
  NAND U1316 ( .A(n718), .B(n717), .Z(n730) );
  XNOR U1317 ( .A(n729), .B(n730), .Z(n731) );
  XOR U1318 ( .A(n732), .B(n731), .Z(n724) );
  XNOR U1319 ( .A(sreg[103]), .B(n724), .Z(n726) );
  NAND U1320 ( .A(n719), .B(sreg[102]), .Z(n723) );
  OR U1321 ( .A(n721), .B(n720), .Z(n722) );
  AND U1322 ( .A(n723), .B(n722), .Z(n725) );
  XOR U1323 ( .A(n726), .B(n725), .Z(c[103]) );
  NAND U1324 ( .A(sreg[103]), .B(n724), .Z(n728) );
  OR U1325 ( .A(n726), .B(n725), .Z(n727) );
  NAND U1326 ( .A(n728), .B(n727), .Z(n803) );
  XNOR U1327 ( .A(n803), .B(sreg[104]), .Z(n805) );
  NANDN U1328 ( .A(n730), .B(n729), .Z(n734) );
  NAND U1329 ( .A(n732), .B(n731), .Z(n733) );
  NAND U1330 ( .A(n734), .B(n733), .Z(n764) );
  NAND U1331 ( .A(n736), .B(n735), .Z(n740) );
  OR U1332 ( .A(n738), .B(n737), .Z(n739) );
  NAND U1333 ( .A(n740), .B(n739), .Z(n761) );
  NANDN U1334 ( .A(n742), .B(n741), .Z(n746) );
  NAND U1335 ( .A(n744), .B(n743), .Z(n745) );
  NAND U1336 ( .A(n746), .B(n745), .Z(n800) );
  NAND U1337 ( .A(n747), .B(n17553), .Z(n749) );
  XOR U1338 ( .A(b[7]), .B(a[2]), .Z(n773) );
  NAND U1339 ( .A(n773), .B(n17555), .Z(n748) );
  NAND U1340 ( .A(n749), .B(n748), .Z(n767) );
  OR U1341 ( .A(n750), .B(n16988), .Z(n752) );
  XNOR U1342 ( .A(b[3]), .B(a[6]), .Z(n785) );
  NANDN U1343 ( .A(n785), .B(n16990), .Z(n751) );
  AND U1344 ( .A(n752), .B(n751), .Z(n768) );
  XNOR U1345 ( .A(n767), .B(n768), .Z(n769) );
  NAND U1346 ( .A(n754), .B(n753), .Z(n770) );
  XOR U1347 ( .A(n769), .B(n770), .Z(n797) );
  XOR U1348 ( .A(b[8]), .B(b[7]), .Z(n17814) );
  NAND U1349 ( .A(a[0]), .B(n17814), .Z(n794) );
  NANDN U1350 ( .A(n577), .B(a[8]), .Z(n755) );
  XOR U1351 ( .A(n17151), .B(n755), .Z(n757) );
  NANDN U1352 ( .A(b[0]), .B(a[7]), .Z(n756) );
  AND U1353 ( .A(n757), .B(n756), .Z(n792) );
  XOR U1354 ( .A(b[5]), .B(a[4]), .Z(n782) );
  NAND U1355 ( .A(n17310), .B(n782), .Z(n760) );
  NAND U1356 ( .A(n17311), .B(n758), .Z(n759) );
  AND U1357 ( .A(n760), .B(n759), .Z(n791) );
  XNOR U1358 ( .A(n792), .B(n791), .Z(n793) );
  XNOR U1359 ( .A(n794), .B(n793), .Z(n798) );
  XNOR U1360 ( .A(n797), .B(n798), .Z(n799) );
  XNOR U1361 ( .A(n800), .B(n799), .Z(n762) );
  XNOR U1362 ( .A(n761), .B(n762), .Z(n763) );
  XNOR U1363 ( .A(n764), .B(n763), .Z(n804) );
  XOR U1364 ( .A(n805), .B(n804), .Z(c[104]) );
  NANDN U1365 ( .A(n762), .B(n761), .Z(n766) );
  NANDN U1366 ( .A(n764), .B(n763), .Z(n765) );
  NAND U1367 ( .A(n766), .B(n765), .Z(n816) );
  NANDN U1368 ( .A(n768), .B(n767), .Z(n772) );
  NANDN U1369 ( .A(n770), .B(n769), .Z(n771) );
  NAND U1370 ( .A(n772), .B(n771), .Z(n820) );
  NAND U1371 ( .A(n773), .B(n17553), .Z(n775) );
  XOR U1372 ( .A(b[7]), .B(a[3]), .Z(n843) );
  NAND U1373 ( .A(n843), .B(n17555), .Z(n774) );
  NAND U1374 ( .A(n775), .B(n774), .Z(n835) );
  XNOR U1375 ( .A(n579), .B(a[0]), .Z(n778) );
  XNOR U1376 ( .A(n579), .B(b[7]), .Z(n777) );
  XNOR U1377 ( .A(n579), .B(b[8]), .Z(n776) );
  AND U1378 ( .A(n777), .B(n776), .Z(n17815) );
  NAND U1379 ( .A(n778), .B(n17815), .Z(n780) );
  XNOR U1380 ( .A(b[9]), .B(a[1]), .Z(n832) );
  ANDN U1381 ( .B(n17814), .A(n832), .Z(n779) );
  ANDN U1382 ( .B(n780), .A(n779), .Z(n836) );
  XOR U1383 ( .A(n835), .B(n836), .Z(n825) );
  NAND U1384 ( .A(b[8]), .B(b[7]), .Z(n17963) );
  ANDN U1385 ( .B(n17963), .A(n579), .Z(n18149) );
  NANDN U1386 ( .A(n2921), .B(n17814), .Z(n781) );
  AND U1387 ( .A(n18149), .B(n781), .Z(n823) );
  XOR U1388 ( .A(b[5]), .B(a[5]), .Z(n829) );
  NAND U1389 ( .A(n829), .B(n17310), .Z(n784) );
  NAND U1390 ( .A(n782), .B(n17311), .Z(n783) );
  NAND U1391 ( .A(n784), .B(n783), .Z(n824) );
  XNOR U1392 ( .A(n823), .B(n824), .Z(n826) );
  XNOR U1393 ( .A(n825), .B(n826), .Z(n849) );
  OR U1394 ( .A(n785), .B(n16988), .Z(n787) );
  XNOR U1395 ( .A(b[3]), .B(a[7]), .Z(n837) );
  NANDN U1396 ( .A(n837), .B(n16990), .Z(n786) );
  AND U1397 ( .A(n787), .B(n786), .Z(n847) );
  NANDN U1398 ( .A(n577), .B(a[9]), .Z(n788) );
  XOR U1399 ( .A(n17151), .B(n788), .Z(n790) );
  NANDN U1400 ( .A(b[0]), .B(a[8]), .Z(n789) );
  AND U1401 ( .A(n790), .B(n789), .Z(n846) );
  XNOR U1402 ( .A(n847), .B(n846), .Z(n848) );
  XNOR U1403 ( .A(n849), .B(n848), .Z(n817) );
  NANDN U1404 ( .A(n792), .B(n791), .Z(n796) );
  NAND U1405 ( .A(n794), .B(n793), .Z(n795) );
  AND U1406 ( .A(n796), .B(n795), .Z(n818) );
  XOR U1407 ( .A(n817), .B(n818), .Z(n819) );
  XNOR U1408 ( .A(n820), .B(n819), .Z(n813) );
  NANDN U1409 ( .A(n798), .B(n797), .Z(n802) );
  NAND U1410 ( .A(n800), .B(n799), .Z(n801) );
  AND U1411 ( .A(n802), .B(n801), .Z(n814) );
  XNOR U1412 ( .A(n813), .B(n814), .Z(n815) );
  XNOR U1413 ( .A(n816), .B(n815), .Z(n808) );
  XNOR U1414 ( .A(n808), .B(sreg[105]), .Z(n810) );
  NAND U1415 ( .A(n803), .B(sreg[104]), .Z(n807) );
  OR U1416 ( .A(n805), .B(n804), .Z(n806) );
  AND U1417 ( .A(n807), .B(n806), .Z(n809) );
  XOR U1418 ( .A(n810), .B(n809), .Z(c[105]) );
  NAND U1419 ( .A(n808), .B(sreg[105]), .Z(n812) );
  OR U1420 ( .A(n810), .B(n809), .Z(n811) );
  NAND U1421 ( .A(n812), .B(n811), .Z(n900) );
  XNOR U1422 ( .A(n900), .B(sreg[106]), .Z(n902) );
  NAND U1423 ( .A(n818), .B(n817), .Z(n822) );
  NAND U1424 ( .A(n820), .B(n819), .Z(n821) );
  NAND U1425 ( .A(n822), .B(n821), .Z(n851) );
  OR U1426 ( .A(n824), .B(n823), .Z(n828) );
  NANDN U1427 ( .A(n826), .B(n825), .Z(n827) );
  NAND U1428 ( .A(n828), .B(n827), .Z(n858) );
  XOR U1429 ( .A(b[5]), .B(a[6]), .Z(n897) );
  NAND U1430 ( .A(n897), .B(n17310), .Z(n831) );
  NAND U1431 ( .A(n829), .B(n17311), .Z(n830) );
  NAND U1432 ( .A(n831), .B(n830), .Z(n874) );
  XNOR U1433 ( .A(b[9]), .B(a[2]), .Z(n886) );
  NANDN U1434 ( .A(n886), .B(n17814), .Z(n834) );
  NANDN U1435 ( .A(n832), .B(n17815), .Z(n833) );
  AND U1436 ( .A(n834), .B(n833), .Z(n875) );
  XNOR U1437 ( .A(n874), .B(n875), .Z(n876) );
  NANDN U1438 ( .A(n836), .B(n835), .Z(n877) );
  XOR U1439 ( .A(n876), .B(n877), .Z(n862) );
  XNOR U1440 ( .A(b[3]), .B(a[8]), .Z(n883) );
  NANDN U1441 ( .A(n883), .B(n16990), .Z(n839) );
  OR U1442 ( .A(n837), .B(n16988), .Z(n838) );
  NAND U1443 ( .A(n839), .B(n838), .Z(n863) );
  XNOR U1444 ( .A(n862), .B(n863), .Z(n864) );
  XOR U1445 ( .A(n579), .B(b[10]), .Z(n18194) );
  NOR U1446 ( .A(n2921), .B(n18194), .Z(n871) );
  NANDN U1447 ( .A(n577), .B(a[10]), .Z(n840) );
  XOR U1448 ( .A(n17151), .B(n840), .Z(n842) );
  NANDN U1449 ( .A(b[0]), .B(a[9]), .Z(n841) );
  AND U1450 ( .A(n842), .B(n841), .Z(n869) );
  XNOR U1451 ( .A(b[7]), .B(a[4]), .Z(n880) );
  NANDN U1452 ( .A(n880), .B(n17555), .Z(n845) );
  NAND U1453 ( .A(n843), .B(n17553), .Z(n844) );
  AND U1454 ( .A(n845), .B(n844), .Z(n868) );
  XNOR U1455 ( .A(n869), .B(n868), .Z(n870) );
  XOR U1456 ( .A(n871), .B(n870), .Z(n865) );
  XNOR U1457 ( .A(n864), .B(n865), .Z(n856) );
  XNOR U1458 ( .A(n856), .B(n857), .Z(n859) );
  XNOR U1459 ( .A(n858), .B(n859), .Z(n850) );
  XNOR U1460 ( .A(n851), .B(n850), .Z(n852) );
  XOR U1461 ( .A(n853), .B(n852), .Z(n901) );
  XOR U1462 ( .A(n902), .B(n901), .Z(c[106]) );
  NANDN U1463 ( .A(n851), .B(n850), .Z(n855) );
  NAND U1464 ( .A(n853), .B(n852), .Z(n854) );
  NAND U1465 ( .A(n855), .B(n854), .Z(n913) );
  NAND U1466 ( .A(n857), .B(n856), .Z(n861) );
  NANDN U1467 ( .A(n859), .B(n858), .Z(n860) );
  NAND U1468 ( .A(n861), .B(n860), .Z(n910) );
  NANDN U1469 ( .A(n863), .B(n862), .Z(n867) );
  NANDN U1470 ( .A(n865), .B(n864), .Z(n866) );
  NAND U1471 ( .A(n867), .B(n866), .Z(n919) );
  NANDN U1472 ( .A(n869), .B(n868), .Z(n873) );
  NANDN U1473 ( .A(n871), .B(n870), .Z(n872) );
  NAND U1474 ( .A(n873), .B(n872), .Z(n916) );
  NANDN U1475 ( .A(n875), .B(n874), .Z(n879) );
  NANDN U1476 ( .A(n877), .B(n876), .Z(n878) );
  NAND U1477 ( .A(n879), .B(n878), .Z(n957) );
  XNOR U1478 ( .A(b[7]), .B(a[5]), .Z(n936) );
  NANDN U1479 ( .A(n936), .B(n17555), .Z(n882) );
  NANDN U1480 ( .A(n880), .B(n17553), .Z(n881) );
  NAND U1481 ( .A(n882), .B(n881), .Z(n925) );
  XNOR U1482 ( .A(b[3]), .B(a[9]), .Z(n939) );
  NANDN U1483 ( .A(n939), .B(n16990), .Z(n885) );
  OR U1484 ( .A(n883), .B(n16988), .Z(n884) );
  NAND U1485 ( .A(n885), .B(n884), .Z(n923) );
  XOR U1486 ( .A(n922), .B(n923), .Z(n924) );
  XNOR U1487 ( .A(n925), .B(n924), .Z(n955) );
  XNOR U1488 ( .A(n579), .B(a[3]), .Z(n945) );
  NAND U1489 ( .A(n17814), .B(n945), .Z(n888) );
  NANDN U1490 ( .A(n886), .B(n17815), .Z(n887) );
  NAND U1491 ( .A(n888), .B(n887), .Z(n935) );
  XNOR U1492 ( .A(b[11]), .B(n2921), .Z(n891) );
  XNOR U1493 ( .A(b[11]), .B(n579), .Z(n890) );
  XOR U1494 ( .A(b[11]), .B(b[10]), .Z(n889) );
  AND U1495 ( .A(n890), .B(n889), .Z(n18104) );
  NAND U1496 ( .A(n891), .B(n18104), .Z(n893) );
  XNOR U1497 ( .A(b[11]), .B(a[1]), .Z(n931) );
  OR U1498 ( .A(n931), .B(n18194), .Z(n892) );
  NAND U1499 ( .A(n893), .B(n892), .Z(n934) );
  XNOR U1500 ( .A(n935), .B(n934), .Z(n951) );
  NANDN U1501 ( .A(n577), .B(a[11]), .Z(n894) );
  XOR U1502 ( .A(n17151), .B(n894), .Z(n896) );
  NANDN U1503 ( .A(b[0]), .B(a[10]), .Z(n895) );
  AND U1504 ( .A(n896), .B(n895), .Z(n949) );
  XNOR U1505 ( .A(b[5]), .B(a[7]), .Z(n928) );
  NANDN U1506 ( .A(n928), .B(n17310), .Z(n899) );
  NAND U1507 ( .A(n17311), .B(n897), .Z(n898) );
  AND U1508 ( .A(n899), .B(n898), .Z(n948) );
  XNOR U1509 ( .A(n949), .B(n948), .Z(n950) );
  XOR U1510 ( .A(n951), .B(n950), .Z(n954) );
  XOR U1511 ( .A(n955), .B(n954), .Z(n956) );
  XOR U1512 ( .A(n957), .B(n956), .Z(n917) );
  XNOR U1513 ( .A(n916), .B(n917), .Z(n918) );
  XNOR U1514 ( .A(n919), .B(n918), .Z(n911) );
  XNOR U1515 ( .A(n910), .B(n911), .Z(n912) );
  XNOR U1516 ( .A(n913), .B(n912), .Z(n905) );
  XNOR U1517 ( .A(n905), .B(sreg[107]), .Z(n907) );
  NAND U1518 ( .A(n900), .B(sreg[106]), .Z(n904) );
  OR U1519 ( .A(n902), .B(n901), .Z(n903) );
  AND U1520 ( .A(n904), .B(n903), .Z(n906) );
  XOR U1521 ( .A(n907), .B(n906), .Z(c[107]) );
  NAND U1522 ( .A(n905), .B(sreg[107]), .Z(n909) );
  OR U1523 ( .A(n907), .B(n906), .Z(n908) );
  NAND U1524 ( .A(n909), .B(n908), .Z(n1019) );
  XNOR U1525 ( .A(n1019), .B(sreg[108]), .Z(n1021) );
  NANDN U1526 ( .A(n911), .B(n910), .Z(n915) );
  NAND U1527 ( .A(n913), .B(n912), .Z(n914) );
  NAND U1528 ( .A(n915), .B(n914), .Z(n963) );
  NANDN U1529 ( .A(n917), .B(n916), .Z(n921) );
  NAND U1530 ( .A(n919), .B(n918), .Z(n920) );
  NAND U1531 ( .A(n921), .B(n920), .Z(n960) );
  OR U1532 ( .A(n923), .B(n922), .Z(n927) );
  NANDN U1533 ( .A(n925), .B(n924), .Z(n926) );
  NAND U1534 ( .A(n927), .B(n926), .Z(n969) );
  XOR U1535 ( .A(b[5]), .B(a[8]), .Z(n998) );
  NAND U1536 ( .A(n17310), .B(n998), .Z(n930) );
  NANDN U1537 ( .A(n928), .B(n17311), .Z(n929) );
  NAND U1538 ( .A(n930), .B(n929), .Z(n979) );
  XOR U1539 ( .A(b[11]), .B(a[2]), .Z(n984) );
  NANDN U1540 ( .A(n18194), .B(n984), .Z(n933) );
  NANDN U1541 ( .A(n931), .B(n18104), .Z(n932) );
  AND U1542 ( .A(n933), .B(n932), .Z(n978) );
  XNOR U1543 ( .A(n979), .B(n978), .Z(n980) );
  NAND U1544 ( .A(n935), .B(n934), .Z(n1010) );
  XNOR U1545 ( .A(b[7]), .B(a[6]), .Z(n995) );
  NANDN U1546 ( .A(n995), .B(n17555), .Z(n938) );
  NANDN U1547 ( .A(n936), .B(n17553), .Z(n937) );
  NAND U1548 ( .A(n938), .B(n937), .Z(n1008) );
  XNOR U1549 ( .A(b[3]), .B(a[10]), .Z(n1001) );
  NANDN U1550 ( .A(n1001), .B(n16990), .Z(n941) );
  OR U1551 ( .A(n939), .B(n16988), .Z(n940) );
  AND U1552 ( .A(n941), .B(n940), .Z(n1007) );
  XNOR U1553 ( .A(n1008), .B(n1007), .Z(n1009) );
  XNOR U1554 ( .A(n1010), .B(n1009), .Z(n981) );
  XOR U1555 ( .A(n980), .B(n981), .Z(n975) );
  NANDN U1556 ( .A(n577), .B(a[12]), .Z(n942) );
  XOR U1557 ( .A(n17151), .B(n942), .Z(n944) );
  IV U1558 ( .A(a[11]), .Z(n4573) );
  NANDN U1559 ( .A(n4573), .B(n577), .Z(n943) );
  AND U1560 ( .A(n944), .B(n943), .Z(n1013) );
  XNOR U1561 ( .A(b[9]), .B(a[4]), .Z(n1004) );
  NANDN U1562 ( .A(n1004), .B(n17814), .Z(n947) );
  NAND U1563 ( .A(n945), .B(n17815), .Z(n946) );
  AND U1564 ( .A(n947), .B(n946), .Z(n1014) );
  XOR U1565 ( .A(n1013), .B(n1014), .Z(n1016) );
  XOR U1566 ( .A(b[11]), .B(b[12]), .Z(n18336) );
  NANDN U1567 ( .A(n2921), .B(n18336), .Z(n1015) );
  XOR U1568 ( .A(n1016), .B(n1015), .Z(n972) );
  NANDN U1569 ( .A(n949), .B(n948), .Z(n953) );
  NAND U1570 ( .A(n951), .B(n950), .Z(n952) );
  AND U1571 ( .A(n953), .B(n952), .Z(n973) );
  XOR U1572 ( .A(n972), .B(n973), .Z(n974) );
  XNOR U1573 ( .A(n975), .B(n974), .Z(n966) );
  OR U1574 ( .A(n955), .B(n954), .Z(n959) );
  NAND U1575 ( .A(n957), .B(n956), .Z(n958) );
  NAND U1576 ( .A(n959), .B(n958), .Z(n967) );
  XNOR U1577 ( .A(n966), .B(n967), .Z(n968) );
  XNOR U1578 ( .A(n969), .B(n968), .Z(n961) );
  XNOR U1579 ( .A(n960), .B(n961), .Z(n962) );
  XOR U1580 ( .A(n963), .B(n962), .Z(n1020) );
  XOR U1581 ( .A(n1021), .B(n1020), .Z(c[108]) );
  NANDN U1582 ( .A(n961), .B(n960), .Z(n965) );
  NAND U1583 ( .A(n963), .B(n962), .Z(n964) );
  NAND U1584 ( .A(n965), .B(n964), .Z(n1032) );
  NANDN U1585 ( .A(n967), .B(n966), .Z(n971) );
  NAND U1586 ( .A(n969), .B(n968), .Z(n970) );
  NAND U1587 ( .A(n971), .B(n970), .Z(n1030) );
  NAND U1588 ( .A(n973), .B(n972), .Z(n977) );
  NAND U1589 ( .A(n975), .B(n974), .Z(n976) );
  NAND U1590 ( .A(n977), .B(n976), .Z(n1037) );
  NANDN U1591 ( .A(n979), .B(n978), .Z(n983) );
  NANDN U1592 ( .A(n981), .B(n980), .Z(n982) );
  NAND U1593 ( .A(n983), .B(n982), .Z(n1036) );
  XOR U1594 ( .A(b[11]), .B(a[3]), .Z(n1062) );
  NANDN U1595 ( .A(n18194), .B(n1062), .Z(n986) );
  NAND U1596 ( .A(n984), .B(n18104), .Z(n985) );
  NAND U1597 ( .A(n986), .B(n985), .Z(n1051) );
  XNOR U1598 ( .A(n580), .B(a[0]), .Z(n989) );
  XNOR U1599 ( .A(n580), .B(b[11]), .Z(n988) );
  XNOR U1600 ( .A(n580), .B(b[12]), .Z(n987) );
  AND U1601 ( .A(n988), .B(n987), .Z(n18337) );
  NAND U1602 ( .A(n989), .B(n18337), .Z(n991) );
  XNOR U1603 ( .A(n580), .B(a[1]), .Z(n1045) );
  NAND U1604 ( .A(n1045), .B(n18336), .Z(n990) );
  NAND U1605 ( .A(n991), .B(n990), .Z(n1052) );
  XNOR U1606 ( .A(n1051), .B(n1052), .Z(n1077) );
  NANDN U1607 ( .A(n577), .B(a[13]), .Z(n992) );
  XOR U1608 ( .A(n17151), .B(n992), .Z(n994) );
  NANDN U1609 ( .A(b[0]), .B(a[12]), .Z(n993) );
  AND U1610 ( .A(n994), .B(n993), .Z(n1075) );
  XNOR U1611 ( .A(b[7]), .B(a[7]), .Z(n1068) );
  NANDN U1612 ( .A(n1068), .B(n17555), .Z(n997) );
  NANDN U1613 ( .A(n995), .B(n17553), .Z(n996) );
  AND U1614 ( .A(n997), .B(n996), .Z(n1074) );
  XNOR U1615 ( .A(n1075), .B(n1074), .Z(n1076) );
  XOR U1616 ( .A(n1077), .B(n1076), .Z(n1082) );
  XOR U1617 ( .A(b[5]), .B(a[9]), .Z(n1065) );
  NAND U1618 ( .A(n1065), .B(n17310), .Z(n1000) );
  NAND U1619 ( .A(n998), .B(n17311), .Z(n999) );
  NAND U1620 ( .A(n1000), .B(n999), .Z(n1081) );
  OR U1621 ( .A(n1001), .B(n16988), .Z(n1003) );
  XOR U1622 ( .A(b[3]), .B(n4573), .Z(n1071) );
  NANDN U1623 ( .A(n1071), .B(n16990), .Z(n1002) );
  NAND U1624 ( .A(n1003), .B(n1002), .Z(n1053) );
  XNOR U1625 ( .A(b[9]), .B(a[5]), .Z(n1048) );
  NANDN U1626 ( .A(n1048), .B(n17814), .Z(n1006) );
  NANDN U1627 ( .A(n1004), .B(n17815), .Z(n1005) );
  AND U1628 ( .A(n1006), .B(n1005), .Z(n1054) );
  XNOR U1629 ( .A(n1053), .B(n1054), .Z(n1055) );
  XNOR U1630 ( .A(n1056), .B(n1055), .Z(n1080) );
  XNOR U1631 ( .A(n1081), .B(n1080), .Z(n1083) );
  XOR U1632 ( .A(n1082), .B(n1083), .Z(n1042) );
  NANDN U1633 ( .A(n1008), .B(n1007), .Z(n1012) );
  NAND U1634 ( .A(n1010), .B(n1009), .Z(n1011) );
  NAND U1635 ( .A(n1012), .B(n1011), .Z(n1039) );
  NANDN U1636 ( .A(n1014), .B(n1013), .Z(n1018) );
  OR U1637 ( .A(n1016), .B(n1015), .Z(n1017) );
  NAND U1638 ( .A(n1018), .B(n1017), .Z(n1040) );
  XNOR U1639 ( .A(n1039), .B(n1040), .Z(n1041) );
  XNOR U1640 ( .A(n1042), .B(n1041), .Z(n1035) );
  XNOR U1641 ( .A(n1036), .B(n1035), .Z(n1038) );
  XOR U1642 ( .A(n1037), .B(n1038), .Z(n1029) );
  XOR U1643 ( .A(n1030), .B(n1029), .Z(n1031) );
  XNOR U1644 ( .A(n1032), .B(n1031), .Z(n1024) );
  XNOR U1645 ( .A(n1024), .B(sreg[109]), .Z(n1026) );
  NAND U1646 ( .A(n1019), .B(sreg[108]), .Z(n1023) );
  OR U1647 ( .A(n1021), .B(n1020), .Z(n1022) );
  AND U1648 ( .A(n1023), .B(n1022), .Z(n1025) );
  XOR U1649 ( .A(n1026), .B(n1025), .Z(c[109]) );
  NAND U1650 ( .A(n1024), .B(sreg[109]), .Z(n1028) );
  OR U1651 ( .A(n1026), .B(n1025), .Z(n1027) );
  NAND U1652 ( .A(n1028), .B(n1027), .Z(n1150) );
  XNOR U1653 ( .A(n1150), .B(sreg[110]), .Z(n1152) );
  NAND U1654 ( .A(n1030), .B(n1029), .Z(n1034) );
  NAND U1655 ( .A(n1032), .B(n1031), .Z(n1033) );
  NAND U1656 ( .A(n1034), .B(n1033), .Z(n1087) );
  NANDN U1657 ( .A(n1040), .B(n1039), .Z(n1044) );
  NANDN U1658 ( .A(n1042), .B(n1041), .Z(n1043) );
  NAND U1659 ( .A(n1044), .B(n1043), .Z(n1092) );
  XNOR U1660 ( .A(b[13]), .B(a[2]), .Z(n1106) );
  NANDN U1661 ( .A(n1106), .B(n18336), .Z(n1047) );
  NAND U1662 ( .A(n1045), .B(n18337), .Z(n1046) );
  NAND U1663 ( .A(n1047), .B(n1046), .Z(n1144) );
  XNOR U1664 ( .A(b[9]), .B(a[6]), .Z(n1103) );
  NANDN U1665 ( .A(n1103), .B(n17814), .Z(n1050) );
  NANDN U1666 ( .A(n1048), .B(n17815), .Z(n1049) );
  AND U1667 ( .A(n1050), .B(n1049), .Z(n1145) );
  XNOR U1668 ( .A(n1144), .B(n1145), .Z(n1146) );
  NAND U1669 ( .A(n1052), .B(n1051), .Z(n1147) );
  XOR U1670 ( .A(n1146), .B(n1147), .Z(n1099) );
  NANDN U1671 ( .A(n1054), .B(n1053), .Z(n1058) );
  NANDN U1672 ( .A(n1056), .B(n1055), .Z(n1057) );
  NAND U1673 ( .A(n1058), .B(n1057), .Z(n1137) );
  XNOR U1674 ( .A(b[13]), .B(b[14]), .Z(n18512) );
  NOR U1675 ( .A(n2921), .B(n18512), .Z(n1141) );
  NANDN U1676 ( .A(n577), .B(a[14]), .Z(n1059) );
  XOR U1677 ( .A(n17151), .B(n1059), .Z(n1061) );
  IV U1678 ( .A(a[13]), .Z(n4875) );
  NANDN U1679 ( .A(n4875), .B(n577), .Z(n1060) );
  AND U1680 ( .A(n1061), .B(n1060), .Z(n1139) );
  XOR U1681 ( .A(b[11]), .B(a[4]), .Z(n1120) );
  NANDN U1682 ( .A(n18194), .B(n1120), .Z(n1064) );
  NAND U1683 ( .A(n18104), .B(n1062), .Z(n1063) );
  AND U1684 ( .A(n1064), .B(n1063), .Z(n1138) );
  XNOR U1685 ( .A(n1139), .B(n1138), .Z(n1140) );
  XOR U1686 ( .A(n1141), .B(n1140), .Z(n1134) );
  XOR U1687 ( .A(b[5]), .B(a[10]), .Z(n1123) );
  NAND U1688 ( .A(n1123), .B(n17310), .Z(n1067) );
  NAND U1689 ( .A(n1065), .B(n17311), .Z(n1066) );
  NAND U1690 ( .A(n1067), .B(n1066), .Z(n1117) );
  NANDN U1691 ( .A(n1068), .B(n17553), .Z(n1070) );
  XOR U1692 ( .A(b[7]), .B(a[8]), .Z(n1131) );
  NAND U1693 ( .A(n1131), .B(n17555), .Z(n1069) );
  NAND U1694 ( .A(n1070), .B(n1069), .Z(n1114) );
  OR U1695 ( .A(n1071), .B(n16988), .Z(n1073) );
  XNOR U1696 ( .A(b[3]), .B(a[12]), .Z(n1126) );
  NANDN U1697 ( .A(n1126), .B(n16990), .Z(n1072) );
  AND U1698 ( .A(n1073), .B(n1072), .Z(n1115) );
  XNOR U1699 ( .A(n1114), .B(n1115), .Z(n1116) );
  XNOR U1700 ( .A(n1117), .B(n1116), .Z(n1135) );
  XNOR U1701 ( .A(n1134), .B(n1135), .Z(n1136) );
  XNOR U1702 ( .A(n1137), .B(n1136), .Z(n1096) );
  NANDN U1703 ( .A(n1075), .B(n1074), .Z(n1079) );
  NAND U1704 ( .A(n1077), .B(n1076), .Z(n1078) );
  AND U1705 ( .A(n1079), .B(n1078), .Z(n1097) );
  XNOR U1706 ( .A(n1096), .B(n1097), .Z(n1098) );
  XNOR U1707 ( .A(n1099), .B(n1098), .Z(n1090) );
  XOR U1708 ( .A(n1090), .B(n1091), .Z(n1093) );
  XOR U1709 ( .A(n1092), .B(n1093), .Z(n1085) );
  XNOR U1710 ( .A(n1084), .B(n1085), .Z(n1086) );
  XOR U1711 ( .A(n1087), .B(n1086), .Z(n1151) );
  XOR U1712 ( .A(n1152), .B(n1151), .Z(c[110]) );
  NANDN U1713 ( .A(n1085), .B(n1084), .Z(n1089) );
  NAND U1714 ( .A(n1087), .B(n1086), .Z(n1088) );
  NAND U1715 ( .A(n1089), .B(n1088), .Z(n1163) );
  NANDN U1716 ( .A(n1091), .B(n1090), .Z(n1095) );
  OR U1717 ( .A(n1093), .B(n1092), .Z(n1094) );
  NAND U1718 ( .A(n1095), .B(n1094), .Z(n1161) );
  NANDN U1719 ( .A(n577), .B(a[15]), .Z(n1100) );
  XOR U1720 ( .A(n17151), .B(n1100), .Z(n1102) );
  NANDN U1721 ( .A(b[0]), .B(a[14]), .Z(n1101) );
  AND U1722 ( .A(n1102), .B(n1101), .Z(n1188) );
  XNOR U1723 ( .A(n579), .B(a[7]), .Z(n1194) );
  NAND U1724 ( .A(n17814), .B(n1194), .Z(n1105) );
  NANDN U1725 ( .A(n1103), .B(n17815), .Z(n1104) );
  AND U1726 ( .A(n1105), .B(n1104), .Z(n1189) );
  XNOR U1727 ( .A(n1188), .B(n1189), .Z(n1190) );
  XNOR U1728 ( .A(b[13]), .B(a[3]), .Z(n1185) );
  NANDN U1729 ( .A(n1185), .B(n18336), .Z(n1108) );
  NANDN U1730 ( .A(n1106), .B(n18337), .Z(n1107) );
  NAND U1731 ( .A(n1108), .B(n1107), .Z(n1192) );
  XNOR U1732 ( .A(b[15]), .B(n2921), .Z(n1111) );
  XNOR U1733 ( .A(b[15]), .B(n580), .Z(n1110) );
  XOR U1734 ( .A(b[15]), .B(b[14]), .Z(n1109) );
  AND U1735 ( .A(n1110), .B(n1109), .Z(n18513) );
  NAND U1736 ( .A(n1111), .B(n18513), .Z(n1113) );
  XOR U1737 ( .A(b[15]), .B(a[1]), .Z(n1206) );
  ANDN U1738 ( .B(n1206), .A(n18512), .Z(n1112) );
  ANDN U1739 ( .B(n1113), .A(n1112), .Z(n1193) );
  XNOR U1740 ( .A(n1192), .B(n1193), .Z(n1191) );
  XOR U1741 ( .A(n1190), .B(n1191), .Z(n1218) );
  NANDN U1742 ( .A(n1115), .B(n1114), .Z(n1119) );
  NAND U1743 ( .A(n1117), .B(n1116), .Z(n1118) );
  NAND U1744 ( .A(n1119), .B(n1118), .Z(n1219) );
  XOR U1745 ( .A(n1218), .B(n1219), .Z(n1220) );
  XOR U1746 ( .A(b[11]), .B(a[5]), .Z(n1203) );
  NANDN U1747 ( .A(n18194), .B(n1203), .Z(n1122) );
  NAND U1748 ( .A(n1120), .B(n18104), .Z(n1121) );
  NAND U1749 ( .A(n1122), .B(n1121), .Z(n1179) );
  XNOR U1750 ( .A(b[5]), .B(a[11]), .Z(n1209) );
  NANDN U1751 ( .A(n1209), .B(n17310), .Z(n1125) );
  NAND U1752 ( .A(n1123), .B(n17311), .Z(n1124) );
  NAND U1753 ( .A(n1125), .B(n1124), .Z(n1176) );
  OR U1754 ( .A(n1126), .B(n16988), .Z(n1128) );
  XOR U1755 ( .A(b[3]), .B(n4875), .Z(n1197) );
  NANDN U1756 ( .A(n1197), .B(n16990), .Z(n1127) );
  AND U1757 ( .A(n1128), .B(n1127), .Z(n1177) );
  XNOR U1758 ( .A(n1176), .B(n1177), .Z(n1178) );
  XNOR U1759 ( .A(n1179), .B(n1178), .Z(n1215) );
  NANDN U1760 ( .A(b[14]), .B(n580), .Z(n1129) );
  NANDN U1761 ( .A(n2921), .B(n1129), .Z(n1130) );
  NANDN U1762 ( .A(n580), .B(b[14]), .Z(n18577) );
  AND U1763 ( .A(n18577), .B(b[15]), .Z(n18768) );
  NAND U1764 ( .A(n1130), .B(n18768), .Z(n1212) );
  XNOR U1765 ( .A(b[7]), .B(a[9]), .Z(n1200) );
  NANDN U1766 ( .A(n1200), .B(n17555), .Z(n1133) );
  NAND U1767 ( .A(n1131), .B(n17553), .Z(n1132) );
  NAND U1768 ( .A(n1133), .B(n1132), .Z(n1213) );
  XNOR U1769 ( .A(n1212), .B(n1213), .Z(n1214) );
  XOR U1770 ( .A(n1215), .B(n1214), .Z(n1221) );
  XOR U1771 ( .A(n1220), .B(n1221), .Z(n1164) );
  XNOR U1772 ( .A(n1165), .B(n1164), .Z(n1166) );
  NANDN U1773 ( .A(n1139), .B(n1138), .Z(n1143) );
  NANDN U1774 ( .A(n1141), .B(n1140), .Z(n1142) );
  NAND U1775 ( .A(n1143), .B(n1142), .Z(n1170) );
  NANDN U1776 ( .A(n1145), .B(n1144), .Z(n1149) );
  NANDN U1777 ( .A(n1147), .B(n1146), .Z(n1148) );
  NAND U1778 ( .A(n1149), .B(n1148), .Z(n1171) );
  XNOR U1779 ( .A(n1170), .B(n1171), .Z(n1172) );
  XOR U1780 ( .A(n1173), .B(n1172), .Z(n1167) );
  XOR U1781 ( .A(n1166), .B(n1167), .Z(n1160) );
  XNOR U1782 ( .A(n1161), .B(n1160), .Z(n1162) );
  XNOR U1783 ( .A(n1163), .B(n1162), .Z(n1155) );
  XNOR U1784 ( .A(n1155), .B(sreg[111]), .Z(n1157) );
  NAND U1785 ( .A(n1150), .B(sreg[110]), .Z(n1154) );
  OR U1786 ( .A(n1152), .B(n1151), .Z(n1153) );
  AND U1787 ( .A(n1154), .B(n1153), .Z(n1156) );
  XOR U1788 ( .A(n1157), .B(n1156), .Z(c[111]) );
  NAND U1789 ( .A(n1155), .B(sreg[111]), .Z(n1159) );
  OR U1790 ( .A(n1157), .B(n1156), .Z(n1158) );
  NAND U1791 ( .A(n1159), .B(n1158), .Z(n1303) );
  XNOR U1792 ( .A(n1303), .B(sreg[112]), .Z(n1305) );
  NAND U1793 ( .A(n1165), .B(n1164), .Z(n1169) );
  OR U1794 ( .A(n1167), .B(n1166), .Z(n1168) );
  NAND U1795 ( .A(n1169), .B(n1168), .Z(n1224) );
  NANDN U1796 ( .A(n1171), .B(n1170), .Z(n1175) );
  NANDN U1797 ( .A(n1173), .B(n1172), .Z(n1174) );
  NAND U1798 ( .A(n1175), .B(n1174), .Z(n1300) );
  NANDN U1799 ( .A(n1177), .B(n1176), .Z(n1181) );
  NAND U1800 ( .A(n1179), .B(n1178), .Z(n1180) );
  NAND U1801 ( .A(n1181), .B(n1180), .Z(n1239) );
  NANDN U1802 ( .A(n577), .B(a[16]), .Z(n1182) );
  XOR U1803 ( .A(n17151), .B(n1182), .Z(n1184) );
  IV U1804 ( .A(a[15]), .Z(n5159) );
  NANDN U1805 ( .A(n5159), .B(n577), .Z(n1183) );
  AND U1806 ( .A(n1184), .B(n1183), .Z(n1269) );
  XNOR U1807 ( .A(b[13]), .B(a[4]), .Z(n1254) );
  NANDN U1808 ( .A(n1254), .B(n18336), .Z(n1187) );
  NANDN U1809 ( .A(n1185), .B(n18337), .Z(n1186) );
  NAND U1810 ( .A(n1187), .B(n1186), .Z(n1267) );
  XOR U1811 ( .A(b[15]), .B(b[16]), .Z(n18673) );
  NANDN U1812 ( .A(n2921), .B(n18673), .Z(n1268) );
  XNOR U1813 ( .A(n1267), .B(n1268), .Z(n1270) );
  XOR U1814 ( .A(n1269), .B(n1270), .Z(n1236) );
  XOR U1815 ( .A(n1236), .B(n1237), .Z(n1238) );
  XOR U1816 ( .A(n1239), .B(n1238), .Z(n1231) );
  NANDN U1817 ( .A(n1193), .B(n1192), .Z(n1244) );
  XOR U1818 ( .A(n579), .B(a[8]), .Z(n1285) );
  NANDN U1819 ( .A(n1285), .B(n17814), .Z(n1196) );
  NAND U1820 ( .A(n17815), .B(n1194), .Z(n1195) );
  NAND U1821 ( .A(n1196), .B(n1195), .Z(n1243) );
  XNOR U1822 ( .A(b[3]), .B(a[14]), .Z(n1291) );
  NANDN U1823 ( .A(n1291), .B(n16990), .Z(n1199) );
  OR U1824 ( .A(n1197), .B(n16988), .Z(n1198) );
  NAND U1825 ( .A(n1199), .B(n1198), .Z(n1242) );
  XNOR U1826 ( .A(n1243), .B(n1242), .Z(n1245) );
  XNOR U1827 ( .A(n1244), .B(n1245), .Z(n1263) );
  NANDN U1828 ( .A(n1200), .B(n17553), .Z(n1202) );
  XOR U1829 ( .A(b[7]), .B(a[10]), .Z(n1248) );
  NAND U1830 ( .A(n1248), .B(n17555), .Z(n1201) );
  NAND U1831 ( .A(n1202), .B(n1201), .Z(n1262) );
  XOR U1832 ( .A(b[11]), .B(a[6]), .Z(n1251) );
  NANDN U1833 ( .A(n18194), .B(n1251), .Z(n1205) );
  NAND U1834 ( .A(n18104), .B(n1203), .Z(n1204) );
  AND U1835 ( .A(n1205), .B(n1204), .Z(n1260) );
  XNOR U1836 ( .A(b[15]), .B(a[2]), .Z(n1273) );
  OR U1837 ( .A(n1273), .B(n18512), .Z(n1208) );
  NAND U1838 ( .A(n1206), .B(n18513), .Z(n1207) );
  NAND U1839 ( .A(n1208), .B(n1207), .Z(n1257) );
  XOR U1840 ( .A(b[5]), .B(a[12]), .Z(n1294) );
  NAND U1841 ( .A(n1294), .B(n17310), .Z(n1211) );
  NANDN U1842 ( .A(n1209), .B(n17311), .Z(n1210) );
  AND U1843 ( .A(n1211), .B(n1210), .Z(n1258) );
  XNOR U1844 ( .A(n1257), .B(n1258), .Z(n1259) );
  XNOR U1845 ( .A(n1260), .B(n1259), .Z(n1261) );
  XNOR U1846 ( .A(n1262), .B(n1261), .Z(n1264) );
  XOR U1847 ( .A(n1263), .B(n1264), .Z(n1230) );
  XNOR U1848 ( .A(n1231), .B(n1230), .Z(n1233) );
  NANDN U1849 ( .A(n1213), .B(n1212), .Z(n1217) );
  NAND U1850 ( .A(n1215), .B(n1214), .Z(n1216) );
  NAND U1851 ( .A(n1217), .B(n1216), .Z(n1232) );
  XNOR U1852 ( .A(n1233), .B(n1232), .Z(n1297) );
  OR U1853 ( .A(n1219), .B(n1218), .Z(n1223) );
  NAND U1854 ( .A(n1221), .B(n1220), .Z(n1222) );
  AND U1855 ( .A(n1223), .B(n1222), .Z(n1298) );
  XNOR U1856 ( .A(n1297), .B(n1298), .Z(n1299) );
  XNOR U1857 ( .A(n1300), .B(n1299), .Z(n1225) );
  XNOR U1858 ( .A(n1224), .B(n1225), .Z(n1226) );
  XOR U1859 ( .A(n1227), .B(n1226), .Z(n1304) );
  XOR U1860 ( .A(n1305), .B(n1304), .Z(c[112]) );
  NANDN U1861 ( .A(n1225), .B(n1224), .Z(n1229) );
  NAND U1862 ( .A(n1227), .B(n1226), .Z(n1228) );
  NAND U1863 ( .A(n1229), .B(n1228), .Z(n1316) );
  NAND U1864 ( .A(n1231), .B(n1230), .Z(n1235) );
  OR U1865 ( .A(n1233), .B(n1232), .Z(n1234) );
  NAND U1866 ( .A(n1235), .B(n1234), .Z(n1319) );
  OR U1867 ( .A(n1237), .B(n1236), .Z(n1241) );
  NANDN U1868 ( .A(n1239), .B(n1238), .Z(n1240) );
  NAND U1869 ( .A(n1241), .B(n1240), .Z(n1320) );
  XNOR U1870 ( .A(n1319), .B(n1320), .Z(n1321) );
  OR U1871 ( .A(n1243), .B(n1242), .Z(n1247) );
  NANDN U1872 ( .A(n1245), .B(n1244), .Z(n1246) );
  NAND U1873 ( .A(n1247), .B(n1246), .Z(n1325) );
  NAND U1874 ( .A(n1248), .B(n17553), .Z(n1250) );
  XNOR U1875 ( .A(b[7]), .B(a[11]), .Z(n1367) );
  NANDN U1876 ( .A(n1367), .B(n17555), .Z(n1249) );
  NAND U1877 ( .A(n1250), .B(n1249), .Z(n1373) );
  XOR U1878 ( .A(b[11]), .B(a[7]), .Z(n1352) );
  NANDN U1879 ( .A(n18194), .B(n1352), .Z(n1253) );
  NAND U1880 ( .A(n1251), .B(n18104), .Z(n1252) );
  NAND U1881 ( .A(n1253), .B(n1252), .Z(n1370) );
  XNOR U1882 ( .A(b[13]), .B(a[5]), .Z(n1361) );
  NANDN U1883 ( .A(n1361), .B(n18336), .Z(n1256) );
  NANDN U1884 ( .A(n1254), .B(n18337), .Z(n1255) );
  AND U1885 ( .A(n1256), .B(n1255), .Z(n1371) );
  XNOR U1886 ( .A(n1370), .B(n1371), .Z(n1372) );
  XOR U1887 ( .A(n1373), .B(n1372), .Z(n1326) );
  XNOR U1888 ( .A(n1325), .B(n1326), .Z(n1327) );
  XNOR U1889 ( .A(n1327), .B(n1328), .Z(n1332) );
  NAND U1890 ( .A(n1262), .B(n1261), .Z(n1266) );
  OR U1891 ( .A(n1264), .B(n1263), .Z(n1265) );
  NAND U1892 ( .A(n1266), .B(n1265), .Z(n1329) );
  NANDN U1893 ( .A(n1268), .B(n1267), .Z(n1272) );
  NAND U1894 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U1895 ( .A(n1272), .B(n1271), .Z(n1379) );
  NANDN U1896 ( .A(n1273), .B(n18513), .Z(n1275) );
  XOR U1897 ( .A(b[15]), .B(a[3]), .Z(n1344) );
  NANDN U1898 ( .A(n18512), .B(n1344), .Z(n1274) );
  NAND U1899 ( .A(n1275), .B(n1274), .Z(n1348) );
  XNOR U1900 ( .A(b[17]), .B(n2921), .Z(n1278) );
  XOR U1901 ( .A(b[17]), .B(b[15]), .Z(n1277) );
  XOR U1902 ( .A(b[17]), .B(b[16]), .Z(n1276) );
  AND U1903 ( .A(n1277), .B(n1276), .Z(n18674) );
  NAND U1904 ( .A(n1278), .B(n18674), .Z(n1280) );
  XOR U1905 ( .A(b[17]), .B(a[1]), .Z(n1349) );
  NAND U1906 ( .A(n1349), .B(n18673), .Z(n1279) );
  NAND U1907 ( .A(n1280), .B(n1279), .Z(n1347) );
  XNOR U1908 ( .A(n1348), .B(n1347), .Z(n1338) );
  ANDN U1909 ( .B(b[15]), .A(n2921), .Z(n1284) );
  OR U1910 ( .A(b[15]), .B(a[0]), .Z(n1281) );
  NAND U1911 ( .A(n1281), .B(b[16]), .Z(n1282) );
  AND U1912 ( .A(b[17]), .B(n1282), .Z(n1283) );
  NANDN U1913 ( .A(n1284), .B(n1283), .Z(n1335) );
  XNOR U1914 ( .A(b[9]), .B(a[9]), .Z(n1358) );
  NANDN U1915 ( .A(n1358), .B(n17814), .Z(n1287) );
  NANDN U1916 ( .A(n1285), .B(n17815), .Z(n1286) );
  NAND U1917 ( .A(n1287), .B(n1286), .Z(n1336) );
  XNOR U1918 ( .A(n1335), .B(n1336), .Z(n1337) );
  XOR U1919 ( .A(n1338), .B(n1337), .Z(n1376) );
  NANDN U1920 ( .A(n577), .B(a[17]), .Z(n1288) );
  XOR U1921 ( .A(n17151), .B(n1288), .Z(n1290) );
  NANDN U1922 ( .A(b[0]), .B(a[16]), .Z(n1289) );
  AND U1923 ( .A(n1290), .B(n1289), .Z(n1384) );
  XOR U1924 ( .A(b[3]), .B(n5159), .Z(n1355) );
  NANDN U1925 ( .A(n1355), .B(n16990), .Z(n1293) );
  OR U1926 ( .A(n1291), .B(n16988), .Z(n1292) );
  NAND U1927 ( .A(n1293), .B(n1292), .Z(n1382) );
  XNOR U1928 ( .A(b[5]), .B(n4875), .Z(n1364) );
  NAND U1929 ( .A(n1364), .B(n17310), .Z(n1296) );
  NAND U1930 ( .A(n1294), .B(n17311), .Z(n1295) );
  AND U1931 ( .A(n1296), .B(n1295), .Z(n1383) );
  XNOR U1932 ( .A(n1382), .B(n1383), .Z(n1385) );
  XNOR U1933 ( .A(n1384), .B(n1385), .Z(n1377) );
  XOR U1934 ( .A(n1376), .B(n1377), .Z(n1378) );
  XNOR U1935 ( .A(n1379), .B(n1378), .Z(n1330) );
  XNOR U1936 ( .A(n1329), .B(n1330), .Z(n1331) );
  XOR U1937 ( .A(n1332), .B(n1331), .Z(n1322) );
  XOR U1938 ( .A(n1321), .B(n1322), .Z(n1313) );
  NANDN U1939 ( .A(n1298), .B(n1297), .Z(n1302) );
  NAND U1940 ( .A(n1300), .B(n1299), .Z(n1301) );
  AND U1941 ( .A(n1302), .B(n1301), .Z(n1314) );
  XNOR U1942 ( .A(n1313), .B(n1314), .Z(n1315) );
  XNOR U1943 ( .A(n1316), .B(n1315), .Z(n1308) );
  XNOR U1944 ( .A(n1308), .B(sreg[113]), .Z(n1310) );
  NAND U1945 ( .A(n1303), .B(sreg[112]), .Z(n1307) );
  OR U1946 ( .A(n1305), .B(n1304), .Z(n1306) );
  AND U1947 ( .A(n1307), .B(n1306), .Z(n1309) );
  XOR U1948 ( .A(n1310), .B(n1309), .Z(c[113]) );
  NAND U1949 ( .A(n1308), .B(sreg[113]), .Z(n1312) );
  OR U1950 ( .A(n1310), .B(n1309), .Z(n1311) );
  NAND U1951 ( .A(n1312), .B(n1311), .Z(n1470) );
  XNOR U1952 ( .A(n1470), .B(sreg[114]), .Z(n1472) );
  NANDN U1953 ( .A(n1314), .B(n1313), .Z(n1318) );
  NAND U1954 ( .A(n1316), .B(n1315), .Z(n1317) );
  NAND U1955 ( .A(n1318), .B(n1317), .Z(n1389) );
  NANDN U1956 ( .A(n1320), .B(n1319), .Z(n1324) );
  NANDN U1957 ( .A(n1322), .B(n1321), .Z(n1323) );
  NAND U1958 ( .A(n1324), .B(n1323), .Z(n1387) );
  NANDN U1959 ( .A(n1330), .B(n1329), .Z(n1334) );
  NANDN U1960 ( .A(n1332), .B(n1331), .Z(n1333) );
  NAND U1961 ( .A(n1334), .B(n1333), .Z(n1393) );
  XNOR U1962 ( .A(n1392), .B(n1393), .Z(n1394) );
  NANDN U1963 ( .A(n1336), .B(n1335), .Z(n1340) );
  NAND U1964 ( .A(n1338), .B(n1337), .Z(n1339) );
  NAND U1965 ( .A(n1340), .B(n1339), .Z(n1407) );
  NANDN U1966 ( .A(n577), .B(a[18]), .Z(n1341) );
  XOR U1967 ( .A(n17151), .B(n1341), .Z(n1343) );
  NANDN U1968 ( .A(b[0]), .B(a[17]), .Z(n1342) );
  AND U1969 ( .A(n1343), .B(n1342), .Z(n1458) );
  NAND U1970 ( .A(n1344), .B(n18513), .Z(n1346) );
  XOR U1971 ( .A(b[15]), .B(a[4]), .Z(n1440) );
  NANDN U1972 ( .A(n18512), .B(n1440), .Z(n1345) );
  AND U1973 ( .A(n1346), .B(n1345), .Z(n1459) );
  XOR U1974 ( .A(n1458), .B(n1459), .Z(n1461) );
  XOR U1975 ( .A(b[17]), .B(b[18]), .Z(n18834) );
  NANDN U1976 ( .A(n2921), .B(n18834), .Z(n1460) );
  XNOR U1977 ( .A(n1461), .B(n1460), .Z(n1404) );
  NAND U1978 ( .A(n1348), .B(n1347), .Z(n1428) );
  XOR U1979 ( .A(b[17]), .B(a[2]), .Z(n1408) );
  NAND U1980 ( .A(n18673), .B(n1408), .Z(n1351) );
  NAND U1981 ( .A(n18674), .B(n1349), .Z(n1350) );
  NAND U1982 ( .A(n1351), .B(n1350), .Z(n1426) );
  XOR U1983 ( .A(b[11]), .B(a[8]), .Z(n1452) );
  NANDN U1984 ( .A(n18194), .B(n1452), .Z(n1354) );
  NAND U1985 ( .A(n18104), .B(n1352), .Z(n1353) );
  AND U1986 ( .A(n1354), .B(n1353), .Z(n1425) );
  XNOR U1987 ( .A(n1426), .B(n1425), .Z(n1427) );
  XNOR U1988 ( .A(n1428), .B(n1427), .Z(n1405) );
  XNOR U1989 ( .A(n1404), .B(n1405), .Z(n1406) );
  XNOR U1990 ( .A(n1407), .B(n1406), .Z(n1467) );
  OR U1991 ( .A(n1355), .B(n16988), .Z(n1357) );
  XNOR U1992 ( .A(b[3]), .B(a[16]), .Z(n1446) );
  NANDN U1993 ( .A(n1446), .B(n16990), .Z(n1356) );
  NAND U1994 ( .A(n1357), .B(n1356), .Z(n1422) );
  XNOR U1995 ( .A(n579), .B(a[10]), .Z(n1416) );
  NAND U1996 ( .A(n17814), .B(n1416), .Z(n1360) );
  NANDN U1997 ( .A(n1358), .B(n17815), .Z(n1359) );
  NAND U1998 ( .A(n1360), .B(n1359), .Z(n1419) );
  XNOR U1999 ( .A(b[13]), .B(a[6]), .Z(n1437) );
  NANDN U2000 ( .A(n1437), .B(n18336), .Z(n1363) );
  NANDN U2001 ( .A(n1361), .B(n18337), .Z(n1362) );
  AND U2002 ( .A(n1363), .B(n1362), .Z(n1420) );
  XNOR U2003 ( .A(n1419), .B(n1420), .Z(n1421) );
  XNOR U2004 ( .A(n1422), .B(n1421), .Z(n1434) );
  XOR U2005 ( .A(b[5]), .B(a[14]), .Z(n1443) );
  NAND U2006 ( .A(n17310), .B(n1443), .Z(n1366) );
  NAND U2007 ( .A(n17311), .B(n1364), .Z(n1365) );
  NAND U2008 ( .A(n1366), .B(n1365), .Z(n1432) );
  XNOR U2009 ( .A(b[7]), .B(a[12]), .Z(n1455) );
  NANDN U2010 ( .A(n1455), .B(n17555), .Z(n1369) );
  NANDN U2011 ( .A(n1367), .B(n17553), .Z(n1368) );
  AND U2012 ( .A(n1369), .B(n1368), .Z(n1431) );
  XNOR U2013 ( .A(n1432), .B(n1431), .Z(n1433) );
  XOR U2014 ( .A(n1434), .B(n1433), .Z(n1465) );
  NANDN U2015 ( .A(n1371), .B(n1370), .Z(n1375) );
  NAND U2016 ( .A(n1373), .B(n1372), .Z(n1374) );
  AND U2017 ( .A(n1375), .B(n1374), .Z(n1464) );
  XOR U2018 ( .A(n1465), .B(n1464), .Z(n1466) );
  XOR U2019 ( .A(n1467), .B(n1466), .Z(n1401) );
  OR U2020 ( .A(n1377), .B(n1376), .Z(n1381) );
  NAND U2021 ( .A(n1379), .B(n1378), .Z(n1380) );
  NAND U2022 ( .A(n1381), .B(n1380), .Z(n1399) );
  XNOR U2023 ( .A(n1399), .B(n1398), .Z(n1400) );
  XOR U2024 ( .A(n1401), .B(n1400), .Z(n1395) );
  XNOR U2025 ( .A(n1394), .B(n1395), .Z(n1386) );
  XNOR U2026 ( .A(n1387), .B(n1386), .Z(n1388) );
  XOR U2027 ( .A(n1389), .B(n1388), .Z(n1471) );
  XOR U2028 ( .A(n1472), .B(n1471), .Z(c[114]) );
  NANDN U2029 ( .A(n1387), .B(n1386), .Z(n1391) );
  NAND U2030 ( .A(n1389), .B(n1388), .Z(n1390) );
  NAND U2031 ( .A(n1391), .B(n1390), .Z(n1483) );
  NANDN U2032 ( .A(n1393), .B(n1392), .Z(n1397) );
  NANDN U2033 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U2034 ( .A(n1397), .B(n1396), .Z(n1480) );
  NANDN U2035 ( .A(n1399), .B(n1398), .Z(n1403) );
  NANDN U2036 ( .A(n1401), .B(n1400), .Z(n1402) );
  NAND U2037 ( .A(n1403), .B(n1402), .Z(n1489) );
  XOR U2038 ( .A(b[17]), .B(a[3]), .Z(n1528) );
  NAND U2039 ( .A(n1528), .B(n18673), .Z(n1410) );
  NAND U2040 ( .A(n1408), .B(n18674), .Z(n1409) );
  NAND U2041 ( .A(n1410), .B(n1409), .Z(n1542) );
  XNOR U2042 ( .A(n581), .B(a[0]), .Z(n1413) );
  XNOR U2043 ( .A(n581), .B(b[17]), .Z(n1412) );
  XNOR U2044 ( .A(n581), .B(b[18]), .Z(n1411) );
  AND U2045 ( .A(n1412), .B(n1411), .Z(n18832) );
  NAND U2046 ( .A(n1413), .B(n18832), .Z(n1415) );
  XNOR U2047 ( .A(n581), .B(a[1]), .Z(n1543) );
  NAND U2048 ( .A(n1543), .B(n18834), .Z(n1414) );
  NAND U2049 ( .A(n1415), .B(n1414), .Z(n1541) );
  XNOR U2050 ( .A(n1542), .B(n1541), .Z(n1534) );
  XOR U2051 ( .A(n579), .B(a[11]), .Z(n1549) );
  NANDN U2052 ( .A(n1549), .B(n17814), .Z(n1418) );
  NAND U2053 ( .A(n17815), .B(n1416), .Z(n1417) );
  AND U2054 ( .A(n1418), .B(n1417), .Z(n1531) );
  XNOR U2055 ( .A(n1532), .B(n1531), .Z(n1533) );
  XOR U2056 ( .A(n1534), .B(n1533), .Z(n1499) );
  NANDN U2057 ( .A(n1420), .B(n1419), .Z(n1424) );
  NAND U2058 ( .A(n1422), .B(n1421), .Z(n1423) );
  AND U2059 ( .A(n1424), .B(n1423), .Z(n1498) );
  XOR U2060 ( .A(n1499), .B(n1498), .Z(n1500) );
  NANDN U2061 ( .A(n1426), .B(n1425), .Z(n1430) );
  NAND U2062 ( .A(n1428), .B(n1427), .Z(n1429) );
  AND U2063 ( .A(n1430), .B(n1429), .Z(n1501) );
  XOR U2064 ( .A(n1500), .B(n1501), .Z(n1558) );
  XNOR U2065 ( .A(n1559), .B(n1558), .Z(n1560) );
  NANDN U2066 ( .A(n1432), .B(n1431), .Z(n1436) );
  NAND U2067 ( .A(n1434), .B(n1433), .Z(n1435) );
  NAND U2068 ( .A(n1436), .B(n1435), .Z(n1493) );
  XNOR U2069 ( .A(b[13]), .B(a[7]), .Z(n1552) );
  NANDN U2070 ( .A(n1552), .B(n18336), .Z(n1439) );
  NANDN U2071 ( .A(n1437), .B(n18337), .Z(n1438) );
  NAND U2072 ( .A(n1439), .B(n1438), .Z(n1513) );
  NAND U2073 ( .A(n1440), .B(n18513), .Z(n1442) );
  XOR U2074 ( .A(b[15]), .B(a[5]), .Z(n1555) );
  NANDN U2075 ( .A(n18512), .B(n1555), .Z(n1441) );
  NAND U2076 ( .A(n1442), .B(n1441), .Z(n1510) );
  XNOR U2077 ( .A(b[5]), .B(n5159), .Z(n1519) );
  NAND U2078 ( .A(n1519), .B(n17310), .Z(n1445) );
  NAND U2079 ( .A(n1443), .B(n17311), .Z(n1444) );
  AND U2080 ( .A(n1445), .B(n1444), .Z(n1511) );
  XNOR U2081 ( .A(n1510), .B(n1511), .Z(n1512) );
  XNOR U2082 ( .A(n1513), .B(n1512), .Z(n1507) );
  OR U2083 ( .A(n1446), .B(n16988), .Z(n1448) );
  XNOR U2084 ( .A(n578), .B(a[17]), .Z(n1516) );
  NAND U2085 ( .A(n1516), .B(n16990), .Z(n1447) );
  NAND U2086 ( .A(n1448), .B(n1447), .Z(n1540) );
  NANDN U2087 ( .A(n577), .B(a[19]), .Z(n1449) );
  XOR U2088 ( .A(n17151), .B(n1449), .Z(n1451) );
  NANDN U2089 ( .A(b[0]), .B(a[18]), .Z(n1450) );
  AND U2090 ( .A(n1451), .B(n1450), .Z(n1537) );
  XOR U2091 ( .A(b[11]), .B(a[9]), .Z(n1546) );
  NANDN U2092 ( .A(n18194), .B(n1546), .Z(n1454) );
  NAND U2093 ( .A(n1452), .B(n18104), .Z(n1453) );
  AND U2094 ( .A(n1454), .B(n1453), .Z(n1538) );
  XNOR U2095 ( .A(n1537), .B(n1538), .Z(n1539) );
  XNOR U2096 ( .A(n1540), .B(n1539), .Z(n1504) );
  XNOR U2097 ( .A(b[7]), .B(a[13]), .Z(n1522) );
  NANDN U2098 ( .A(n1522), .B(n17555), .Z(n1457) );
  NANDN U2099 ( .A(n1455), .B(n17553), .Z(n1456) );
  NAND U2100 ( .A(n1457), .B(n1456), .Z(n1505) );
  XNOR U2101 ( .A(n1504), .B(n1505), .Z(n1506) );
  XOR U2102 ( .A(n1507), .B(n1506), .Z(n1492) );
  XNOR U2103 ( .A(n1493), .B(n1492), .Z(n1495) );
  NANDN U2104 ( .A(n1459), .B(n1458), .Z(n1463) );
  OR U2105 ( .A(n1461), .B(n1460), .Z(n1462) );
  AND U2106 ( .A(n1463), .B(n1462), .Z(n1494) );
  XOR U2107 ( .A(n1495), .B(n1494), .Z(n1561) );
  XOR U2108 ( .A(n1560), .B(n1561), .Z(n1486) );
  OR U2109 ( .A(n1465), .B(n1464), .Z(n1469) );
  NAND U2110 ( .A(n1467), .B(n1466), .Z(n1468) );
  NAND U2111 ( .A(n1469), .B(n1468), .Z(n1487) );
  XOR U2112 ( .A(n1486), .B(n1487), .Z(n1488) );
  XNOR U2113 ( .A(n1489), .B(n1488), .Z(n1481) );
  XNOR U2114 ( .A(n1480), .B(n1481), .Z(n1482) );
  XNOR U2115 ( .A(n1483), .B(n1482), .Z(n1475) );
  XNOR U2116 ( .A(n1475), .B(sreg[115]), .Z(n1477) );
  NAND U2117 ( .A(n1470), .B(sreg[114]), .Z(n1474) );
  OR U2118 ( .A(n1472), .B(n1471), .Z(n1473) );
  AND U2119 ( .A(n1474), .B(n1473), .Z(n1476) );
  XOR U2120 ( .A(n1477), .B(n1476), .Z(c[115]) );
  NAND U2121 ( .A(n1475), .B(sreg[115]), .Z(n1479) );
  OR U2122 ( .A(n1477), .B(n1476), .Z(n1478) );
  NAND U2123 ( .A(n1479), .B(n1478), .Z(n1647) );
  XNOR U2124 ( .A(n1647), .B(sreg[116]), .Z(n1649) );
  NANDN U2125 ( .A(n1481), .B(n1480), .Z(n1485) );
  NAND U2126 ( .A(n1483), .B(n1482), .Z(n1484) );
  NAND U2127 ( .A(n1485), .B(n1484), .Z(n1565) );
  OR U2128 ( .A(n1487), .B(n1486), .Z(n1491) );
  NAND U2129 ( .A(n1489), .B(n1488), .Z(n1490) );
  NAND U2130 ( .A(n1491), .B(n1490), .Z(n1562) );
  OR U2131 ( .A(n1493), .B(n1492), .Z(n1497) );
  OR U2132 ( .A(n1495), .B(n1494), .Z(n1496) );
  NAND U2133 ( .A(n1497), .B(n1496), .Z(n1571) );
  OR U2134 ( .A(n1499), .B(n1498), .Z(n1503) );
  NAND U2135 ( .A(n1501), .B(n1500), .Z(n1502) );
  NAND U2136 ( .A(n1503), .B(n1502), .Z(n1572) );
  NANDN U2137 ( .A(n1505), .B(n1504), .Z(n1509) );
  NAND U2138 ( .A(n1507), .B(n1506), .Z(n1508) );
  NAND U2139 ( .A(n1509), .B(n1508), .Z(n1573) );
  XNOR U2140 ( .A(n1572), .B(n1573), .Z(n1574) );
  NANDN U2141 ( .A(n1511), .B(n1510), .Z(n1515) );
  NAND U2142 ( .A(n1513), .B(n1512), .Z(n1514) );
  NAND U2143 ( .A(n1515), .B(n1514), .Z(n1591) );
  XNOR U2144 ( .A(b[3]), .B(a[18]), .Z(n1622) );
  NANDN U2145 ( .A(n1622), .B(n16990), .Z(n1518) );
  NANDN U2146 ( .A(n16988), .B(n1516), .Z(n1517) );
  NAND U2147 ( .A(n1518), .B(n1517), .Z(n1596) );
  XOR U2148 ( .A(b[5]), .B(a[16]), .Z(n1631) );
  NAND U2149 ( .A(n17310), .B(n1631), .Z(n1521) );
  NAND U2150 ( .A(n17311), .B(n1519), .Z(n1520) );
  NAND U2151 ( .A(n1521), .B(n1520), .Z(n1594) );
  XNOR U2152 ( .A(b[7]), .B(a[14]), .Z(n1628) );
  NANDN U2153 ( .A(n1628), .B(n17555), .Z(n1524) );
  NANDN U2154 ( .A(n1522), .B(n17553), .Z(n1523) );
  NAND U2155 ( .A(n1524), .B(n1523), .Z(n1595) );
  XNOR U2156 ( .A(n1594), .B(n1595), .Z(n1597) );
  XOR U2157 ( .A(n1596), .B(n1597), .Z(n1588) );
  NANDN U2158 ( .A(n577), .B(a[20]), .Z(n1525) );
  XOR U2159 ( .A(n17151), .B(n1525), .Z(n1527) );
  NANDN U2160 ( .A(b[0]), .B(a[19]), .Z(n1526) );
  AND U2161 ( .A(n1527), .B(n1526), .Z(n1613) );
  XOR U2162 ( .A(b[17]), .B(a[4]), .Z(n1637) );
  NAND U2163 ( .A(n1637), .B(n18673), .Z(n1530) );
  NAND U2164 ( .A(n1528), .B(n18674), .Z(n1529) );
  AND U2165 ( .A(n1530), .B(n1529), .Z(n1614) );
  XOR U2166 ( .A(n1613), .B(n1614), .Z(n1616) );
  XNOR U2167 ( .A(n581), .B(b[20]), .Z(n19015) );
  NANDN U2168 ( .A(n2921), .B(n19015), .Z(n1615) );
  XOR U2169 ( .A(n1616), .B(n1615), .Z(n1589) );
  XNOR U2170 ( .A(n1588), .B(n1589), .Z(n1590) );
  XOR U2171 ( .A(n1591), .B(n1590), .Z(n1578) );
  NANDN U2172 ( .A(n1532), .B(n1531), .Z(n1536) );
  NAND U2173 ( .A(n1534), .B(n1533), .Z(n1535) );
  NAND U2174 ( .A(n1536), .B(n1535), .Z(n1579) );
  XNOR U2175 ( .A(n1578), .B(n1579), .Z(n1580) );
  NAND U2176 ( .A(n1542), .B(n1541), .Z(n1645) );
  XNOR U2177 ( .A(b[19]), .B(a[2]), .Z(n1602) );
  NANDN U2178 ( .A(n1602), .B(n18834), .Z(n1545) );
  NAND U2179 ( .A(n18832), .B(n1543), .Z(n1544) );
  NAND U2180 ( .A(n1545), .B(n1544), .Z(n1644) );
  XNOR U2181 ( .A(b[11]), .B(a[10]), .Z(n1610) );
  OR U2182 ( .A(n1610), .B(n18194), .Z(n1548) );
  NAND U2183 ( .A(n18104), .B(n1546), .Z(n1547) );
  AND U2184 ( .A(n1548), .B(n1547), .Z(n1643) );
  XNOR U2185 ( .A(n1644), .B(n1643), .Z(n1646) );
  XNOR U2186 ( .A(n1645), .B(n1646), .Z(n1599) );
  XOR U2187 ( .A(n579), .B(a[12]), .Z(n1625) );
  NANDN U2188 ( .A(n1625), .B(n17814), .Z(n1551) );
  NANDN U2189 ( .A(n1549), .B(n17815), .Z(n1550) );
  NAND U2190 ( .A(n1551), .B(n1550), .Z(n1586) );
  XNOR U2191 ( .A(b[13]), .B(a[8]), .Z(n1634) );
  NANDN U2192 ( .A(n1634), .B(n18336), .Z(n1554) );
  NANDN U2193 ( .A(n1552), .B(n18337), .Z(n1553) );
  NAND U2194 ( .A(n1554), .B(n1553), .Z(n1584) );
  NAND U2195 ( .A(n1555), .B(n18513), .Z(n1557) );
  XOR U2196 ( .A(b[15]), .B(a[6]), .Z(n1640) );
  NANDN U2197 ( .A(n18512), .B(n1640), .Z(n1556) );
  AND U2198 ( .A(n1557), .B(n1556), .Z(n1585) );
  XNOR U2199 ( .A(n1584), .B(n1585), .Z(n1587) );
  XOR U2200 ( .A(n1586), .B(n1587), .Z(n1598) );
  XOR U2201 ( .A(n1599), .B(n1598), .Z(n1600) );
  XOR U2202 ( .A(n1601), .B(n1600), .Z(n1581) );
  XOR U2203 ( .A(n1580), .B(n1581), .Z(n1575) );
  XNOR U2204 ( .A(n1574), .B(n1575), .Z(n1568) );
  XNOR U2205 ( .A(n1568), .B(n1569), .Z(n1570) );
  XOR U2206 ( .A(n1571), .B(n1570), .Z(n1563) );
  XNOR U2207 ( .A(n1562), .B(n1563), .Z(n1564) );
  XOR U2208 ( .A(n1565), .B(n1564), .Z(n1648) );
  XOR U2209 ( .A(n1649), .B(n1648), .Z(c[116]) );
  NANDN U2210 ( .A(n1563), .B(n1562), .Z(n1567) );
  NAND U2211 ( .A(n1565), .B(n1564), .Z(n1566) );
  NAND U2212 ( .A(n1567), .B(n1566), .Z(n1660) );
  NANDN U2213 ( .A(n1573), .B(n1572), .Z(n1577) );
  NAND U2214 ( .A(n1575), .B(n1574), .Z(n1576) );
  NAND U2215 ( .A(n1577), .B(n1576), .Z(n1747) );
  NANDN U2216 ( .A(n1579), .B(n1578), .Z(n1583) );
  NAND U2217 ( .A(n1581), .B(n1580), .Z(n1582) );
  NAND U2218 ( .A(n1583), .B(n1582), .Z(n1745) );
  NANDN U2219 ( .A(n1589), .B(n1588), .Z(n1593) );
  NANDN U2220 ( .A(n1591), .B(n1590), .Z(n1592) );
  NAND U2221 ( .A(n1593), .B(n1592), .Z(n1663) );
  XNOR U2222 ( .A(n1663), .B(n1664), .Z(n1665) );
  XNOR U2223 ( .A(n1666), .B(n1665), .Z(n1669) );
  NANDN U2224 ( .A(n1602), .B(n18832), .Z(n1604) );
  XNOR U2225 ( .A(b[19]), .B(a[3]), .Z(n1735) );
  NANDN U2226 ( .A(n1735), .B(n18834), .Z(n1603) );
  NAND U2227 ( .A(n1604), .B(n1603), .Z(n1725) );
  XNOR U2228 ( .A(b[21]), .B(a[1]), .Z(n1694) );
  ANDN U2229 ( .B(n19015), .A(n1694), .Z(n1609) );
  XNOR U2230 ( .A(n582), .B(a[0]), .Z(n1607) );
  XNOR U2231 ( .A(n582), .B(b[19]), .Z(n1606) );
  XNOR U2232 ( .A(n582), .B(b[20]), .Z(n1605) );
  AND U2233 ( .A(n1606), .B(n1605), .Z(n19013) );
  NAND U2234 ( .A(n1607), .B(n19013), .Z(n1608) );
  NANDN U2235 ( .A(n1609), .B(n1608), .Z(n1724) );
  XNOR U2236 ( .A(n1725), .B(n1724), .Z(n1721) );
  XOR U2237 ( .A(b[11]), .B(n4573), .Z(n1697) );
  OR U2238 ( .A(n1697), .B(n18194), .Z(n1612) );
  NANDN U2239 ( .A(n1610), .B(n18104), .Z(n1611) );
  AND U2240 ( .A(n1612), .B(n1611), .Z(n1718) );
  XNOR U2241 ( .A(n1719), .B(n1718), .Z(n1720) );
  XOR U2242 ( .A(n1721), .B(n1720), .Z(n1676) );
  NANDN U2243 ( .A(n1614), .B(n1613), .Z(n1618) );
  OR U2244 ( .A(n1616), .B(n1615), .Z(n1617) );
  NAND U2245 ( .A(n1618), .B(n1617), .Z(n1674) );
  NANDN U2246 ( .A(n577), .B(a[21]), .Z(n1619) );
  XOR U2247 ( .A(n17151), .B(n1619), .Z(n1621) );
  NANDN U2248 ( .A(b[0]), .B(a[20]), .Z(n1620) );
  AND U2249 ( .A(n1621), .B(n1620), .Z(n1707) );
  XNOR U2250 ( .A(b[3]), .B(a[19]), .Z(n1729) );
  NANDN U2251 ( .A(n1729), .B(n16990), .Z(n1624) );
  OR U2252 ( .A(n1622), .B(n16988), .Z(n1623) );
  AND U2253 ( .A(n1624), .B(n1623), .Z(n1706) );
  XNOR U2254 ( .A(n1707), .B(n1706), .Z(n1708) );
  XOR U2255 ( .A(b[9]), .B(n4875), .Z(n1688) );
  NANDN U2256 ( .A(n1688), .B(n17814), .Z(n1627) );
  NANDN U2257 ( .A(n1625), .B(n17815), .Z(n1626) );
  NAND U2258 ( .A(n1627), .B(n1626), .Z(n1709) );
  XOR U2259 ( .A(n1708), .B(n1709), .Z(n1673) );
  XOR U2260 ( .A(n1674), .B(n1673), .Z(n1675) );
  XOR U2261 ( .A(n1676), .B(n1675), .Z(n1740) );
  NANDN U2262 ( .A(n1628), .B(n17553), .Z(n1630) );
  XNOR U2263 ( .A(b[7]), .B(a[15]), .Z(n1679) );
  NANDN U2264 ( .A(n1679), .B(n17555), .Z(n1629) );
  NAND U2265 ( .A(n1630), .B(n1629), .Z(n1712) );
  XOR U2266 ( .A(b[5]), .B(a[17]), .Z(n1682) );
  NAND U2267 ( .A(n1682), .B(n17310), .Z(n1633) );
  NAND U2268 ( .A(n1631), .B(n17311), .Z(n1632) );
  AND U2269 ( .A(n1633), .B(n1632), .Z(n1713) );
  XNOR U2270 ( .A(n1712), .B(n1713), .Z(n1714) );
  XNOR U2271 ( .A(n580), .B(a[9]), .Z(n1726) );
  NAND U2272 ( .A(n1726), .B(n18336), .Z(n1636) );
  NANDN U2273 ( .A(n1634), .B(n18337), .Z(n1635) );
  NAND U2274 ( .A(n1636), .B(n1635), .Z(n1703) );
  XOR U2275 ( .A(b[17]), .B(a[5]), .Z(n1691) );
  NAND U2276 ( .A(n1691), .B(n18673), .Z(n1639) );
  NAND U2277 ( .A(n1637), .B(n18674), .Z(n1638) );
  NAND U2278 ( .A(n1639), .B(n1638), .Z(n1700) );
  NAND U2279 ( .A(n1640), .B(n18513), .Z(n1642) );
  XOR U2280 ( .A(b[15]), .B(a[7]), .Z(n1685) );
  NANDN U2281 ( .A(n18512), .B(n1685), .Z(n1641) );
  AND U2282 ( .A(n1642), .B(n1641), .Z(n1701) );
  XNOR U2283 ( .A(n1700), .B(n1701), .Z(n1702) );
  XOR U2284 ( .A(n1703), .B(n1702), .Z(n1715) );
  XOR U2285 ( .A(n1714), .B(n1715), .Z(n1738) );
  XNOR U2286 ( .A(n1738), .B(n1739), .Z(n1741) );
  XOR U2287 ( .A(n1740), .B(n1741), .Z(n1667) );
  XNOR U2288 ( .A(n1668), .B(n1667), .Z(n1670) );
  XOR U2289 ( .A(n1669), .B(n1670), .Z(n1744) );
  XOR U2290 ( .A(n1745), .B(n1744), .Z(n1746) );
  XOR U2291 ( .A(n1747), .B(n1746), .Z(n1658) );
  XNOR U2292 ( .A(n1657), .B(n1658), .Z(n1659) );
  XNOR U2293 ( .A(n1660), .B(n1659), .Z(n1652) );
  XNOR U2294 ( .A(n1652), .B(sreg[117]), .Z(n1654) );
  NAND U2295 ( .A(n1647), .B(sreg[116]), .Z(n1651) );
  OR U2296 ( .A(n1649), .B(n1648), .Z(n1650) );
  AND U2297 ( .A(n1651), .B(n1650), .Z(n1653) );
  XOR U2298 ( .A(n1654), .B(n1653), .Z(c[117]) );
  NAND U2299 ( .A(n1652), .B(sreg[117]), .Z(n1656) );
  OR U2300 ( .A(n1654), .B(n1653), .Z(n1655) );
  NAND U2301 ( .A(n1656), .B(n1655), .Z(n1856) );
  XNOR U2302 ( .A(n1856), .B(sreg[118]), .Z(n1858) );
  NANDN U2303 ( .A(n1658), .B(n1657), .Z(n1662) );
  NAND U2304 ( .A(n1660), .B(n1659), .Z(n1661) );
  NAND U2305 ( .A(n1662), .B(n1661), .Z(n1753) );
  NAND U2306 ( .A(n1668), .B(n1667), .Z(n1672) );
  OR U2307 ( .A(n1670), .B(n1669), .Z(n1671) );
  NAND U2308 ( .A(n1672), .B(n1671), .Z(n1757) );
  XNOR U2309 ( .A(n1756), .B(n1757), .Z(n1758) );
  OR U2310 ( .A(n1674), .B(n1673), .Z(n1678) );
  NAND U2311 ( .A(n1676), .B(n1675), .Z(n1677) );
  NAND U2312 ( .A(n1678), .B(n1677), .Z(n1764) );
  NANDN U2313 ( .A(n1679), .B(n17553), .Z(n1681) );
  XOR U2314 ( .A(b[7]), .B(a[16]), .Z(n1774) );
  NAND U2315 ( .A(n1774), .B(n17555), .Z(n1680) );
  NAND U2316 ( .A(n1681), .B(n1680), .Z(n1800) );
  XOR U2317 ( .A(b[5]), .B(a[18]), .Z(n1780) );
  NAND U2318 ( .A(n1780), .B(n17310), .Z(n1684) );
  NAND U2319 ( .A(n1682), .B(n17311), .Z(n1683) );
  NAND U2320 ( .A(n1684), .B(n1683), .Z(n1797) );
  NAND U2321 ( .A(n1685), .B(n18513), .Z(n1687) );
  XOR U2322 ( .A(b[15]), .B(a[8]), .Z(n1829) );
  NANDN U2323 ( .A(n18512), .B(n1829), .Z(n1686) );
  AND U2324 ( .A(n1687), .B(n1686), .Z(n1798) );
  XNOR U2325 ( .A(n1797), .B(n1798), .Z(n1799) );
  XNOR U2326 ( .A(n1800), .B(n1799), .Z(n1834) );
  XNOR U2327 ( .A(b[9]), .B(a[14]), .Z(n1777) );
  NANDN U2328 ( .A(n1777), .B(n17814), .Z(n1690) );
  NANDN U2329 ( .A(n1688), .B(n17815), .Z(n1689) );
  NAND U2330 ( .A(n1690), .B(n1689), .Z(n1806) );
  XOR U2331 ( .A(b[17]), .B(a[6]), .Z(n1815) );
  NAND U2332 ( .A(n1815), .B(n18673), .Z(n1693) );
  NAND U2333 ( .A(n1691), .B(n18674), .Z(n1692) );
  NAND U2334 ( .A(n1693), .B(n1692), .Z(n1803) );
  NANDN U2335 ( .A(n1694), .B(n19013), .Z(n1696) );
  XNOR U2336 ( .A(b[21]), .B(a[2]), .Z(n1789) );
  NANDN U2337 ( .A(n1789), .B(n19015), .Z(n1695) );
  AND U2338 ( .A(n1696), .B(n1695), .Z(n1804) );
  XNOR U2339 ( .A(n1803), .B(n1804), .Z(n1805) );
  XNOR U2340 ( .A(n1806), .B(n1805), .Z(n1832) );
  XOR U2341 ( .A(b[11]), .B(a[12]), .Z(n1786) );
  NANDN U2342 ( .A(n18194), .B(n1786), .Z(n1699) );
  NANDN U2343 ( .A(n1697), .B(n18104), .Z(n1698) );
  NAND U2344 ( .A(n1699), .B(n1698), .Z(n1833) );
  XOR U2345 ( .A(n1832), .B(n1833), .Z(n1835) );
  XNOR U2346 ( .A(n1834), .B(n1835), .Z(n1853) );
  NANDN U2347 ( .A(n1701), .B(n1700), .Z(n1705) );
  NAND U2348 ( .A(n1703), .B(n1702), .Z(n1704) );
  NAND U2349 ( .A(n1705), .B(n1704), .Z(n1850) );
  NANDN U2350 ( .A(n1707), .B(n1706), .Z(n1711) );
  NANDN U2351 ( .A(n1709), .B(n1708), .Z(n1710) );
  NAND U2352 ( .A(n1711), .B(n1710), .Z(n1851) );
  XNOR U2353 ( .A(n1850), .B(n1851), .Z(n1852) );
  XNOR U2354 ( .A(n1853), .B(n1852), .Z(n1840) );
  NANDN U2355 ( .A(n1713), .B(n1712), .Z(n1717) );
  NAND U2356 ( .A(n1715), .B(n1714), .Z(n1716) );
  NAND U2357 ( .A(n1717), .B(n1716), .Z(n1839) );
  NANDN U2358 ( .A(n1719), .B(n1718), .Z(n1723) );
  NAND U2359 ( .A(n1721), .B(n1720), .Z(n1722) );
  NAND U2360 ( .A(n1723), .B(n1722), .Z(n1844) );
  NAND U2361 ( .A(n1725), .B(n1724), .Z(n1771) );
  XNOR U2362 ( .A(b[13]), .B(a[10]), .Z(n1821) );
  NANDN U2363 ( .A(n1821), .B(n18336), .Z(n1728) );
  NAND U2364 ( .A(n18337), .B(n1726), .Z(n1727) );
  NAND U2365 ( .A(n1728), .B(n1727), .Z(n1769) );
  XNOR U2366 ( .A(b[3]), .B(a[20]), .Z(n1826) );
  NANDN U2367 ( .A(n1826), .B(n16990), .Z(n1731) );
  OR U2368 ( .A(n1729), .B(n16988), .Z(n1730) );
  AND U2369 ( .A(n1731), .B(n1730), .Z(n1768) );
  XNOR U2370 ( .A(n1769), .B(n1768), .Z(n1770) );
  XNOR U2371 ( .A(n1771), .B(n1770), .Z(n1845) );
  XNOR U2372 ( .A(n1844), .B(n1845), .Z(n1846) );
  XNOR U2373 ( .A(b[21]), .B(b[22]), .Z(n19127) );
  NOR U2374 ( .A(n2921), .B(n19127), .Z(n1812) );
  NANDN U2375 ( .A(n577), .B(a[22]), .Z(n1732) );
  XOR U2376 ( .A(n17151), .B(n1732), .Z(n1734) );
  NANDN U2377 ( .A(b[0]), .B(a[21]), .Z(n1733) );
  AND U2378 ( .A(n1734), .B(n1733), .Z(n1810) );
  XNOR U2379 ( .A(b[19]), .B(a[4]), .Z(n1818) );
  NANDN U2380 ( .A(n1818), .B(n18834), .Z(n1737) );
  NANDN U2381 ( .A(n1735), .B(n18832), .Z(n1736) );
  AND U2382 ( .A(n1737), .B(n1736), .Z(n1809) );
  XNOR U2383 ( .A(n1810), .B(n1809), .Z(n1811) );
  XOR U2384 ( .A(n1812), .B(n1811), .Z(n1847) );
  XNOR U2385 ( .A(n1846), .B(n1847), .Z(n1838) );
  XOR U2386 ( .A(n1839), .B(n1838), .Z(n1841) );
  XOR U2387 ( .A(n1840), .B(n1841), .Z(n1762) );
  NAND U2388 ( .A(n1739), .B(n1738), .Z(n1743) );
  OR U2389 ( .A(n1741), .B(n1740), .Z(n1742) );
  AND U2390 ( .A(n1743), .B(n1742), .Z(n1763) );
  XNOR U2391 ( .A(n1762), .B(n1763), .Z(n1765) );
  XNOR U2392 ( .A(n1764), .B(n1765), .Z(n1759) );
  XOR U2393 ( .A(n1758), .B(n1759), .Z(n1750) );
  NAND U2394 ( .A(n1745), .B(n1744), .Z(n1749) );
  NAND U2395 ( .A(n1747), .B(n1746), .Z(n1748) );
  AND U2396 ( .A(n1749), .B(n1748), .Z(n1751) );
  XOR U2397 ( .A(n1750), .B(n1751), .Z(n1752) );
  XOR U2398 ( .A(n1753), .B(n1752), .Z(n1857) );
  XOR U2399 ( .A(n1858), .B(n1857), .Z(c[118]) );
  NAND U2400 ( .A(n1751), .B(n1750), .Z(n1755) );
  NAND U2401 ( .A(n1753), .B(n1752), .Z(n1754) );
  NAND U2402 ( .A(n1755), .B(n1754), .Z(n1869) );
  NANDN U2403 ( .A(n1757), .B(n1756), .Z(n1761) );
  NAND U2404 ( .A(n1759), .B(n1758), .Z(n1760) );
  NAND U2405 ( .A(n1761), .B(n1760), .Z(n1866) );
  NAND U2406 ( .A(n1763), .B(n1762), .Z(n1767) );
  NANDN U2407 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U2408 ( .A(n1767), .B(n1766), .Z(n1875) );
  NANDN U2409 ( .A(n1769), .B(n1768), .Z(n1773) );
  NAND U2410 ( .A(n1771), .B(n1770), .Z(n1772) );
  NAND U2411 ( .A(n1773), .B(n1772), .Z(n1953) );
  NAND U2412 ( .A(n1774), .B(n17553), .Z(n1776) );
  XOR U2413 ( .A(b[7]), .B(a[17]), .Z(n1929) );
  NAND U2414 ( .A(n1929), .B(n17555), .Z(n1775) );
  NAND U2415 ( .A(n1776), .B(n1775), .Z(n1947) );
  XOR U2416 ( .A(b[9]), .B(n5159), .Z(n1914) );
  NANDN U2417 ( .A(n1914), .B(n17814), .Z(n1779) );
  NANDN U2418 ( .A(n1777), .B(n17815), .Z(n1778) );
  NAND U2419 ( .A(n1779), .B(n1778), .Z(n1944) );
  XOR U2420 ( .A(b[5]), .B(a[19]), .Z(n1932) );
  NAND U2421 ( .A(n1932), .B(n17310), .Z(n1782) );
  NAND U2422 ( .A(n1780), .B(n17311), .Z(n1781) );
  AND U2423 ( .A(n1782), .B(n1781), .Z(n1945) );
  XNOR U2424 ( .A(n1944), .B(n1945), .Z(n1946) );
  XNOR U2425 ( .A(n1947), .B(n1946), .Z(n1951) );
  NANDN U2426 ( .A(n577), .B(a[23]), .Z(n1783) );
  XOR U2427 ( .A(n17151), .B(n1783), .Z(n1785) );
  NANDN U2428 ( .A(b[0]), .B(a[22]), .Z(n1784) );
  AND U2429 ( .A(n1785), .B(n1784), .Z(n1896) );
  XNOR U2430 ( .A(b[11]), .B(a[13]), .Z(n1908) );
  OR U2431 ( .A(n1908), .B(n18194), .Z(n1788) );
  NAND U2432 ( .A(n1786), .B(n18104), .Z(n1787) );
  AND U2433 ( .A(n1788), .B(n1787), .Z(n1897) );
  XNOR U2434 ( .A(n1896), .B(n1897), .Z(n1898) );
  NANDN U2435 ( .A(n1789), .B(n19013), .Z(n1791) );
  XNOR U2436 ( .A(b[21]), .B(a[3]), .Z(n1923) );
  NANDN U2437 ( .A(n1923), .B(n19015), .Z(n1790) );
  NAND U2438 ( .A(n1791), .B(n1790), .Z(n1900) );
  XNOR U2439 ( .A(b[23]), .B(n2921), .Z(n1794) );
  XNOR U2440 ( .A(b[23]), .B(n582), .Z(n1793) );
  XOR U2441 ( .A(b[23]), .B(b[22]), .Z(n1792) );
  AND U2442 ( .A(n1793), .B(n1792), .Z(n19128) );
  NAND U2443 ( .A(n1794), .B(n19128), .Z(n1796) );
  XOR U2444 ( .A(b[23]), .B(a[1]), .Z(n1920) );
  ANDN U2445 ( .B(n1920), .A(n19127), .Z(n1795) );
  ANDN U2446 ( .B(n1796), .A(n1795), .Z(n1901) );
  XNOR U2447 ( .A(n1900), .B(n1901), .Z(n1899) );
  XOR U2448 ( .A(n1898), .B(n1899), .Z(n1950) );
  XNOR U2449 ( .A(n1951), .B(n1950), .Z(n1952) );
  XNOR U2450 ( .A(n1953), .B(n1952), .Z(n1887) );
  NANDN U2451 ( .A(n1798), .B(n1797), .Z(n1802) );
  NAND U2452 ( .A(n1800), .B(n1799), .Z(n1801) );
  NAND U2453 ( .A(n1802), .B(n1801), .Z(n1885) );
  NANDN U2454 ( .A(n1804), .B(n1803), .Z(n1808) );
  NAND U2455 ( .A(n1806), .B(n1805), .Z(n1807) );
  AND U2456 ( .A(n1808), .B(n1807), .Z(n1884) );
  XNOR U2457 ( .A(n1885), .B(n1884), .Z(n1886) );
  XNOR U2458 ( .A(n1887), .B(n1886), .Z(n1965) );
  NANDN U2459 ( .A(n1810), .B(n1809), .Z(n1814) );
  NANDN U2460 ( .A(n1812), .B(n1811), .Z(n1813) );
  NAND U2461 ( .A(n1814), .B(n1813), .Z(n1878) );
  XOR U2462 ( .A(b[17]), .B(a[7]), .Z(n1935) );
  NAND U2463 ( .A(n1935), .B(n18673), .Z(n1817) );
  NAND U2464 ( .A(n1815), .B(n18674), .Z(n1816) );
  NAND U2465 ( .A(n1817), .B(n1816), .Z(n1893) );
  NANDN U2466 ( .A(n1818), .B(n18832), .Z(n1820) );
  XNOR U2467 ( .A(b[19]), .B(a[5]), .Z(n1917) );
  NANDN U2468 ( .A(n1917), .B(n18834), .Z(n1819) );
  NAND U2469 ( .A(n1820), .B(n1819), .Z(n1890) );
  XOR U2470 ( .A(n580), .B(n4573), .Z(n1905) );
  NAND U2471 ( .A(n1905), .B(n18336), .Z(n1823) );
  NANDN U2472 ( .A(n1821), .B(n18337), .Z(n1822) );
  AND U2473 ( .A(n1823), .B(n1822), .Z(n1891) );
  XNOR U2474 ( .A(n1890), .B(n1891), .Z(n1892) );
  XOR U2475 ( .A(n1893), .B(n1892), .Z(n1879) );
  XNOR U2476 ( .A(n1878), .B(n1879), .Z(n1880) );
  NANDN U2477 ( .A(n582), .B(b[22]), .Z(n19183) );
  AND U2478 ( .A(n19183), .B(b[23]), .Z(n19287) );
  XNOR U2479 ( .A(b[22]), .B(n582), .Z(n1824) );
  NANDN U2480 ( .A(n2921), .B(n1824), .Z(n1825) );
  AND U2481 ( .A(n19287), .B(n1825), .Z(n1939) );
  XNOR U2482 ( .A(b[3]), .B(a[21]), .Z(n1902) );
  NANDN U2483 ( .A(n1902), .B(n16990), .Z(n1828) );
  OR U2484 ( .A(n1826), .B(n16988), .Z(n1827) );
  AND U2485 ( .A(n1828), .B(n1827), .Z(n1938) );
  XNOR U2486 ( .A(n1939), .B(n1938), .Z(n1940) );
  XNOR U2487 ( .A(b[15]), .B(a[9]), .Z(n1911) );
  OR U2488 ( .A(n1911), .B(n18512), .Z(n1831) );
  NAND U2489 ( .A(n1829), .B(n18513), .Z(n1830) );
  AND U2490 ( .A(n1831), .B(n1830), .Z(n1941) );
  XNOR U2491 ( .A(n1940), .B(n1941), .Z(n1881) );
  XOR U2492 ( .A(n1880), .B(n1881), .Z(n1962) );
  NANDN U2493 ( .A(n1833), .B(n1832), .Z(n1837) );
  NANDN U2494 ( .A(n1835), .B(n1834), .Z(n1836) );
  NAND U2495 ( .A(n1837), .B(n1836), .Z(n1963) );
  XNOR U2496 ( .A(n1962), .B(n1963), .Z(n1964) );
  XNOR U2497 ( .A(n1965), .B(n1964), .Z(n1872) );
  NANDN U2498 ( .A(n1839), .B(n1838), .Z(n1843) );
  OR U2499 ( .A(n1841), .B(n1840), .Z(n1842) );
  NAND U2500 ( .A(n1843), .B(n1842), .Z(n1959) );
  NANDN U2501 ( .A(n1845), .B(n1844), .Z(n1849) );
  NANDN U2502 ( .A(n1847), .B(n1846), .Z(n1848) );
  NAND U2503 ( .A(n1849), .B(n1848), .Z(n1956) );
  NANDN U2504 ( .A(n1851), .B(n1850), .Z(n1855) );
  NANDN U2505 ( .A(n1853), .B(n1852), .Z(n1854) );
  NAND U2506 ( .A(n1855), .B(n1854), .Z(n1957) );
  XNOR U2507 ( .A(n1956), .B(n1957), .Z(n1958) );
  XNOR U2508 ( .A(n1959), .B(n1958), .Z(n1873) );
  XOR U2509 ( .A(n1872), .B(n1873), .Z(n1874) );
  XNOR U2510 ( .A(n1875), .B(n1874), .Z(n1867) );
  XNOR U2511 ( .A(n1866), .B(n1867), .Z(n1868) );
  XNOR U2512 ( .A(n1869), .B(n1868), .Z(n1861) );
  XNOR U2513 ( .A(n1861), .B(sreg[119]), .Z(n1863) );
  NAND U2514 ( .A(n1856), .B(sreg[118]), .Z(n1860) );
  OR U2515 ( .A(n1858), .B(n1857), .Z(n1859) );
  AND U2516 ( .A(n1860), .B(n1859), .Z(n1862) );
  XOR U2517 ( .A(n1863), .B(n1862), .Z(c[119]) );
  NAND U2518 ( .A(n1861), .B(sreg[119]), .Z(n1865) );
  OR U2519 ( .A(n1863), .B(n1862), .Z(n1864) );
  NAND U2520 ( .A(n1865), .B(n1864), .Z(n2079) );
  XNOR U2521 ( .A(n2079), .B(sreg[120]), .Z(n2081) );
  NANDN U2522 ( .A(n1867), .B(n1866), .Z(n1871) );
  NAND U2523 ( .A(n1869), .B(n1868), .Z(n1870) );
  NAND U2524 ( .A(n1871), .B(n1870), .Z(n1971) );
  OR U2525 ( .A(n1873), .B(n1872), .Z(n1877) );
  NAND U2526 ( .A(n1875), .B(n1874), .Z(n1876) );
  NAND U2527 ( .A(n1877), .B(n1876), .Z(n1968) );
  NANDN U2528 ( .A(n1879), .B(n1878), .Z(n1883) );
  NANDN U2529 ( .A(n1881), .B(n1880), .Z(n1882) );
  NAND U2530 ( .A(n1883), .B(n1882), .Z(n2076) );
  NANDN U2531 ( .A(n1885), .B(n1884), .Z(n1889) );
  NANDN U2532 ( .A(n1887), .B(n1886), .Z(n1888) );
  NAND U2533 ( .A(n1889), .B(n1888), .Z(n2070) );
  NANDN U2534 ( .A(n1891), .B(n1890), .Z(n1895) );
  NAND U2535 ( .A(n1893), .B(n1892), .Z(n1894) );
  NAND U2536 ( .A(n1895), .B(n1894), .Z(n1981) );
  XNOR U2537 ( .A(n1981), .B(n1980), .Z(n1982) );
  NANDN U2538 ( .A(n1901), .B(n1900), .Z(n2020) );
  XNOR U2539 ( .A(b[3]), .B(a[22]), .Z(n1998) );
  NANDN U2540 ( .A(n1998), .B(n16990), .Z(n1904) );
  OR U2541 ( .A(n1902), .B(n16988), .Z(n1903) );
  NAND U2542 ( .A(n1904), .B(n1903), .Z(n2019) );
  XNOR U2543 ( .A(b[13]), .B(a[12]), .Z(n2007) );
  NANDN U2544 ( .A(n2007), .B(n18336), .Z(n1907) );
  NAND U2545 ( .A(n18337), .B(n1905), .Z(n1906) );
  AND U2546 ( .A(n1907), .B(n1906), .Z(n2018) );
  XNOR U2547 ( .A(n2019), .B(n2018), .Z(n2021) );
  XNOR U2548 ( .A(n2020), .B(n2021), .Z(n1983) );
  XNOR U2549 ( .A(n1982), .B(n1983), .Z(n2067) );
  XOR U2550 ( .A(b[11]), .B(a[14]), .Z(n2052) );
  NANDN U2551 ( .A(n18194), .B(n2052), .Z(n1910) );
  NANDN U2552 ( .A(n1908), .B(n18104), .Z(n1909) );
  NAND U2553 ( .A(n1910), .B(n1909), .Z(n2028) );
  NANDN U2554 ( .A(n1911), .B(n18513), .Z(n1913) );
  XOR U2555 ( .A(b[15]), .B(a[10]), .Z(n2001) );
  NANDN U2556 ( .A(n18512), .B(n2001), .Z(n1912) );
  AND U2557 ( .A(n1913), .B(n1912), .Z(n2029) );
  XNOR U2558 ( .A(n2028), .B(n2029), .Z(n2030) );
  XNOR U2559 ( .A(b[9]), .B(a[16]), .Z(n2040) );
  NANDN U2560 ( .A(n2040), .B(n17814), .Z(n1916) );
  NANDN U2561 ( .A(n1914), .B(n17815), .Z(n1915) );
  NAND U2562 ( .A(n1916), .B(n1915), .Z(n2024) );
  NANDN U2563 ( .A(n1917), .B(n18832), .Z(n1919) );
  XNOR U2564 ( .A(b[19]), .B(a[6]), .Z(n2034) );
  NANDN U2565 ( .A(n2034), .B(n18834), .Z(n1918) );
  AND U2566 ( .A(n1919), .B(n1918), .Z(n2022) );
  XOR U2567 ( .A(b[23]), .B(a[2]), .Z(n2010) );
  NANDN U2568 ( .A(n19127), .B(n2010), .Z(n1922) );
  NAND U2569 ( .A(n1920), .B(n19128), .Z(n1921) );
  AND U2570 ( .A(n1922), .B(n1921), .Z(n2023) );
  XOR U2571 ( .A(n2024), .B(n2025), .Z(n2031) );
  XNOR U2572 ( .A(n2030), .B(n2031), .Z(n2063) );
  NANDN U2573 ( .A(n1923), .B(n19013), .Z(n1925) );
  XNOR U2574 ( .A(b[21]), .B(a[4]), .Z(n2037) );
  NANDN U2575 ( .A(n2037), .B(n19015), .Z(n1924) );
  NAND U2576 ( .A(n1925), .B(n1924), .Z(n1992) );
  XOR U2577 ( .A(b[24]), .B(b[23]), .Z(n19240) );
  NANDN U2578 ( .A(n2921), .B(n19240), .Z(n1997) );
  XNOR U2579 ( .A(n1992), .B(n1997), .Z(n1994) );
  NANDN U2580 ( .A(n577), .B(a[24]), .Z(n1926) );
  XOR U2581 ( .A(n17151), .B(n1926), .Z(n1928) );
  NANDN U2582 ( .A(b[0]), .B(a[23]), .Z(n1927) );
  AND U2583 ( .A(n1928), .B(n1927), .Z(n1993) );
  XOR U2584 ( .A(n1994), .B(n1993), .Z(n2061) );
  NAND U2585 ( .A(n1929), .B(n17553), .Z(n1931) );
  XOR U2586 ( .A(b[7]), .B(a[18]), .Z(n2043) );
  NAND U2587 ( .A(n2043), .B(n17555), .Z(n1930) );
  NAND U2588 ( .A(n1931), .B(n1930), .Z(n2058) );
  XOR U2589 ( .A(b[5]), .B(a[20]), .Z(n2046) );
  NAND U2590 ( .A(n2046), .B(n17310), .Z(n1934) );
  NAND U2591 ( .A(n1932), .B(n17311), .Z(n1933) );
  NAND U2592 ( .A(n1934), .B(n1933), .Z(n2055) );
  XOR U2593 ( .A(b[17]), .B(a[8]), .Z(n2049) );
  NAND U2594 ( .A(n2049), .B(n18673), .Z(n1937) );
  NAND U2595 ( .A(n1935), .B(n18674), .Z(n1936) );
  AND U2596 ( .A(n1937), .B(n1936), .Z(n2056) );
  XNOR U2597 ( .A(n2055), .B(n2056), .Z(n2057) );
  XOR U2598 ( .A(n2058), .B(n2057), .Z(n2062) );
  XNOR U2599 ( .A(n2061), .B(n2062), .Z(n2064) );
  XNOR U2600 ( .A(n2063), .B(n2064), .Z(n1989) );
  NANDN U2601 ( .A(n1939), .B(n1938), .Z(n1943) );
  NAND U2602 ( .A(n1941), .B(n1940), .Z(n1942) );
  NAND U2603 ( .A(n1943), .B(n1942), .Z(n1986) );
  NANDN U2604 ( .A(n1945), .B(n1944), .Z(n1949) );
  NAND U2605 ( .A(n1947), .B(n1946), .Z(n1948) );
  NAND U2606 ( .A(n1949), .B(n1948), .Z(n1987) );
  XNOR U2607 ( .A(n1986), .B(n1987), .Z(n1988) );
  XOR U2608 ( .A(n1989), .B(n1988), .Z(n2068) );
  XNOR U2609 ( .A(n2067), .B(n2068), .Z(n2069) );
  XNOR U2610 ( .A(n2070), .B(n2069), .Z(n2074) );
  NANDN U2611 ( .A(n1951), .B(n1950), .Z(n1955) );
  NANDN U2612 ( .A(n1953), .B(n1952), .Z(n1954) );
  AND U2613 ( .A(n1955), .B(n1954), .Z(n2073) );
  XNOR U2614 ( .A(n2074), .B(n2073), .Z(n2075) );
  XNOR U2615 ( .A(n2076), .B(n2075), .Z(n1977) );
  NANDN U2616 ( .A(n1957), .B(n1956), .Z(n1961) );
  NAND U2617 ( .A(n1959), .B(n1958), .Z(n1960) );
  NAND U2618 ( .A(n1961), .B(n1960), .Z(n1974) );
  NANDN U2619 ( .A(n1963), .B(n1962), .Z(n1967) );
  NANDN U2620 ( .A(n1965), .B(n1964), .Z(n1966) );
  NAND U2621 ( .A(n1967), .B(n1966), .Z(n1975) );
  XNOR U2622 ( .A(n1974), .B(n1975), .Z(n1976) );
  XOR U2623 ( .A(n1977), .B(n1976), .Z(n1969) );
  XNOR U2624 ( .A(n1968), .B(n1969), .Z(n1970) );
  XOR U2625 ( .A(n1971), .B(n1970), .Z(n2080) );
  XOR U2626 ( .A(n2081), .B(n2080), .Z(c[120]) );
  NANDN U2627 ( .A(n1969), .B(n1968), .Z(n1973) );
  NAND U2628 ( .A(n1971), .B(n1970), .Z(n1972) );
  NAND U2629 ( .A(n1973), .B(n1972), .Z(n2092) );
  NANDN U2630 ( .A(n1975), .B(n1974), .Z(n1979) );
  NANDN U2631 ( .A(n1977), .B(n1976), .Z(n1978) );
  NAND U2632 ( .A(n1979), .B(n1978), .Z(n2089) );
  NANDN U2633 ( .A(n1981), .B(n1980), .Z(n1985) );
  NANDN U2634 ( .A(n1983), .B(n1982), .Z(n1984) );
  NAND U2635 ( .A(n1985), .B(n1984), .Z(n2194) );
  NANDN U2636 ( .A(n1987), .B(n1986), .Z(n1991) );
  NANDN U2637 ( .A(n1989), .B(n1988), .Z(n1990) );
  AND U2638 ( .A(n1991), .B(n1990), .Z(n2195) );
  XNOR U2639 ( .A(n2194), .B(n2195), .Z(n2196) );
  NANDN U2640 ( .A(n1997), .B(n1992), .Z(n1996) );
  NAND U2641 ( .A(n1994), .B(n1993), .Z(n1995) );
  NAND U2642 ( .A(n1996), .B(n1995), .Z(n2191) );
  NAND U2643 ( .A(b[24]), .B(b[23]), .Z(n19271) );
  AND U2644 ( .A(n19271), .B(b[25]), .Z(n19381) );
  AND U2645 ( .A(n19381), .B(n1997), .Z(n2170) );
  XNOR U2646 ( .A(b[3]), .B(a[23]), .Z(n2136) );
  NANDN U2647 ( .A(n2136), .B(n16990), .Z(n2000) );
  OR U2648 ( .A(n1998), .B(n16988), .Z(n1999) );
  AND U2649 ( .A(n2000), .B(n1999), .Z(n2169) );
  XNOR U2650 ( .A(n2170), .B(n2169), .Z(n2171) );
  XNOR U2651 ( .A(b[15]), .B(a[11]), .Z(n2133) );
  OR U2652 ( .A(n2133), .B(n18512), .Z(n2003) );
  NAND U2653 ( .A(n2001), .B(n18513), .Z(n2002) );
  NAND U2654 ( .A(n2003), .B(n2002), .Z(n2172) );
  XOR U2655 ( .A(n2171), .B(n2172), .Z(n2189) );
  NANDN U2656 ( .A(n577), .B(a[25]), .Z(n2004) );
  XOR U2657 ( .A(n17151), .B(n2004), .Z(n2006) );
  NANDN U2658 ( .A(b[0]), .B(a[24]), .Z(n2005) );
  AND U2659 ( .A(n2006), .B(n2005), .Z(n2184) );
  XOR U2660 ( .A(b[13]), .B(n4875), .Z(n2142) );
  NANDN U2661 ( .A(n2142), .B(n18336), .Z(n2009) );
  NANDN U2662 ( .A(n2007), .B(n18337), .Z(n2008) );
  AND U2663 ( .A(n2009), .B(n2008), .Z(n2185) );
  XNOR U2664 ( .A(n2184), .B(n2185), .Z(n2186) );
  XOR U2665 ( .A(b[23]), .B(a[3]), .Z(n2166) );
  NANDN U2666 ( .A(n19127), .B(n2166), .Z(n2012) );
  NAND U2667 ( .A(n2010), .B(n19128), .Z(n2011) );
  NAND U2668 ( .A(n2012), .B(n2011), .Z(n2131) );
  XNOR U2669 ( .A(b[25]), .B(n2921), .Z(n2015) );
  XOR U2670 ( .A(b[25]), .B(b[23]), .Z(n2014) );
  XOR U2671 ( .A(b[25]), .B(b[24]), .Z(n2013) );
  AND U2672 ( .A(n2014), .B(n2013), .Z(n19242) );
  NAND U2673 ( .A(n2015), .B(n19242), .Z(n2017) );
  XOR U2674 ( .A(b[25]), .B(a[1]), .Z(n2181) );
  AND U2675 ( .A(n19240), .B(n2181), .Z(n2016) );
  ANDN U2676 ( .B(n2017), .A(n2016), .Z(n2132) );
  XNOR U2677 ( .A(n2131), .B(n2132), .Z(n2187) );
  XOR U2678 ( .A(n2186), .B(n2187), .Z(n2188) );
  XOR U2679 ( .A(n2189), .B(n2188), .Z(n2190) );
  XNOR U2680 ( .A(n2191), .B(n2190), .Z(n2116) );
  OR U2681 ( .A(n2023), .B(n2022), .Z(n2027) );
  NANDN U2682 ( .A(n2025), .B(n2024), .Z(n2026) );
  NAND U2683 ( .A(n2027), .B(n2026), .Z(n2114) );
  XNOR U2684 ( .A(n2113), .B(n2114), .Z(n2115) );
  XOR U2685 ( .A(n2116), .B(n2115), .Z(n2103) );
  NANDN U2686 ( .A(n2029), .B(n2028), .Z(n2033) );
  NANDN U2687 ( .A(n2031), .B(n2030), .Z(n2032) );
  NAND U2688 ( .A(n2033), .B(n2032), .Z(n2110) );
  NANDN U2689 ( .A(n2034), .B(n18832), .Z(n2036) );
  XNOR U2690 ( .A(b[19]), .B(a[7]), .Z(n2145) );
  NANDN U2691 ( .A(n2145), .B(n18834), .Z(n2035) );
  NAND U2692 ( .A(n2036), .B(n2035), .Z(n2151) );
  NANDN U2693 ( .A(n2037), .B(n19013), .Z(n2039) );
  XNOR U2694 ( .A(b[21]), .B(a[5]), .Z(n2178) );
  NANDN U2695 ( .A(n2178), .B(n19015), .Z(n2038) );
  NAND U2696 ( .A(n2039), .B(n2038), .Z(n2148) );
  XNOR U2697 ( .A(b[9]), .B(a[17]), .Z(n2157) );
  NANDN U2698 ( .A(n2157), .B(n17814), .Z(n2042) );
  NANDN U2699 ( .A(n2040), .B(n17815), .Z(n2041) );
  AND U2700 ( .A(n2042), .B(n2041), .Z(n2149) );
  XNOR U2701 ( .A(n2148), .B(n2149), .Z(n2150) );
  XNOR U2702 ( .A(n2151), .B(n2150), .Z(n2122) );
  NAND U2703 ( .A(n2043), .B(n17553), .Z(n2045) );
  XOR U2704 ( .A(b[7]), .B(a[19]), .Z(n2154) );
  NAND U2705 ( .A(n2154), .B(n17555), .Z(n2044) );
  NAND U2706 ( .A(n2045), .B(n2044), .Z(n2128) );
  XOR U2707 ( .A(b[5]), .B(a[21]), .Z(n2139) );
  NAND U2708 ( .A(n2139), .B(n17310), .Z(n2048) );
  NAND U2709 ( .A(n2046), .B(n17311), .Z(n2047) );
  NAND U2710 ( .A(n2048), .B(n2047), .Z(n2125) );
  XOR U2711 ( .A(b[17]), .B(a[9]), .Z(n2175) );
  NAND U2712 ( .A(n2175), .B(n18673), .Z(n2051) );
  NAND U2713 ( .A(n2049), .B(n18674), .Z(n2050) );
  AND U2714 ( .A(n2051), .B(n2050), .Z(n2126) );
  XNOR U2715 ( .A(n2125), .B(n2126), .Z(n2127) );
  XNOR U2716 ( .A(n2128), .B(n2127), .Z(n2119) );
  XNOR U2717 ( .A(b[11]), .B(a[15]), .Z(n2160) );
  OR U2718 ( .A(n2160), .B(n18194), .Z(n2054) );
  NAND U2719 ( .A(n18104), .B(n2052), .Z(n2053) );
  NAND U2720 ( .A(n2054), .B(n2053), .Z(n2120) );
  XNOR U2721 ( .A(n2119), .B(n2120), .Z(n2121) );
  XOR U2722 ( .A(n2122), .B(n2121), .Z(n2108) );
  NANDN U2723 ( .A(n2056), .B(n2055), .Z(n2060) );
  NAND U2724 ( .A(n2058), .B(n2057), .Z(n2059) );
  AND U2725 ( .A(n2060), .B(n2059), .Z(n2107) );
  XOR U2726 ( .A(n2108), .B(n2107), .Z(n2109) );
  XOR U2727 ( .A(n2110), .B(n2109), .Z(n2102) );
  OR U2728 ( .A(n2062), .B(n2061), .Z(n2066) );
  OR U2729 ( .A(n2064), .B(n2063), .Z(n2065) );
  AND U2730 ( .A(n2066), .B(n2065), .Z(n2101) );
  XNOR U2731 ( .A(n2102), .B(n2101), .Z(n2104) );
  XOR U2732 ( .A(n2103), .B(n2104), .Z(n2197) );
  XOR U2733 ( .A(n2196), .B(n2197), .Z(n2095) );
  NANDN U2734 ( .A(n2068), .B(n2067), .Z(n2072) );
  NAND U2735 ( .A(n2070), .B(n2069), .Z(n2071) );
  NAND U2736 ( .A(n2072), .B(n2071), .Z(n2096) );
  XNOR U2737 ( .A(n2095), .B(n2096), .Z(n2097) );
  NANDN U2738 ( .A(n2074), .B(n2073), .Z(n2078) );
  NAND U2739 ( .A(n2076), .B(n2075), .Z(n2077) );
  NAND U2740 ( .A(n2078), .B(n2077), .Z(n2098) );
  XNOR U2741 ( .A(n2097), .B(n2098), .Z(n2090) );
  XNOR U2742 ( .A(n2089), .B(n2090), .Z(n2091) );
  XNOR U2743 ( .A(n2092), .B(n2091), .Z(n2084) );
  XNOR U2744 ( .A(n2084), .B(sreg[121]), .Z(n2086) );
  NAND U2745 ( .A(n2079), .B(sreg[120]), .Z(n2083) );
  OR U2746 ( .A(n2081), .B(n2080), .Z(n2082) );
  AND U2747 ( .A(n2083), .B(n2082), .Z(n2085) );
  XOR U2748 ( .A(n2086), .B(n2085), .Z(c[121]) );
  NAND U2749 ( .A(n2084), .B(sreg[121]), .Z(n2088) );
  OR U2750 ( .A(n2086), .B(n2085), .Z(n2087) );
  NAND U2751 ( .A(n2088), .B(n2087), .Z(n2317) );
  XNOR U2752 ( .A(n2317), .B(sreg[122]), .Z(n2319) );
  NANDN U2753 ( .A(n2090), .B(n2089), .Z(n2094) );
  NAND U2754 ( .A(n2092), .B(n2091), .Z(n2093) );
  NAND U2755 ( .A(n2094), .B(n2093), .Z(n2203) );
  NANDN U2756 ( .A(n2096), .B(n2095), .Z(n2100) );
  NANDN U2757 ( .A(n2098), .B(n2097), .Z(n2099) );
  NAND U2758 ( .A(n2100), .B(n2099), .Z(n2201) );
  OR U2759 ( .A(n2102), .B(n2101), .Z(n2106) );
  NANDN U2760 ( .A(n2104), .B(n2103), .Z(n2105) );
  NAND U2761 ( .A(n2106), .B(n2105), .Z(n2209) );
  OR U2762 ( .A(n2108), .B(n2107), .Z(n2112) );
  NAND U2763 ( .A(n2110), .B(n2109), .Z(n2111) );
  NAND U2764 ( .A(n2112), .B(n2111), .Z(n2210) );
  NANDN U2765 ( .A(n2114), .B(n2113), .Z(n2118) );
  NAND U2766 ( .A(n2116), .B(n2115), .Z(n2117) );
  NAND U2767 ( .A(n2118), .B(n2117), .Z(n2211) );
  XNOR U2768 ( .A(n2210), .B(n2211), .Z(n2212) );
  NANDN U2769 ( .A(n2120), .B(n2119), .Z(n2124) );
  NAND U2770 ( .A(n2122), .B(n2121), .Z(n2123) );
  AND U2771 ( .A(n2124), .B(n2123), .Z(n2216) );
  NANDN U2772 ( .A(n2126), .B(n2125), .Z(n2130) );
  NAND U2773 ( .A(n2128), .B(n2127), .Z(n2129) );
  NAND U2774 ( .A(n2130), .B(n2129), .Z(n2241) );
  NANDN U2775 ( .A(n2132), .B(n2131), .Z(n2303) );
  XOR U2776 ( .A(b[15]), .B(a[12]), .Z(n2275) );
  NANDN U2777 ( .A(n18512), .B(n2275), .Z(n2135) );
  NANDN U2778 ( .A(n2133), .B(n18513), .Z(n2134) );
  NAND U2779 ( .A(n2135), .B(n2134), .Z(n2302) );
  XNOR U2780 ( .A(n578), .B(a[24]), .Z(n2272) );
  NAND U2781 ( .A(n16990), .B(n2272), .Z(n2138) );
  OR U2782 ( .A(n2136), .B(n16988), .Z(n2137) );
  AND U2783 ( .A(n2138), .B(n2137), .Z(n2301) );
  XNOR U2784 ( .A(n2302), .B(n2301), .Z(n2304) );
  XNOR U2785 ( .A(n2303), .B(n2304), .Z(n2238) );
  XOR U2786 ( .A(b[5]), .B(a[22]), .Z(n2295) );
  NAND U2787 ( .A(n2295), .B(n17310), .Z(n2141) );
  NAND U2788 ( .A(n2139), .B(n17311), .Z(n2140) );
  NAND U2789 ( .A(n2141), .B(n2140), .Z(n2247) );
  XNOR U2790 ( .A(n580), .B(a[14]), .Z(n2289) );
  NAND U2791 ( .A(n2289), .B(n18336), .Z(n2144) );
  NANDN U2792 ( .A(n2142), .B(n18337), .Z(n2143) );
  NAND U2793 ( .A(n2144), .B(n2143), .Z(n2244) );
  NANDN U2794 ( .A(n2145), .B(n18832), .Z(n2147) );
  XNOR U2795 ( .A(b[19]), .B(a[8]), .Z(n2298) );
  NANDN U2796 ( .A(n2298), .B(n18834), .Z(n2146) );
  AND U2797 ( .A(n2147), .B(n2146), .Z(n2245) );
  XNOR U2798 ( .A(n2244), .B(n2245), .Z(n2246) );
  XNOR U2799 ( .A(n2247), .B(n2246), .Z(n2239) );
  XNOR U2800 ( .A(n2238), .B(n2239), .Z(n2240) );
  XOR U2801 ( .A(n2241), .B(n2240), .Z(n2217) );
  XOR U2802 ( .A(n2216), .B(n2217), .Z(n2219) );
  NANDN U2803 ( .A(n2149), .B(n2148), .Z(n2153) );
  NAND U2804 ( .A(n2151), .B(n2150), .Z(n2152) );
  NAND U2805 ( .A(n2153), .B(n2152), .Z(n2234) );
  NAND U2806 ( .A(n2154), .B(n17553), .Z(n2156) );
  XOR U2807 ( .A(b[7]), .B(a[20]), .Z(n2292) );
  NAND U2808 ( .A(n2292), .B(n17555), .Z(n2155) );
  NAND U2809 ( .A(n2156), .B(n2155), .Z(n2308) );
  XNOR U2810 ( .A(b[9]), .B(a[18]), .Z(n2256) );
  NANDN U2811 ( .A(n2256), .B(n17814), .Z(n2159) );
  NANDN U2812 ( .A(n2157), .B(n17815), .Z(n2158) );
  NAND U2813 ( .A(n2159), .B(n2158), .Z(n2305) );
  XOR U2814 ( .A(b[11]), .B(a[16]), .Z(n2253) );
  NANDN U2815 ( .A(n18194), .B(n2253), .Z(n2162) );
  NANDN U2816 ( .A(n2160), .B(n18104), .Z(n2161) );
  AND U2817 ( .A(n2162), .B(n2161), .Z(n2306) );
  XNOR U2818 ( .A(n2305), .B(n2306), .Z(n2307) );
  XNOR U2819 ( .A(n2308), .B(n2307), .Z(n2232) );
  XOR U2820 ( .A(b[26]), .B(b[25]), .Z(n19336) );
  NAND U2821 ( .A(a[0]), .B(n19336), .Z(n2268) );
  NANDN U2822 ( .A(n577), .B(a[26]), .Z(n2163) );
  XOR U2823 ( .A(n17151), .B(n2163), .Z(n2165) );
  NANDN U2824 ( .A(b[0]), .B(a[25]), .Z(n2164) );
  AND U2825 ( .A(n2165), .B(n2164), .Z(n2266) );
  XOR U2826 ( .A(b[23]), .B(a[4]), .Z(n2262) );
  NANDN U2827 ( .A(n19127), .B(n2262), .Z(n2168) );
  NAND U2828 ( .A(n19128), .B(n2166), .Z(n2167) );
  AND U2829 ( .A(n2168), .B(n2167), .Z(n2265) );
  XNOR U2830 ( .A(n2266), .B(n2265), .Z(n2267) );
  XNOR U2831 ( .A(n2268), .B(n2267), .Z(n2233) );
  XOR U2832 ( .A(n2232), .B(n2233), .Z(n2235) );
  XOR U2833 ( .A(n2234), .B(n2235), .Z(n2218) );
  XOR U2834 ( .A(n2219), .B(n2218), .Z(n2224) );
  NANDN U2835 ( .A(n2170), .B(n2169), .Z(n2174) );
  NANDN U2836 ( .A(n2172), .B(n2171), .Z(n2173) );
  NAND U2837 ( .A(n2174), .B(n2173), .Z(n2231) );
  XOR U2838 ( .A(b[17]), .B(a[10]), .Z(n2250) );
  NAND U2839 ( .A(n2250), .B(n18673), .Z(n2177) );
  NAND U2840 ( .A(n2175), .B(n18674), .Z(n2176) );
  NAND U2841 ( .A(n2177), .B(n2176), .Z(n2314) );
  NANDN U2842 ( .A(n2178), .B(n19013), .Z(n2180) );
  XNOR U2843 ( .A(b[21]), .B(a[6]), .Z(n2259) );
  NANDN U2844 ( .A(n2259), .B(n19015), .Z(n2179) );
  NAND U2845 ( .A(n2180), .B(n2179), .Z(n2311) );
  XOR U2846 ( .A(b[25]), .B(a[2]), .Z(n2278) );
  NAND U2847 ( .A(n2278), .B(n19240), .Z(n2183) );
  NAND U2848 ( .A(n2181), .B(n19242), .Z(n2182) );
  AND U2849 ( .A(n2183), .B(n2182), .Z(n2312) );
  XNOR U2850 ( .A(n2311), .B(n2312), .Z(n2313) );
  XNOR U2851 ( .A(n2314), .B(n2313), .Z(n2228) );
  XNOR U2852 ( .A(n2228), .B(n2229), .Z(n2230) );
  XNOR U2853 ( .A(n2231), .B(n2230), .Z(n2222) );
  NAND U2854 ( .A(n2189), .B(n2188), .Z(n2193) );
  NAND U2855 ( .A(n2191), .B(n2190), .Z(n2192) );
  AND U2856 ( .A(n2193), .B(n2192), .Z(n2223) );
  XOR U2857 ( .A(n2222), .B(n2223), .Z(n2225) );
  XOR U2858 ( .A(n2224), .B(n2225), .Z(n2213) );
  XNOR U2859 ( .A(n2212), .B(n2213), .Z(n2206) );
  NANDN U2860 ( .A(n2195), .B(n2194), .Z(n2199) );
  NANDN U2861 ( .A(n2197), .B(n2196), .Z(n2198) );
  AND U2862 ( .A(n2199), .B(n2198), .Z(n2207) );
  XNOR U2863 ( .A(n2206), .B(n2207), .Z(n2208) );
  XOR U2864 ( .A(n2209), .B(n2208), .Z(n2200) );
  XNOR U2865 ( .A(n2201), .B(n2200), .Z(n2202) );
  XOR U2866 ( .A(n2203), .B(n2202), .Z(n2318) );
  XOR U2867 ( .A(n2319), .B(n2318), .Z(c[122]) );
  NANDN U2868 ( .A(n2201), .B(n2200), .Z(n2205) );
  NAND U2869 ( .A(n2203), .B(n2202), .Z(n2204) );
  NAND U2870 ( .A(n2205), .B(n2204), .Z(n2330) );
  NANDN U2871 ( .A(n2211), .B(n2210), .Z(n2215) );
  NAND U2872 ( .A(n2213), .B(n2212), .Z(n2214) );
  NAND U2873 ( .A(n2215), .B(n2214), .Z(n2334) );
  OR U2874 ( .A(n2217), .B(n2216), .Z(n2221) );
  NAND U2875 ( .A(n2219), .B(n2218), .Z(n2220) );
  NAND U2876 ( .A(n2221), .B(n2220), .Z(n2331) );
  NANDN U2877 ( .A(n2223), .B(n2222), .Z(n2227) );
  OR U2878 ( .A(n2225), .B(n2224), .Z(n2226) );
  NAND U2879 ( .A(n2227), .B(n2226), .Z(n2442) );
  NANDN U2880 ( .A(n2233), .B(n2232), .Z(n2237) );
  OR U2881 ( .A(n2235), .B(n2234), .Z(n2236) );
  NAND U2882 ( .A(n2237), .B(n2236), .Z(n2423) );
  NANDN U2883 ( .A(n2239), .B(n2238), .Z(n2243) );
  NAND U2884 ( .A(n2241), .B(n2240), .Z(n2242) );
  NAND U2885 ( .A(n2243), .B(n2242), .Z(n2424) );
  XNOR U2886 ( .A(n2423), .B(n2424), .Z(n2425) );
  XNOR U2887 ( .A(n2426), .B(n2425), .Z(n2439) );
  NANDN U2888 ( .A(n2245), .B(n2244), .Z(n2249) );
  NAND U2889 ( .A(n2247), .B(n2246), .Z(n2248) );
  NAND U2890 ( .A(n2249), .B(n2248), .Z(n2430) );
  XNOR U2891 ( .A(b[17]), .B(a[11]), .Z(n2417) );
  NANDN U2892 ( .A(n2417), .B(n18673), .Z(n2252) );
  NAND U2893 ( .A(n2250), .B(n18674), .Z(n2251) );
  NAND U2894 ( .A(n2252), .B(n2251), .Z(n2343) );
  XOR U2895 ( .A(b[11]), .B(a[17]), .Z(n2414) );
  NANDN U2896 ( .A(n18194), .B(n2414), .Z(n2255) );
  NAND U2897 ( .A(n2253), .B(n18104), .Z(n2254) );
  AND U2898 ( .A(n2255), .B(n2254), .Z(n2344) );
  XNOR U2899 ( .A(n2343), .B(n2344), .Z(n2345) );
  XNOR U2900 ( .A(b[9]), .B(a[19]), .Z(n2420) );
  NANDN U2901 ( .A(n2420), .B(n17814), .Z(n2258) );
  NANDN U2902 ( .A(n2256), .B(n17815), .Z(n2257) );
  NAND U2903 ( .A(n2258), .B(n2257), .Z(n2384) );
  NANDN U2904 ( .A(n2259), .B(n19013), .Z(n2261) );
  XNOR U2905 ( .A(b[21]), .B(a[7]), .Z(n2408) );
  NANDN U2906 ( .A(n2408), .B(n19015), .Z(n2260) );
  NAND U2907 ( .A(n2261), .B(n2260), .Z(n2381) );
  XOR U2908 ( .A(b[23]), .B(a[5]), .Z(n2399) );
  NANDN U2909 ( .A(n19127), .B(n2399), .Z(n2264) );
  NAND U2910 ( .A(n2262), .B(n19128), .Z(n2263) );
  AND U2911 ( .A(n2264), .B(n2263), .Z(n2382) );
  XNOR U2912 ( .A(n2381), .B(n2382), .Z(n2383) );
  XNOR U2913 ( .A(n2384), .B(n2383), .Z(n2346) );
  XOR U2914 ( .A(n2345), .B(n2346), .Z(n2340) );
  NANDN U2915 ( .A(n2266), .B(n2265), .Z(n2270) );
  NAND U2916 ( .A(n2268), .B(n2267), .Z(n2269) );
  NAND U2917 ( .A(n2270), .B(n2269), .Z(n2337) );
  NAND U2918 ( .A(b[26]), .B(b[25]), .Z(n19368) );
  ANDN U2919 ( .B(n19368), .A(n583), .Z(n19450) );
  NANDN U2920 ( .A(n2921), .B(n19336), .Z(n2271) );
  NAND U2921 ( .A(n19450), .B(n2271), .Z(n2372) );
  NANDN U2922 ( .A(n16988), .B(n2272), .Z(n2274) );
  XNOR U2923 ( .A(b[3]), .B(a[25]), .Z(n2396) );
  NANDN U2924 ( .A(n2396), .B(n16990), .Z(n2273) );
  NAND U2925 ( .A(n2274), .B(n2273), .Z(n2369) );
  NAND U2926 ( .A(n2275), .B(n18513), .Z(n2277) );
  XNOR U2927 ( .A(b[15]), .B(a[13]), .Z(n2364) );
  OR U2928 ( .A(n2364), .B(n18512), .Z(n2276) );
  AND U2929 ( .A(n2277), .B(n2276), .Z(n2370) );
  XNOR U2930 ( .A(n2369), .B(n2370), .Z(n2371) );
  XNOR U2931 ( .A(n2372), .B(n2371), .Z(n2338) );
  XNOR U2932 ( .A(n2337), .B(n2338), .Z(n2339) );
  XOR U2933 ( .A(n2340), .B(n2339), .Z(n2429) );
  XOR U2934 ( .A(n2430), .B(n2429), .Z(n2432) );
  XOR U2935 ( .A(b[25]), .B(a[3]), .Z(n2358) );
  NAND U2936 ( .A(n2358), .B(n19240), .Z(n2280) );
  NAND U2937 ( .A(n2278), .B(n19242), .Z(n2279) );
  NAND U2938 ( .A(n2280), .B(n2279), .Z(n2368) );
  XNOR U2939 ( .A(b[27]), .B(a[1]), .Z(n2361) );
  ANDN U2940 ( .B(n19336), .A(n2361), .Z(n2285) );
  XNOR U2941 ( .A(n583), .B(a[0]), .Z(n2283) );
  XNOR U2942 ( .A(n583), .B(b[25]), .Z(n2282) );
  XNOR U2943 ( .A(n583), .B(b[26]), .Z(n2281) );
  AND U2944 ( .A(n2282), .B(n2281), .Z(n19337) );
  NAND U2945 ( .A(n2283), .B(n19337), .Z(n2284) );
  NANDN U2946 ( .A(n2285), .B(n2284), .Z(n2367) );
  XNOR U2947 ( .A(n2368), .B(n2367), .Z(n2390) );
  NANDN U2948 ( .A(n577), .B(a[27]), .Z(n2286) );
  XOR U2949 ( .A(n17151), .B(n2286), .Z(n2288) );
  NANDN U2950 ( .A(b[0]), .B(a[26]), .Z(n2287) );
  AND U2951 ( .A(n2288), .B(n2287), .Z(n2388) );
  XOR U2952 ( .A(b[13]), .B(n5159), .Z(n2393) );
  NANDN U2953 ( .A(n2393), .B(n18336), .Z(n2291) );
  NAND U2954 ( .A(n18337), .B(n2289), .Z(n2290) );
  AND U2955 ( .A(n2291), .B(n2290), .Z(n2387) );
  XNOR U2956 ( .A(n2388), .B(n2387), .Z(n2389) );
  XOR U2957 ( .A(n2390), .B(n2389), .Z(n2375) );
  NAND U2958 ( .A(n2292), .B(n17553), .Z(n2294) );
  XOR U2959 ( .A(b[7]), .B(a[21]), .Z(n2411) );
  NAND U2960 ( .A(n2411), .B(n17555), .Z(n2293) );
  NAND U2961 ( .A(n2294), .B(n2293), .Z(n2352) );
  XOR U2962 ( .A(b[5]), .B(a[23]), .Z(n2402) );
  NAND U2963 ( .A(n2402), .B(n17310), .Z(n2297) );
  NAND U2964 ( .A(n2295), .B(n17311), .Z(n2296) );
  NAND U2965 ( .A(n2297), .B(n2296), .Z(n2349) );
  NANDN U2966 ( .A(n2298), .B(n18832), .Z(n2300) );
  XNOR U2967 ( .A(b[19]), .B(a[9]), .Z(n2405) );
  NANDN U2968 ( .A(n2405), .B(n18834), .Z(n2299) );
  AND U2969 ( .A(n2300), .B(n2299), .Z(n2350) );
  XNOR U2970 ( .A(n2349), .B(n2350), .Z(n2351) );
  XNOR U2971 ( .A(n2352), .B(n2351), .Z(n2376) );
  XOR U2972 ( .A(n2375), .B(n2376), .Z(n2377) );
  XOR U2973 ( .A(n2377), .B(n2378), .Z(n2438) );
  NANDN U2974 ( .A(n2306), .B(n2305), .Z(n2310) );
  NAND U2975 ( .A(n2308), .B(n2307), .Z(n2309) );
  NAND U2976 ( .A(n2310), .B(n2309), .Z(n2436) );
  NANDN U2977 ( .A(n2312), .B(n2311), .Z(n2316) );
  NAND U2978 ( .A(n2314), .B(n2313), .Z(n2315) );
  AND U2979 ( .A(n2316), .B(n2315), .Z(n2435) );
  XNOR U2980 ( .A(n2436), .B(n2435), .Z(n2437) );
  XOR U2981 ( .A(n2438), .B(n2437), .Z(n2431) );
  XOR U2982 ( .A(n2432), .B(n2431), .Z(n2440) );
  XNOR U2983 ( .A(n2439), .B(n2440), .Z(n2441) );
  XOR U2984 ( .A(n2442), .B(n2441), .Z(n2332) );
  XNOR U2985 ( .A(n2331), .B(n2332), .Z(n2333) );
  XNOR U2986 ( .A(n2334), .B(n2333), .Z(n2327) );
  XOR U2987 ( .A(n2328), .B(n2327), .Z(n2329) );
  XNOR U2988 ( .A(n2330), .B(n2329), .Z(n2322) );
  XNOR U2989 ( .A(n2322), .B(sreg[123]), .Z(n2324) );
  NAND U2990 ( .A(n2317), .B(sreg[122]), .Z(n2321) );
  OR U2991 ( .A(n2319), .B(n2318), .Z(n2320) );
  AND U2992 ( .A(n2321), .B(n2320), .Z(n2323) );
  XOR U2993 ( .A(n2324), .B(n2323), .Z(c[123]) );
  NAND U2994 ( .A(n2322), .B(sreg[123]), .Z(n2326) );
  OR U2995 ( .A(n2324), .B(n2323), .Z(n2325) );
  NAND U2996 ( .A(n2326), .B(n2325), .Z(n2576) );
  XNOR U2997 ( .A(n2576), .B(sreg[124]), .Z(n2578) );
  NANDN U2998 ( .A(n2332), .B(n2331), .Z(n2336) );
  NANDN U2999 ( .A(n2334), .B(n2333), .Z(n2335) );
  NAND U3000 ( .A(n2336), .B(n2335), .Z(n2445) );
  NANDN U3001 ( .A(n2338), .B(n2337), .Z(n2342) );
  NAND U3002 ( .A(n2340), .B(n2339), .Z(n2341) );
  NAND U3003 ( .A(n2342), .B(n2341), .Z(n2464) );
  NANDN U3004 ( .A(n2344), .B(n2343), .Z(n2348) );
  NANDN U3005 ( .A(n2346), .B(n2345), .Z(n2347) );
  NAND U3006 ( .A(n2348), .B(n2347), .Z(n2472) );
  NANDN U3007 ( .A(n2350), .B(n2349), .Z(n2354) );
  NAND U3008 ( .A(n2352), .B(n2351), .Z(n2353) );
  NAND U3009 ( .A(n2354), .B(n2353), .Z(n2567) );
  NANDN U3010 ( .A(n577), .B(a[28]), .Z(n2355) );
  XOR U3011 ( .A(n17151), .B(n2355), .Z(n2357) );
  NANDN U3012 ( .A(b[0]), .B(a[27]), .Z(n2356) );
  AND U3013 ( .A(n2357), .B(n2356), .Z(n2485) );
  AND U3014 ( .A(a[0]), .B(n575), .Z(n2539) );
  XOR U3015 ( .A(b[25]), .B(a[4]), .Z(n2478) );
  NAND U3016 ( .A(n2478), .B(n19240), .Z(n2360) );
  NAND U3017 ( .A(n2358), .B(n19242), .Z(n2359) );
  NAND U3018 ( .A(n2360), .B(n2359), .Z(n2484) );
  XNOR U3019 ( .A(n2539), .B(n2484), .Z(n2486) );
  XNOR U3020 ( .A(n2485), .B(n2486), .Z(n2565) );
  XNOR U3021 ( .A(b[27]), .B(a[2]), .Z(n2501) );
  NANDN U3022 ( .A(n2501), .B(n19336), .Z(n2363) );
  NANDN U3023 ( .A(n2361), .B(n19337), .Z(n2362) );
  NAND U3024 ( .A(n2363), .B(n2362), .Z(n2495) );
  NANDN U3025 ( .A(n2364), .B(n18513), .Z(n2366) );
  XOR U3026 ( .A(b[15]), .B(a[14]), .Z(n2511) );
  NANDN U3027 ( .A(n18512), .B(n2511), .Z(n2365) );
  AND U3028 ( .A(n2366), .B(n2365), .Z(n2496) );
  XNOR U3029 ( .A(n2495), .B(n2496), .Z(n2497) );
  NAND U3030 ( .A(n2368), .B(n2367), .Z(n2498) );
  XNOR U3031 ( .A(n2497), .B(n2498), .Z(n2564) );
  XOR U3032 ( .A(n2565), .B(n2564), .Z(n2566) );
  XOR U3033 ( .A(n2567), .B(n2566), .Z(n2469) );
  NANDN U3034 ( .A(n2370), .B(n2369), .Z(n2374) );
  NANDN U3035 ( .A(n2372), .B(n2371), .Z(n2373) );
  AND U3036 ( .A(n2374), .B(n2373), .Z(n2470) );
  XNOR U3037 ( .A(n2469), .B(n2470), .Z(n2471) );
  XOR U3038 ( .A(n2472), .B(n2471), .Z(n2463) );
  XOR U3039 ( .A(n2464), .B(n2463), .Z(n2466) );
  OR U3040 ( .A(n2376), .B(n2375), .Z(n2380) );
  NAND U3041 ( .A(n2378), .B(n2377), .Z(n2379) );
  NAND U3042 ( .A(n2380), .B(n2379), .Z(n2573) );
  NANDN U3043 ( .A(n2382), .B(n2381), .Z(n2386) );
  NAND U3044 ( .A(n2384), .B(n2383), .Z(n2385) );
  NAND U3045 ( .A(n2386), .B(n2385), .Z(n2561) );
  NANDN U3046 ( .A(n2388), .B(n2387), .Z(n2392) );
  NAND U3047 ( .A(n2390), .B(n2389), .Z(n2391) );
  NAND U3048 ( .A(n2392), .B(n2391), .Z(n2558) );
  XNOR U3049 ( .A(b[13]), .B(a[16]), .Z(n2514) );
  NANDN U3050 ( .A(n2514), .B(n18336), .Z(n2395) );
  NANDN U3051 ( .A(n2393), .B(n18337), .Z(n2394) );
  NAND U3052 ( .A(n2395), .B(n2394), .Z(n2526) );
  OR U3053 ( .A(n2396), .B(n16988), .Z(n2398) );
  XNOR U3054 ( .A(b[3]), .B(a[26]), .Z(n2532) );
  NANDN U3055 ( .A(n2532), .B(n16990), .Z(n2397) );
  NAND U3056 ( .A(n2398), .B(n2397), .Z(n2523) );
  XOR U3057 ( .A(b[23]), .B(a[6]), .Z(n2475) );
  NANDN U3058 ( .A(n19127), .B(n2475), .Z(n2401) );
  NAND U3059 ( .A(n2399), .B(n19128), .Z(n2400) );
  AND U3060 ( .A(n2401), .B(n2400), .Z(n2524) );
  XNOR U3061 ( .A(n2523), .B(n2524), .Z(n2525) );
  XOR U3062 ( .A(n2526), .B(n2525), .Z(n2559) );
  XNOR U3063 ( .A(n2558), .B(n2559), .Z(n2560) );
  XOR U3064 ( .A(n2561), .B(n2560), .Z(n2570) );
  XOR U3065 ( .A(b[5]), .B(a[24]), .Z(n2529) );
  NAND U3066 ( .A(n2529), .B(n17310), .Z(n2404) );
  NAND U3067 ( .A(n2402), .B(n17311), .Z(n2403) );
  NAND U3068 ( .A(n2404), .B(n2403), .Z(n2549) );
  NANDN U3069 ( .A(n2405), .B(n18832), .Z(n2407) );
  XNOR U3070 ( .A(b[19]), .B(a[10]), .Z(n2517) );
  NANDN U3071 ( .A(n2517), .B(n18834), .Z(n2406) );
  NAND U3072 ( .A(n2407), .B(n2406), .Z(n2546) );
  NANDN U3073 ( .A(n2408), .B(n19013), .Z(n2410) );
  XNOR U3074 ( .A(n582), .B(a[8]), .Z(n2543) );
  NAND U3075 ( .A(n2543), .B(n19015), .Z(n2409) );
  AND U3076 ( .A(n2410), .B(n2409), .Z(n2547) );
  XNOR U3077 ( .A(n2546), .B(n2547), .Z(n2548) );
  XNOR U3078 ( .A(n2549), .B(n2548), .Z(n2555) );
  NAND U3079 ( .A(n2411), .B(n17553), .Z(n2413) );
  XOR U3080 ( .A(b[7]), .B(a[22]), .Z(n2540) );
  NAND U3081 ( .A(n2540), .B(n17555), .Z(n2412) );
  NAND U3082 ( .A(n2413), .B(n2412), .Z(n2492) );
  XOR U3083 ( .A(b[11]), .B(a[18]), .Z(n2520) );
  NANDN U3084 ( .A(n18194), .B(n2520), .Z(n2416) );
  NAND U3085 ( .A(n2414), .B(n18104), .Z(n2415) );
  NAND U3086 ( .A(n2416), .B(n2415), .Z(n2489) );
  XOR U3087 ( .A(b[17]), .B(a[12]), .Z(n2535) );
  NAND U3088 ( .A(n2535), .B(n18673), .Z(n2419) );
  NANDN U3089 ( .A(n2417), .B(n18674), .Z(n2418) );
  AND U3090 ( .A(n2419), .B(n2418), .Z(n2490) );
  XNOR U3091 ( .A(n2489), .B(n2490), .Z(n2491) );
  XNOR U3092 ( .A(n2492), .B(n2491), .Z(n2552) );
  XNOR U3093 ( .A(b[9]), .B(a[20]), .Z(n2481) );
  NANDN U3094 ( .A(n2481), .B(n17814), .Z(n2422) );
  NANDN U3095 ( .A(n2420), .B(n17815), .Z(n2421) );
  NAND U3096 ( .A(n2422), .B(n2421), .Z(n2553) );
  XNOR U3097 ( .A(n2552), .B(n2553), .Z(n2554) );
  XOR U3098 ( .A(n2555), .B(n2554), .Z(n2571) );
  XNOR U3099 ( .A(n2570), .B(n2571), .Z(n2572) );
  XNOR U3100 ( .A(n2573), .B(n2572), .Z(n2465) );
  XNOR U3101 ( .A(n2466), .B(n2465), .Z(n2454) );
  NANDN U3102 ( .A(n2424), .B(n2423), .Z(n2428) );
  NAND U3103 ( .A(n2426), .B(n2425), .Z(n2427) );
  NAND U3104 ( .A(n2428), .B(n2427), .Z(n2460) );
  NANDN U3105 ( .A(n2430), .B(n2429), .Z(n2434) );
  OR U3106 ( .A(n2432), .B(n2431), .Z(n2433) );
  NAND U3107 ( .A(n2434), .B(n2433), .Z(n2458) );
  XNOR U3108 ( .A(n2458), .B(n2457), .Z(n2459) );
  XOR U3109 ( .A(n2460), .B(n2459), .Z(n2451) );
  NANDN U3110 ( .A(n2440), .B(n2439), .Z(n2444) );
  NAND U3111 ( .A(n2442), .B(n2441), .Z(n2443) );
  NAND U3112 ( .A(n2444), .B(n2443), .Z(n2452) );
  XNOR U3113 ( .A(n2451), .B(n2452), .Z(n2453) );
  XNOR U3114 ( .A(n2454), .B(n2453), .Z(n2446) );
  XNOR U3115 ( .A(n2445), .B(n2446), .Z(n2447) );
  XOR U3116 ( .A(n2448), .B(n2447), .Z(n2577) );
  XOR U3117 ( .A(n2578), .B(n2577), .Z(c[124]) );
  NANDN U3118 ( .A(n2446), .B(n2445), .Z(n2450) );
  NAND U3119 ( .A(n2448), .B(n2447), .Z(n2449) );
  NAND U3120 ( .A(n2450), .B(n2449), .Z(n2589) );
  NANDN U3121 ( .A(n2452), .B(n2451), .Z(n2456) );
  NAND U3122 ( .A(n2454), .B(n2453), .Z(n2455) );
  NAND U3123 ( .A(n2456), .B(n2455), .Z(n2586) );
  NANDN U3124 ( .A(n2458), .B(n2457), .Z(n2462) );
  NANDN U3125 ( .A(n2460), .B(n2459), .Z(n2461) );
  NAND U3126 ( .A(n2462), .B(n2461), .Z(n2712) );
  NANDN U3127 ( .A(n2464), .B(n2463), .Z(n2468) );
  OR U3128 ( .A(n2466), .B(n2465), .Z(n2467) );
  NAND U3129 ( .A(n2468), .B(n2467), .Z(n2709) );
  NANDN U3130 ( .A(n2470), .B(n2469), .Z(n2474) );
  NAND U3131 ( .A(n2472), .B(n2471), .Z(n2473) );
  NAND U3132 ( .A(n2474), .B(n2473), .Z(n2706) );
  XOR U3133 ( .A(b[23]), .B(a[7]), .Z(n2602) );
  NANDN U3134 ( .A(n19127), .B(n2602), .Z(n2477) );
  NAND U3135 ( .A(n2475), .B(n19128), .Z(n2476) );
  NAND U3136 ( .A(n2477), .B(n2476), .Z(n2620) );
  XOR U3137 ( .A(b[25]), .B(a[5]), .Z(n2605) );
  NAND U3138 ( .A(n2605), .B(n19240), .Z(n2480) );
  NAND U3139 ( .A(n2478), .B(n19242), .Z(n2479) );
  NAND U3140 ( .A(n2480), .B(n2479), .Z(n2617) );
  XNOR U3141 ( .A(b[9]), .B(a[21]), .Z(n2670) );
  NANDN U3142 ( .A(n2670), .B(n17814), .Z(n2483) );
  NANDN U3143 ( .A(n2481), .B(n17815), .Z(n2482) );
  AND U3144 ( .A(n2483), .B(n2482), .Z(n2618) );
  XNOR U3145 ( .A(n2617), .B(n2618), .Z(n2619) );
  XNOR U3146 ( .A(n2620), .B(n2619), .Z(n2641) );
  NAND U3147 ( .A(n2484), .B(n2539), .Z(n2488) );
  NANDN U3148 ( .A(n2486), .B(n2485), .Z(n2487) );
  NAND U3149 ( .A(n2488), .B(n2487), .Z(n2642) );
  XNOR U3150 ( .A(n2641), .B(n2642), .Z(n2643) );
  NANDN U3151 ( .A(n2490), .B(n2489), .Z(n2494) );
  NAND U3152 ( .A(n2492), .B(n2491), .Z(n2493) );
  AND U3153 ( .A(n2494), .B(n2493), .Z(n2644) );
  XNOR U3154 ( .A(n2643), .B(n2644), .Z(n2704) );
  NANDN U3155 ( .A(n2496), .B(n2495), .Z(n2500) );
  NANDN U3156 ( .A(n2498), .B(n2497), .Z(n2499) );
  NAND U3157 ( .A(n2500), .B(n2499), .Z(n2650) );
  XNOR U3158 ( .A(b[27]), .B(a[3]), .Z(n2599) );
  NANDN U3159 ( .A(n2599), .B(n19336), .Z(n2503) );
  NANDN U3160 ( .A(n2501), .B(n19337), .Z(n2502) );
  NAND U3161 ( .A(n2503), .B(n2502), .Z(n2654) );
  XNOR U3162 ( .A(b[29]), .B(a[1]), .Z(n2658) );
  NOR U3163 ( .A(n576), .B(n2658), .Z(n2507) );
  XNOR U3164 ( .A(n2921), .B(b[29]), .Z(n2505) );
  XOR U3165 ( .A(b[28]), .B(b[29]), .Z(n2504) );
  AND U3166 ( .A(n2504), .B(n576), .Z(n19406) );
  NAND U3167 ( .A(n2505), .B(n19406), .Z(n2506) );
  NANDN U3168 ( .A(n2507), .B(n2506), .Z(n2653) );
  XNOR U3169 ( .A(n2654), .B(n2653), .Z(n2688) );
  ANDN U3170 ( .B(a[29]), .A(n577), .Z(n2508) );
  XNOR U3171 ( .A(n17151), .B(n2508), .Z(n2510) );
  NANDN U3172 ( .A(b[0]), .B(a[28]), .Z(n2509) );
  NAND U3173 ( .A(n2510), .B(n2509), .Z(n2685) );
  XNOR U3174 ( .A(b[15]), .B(a[15]), .Z(n2661) );
  OR U3175 ( .A(n2661), .B(n18512), .Z(n2513) );
  NAND U3176 ( .A(n2511), .B(n18513), .Z(n2512) );
  NAND U3177 ( .A(n2513), .B(n2512), .Z(n2686) );
  XNOR U3178 ( .A(n2685), .B(n2686), .Z(n2687) );
  XOR U3179 ( .A(n2688), .B(n2687), .Z(n2647) );
  XNOR U3180 ( .A(b[13]), .B(a[17]), .Z(n2676) );
  NANDN U3181 ( .A(n2676), .B(n18336), .Z(n2516) );
  NANDN U3182 ( .A(n2514), .B(n18337), .Z(n2515) );
  NAND U3183 ( .A(n2516), .B(n2515), .Z(n2694) );
  NANDN U3184 ( .A(n2517), .B(n18832), .Z(n2519) );
  XOR U3185 ( .A(b[19]), .B(n4573), .Z(n2679) );
  NANDN U3186 ( .A(n2679), .B(n18834), .Z(n2518) );
  NAND U3187 ( .A(n2519), .B(n2518), .Z(n2691) );
  XOR U3188 ( .A(b[11]), .B(a[19]), .Z(n2673) );
  NANDN U3189 ( .A(n18194), .B(n2673), .Z(n2522) );
  NAND U3190 ( .A(n2520), .B(n18104), .Z(n2521) );
  AND U3191 ( .A(n2522), .B(n2521), .Z(n2692) );
  XNOR U3192 ( .A(n2691), .B(n2692), .Z(n2693) );
  XNOR U3193 ( .A(n2694), .B(n2693), .Z(n2648) );
  XOR U3194 ( .A(n2647), .B(n2648), .Z(n2649) );
  XNOR U3195 ( .A(n2650), .B(n2649), .Z(n2632) );
  NANDN U3196 ( .A(n2524), .B(n2523), .Z(n2528) );
  NAND U3197 ( .A(n2526), .B(n2525), .Z(n2527) );
  NAND U3198 ( .A(n2528), .B(n2527), .Z(n2629) );
  XOR U3199 ( .A(b[5]), .B(a[25]), .Z(n2664) );
  NAND U3200 ( .A(n2664), .B(n17310), .Z(n2531) );
  NAND U3201 ( .A(n2529), .B(n17311), .Z(n2530) );
  NAND U3202 ( .A(n2531), .B(n2530), .Z(n2614) );
  OR U3203 ( .A(n2532), .B(n16988), .Z(n2534) );
  XNOR U3204 ( .A(b[3]), .B(a[27]), .Z(n2667) );
  NANDN U3205 ( .A(n2667), .B(n16990), .Z(n2533) );
  NAND U3206 ( .A(n2534), .B(n2533), .Z(n2611) );
  XNOR U3207 ( .A(b[17]), .B(n4875), .Z(n2655) );
  NAND U3208 ( .A(n2655), .B(n18673), .Z(n2537) );
  NAND U3209 ( .A(n2535), .B(n18674), .Z(n2536) );
  AND U3210 ( .A(n2537), .B(n2536), .Z(n2612) );
  XNOR U3211 ( .A(n2611), .B(n2612), .Z(n2613) );
  XNOR U3212 ( .A(n2614), .B(n2613), .Z(n2592) );
  IV U3213 ( .A(b[28]), .Z(n19441) );
  NANDN U3214 ( .A(n19441), .B(b[27]), .Z(n2538) );
  AND U3215 ( .A(n2538), .B(b[29]), .Z(n19483) );
  XNOR U3216 ( .A(b[7]), .B(a[23]), .Z(n2682) );
  NANDN U3217 ( .A(n2682), .B(n17555), .Z(n2542) );
  NAND U3218 ( .A(n2540), .B(n17553), .Z(n2541) );
  NAND U3219 ( .A(n2542), .B(n2541), .Z(n2624) );
  XOR U3220 ( .A(n2623), .B(n2624), .Z(n2625) );
  XNOR U3221 ( .A(b[21]), .B(a[9]), .Z(n2608) );
  NANDN U3222 ( .A(n2608), .B(n19015), .Z(n2545) );
  NAND U3223 ( .A(n19013), .B(n2543), .Z(n2544) );
  AND U3224 ( .A(n2545), .B(n2544), .Z(n2626) );
  XNOR U3225 ( .A(n2625), .B(n2626), .Z(n2593) );
  XNOR U3226 ( .A(n2592), .B(n2593), .Z(n2594) );
  NANDN U3227 ( .A(n2547), .B(n2546), .Z(n2551) );
  NAND U3228 ( .A(n2549), .B(n2548), .Z(n2550) );
  AND U3229 ( .A(n2551), .B(n2550), .Z(n2595) );
  XNOR U3230 ( .A(n2594), .B(n2595), .Z(n2630) );
  XOR U3231 ( .A(n2629), .B(n2630), .Z(n2631) );
  XOR U3232 ( .A(n2632), .B(n2631), .Z(n2703) );
  XNOR U3233 ( .A(n2704), .B(n2703), .Z(n2705) );
  XOR U3234 ( .A(n2706), .B(n2705), .Z(n2700) );
  NANDN U3235 ( .A(n2553), .B(n2552), .Z(n2557) );
  NAND U3236 ( .A(n2555), .B(n2554), .Z(n2556) );
  NAND U3237 ( .A(n2557), .B(n2556), .Z(n2638) );
  NANDN U3238 ( .A(n2559), .B(n2558), .Z(n2563) );
  NANDN U3239 ( .A(n2561), .B(n2560), .Z(n2562) );
  NAND U3240 ( .A(n2563), .B(n2562), .Z(n2635) );
  OR U3241 ( .A(n2565), .B(n2564), .Z(n2569) );
  NANDN U3242 ( .A(n2567), .B(n2566), .Z(n2568) );
  AND U3243 ( .A(n2569), .B(n2568), .Z(n2636) );
  XNOR U3244 ( .A(n2635), .B(n2636), .Z(n2637) );
  XNOR U3245 ( .A(n2638), .B(n2637), .Z(n2697) );
  NANDN U3246 ( .A(n2571), .B(n2570), .Z(n2575) );
  NAND U3247 ( .A(n2573), .B(n2572), .Z(n2574) );
  AND U3248 ( .A(n2575), .B(n2574), .Z(n2698) );
  XNOR U3249 ( .A(n2697), .B(n2698), .Z(n2699) );
  XNOR U3250 ( .A(n2700), .B(n2699), .Z(n2710) );
  XNOR U3251 ( .A(n2709), .B(n2710), .Z(n2711) );
  XOR U3252 ( .A(n2712), .B(n2711), .Z(n2587) );
  XNOR U3253 ( .A(n2586), .B(n2587), .Z(n2588) );
  XNOR U3254 ( .A(n2589), .B(n2588), .Z(n2581) );
  XNOR U3255 ( .A(n2581), .B(sreg[125]), .Z(n2583) );
  NAND U3256 ( .A(n2576), .B(sreg[124]), .Z(n2580) );
  OR U3257 ( .A(n2578), .B(n2577), .Z(n2579) );
  AND U3258 ( .A(n2580), .B(n2579), .Z(n2582) );
  XOR U3259 ( .A(n2583), .B(n2582), .Z(c[125]) );
  NAND U3260 ( .A(n2581), .B(sreg[125]), .Z(n2585) );
  OR U3261 ( .A(n2583), .B(n2582), .Z(n2584) );
  NAND U3262 ( .A(n2585), .B(n2584), .Z(n2851) );
  XNOR U3263 ( .A(n2851), .B(sreg[126]), .Z(n2853) );
  NANDN U3264 ( .A(n2587), .B(n2586), .Z(n2591) );
  NAND U3265 ( .A(n2589), .B(n2588), .Z(n2590) );
  NAND U3266 ( .A(n2591), .B(n2590), .Z(n2718) );
  NANDN U3267 ( .A(n577), .B(a[30]), .Z(n2596) );
  XOR U3268 ( .A(n17151), .B(n2596), .Z(n2598) );
  IV U3269 ( .A(a[29]), .Z(n6835) );
  NANDN U3270 ( .A(n6835), .B(n577), .Z(n2597) );
  AND U3271 ( .A(n2598), .B(n2597), .Z(n2767) );
  XNOR U3272 ( .A(b[27]), .B(a[4]), .Z(n2839) );
  NANDN U3273 ( .A(n2839), .B(n19336), .Z(n2601) );
  NANDN U3274 ( .A(n2599), .B(n19337), .Z(n2600) );
  NAND U3275 ( .A(n2601), .B(n2600), .Z(n2765) );
  XNOR U3276 ( .A(n584), .B(b[30]), .Z(n19472) );
  NANDN U3277 ( .A(n2921), .B(n19472), .Z(n2766) );
  XNOR U3278 ( .A(n2765), .B(n2766), .Z(n2768) );
  XOR U3279 ( .A(n2767), .B(n2768), .Z(n2783) );
  XOR U3280 ( .A(b[23]), .B(a[8]), .Z(n2833) );
  NANDN U3281 ( .A(n19127), .B(n2833), .Z(n2604) );
  NAND U3282 ( .A(n2602), .B(n19128), .Z(n2603) );
  NAND U3283 ( .A(n2604), .B(n2603), .Z(n2815) );
  XOR U3284 ( .A(b[25]), .B(a[6]), .Z(n2836) );
  NAND U3285 ( .A(n2836), .B(n19240), .Z(n2607) );
  NAND U3286 ( .A(n2605), .B(n19242), .Z(n2606) );
  NAND U3287 ( .A(n2607), .B(n2606), .Z(n2812) );
  NANDN U3288 ( .A(n2608), .B(n19013), .Z(n2610) );
  XNOR U3289 ( .A(b[21]), .B(a[10]), .Z(n2830) );
  NANDN U3290 ( .A(n2830), .B(n19015), .Z(n2609) );
  AND U3291 ( .A(n2610), .B(n2609), .Z(n2813) );
  XNOR U3292 ( .A(n2812), .B(n2813), .Z(n2814) );
  XNOR U3293 ( .A(n2815), .B(n2814), .Z(n2781) );
  NANDN U3294 ( .A(n2612), .B(n2611), .Z(n2616) );
  NAND U3295 ( .A(n2614), .B(n2613), .Z(n2615) );
  NAND U3296 ( .A(n2616), .B(n2615), .Z(n2782) );
  XOR U3297 ( .A(n2781), .B(n2782), .Z(n2784) );
  XOR U3298 ( .A(n2783), .B(n2784), .Z(n2736) );
  NANDN U3299 ( .A(n2618), .B(n2617), .Z(n2622) );
  NAND U3300 ( .A(n2620), .B(n2619), .Z(n2621) );
  NAND U3301 ( .A(n2622), .B(n2621), .Z(n2733) );
  OR U3302 ( .A(n2624), .B(n2623), .Z(n2628) );
  NAND U3303 ( .A(n2626), .B(n2625), .Z(n2627) );
  NAND U3304 ( .A(n2628), .B(n2627), .Z(n2734) );
  XNOR U3305 ( .A(n2733), .B(n2734), .Z(n2735) );
  XOR U3306 ( .A(n2736), .B(n2735), .Z(n2728) );
  XOR U3307 ( .A(n2727), .B(n2728), .Z(n2729) );
  OR U3308 ( .A(n2630), .B(n2629), .Z(n2634) );
  NAND U3309 ( .A(n2632), .B(n2631), .Z(n2633) );
  NAND U3310 ( .A(n2634), .B(n2633), .Z(n2730) );
  XOR U3311 ( .A(n2729), .B(n2730), .Z(n2724) );
  NANDN U3312 ( .A(n2636), .B(n2635), .Z(n2640) );
  NAND U3313 ( .A(n2638), .B(n2637), .Z(n2639) );
  NAND U3314 ( .A(n2640), .B(n2639), .Z(n2721) );
  NANDN U3315 ( .A(n2642), .B(n2641), .Z(n2646) );
  NAND U3316 ( .A(n2644), .B(n2643), .Z(n2645) );
  NAND U3317 ( .A(n2646), .B(n2645), .Z(n2774) );
  OR U3318 ( .A(n2648), .B(n2647), .Z(n2652) );
  NAND U3319 ( .A(n2650), .B(n2649), .Z(n2651) );
  NAND U3320 ( .A(n2652), .B(n2651), .Z(n2771) );
  NAND U3321 ( .A(n2654), .B(n2653), .Z(n2804) );
  XOR U3322 ( .A(b[17]), .B(a[14]), .Z(n2799) );
  NAND U3323 ( .A(n18673), .B(n2799), .Z(n2657) );
  NAND U3324 ( .A(n18674), .B(n2655), .Z(n2656) );
  NAND U3325 ( .A(n2657), .B(n2656), .Z(n2803) );
  NANDN U3326 ( .A(n2658), .B(n19406), .Z(n2660) );
  XNOR U3327 ( .A(n584), .B(a[2]), .Z(n2751) );
  NANDN U3328 ( .A(n576), .B(n2751), .Z(n2659) );
  AND U3329 ( .A(n2660), .B(n2659), .Z(n2802) );
  XNOR U3330 ( .A(n2803), .B(n2802), .Z(n2805) );
  XNOR U3331 ( .A(n2804), .B(n2805), .Z(n2777) );
  NANDN U3332 ( .A(n2661), .B(n18513), .Z(n2663) );
  XOR U3333 ( .A(b[15]), .B(a[16]), .Z(n2762) );
  NANDN U3334 ( .A(n18512), .B(n2762), .Z(n2662) );
  NAND U3335 ( .A(n2663), .B(n2662), .Z(n2821) );
  XOR U3336 ( .A(b[5]), .B(a[26]), .Z(n2790) );
  NAND U3337 ( .A(n2790), .B(n17310), .Z(n2666) );
  NAND U3338 ( .A(n2664), .B(n17311), .Z(n2665) );
  NAND U3339 ( .A(n2666), .B(n2665), .Z(n2818) );
  OR U3340 ( .A(n2667), .B(n16988), .Z(n2669) );
  XNOR U3341 ( .A(b[3]), .B(a[28]), .Z(n2796) );
  NANDN U3342 ( .A(n2796), .B(n16990), .Z(n2668) );
  AND U3343 ( .A(n2669), .B(n2668), .Z(n2819) );
  XNOR U3344 ( .A(n2818), .B(n2819), .Z(n2820) );
  XNOR U3345 ( .A(n2821), .B(n2820), .Z(n2778) );
  XNOR U3346 ( .A(n2777), .B(n2778), .Z(n2779) );
  XNOR U3347 ( .A(b[9]), .B(a[22]), .Z(n2824) );
  NANDN U3348 ( .A(n2824), .B(n17814), .Z(n2672) );
  NANDN U3349 ( .A(n2670), .B(n17815), .Z(n2671) );
  NAND U3350 ( .A(n2672), .B(n2671), .Z(n2806) );
  XOR U3351 ( .A(b[11]), .B(a[20]), .Z(n2842) );
  NANDN U3352 ( .A(n18194), .B(n2842), .Z(n2675) );
  NAND U3353 ( .A(n2673), .B(n18104), .Z(n2674) );
  AND U3354 ( .A(n2675), .B(n2674), .Z(n2807) );
  XNOR U3355 ( .A(n2806), .B(n2807), .Z(n2808) );
  XNOR U3356 ( .A(b[13]), .B(a[18]), .Z(n2827) );
  NANDN U3357 ( .A(n2827), .B(n18336), .Z(n2678) );
  NANDN U3358 ( .A(n2676), .B(n18337), .Z(n2677) );
  NAND U3359 ( .A(n2678), .B(n2677), .Z(n2748) );
  NANDN U3360 ( .A(n2679), .B(n18832), .Z(n2681) );
  XNOR U3361 ( .A(b[19]), .B(a[12]), .Z(n2793) );
  NANDN U3362 ( .A(n2793), .B(n18834), .Z(n2680) );
  NAND U3363 ( .A(n2681), .B(n2680), .Z(n2745) );
  NANDN U3364 ( .A(n2682), .B(n17553), .Z(n2684) );
  XOR U3365 ( .A(b[7]), .B(a[24]), .Z(n2787) );
  NAND U3366 ( .A(n2787), .B(n17555), .Z(n2683) );
  AND U3367 ( .A(n2684), .B(n2683), .Z(n2746) );
  XNOR U3368 ( .A(n2745), .B(n2746), .Z(n2747) );
  XOR U3369 ( .A(n2748), .B(n2747), .Z(n2809) );
  XOR U3370 ( .A(n2808), .B(n2809), .Z(n2780) );
  XOR U3371 ( .A(n2779), .B(n2780), .Z(n2742) );
  NANDN U3372 ( .A(n2686), .B(n2685), .Z(n2690) );
  NAND U3373 ( .A(n2688), .B(n2687), .Z(n2689) );
  NAND U3374 ( .A(n2690), .B(n2689), .Z(n2739) );
  NANDN U3375 ( .A(n2692), .B(n2691), .Z(n2696) );
  NAND U3376 ( .A(n2694), .B(n2693), .Z(n2695) );
  NAND U3377 ( .A(n2696), .B(n2695), .Z(n2740) );
  XNOR U3378 ( .A(n2739), .B(n2740), .Z(n2741) );
  XOR U3379 ( .A(n2742), .B(n2741), .Z(n2772) );
  XOR U3380 ( .A(n2771), .B(n2772), .Z(n2773) );
  XNOR U3381 ( .A(n2774), .B(n2773), .Z(n2722) );
  XNOR U3382 ( .A(n2721), .B(n2722), .Z(n2723) );
  XNOR U3383 ( .A(n2724), .B(n2723), .Z(n2848) );
  NANDN U3384 ( .A(n2698), .B(n2697), .Z(n2702) );
  NAND U3385 ( .A(n2700), .B(n2699), .Z(n2701) );
  NAND U3386 ( .A(n2702), .B(n2701), .Z(n2845) );
  NANDN U3387 ( .A(n2704), .B(n2703), .Z(n2708) );
  NANDN U3388 ( .A(n2706), .B(n2705), .Z(n2707) );
  NAND U3389 ( .A(n2708), .B(n2707), .Z(n2846) );
  XNOR U3390 ( .A(n2845), .B(n2846), .Z(n2847) );
  XOR U3391 ( .A(n2848), .B(n2847), .Z(n2715) );
  NANDN U3392 ( .A(n2710), .B(n2709), .Z(n2714) );
  NAND U3393 ( .A(n2712), .B(n2711), .Z(n2713) );
  NAND U3394 ( .A(n2714), .B(n2713), .Z(n2716) );
  XOR U3395 ( .A(n2715), .B(n2716), .Z(n2717) );
  XOR U3396 ( .A(n2718), .B(n2717), .Z(n2852) );
  XOR U3397 ( .A(n2853), .B(n2852), .Z(c[126]) );
  OR U3398 ( .A(n2716), .B(n2715), .Z(n2720) );
  NAND U3399 ( .A(n2718), .B(n2717), .Z(n2719) );
  NAND U3400 ( .A(n2720), .B(n2719), .Z(n2864) );
  NANDN U3401 ( .A(n2722), .B(n2721), .Z(n2726) );
  NAND U3402 ( .A(n2724), .B(n2723), .Z(n2725) );
  NAND U3403 ( .A(n2726), .B(n2725), .Z(n2999) );
  OR U3404 ( .A(n2728), .B(n2727), .Z(n2732) );
  NANDN U3405 ( .A(n2730), .B(n2729), .Z(n2731) );
  NAND U3406 ( .A(n2732), .B(n2731), .Z(n2997) );
  NANDN U3407 ( .A(n2734), .B(n2733), .Z(n2738) );
  NANDN U3408 ( .A(n2736), .B(n2735), .Z(n2737) );
  NAND U3409 ( .A(n2738), .B(n2737), .Z(n2876) );
  NANDN U3410 ( .A(n2740), .B(n2739), .Z(n2744) );
  NANDN U3411 ( .A(n2742), .B(n2741), .Z(n2743) );
  NAND U3412 ( .A(n2744), .B(n2743), .Z(n2874) );
  NANDN U3413 ( .A(n2746), .B(n2745), .Z(n2750) );
  NAND U3414 ( .A(n2748), .B(n2747), .Z(n2749) );
  NAND U3415 ( .A(n2750), .B(n2749), .Z(n2894) );
  NAND U3416 ( .A(n2751), .B(n19406), .Z(n2753) );
  XNOR U3417 ( .A(n584), .B(a[3]), .Z(n2915) );
  NANDN U3418 ( .A(n576), .B(n2915), .Z(n2752) );
  NAND U3419 ( .A(n2753), .B(n2752), .Z(n2980) );
  XNOR U3420 ( .A(n585), .B(a[0]), .Z(n2756) );
  XNOR U3421 ( .A(n585), .B(b[29]), .Z(n2755) );
  XNOR U3422 ( .A(n585), .B(b[30]), .Z(n2754) );
  AND U3423 ( .A(n2755), .B(n2754), .Z(n19473) );
  NAND U3424 ( .A(n2756), .B(n19473), .Z(n2758) );
  XNOR U3425 ( .A(n585), .B(a[1]), .Z(n2990) );
  NAND U3426 ( .A(n2990), .B(n19472), .Z(n2757) );
  NAND U3427 ( .A(n2758), .B(n2757), .Z(n2979) );
  XNOR U3428 ( .A(n2980), .B(n2979), .Z(n2912) );
  NANDN U3429 ( .A(n577), .B(a[31]), .Z(n2759) );
  XOR U3430 ( .A(n17151), .B(n2759), .Z(n2761) );
  IV U3431 ( .A(a[30]), .Z(n7336) );
  NANDN U3432 ( .A(n7336), .B(n577), .Z(n2760) );
  AND U3433 ( .A(n2761), .B(n2760), .Z(n2910) );
  XNOR U3434 ( .A(b[15]), .B(a[17]), .Z(n2928) );
  OR U3435 ( .A(n2928), .B(n18512), .Z(n2764) );
  NAND U3436 ( .A(n2762), .B(n18513), .Z(n2763) );
  AND U3437 ( .A(n2764), .B(n2763), .Z(n2909) );
  XNOR U3438 ( .A(n2910), .B(n2909), .Z(n2911) );
  XOR U3439 ( .A(n2912), .B(n2911), .Z(n2892) );
  NANDN U3440 ( .A(n2766), .B(n2765), .Z(n2770) );
  NAND U3441 ( .A(n2768), .B(n2767), .Z(n2769) );
  AND U3442 ( .A(n2770), .B(n2769), .Z(n2891) );
  XOR U3443 ( .A(n2892), .B(n2891), .Z(n2893) );
  XOR U3444 ( .A(n2894), .B(n2893), .Z(n2873) );
  XNOR U3445 ( .A(n2874), .B(n2873), .Z(n2875) );
  XNOR U3446 ( .A(n2876), .B(n2875), .Z(n2870) );
  OR U3447 ( .A(n2772), .B(n2771), .Z(n2776) );
  NAND U3448 ( .A(n2774), .B(n2773), .Z(n2775) );
  NAND U3449 ( .A(n2776), .B(n2775), .Z(n2867) );
  NANDN U3450 ( .A(n2782), .B(n2781), .Z(n2786) );
  OR U3451 ( .A(n2784), .B(n2783), .Z(n2785) );
  NAND U3452 ( .A(n2786), .B(n2785), .Z(n2880) );
  XNOR U3453 ( .A(n2879), .B(n2880), .Z(n2881) );
  NAND U3454 ( .A(n2787), .B(n17553), .Z(n2789) );
  XOR U3455 ( .A(b[7]), .B(a[25]), .Z(n2958) );
  NAND U3456 ( .A(n2958), .B(n17555), .Z(n2788) );
  NAND U3457 ( .A(n2789), .B(n2788), .Z(n2976) );
  XOR U3458 ( .A(b[5]), .B(a[27]), .Z(n2961) );
  NAND U3459 ( .A(n2961), .B(n17310), .Z(n2792) );
  NAND U3460 ( .A(n2790), .B(n17311), .Z(n2791) );
  NAND U3461 ( .A(n2792), .B(n2791), .Z(n2973) );
  NANDN U3462 ( .A(n2793), .B(n18832), .Z(n2795) );
  XOR U3463 ( .A(b[19]), .B(n4875), .Z(n2964) );
  NANDN U3464 ( .A(n2964), .B(n18834), .Z(n2794) );
  AND U3465 ( .A(n2795), .B(n2794), .Z(n2974) );
  XNOR U3466 ( .A(n2973), .B(n2974), .Z(n2975) );
  XNOR U3467 ( .A(n2976), .B(n2975), .Z(n2898) );
  OR U3468 ( .A(n2796), .B(n16988), .Z(n2798) );
  XOR U3469 ( .A(b[3]), .B(n6835), .Z(n2984) );
  NANDN U3470 ( .A(n2984), .B(n16990), .Z(n2797) );
  NAND U3471 ( .A(n2798), .B(n2797), .Z(n2906) );
  XNOR U3472 ( .A(b[17]), .B(n5159), .Z(n2981) );
  NAND U3473 ( .A(n2981), .B(n18673), .Z(n2801) );
  NAND U3474 ( .A(n2799), .B(n18674), .Z(n2800) );
  NAND U3475 ( .A(n2801), .B(n2800), .Z(n2903) );
  XNOR U3476 ( .A(n2903), .B(n2904), .Z(n2905) );
  XOR U3477 ( .A(n2906), .B(n2905), .Z(n2897) );
  XNOR U3478 ( .A(n2898), .B(n2897), .Z(n2899) );
  XNOR U3479 ( .A(n2899), .B(n2900), .Z(n2886) );
  NANDN U3480 ( .A(n2807), .B(n2806), .Z(n2811) );
  NAND U3481 ( .A(n2809), .B(n2808), .Z(n2810) );
  NAND U3482 ( .A(n2811), .B(n2810), .Z(n2940) );
  NANDN U3483 ( .A(n2813), .B(n2812), .Z(n2817) );
  NAND U3484 ( .A(n2815), .B(n2814), .Z(n2816) );
  NAND U3485 ( .A(n2817), .B(n2816), .Z(n2937) );
  NANDN U3486 ( .A(n2819), .B(n2818), .Z(n2823) );
  NAND U3487 ( .A(n2821), .B(n2820), .Z(n2822) );
  AND U3488 ( .A(n2823), .B(n2822), .Z(n2938) );
  XNOR U3489 ( .A(n2937), .B(n2938), .Z(n2939) );
  XNOR U3490 ( .A(n2940), .B(n2939), .Z(n2885) );
  XNOR U3491 ( .A(n2886), .B(n2885), .Z(n2888) );
  XNOR U3492 ( .A(b[9]), .B(a[23]), .Z(n2987) );
  NANDN U3493 ( .A(n2987), .B(n17814), .Z(n2826) );
  NANDN U3494 ( .A(n2824), .B(n17815), .Z(n2825) );
  NAND U3495 ( .A(n2826), .B(n2825), .Z(n2934) );
  XNOR U3496 ( .A(b[13]), .B(a[19]), .Z(n2922) );
  NANDN U3497 ( .A(n2922), .B(n18336), .Z(n2829) );
  NANDN U3498 ( .A(n2827), .B(n18337), .Z(n2828) );
  NAND U3499 ( .A(n2829), .B(n2828), .Z(n2931) );
  NANDN U3500 ( .A(n2830), .B(n19013), .Z(n2832) );
  XOR U3501 ( .A(b[21]), .B(n4573), .Z(n2925) );
  NANDN U3502 ( .A(n2925), .B(n19015), .Z(n2831) );
  AND U3503 ( .A(n2832), .B(n2831), .Z(n2932) );
  XNOR U3504 ( .A(n2931), .B(n2932), .Z(n2933) );
  XNOR U3505 ( .A(n2934), .B(n2933), .Z(n2946) );
  XOR U3506 ( .A(b[23]), .B(a[9]), .Z(n2993) );
  NANDN U3507 ( .A(n19127), .B(n2993), .Z(n2835) );
  NAND U3508 ( .A(n2833), .B(n19128), .Z(n2834) );
  NAND U3509 ( .A(n2835), .B(n2834), .Z(n2970) );
  XOR U3510 ( .A(b[25]), .B(a[7]), .Z(n2952) );
  NAND U3511 ( .A(n2952), .B(n19240), .Z(n2838) );
  NAND U3512 ( .A(n2836), .B(n19242), .Z(n2837) );
  NAND U3513 ( .A(n2838), .B(n2837), .Z(n2967) );
  XNOR U3514 ( .A(b[27]), .B(a[5]), .Z(n2955) );
  NANDN U3515 ( .A(n2955), .B(n19336), .Z(n2841) );
  NANDN U3516 ( .A(n2839), .B(n19337), .Z(n2840) );
  AND U3517 ( .A(n2841), .B(n2840), .Z(n2968) );
  XNOR U3518 ( .A(n2967), .B(n2968), .Z(n2969) );
  XNOR U3519 ( .A(n2970), .B(n2969), .Z(n2943) );
  XOR U3520 ( .A(b[11]), .B(a[21]), .Z(n2949) );
  NANDN U3521 ( .A(n18194), .B(n2949), .Z(n2844) );
  NAND U3522 ( .A(n18104), .B(n2842), .Z(n2843) );
  NAND U3523 ( .A(n2844), .B(n2843), .Z(n2944) );
  XNOR U3524 ( .A(n2943), .B(n2944), .Z(n2945) );
  XOR U3525 ( .A(n2946), .B(n2945), .Z(n2887) );
  XNOR U3526 ( .A(n2888), .B(n2887), .Z(n2882) );
  XOR U3527 ( .A(n2881), .B(n2882), .Z(n2868) );
  XOR U3528 ( .A(n2867), .B(n2868), .Z(n2869) );
  XNOR U3529 ( .A(n2870), .B(n2869), .Z(n2996) );
  XNOR U3530 ( .A(n2997), .B(n2996), .Z(n2998) );
  XNOR U3531 ( .A(n2999), .B(n2998), .Z(n2861) );
  NANDN U3532 ( .A(n2846), .B(n2845), .Z(n2850) );
  NAND U3533 ( .A(n2848), .B(n2847), .Z(n2849) );
  NAND U3534 ( .A(n2850), .B(n2849), .Z(n2862) );
  XNOR U3535 ( .A(n2861), .B(n2862), .Z(n2863) );
  XNOR U3536 ( .A(n2864), .B(n2863), .Z(n2856) );
  XNOR U3537 ( .A(n2856), .B(sreg[127]), .Z(n2858) );
  NAND U3538 ( .A(n2851), .B(sreg[126]), .Z(n2855) );
  OR U3539 ( .A(n2853), .B(n2852), .Z(n2854) );
  AND U3540 ( .A(n2855), .B(n2854), .Z(n2857) );
  XOR U3541 ( .A(n2858), .B(n2857), .Z(c[127]) );
  NAND U3542 ( .A(n2856), .B(sreg[127]), .Z(n2860) );
  OR U3543 ( .A(n2858), .B(n2857), .Z(n2859) );
  NAND U3544 ( .A(n2860), .B(n2859), .Z(n3143) );
  XNOR U3545 ( .A(n3143), .B(sreg[128]), .Z(n3145) );
  NANDN U3546 ( .A(n2862), .B(n2861), .Z(n2866) );
  NAND U3547 ( .A(n2864), .B(n2863), .Z(n2865) );
  NAND U3548 ( .A(n2866), .B(n2865), .Z(n3005) );
  OR U3549 ( .A(n2868), .B(n2867), .Z(n2872) );
  NANDN U3550 ( .A(n2870), .B(n2869), .Z(n2871) );
  NAND U3551 ( .A(n2872), .B(n2871), .Z(n3140) );
  NANDN U3552 ( .A(n2874), .B(n2873), .Z(n2878) );
  NAND U3553 ( .A(n2876), .B(n2875), .Z(n2877) );
  NAND U3554 ( .A(n2878), .B(n2877), .Z(n3138) );
  NANDN U3555 ( .A(n2880), .B(n2879), .Z(n2884) );
  NANDN U3556 ( .A(n2882), .B(n2881), .Z(n2883) );
  NAND U3557 ( .A(n2884), .B(n2883), .Z(n3102) );
  OR U3558 ( .A(n2886), .B(n2885), .Z(n2890) );
  OR U3559 ( .A(n2888), .B(n2887), .Z(n2889) );
  AND U3560 ( .A(n2890), .B(n2889), .Z(n3103) );
  XNOR U3561 ( .A(n3102), .B(n3103), .Z(n3104) );
  OR U3562 ( .A(n2892), .B(n2891), .Z(n2896) );
  NAND U3563 ( .A(n2894), .B(n2893), .Z(n2895) );
  NAND U3564 ( .A(n2896), .B(n2895), .Z(n3132) );
  NANDN U3565 ( .A(n2898), .B(n2897), .Z(n2902) );
  NAND U3566 ( .A(n2900), .B(n2899), .Z(n2901) );
  NAND U3567 ( .A(n2902), .B(n2901), .Z(n3131) );
  NANDN U3568 ( .A(n2904), .B(n2903), .Z(n2908) );
  NAND U3569 ( .A(n2906), .B(n2905), .Z(n2907) );
  NAND U3570 ( .A(n2908), .B(n2907), .Z(n3114) );
  NANDN U3571 ( .A(n2910), .B(n2909), .Z(n2914) );
  NAND U3572 ( .A(n2912), .B(n2911), .Z(n2913) );
  NAND U3573 ( .A(n2914), .B(n2913), .Z(n3115) );
  XNOR U3574 ( .A(n3114), .B(n3115), .Z(n3116) );
  NAND U3575 ( .A(n19406), .B(n2915), .Z(n2917) );
  XNOR U3576 ( .A(n584), .B(a[4]), .Z(n3026) );
  NANDN U3577 ( .A(n576), .B(n3026), .Z(n2916) );
  AND U3578 ( .A(n2917), .B(n2916), .Z(n3042) );
  NANDN U3579 ( .A(n577), .B(a[32]), .Z(n2918) );
  XOR U3580 ( .A(n17151), .B(n2918), .Z(n2920) );
  NANDN U3581 ( .A(b[0]), .B(a[31]), .Z(n2919) );
  AND U3582 ( .A(n2920), .B(n2919), .Z(n3041) );
  XOR U3583 ( .A(n3042), .B(n3041), .Z(n3044) );
  NANDN U3584 ( .A(n2921), .B(b[31]), .Z(n3043) );
  XOR U3585 ( .A(n3044), .B(n3043), .Z(n3008) );
  XNOR U3586 ( .A(n580), .B(a[20]), .Z(n3087) );
  NAND U3587 ( .A(n3087), .B(n18336), .Z(n2924) );
  NANDN U3588 ( .A(n2922), .B(n18337), .Z(n2923) );
  NAND U3589 ( .A(n2924), .B(n2923), .Z(n3054) );
  NANDN U3590 ( .A(n2925), .B(n19013), .Z(n2927) );
  XNOR U3591 ( .A(b[21]), .B(a[12]), .Z(n3014) );
  NANDN U3592 ( .A(n3014), .B(n19015), .Z(n2926) );
  NAND U3593 ( .A(n2927), .B(n2926), .Z(n3051) );
  NANDN U3594 ( .A(n2928), .B(n18513), .Z(n2930) );
  XOR U3595 ( .A(b[15]), .B(a[18]), .Z(n3023) );
  NANDN U3596 ( .A(n18512), .B(n3023), .Z(n2929) );
  AND U3597 ( .A(n2930), .B(n2929), .Z(n3052) );
  XNOR U3598 ( .A(n3051), .B(n3052), .Z(n3053) );
  XNOR U3599 ( .A(n3054), .B(n3053), .Z(n3009) );
  XOR U3600 ( .A(n3008), .B(n3009), .Z(n3011) );
  NANDN U3601 ( .A(n2932), .B(n2931), .Z(n2936) );
  NAND U3602 ( .A(n2934), .B(n2933), .Z(n2935) );
  AND U3603 ( .A(n2936), .B(n2935), .Z(n3010) );
  XOR U3604 ( .A(n3011), .B(n3010), .Z(n3117) );
  XOR U3605 ( .A(n3116), .B(n3117), .Z(n3130) );
  XNOR U3606 ( .A(n3131), .B(n3130), .Z(n3133) );
  XNOR U3607 ( .A(n3132), .B(n3133), .Z(n3110) );
  NANDN U3608 ( .A(n2938), .B(n2937), .Z(n2942) );
  NAND U3609 ( .A(n2940), .B(n2939), .Z(n2941) );
  NAND U3610 ( .A(n2942), .B(n2941), .Z(n3108) );
  NANDN U3611 ( .A(n2944), .B(n2943), .Z(n2948) );
  NAND U3612 ( .A(n2946), .B(n2945), .Z(n2947) );
  NAND U3613 ( .A(n2948), .B(n2947), .Z(n3099) );
  XOR U3614 ( .A(b[11]), .B(a[22]), .Z(n3063) );
  NANDN U3615 ( .A(n18194), .B(n3063), .Z(n2951) );
  NAND U3616 ( .A(n2949), .B(n18104), .Z(n2950) );
  NAND U3617 ( .A(n2951), .B(n2950), .Z(n3093) );
  XOR U3618 ( .A(b[25]), .B(a[8]), .Z(n3084) );
  NAND U3619 ( .A(n3084), .B(n19240), .Z(n2954) );
  NAND U3620 ( .A(n2952), .B(n19242), .Z(n2953) );
  NAND U3621 ( .A(n2954), .B(n2953), .Z(n3090) );
  XNOR U3622 ( .A(b[27]), .B(a[6]), .Z(n3075) );
  NANDN U3623 ( .A(n3075), .B(n19336), .Z(n2957) );
  NANDN U3624 ( .A(n2955), .B(n19337), .Z(n2956) );
  AND U3625 ( .A(n2957), .B(n2956), .Z(n3091) );
  XNOR U3626 ( .A(n3090), .B(n3091), .Z(n3092) );
  XNOR U3627 ( .A(n3093), .B(n3092), .Z(n3120) );
  NAND U3628 ( .A(n2958), .B(n17553), .Z(n2960) );
  XOR U3629 ( .A(b[7]), .B(a[26]), .Z(n3066) );
  NAND U3630 ( .A(n3066), .B(n17555), .Z(n2959) );
  NAND U3631 ( .A(n2960), .B(n2959), .Z(n3032) );
  XOR U3632 ( .A(b[5]), .B(a[28]), .Z(n3069) );
  NAND U3633 ( .A(n3069), .B(n17310), .Z(n2963) );
  NAND U3634 ( .A(n2961), .B(n17311), .Z(n2962) );
  NAND U3635 ( .A(n2963), .B(n2962), .Z(n3029) );
  NANDN U3636 ( .A(n2964), .B(n18832), .Z(n2966) );
  XNOR U3637 ( .A(b[19]), .B(a[14]), .Z(n3020) );
  NANDN U3638 ( .A(n3020), .B(n18834), .Z(n2965) );
  AND U3639 ( .A(n2966), .B(n2965), .Z(n3030) );
  XNOR U3640 ( .A(n3029), .B(n3030), .Z(n3031) );
  XOR U3641 ( .A(n3032), .B(n3031), .Z(n3121) );
  XNOR U3642 ( .A(n3120), .B(n3121), .Z(n3122) );
  NANDN U3643 ( .A(n2968), .B(n2967), .Z(n2972) );
  NAND U3644 ( .A(n2970), .B(n2969), .Z(n2971) );
  AND U3645 ( .A(n2972), .B(n2971), .Z(n3123) );
  XNOR U3646 ( .A(n3122), .B(n3123), .Z(n3096) );
  NANDN U3647 ( .A(n2974), .B(n2973), .Z(n2978) );
  NAND U3648 ( .A(n2976), .B(n2975), .Z(n2977) );
  NAND U3649 ( .A(n2978), .B(n2977), .Z(n3127) );
  NAND U3650 ( .A(n2980), .B(n2979), .Z(n3049) );
  XOR U3651 ( .A(b[17]), .B(a[16]), .Z(n3072) );
  NAND U3652 ( .A(n18673), .B(n3072), .Z(n2983) );
  NAND U3653 ( .A(n18674), .B(n2981), .Z(n2982) );
  NAND U3654 ( .A(n2983), .B(n2982), .Z(n3048) );
  XOR U3655 ( .A(b[3]), .B(n7336), .Z(n3057) );
  NANDN U3656 ( .A(n3057), .B(n16990), .Z(n2986) );
  OR U3657 ( .A(n2984), .B(n16988), .Z(n2985) );
  AND U3658 ( .A(n2986), .B(n2985), .Z(n3047) );
  XNOR U3659 ( .A(n3048), .B(n3047), .Z(n3050) );
  XNOR U3660 ( .A(n3049), .B(n3050), .Z(n3124) );
  XNOR U3661 ( .A(n579), .B(a[24]), .Z(n3060) );
  NAND U3662 ( .A(n17814), .B(n3060), .Z(n2989) );
  NANDN U3663 ( .A(n2987), .B(n17815), .Z(n2988) );
  NAND U3664 ( .A(n2989), .B(n2988), .Z(n3038) );
  XNOR U3665 ( .A(b[31]), .B(a[2]), .Z(n3078) );
  NANDN U3666 ( .A(n3078), .B(n19472), .Z(n2992) );
  NAND U3667 ( .A(n2990), .B(n19473), .Z(n2991) );
  NAND U3668 ( .A(n2992), .B(n2991), .Z(n3035) );
  XOR U3669 ( .A(b[23]), .B(a[10]), .Z(n3017) );
  NANDN U3670 ( .A(n19127), .B(n3017), .Z(n2995) );
  NAND U3671 ( .A(n2993), .B(n19128), .Z(n2994) );
  AND U3672 ( .A(n2995), .B(n2994), .Z(n3036) );
  XNOR U3673 ( .A(n3035), .B(n3036), .Z(n3037) );
  XNOR U3674 ( .A(n3038), .B(n3037), .Z(n3125) );
  XNOR U3675 ( .A(n3124), .B(n3125), .Z(n3126) );
  XNOR U3676 ( .A(n3127), .B(n3126), .Z(n3097) );
  XNOR U3677 ( .A(n3096), .B(n3097), .Z(n3098) );
  XOR U3678 ( .A(n3099), .B(n3098), .Z(n3109) );
  XNOR U3679 ( .A(n3108), .B(n3109), .Z(n3111) );
  XOR U3680 ( .A(n3110), .B(n3111), .Z(n3105) );
  XOR U3681 ( .A(n3104), .B(n3105), .Z(n3137) );
  XOR U3682 ( .A(n3138), .B(n3137), .Z(n3139) );
  XNOR U3683 ( .A(n3140), .B(n3139), .Z(n3002) );
  NAND U3684 ( .A(n2997), .B(n2996), .Z(n3001) );
  OR U3685 ( .A(n2999), .B(n2998), .Z(n3000) );
  NAND U3686 ( .A(n3001), .B(n3000), .Z(n3003) );
  XNOR U3687 ( .A(n3002), .B(n3003), .Z(n3004) );
  XOR U3688 ( .A(n3005), .B(n3004), .Z(n3144) );
  XOR U3689 ( .A(n3145), .B(n3144), .Z(c[128]) );
  NANDN U3690 ( .A(n3003), .B(n3002), .Z(n3007) );
  NAND U3691 ( .A(n3005), .B(n3004), .Z(n3006) );
  NAND U3692 ( .A(n3007), .B(n3006), .Z(n3151) );
  NANDN U3693 ( .A(n3009), .B(n3008), .Z(n3013) );
  OR U3694 ( .A(n3011), .B(n3010), .Z(n3012) );
  NAND U3695 ( .A(n3013), .B(n3012), .Z(n3159) );
  NANDN U3696 ( .A(n3014), .B(n19013), .Z(n3016) );
  XOR U3697 ( .A(n582), .B(n4875), .Z(n3231) );
  NAND U3698 ( .A(n3231), .B(n19015), .Z(n3015) );
  NAND U3699 ( .A(n3016), .B(n3015), .Z(n3264) );
  XNOR U3700 ( .A(b[23]), .B(a[11]), .Z(n3246) );
  OR U3701 ( .A(n3246), .B(n19127), .Z(n3019) );
  NAND U3702 ( .A(n3017), .B(n19128), .Z(n3018) );
  NAND U3703 ( .A(n3019), .B(n3018), .Z(n3261) );
  NANDN U3704 ( .A(n3020), .B(n18832), .Z(n3022) );
  XOR U3705 ( .A(b[19]), .B(n5159), .Z(n3204) );
  NANDN U3706 ( .A(n3204), .B(n18834), .Z(n3021) );
  AND U3707 ( .A(n3022), .B(n3021), .Z(n3262) );
  XNOR U3708 ( .A(n3261), .B(n3262), .Z(n3263) );
  XNOR U3709 ( .A(n3264), .B(n3263), .Z(n3167) );
  NAND U3710 ( .A(n3023), .B(n18513), .Z(n3025) );
  XOR U3711 ( .A(b[15]), .B(a[19]), .Z(n3228) );
  NANDN U3712 ( .A(n18512), .B(n3228), .Z(n3024) );
  NAND U3713 ( .A(n3025), .B(n3024), .Z(n3192) );
  NAND U3714 ( .A(n19406), .B(n3026), .Z(n3028) );
  XNOR U3715 ( .A(n584), .B(a[5]), .Z(n3243) );
  NANDN U3716 ( .A(n576), .B(n3243), .Z(n3027) );
  NAND U3717 ( .A(n3028), .B(n3027), .Z(n3189) );
  NANDN U3718 ( .A(n585), .B(a[1]), .Z(n3190) );
  XNOR U3719 ( .A(n3189), .B(n3190), .Z(n3191) );
  XOR U3720 ( .A(n3192), .B(n3191), .Z(n3168) );
  XNOR U3721 ( .A(n3167), .B(n3168), .Z(n3169) );
  NANDN U3722 ( .A(n3030), .B(n3029), .Z(n3034) );
  NAND U3723 ( .A(n3032), .B(n3031), .Z(n3033) );
  NAND U3724 ( .A(n3034), .B(n3033), .Z(n3170) );
  XOR U3725 ( .A(n3169), .B(n3170), .Z(n3222) );
  NANDN U3726 ( .A(n3036), .B(n3035), .Z(n3040) );
  NAND U3727 ( .A(n3038), .B(n3037), .Z(n3039) );
  NAND U3728 ( .A(n3040), .B(n3039), .Z(n3219) );
  NANDN U3729 ( .A(n3042), .B(n3041), .Z(n3046) );
  OR U3730 ( .A(n3044), .B(n3043), .Z(n3045) );
  AND U3731 ( .A(n3046), .B(n3045), .Z(n3220) );
  XNOR U3732 ( .A(n3219), .B(n3220), .Z(n3221) );
  XNOR U3733 ( .A(n3222), .B(n3221), .Z(n3276) );
  NANDN U3734 ( .A(n3052), .B(n3051), .Z(n3056) );
  NAND U3735 ( .A(n3054), .B(n3053), .Z(n3055) );
  NAND U3736 ( .A(n3056), .B(n3055), .Z(n3216) );
  XNOR U3737 ( .A(b[3]), .B(a[31]), .Z(n3201) );
  NANDN U3738 ( .A(n3201), .B(n16990), .Z(n3059) );
  OR U3739 ( .A(n3057), .B(n16988), .Z(n3058) );
  NAND U3740 ( .A(n3059), .B(n3058), .Z(n3187) );
  XNOR U3741 ( .A(b[9]), .B(a[25]), .Z(n3225) );
  NANDN U3742 ( .A(n3225), .B(n17814), .Z(n3062) );
  NAND U3743 ( .A(n17815), .B(n3060), .Z(n3061) );
  NAND U3744 ( .A(n3062), .B(n3061), .Z(n3185) );
  XNOR U3745 ( .A(b[11]), .B(a[23]), .Z(n3234) );
  OR U3746 ( .A(n3234), .B(n18194), .Z(n3065) );
  NAND U3747 ( .A(n18104), .B(n3063), .Z(n3064) );
  NAND U3748 ( .A(n3065), .B(n3064), .Z(n3186) );
  XNOR U3749 ( .A(n3185), .B(n3186), .Z(n3188) );
  XOR U3750 ( .A(n3187), .B(n3188), .Z(n3176) );
  XNOR U3751 ( .A(b[7]), .B(a[27]), .Z(n3249) );
  NANDN U3752 ( .A(n3249), .B(n17555), .Z(n3068) );
  NAND U3753 ( .A(n3066), .B(n17553), .Z(n3067) );
  NAND U3754 ( .A(n3068), .B(n3067), .Z(n3174) );
  XNOR U3755 ( .A(b[5]), .B(a[29]), .Z(n3210) );
  NANDN U3756 ( .A(n3210), .B(n17310), .Z(n3071) );
  NAND U3757 ( .A(n17311), .B(n3069), .Z(n3070) );
  AND U3758 ( .A(n3071), .B(n3070), .Z(n3173) );
  XNOR U3759 ( .A(n3174), .B(n3173), .Z(n3175) );
  XNOR U3760 ( .A(n3176), .B(n3175), .Z(n3269) );
  XOR U3761 ( .A(b[17]), .B(a[17]), .Z(n3195) );
  NAND U3762 ( .A(n3195), .B(n18673), .Z(n3074) );
  NAND U3763 ( .A(n3072), .B(n18674), .Z(n3073) );
  NAND U3764 ( .A(n3074), .B(n3073), .Z(n3182) );
  XNOR U3765 ( .A(b[27]), .B(a[7]), .Z(n3207) );
  NANDN U3766 ( .A(n3207), .B(n19336), .Z(n3077) );
  NANDN U3767 ( .A(n3075), .B(n19337), .Z(n3076) );
  NAND U3768 ( .A(n3077), .B(n3076), .Z(n3179) );
  XNOR U3769 ( .A(b[31]), .B(a[3]), .Z(n3198) );
  NANDN U3770 ( .A(n3198), .B(n19472), .Z(n3080) );
  NANDN U3771 ( .A(n3078), .B(n19473), .Z(n3079) );
  AND U3772 ( .A(n3080), .B(n3079), .Z(n3180) );
  XNOR U3773 ( .A(n3179), .B(n3180), .Z(n3181) );
  XNOR U3774 ( .A(n3182), .B(n3181), .Z(n3267) );
  NANDN U3775 ( .A(n577), .B(a[33]), .Z(n3081) );
  XOR U3776 ( .A(n17151), .B(n3081), .Z(n3083) );
  NANDN U3777 ( .A(b[0]), .B(a[32]), .Z(n3082) );
  AND U3778 ( .A(n3083), .B(n3082), .Z(n3256) );
  XOR U3779 ( .A(b[25]), .B(a[9]), .Z(n3252) );
  NAND U3780 ( .A(n19240), .B(n3252), .Z(n3086) );
  NAND U3781 ( .A(n19242), .B(n3084), .Z(n3085) );
  AND U3782 ( .A(n3086), .B(n3085), .Z(n3255) );
  XNOR U3783 ( .A(n3256), .B(n3255), .Z(n3257) );
  XOR U3784 ( .A(n580), .B(a[21]), .Z(n3237) );
  NANDN U3785 ( .A(n3237), .B(n18336), .Z(n3089) );
  NAND U3786 ( .A(n18337), .B(n3087), .Z(n3088) );
  AND U3787 ( .A(n3089), .B(n3088), .Z(n3258) );
  XNOR U3788 ( .A(n3257), .B(n3258), .Z(n3268) );
  XOR U3789 ( .A(n3267), .B(n3268), .Z(n3270) );
  XOR U3790 ( .A(n3269), .B(n3270), .Z(n3213) );
  NANDN U3791 ( .A(n3091), .B(n3090), .Z(n3095) );
  NAND U3792 ( .A(n3093), .B(n3092), .Z(n3094) );
  AND U3793 ( .A(n3095), .B(n3094), .Z(n3214) );
  XOR U3794 ( .A(n3216), .B(n3215), .Z(n3274) );
  XNOR U3795 ( .A(n3273), .B(n3274), .Z(n3275) );
  XOR U3796 ( .A(n3276), .B(n3275), .Z(n3158) );
  XOR U3797 ( .A(n3159), .B(n3158), .Z(n3161) );
  NANDN U3798 ( .A(n3097), .B(n3096), .Z(n3101) );
  NANDN U3799 ( .A(n3099), .B(n3098), .Z(n3100) );
  NAND U3800 ( .A(n3101), .B(n3100), .Z(n3160) );
  XNOR U3801 ( .A(n3161), .B(n3160), .Z(n3155) );
  NANDN U3802 ( .A(n3103), .B(n3102), .Z(n3107) );
  NAND U3803 ( .A(n3105), .B(n3104), .Z(n3106) );
  NAND U3804 ( .A(n3107), .B(n3106), .Z(n3152) );
  NANDN U3805 ( .A(n3109), .B(n3108), .Z(n3113) );
  NAND U3806 ( .A(n3111), .B(n3110), .Z(n3112) );
  AND U3807 ( .A(n3113), .B(n3112), .Z(n3166) );
  NANDN U3808 ( .A(n3115), .B(n3114), .Z(n3119) );
  NAND U3809 ( .A(n3117), .B(n3116), .Z(n3118) );
  NAND U3810 ( .A(n3119), .B(n3118), .Z(n3282) );
  NANDN U3811 ( .A(n3125), .B(n3124), .Z(n3129) );
  NAND U3812 ( .A(n3127), .B(n3126), .Z(n3128) );
  NAND U3813 ( .A(n3129), .B(n3128), .Z(n3280) );
  XNOR U3814 ( .A(n3279), .B(n3280), .Z(n3281) );
  XOR U3815 ( .A(n3282), .B(n3281), .Z(n3164) );
  NAND U3816 ( .A(n3131), .B(n3130), .Z(n3135) );
  NANDN U3817 ( .A(n3133), .B(n3132), .Z(n3134) );
  AND U3818 ( .A(n3135), .B(n3134), .Z(n3165) );
  XOR U3819 ( .A(n3164), .B(n3165), .Z(n3136) );
  XNOR U3820 ( .A(n3166), .B(n3136), .Z(n3153) );
  XNOR U3821 ( .A(n3152), .B(n3153), .Z(n3154) );
  XNOR U3822 ( .A(n3155), .B(n3154), .Z(n3148) );
  NAND U3823 ( .A(n3138), .B(n3137), .Z(n3142) );
  NAND U3824 ( .A(n3140), .B(n3139), .Z(n3141) );
  NAND U3825 ( .A(n3142), .B(n3141), .Z(n3149) );
  XNOR U3826 ( .A(n3148), .B(n3149), .Z(n3150) );
  XNOR U3827 ( .A(n3151), .B(n3150), .Z(n3285) );
  XNOR U3828 ( .A(n3285), .B(sreg[129]), .Z(n3287) );
  NAND U3829 ( .A(n3143), .B(sreg[128]), .Z(n3147) );
  OR U3830 ( .A(n3145), .B(n3144), .Z(n3146) );
  AND U3831 ( .A(n3147), .B(n3146), .Z(n3286) );
  XOR U3832 ( .A(n3287), .B(n3286), .Z(c[129]) );
  NANDN U3833 ( .A(n3153), .B(n3152), .Z(n3157) );
  NAND U3834 ( .A(n3155), .B(n3154), .Z(n3156) );
  NAND U3835 ( .A(n3157), .B(n3156), .Z(n3291) );
  NANDN U3836 ( .A(n3159), .B(n3158), .Z(n3163) );
  OR U3837 ( .A(n3161), .B(n3160), .Z(n3162) );
  NAND U3838 ( .A(n3163), .B(n3162), .Z(n3294) );
  XNOR U3839 ( .A(n3294), .B(n3295), .Z(n3296) );
  NANDN U3840 ( .A(n3168), .B(n3167), .Z(n3172) );
  NANDN U3841 ( .A(n3170), .B(n3169), .Z(n3171) );
  NAND U3842 ( .A(n3172), .B(n3171), .Z(n3309) );
  NANDN U3843 ( .A(n3174), .B(n3173), .Z(n3178) );
  NAND U3844 ( .A(n3176), .B(n3175), .Z(n3177) );
  NAND U3845 ( .A(n3178), .B(n3177), .Z(n3414) );
  NANDN U3846 ( .A(n3180), .B(n3179), .Z(n3184) );
  NAND U3847 ( .A(n3182), .B(n3181), .Z(n3183) );
  NAND U3848 ( .A(n3184), .B(n3183), .Z(n3413) );
  XNOR U3849 ( .A(n3413), .B(n3412), .Z(n3415) );
  XOR U3850 ( .A(n3414), .B(n3415), .Z(n3306) );
  NANDN U3851 ( .A(n3190), .B(n3189), .Z(n3194) );
  NAND U3852 ( .A(n3192), .B(n3191), .Z(n3193) );
  NAND U3853 ( .A(n3194), .B(n3193), .Z(n3408) );
  XOR U3854 ( .A(b[17]), .B(a[18]), .Z(n3349) );
  NAND U3855 ( .A(n3349), .B(n18673), .Z(n3197) );
  NAND U3856 ( .A(n3195), .B(n18674), .Z(n3196) );
  NAND U3857 ( .A(n3197), .B(n3196), .Z(n3324) );
  XNOR U3858 ( .A(b[31]), .B(a[4]), .Z(n3352) );
  NANDN U3859 ( .A(n3352), .B(n19472), .Z(n3200) );
  NANDN U3860 ( .A(n3198), .B(n19473), .Z(n3199) );
  AND U3861 ( .A(n3200), .B(n3199), .Z(n3322) );
  OR U3862 ( .A(n3201), .B(n16988), .Z(n3203) );
  XNOR U3863 ( .A(b[3]), .B(a[32]), .Z(n3355) );
  NANDN U3864 ( .A(n3355), .B(n16990), .Z(n3202) );
  AND U3865 ( .A(n3203), .B(n3202), .Z(n3323) );
  XOR U3866 ( .A(n3324), .B(n3325), .Z(n3406) );
  NANDN U3867 ( .A(n3204), .B(n18832), .Z(n3206) );
  XNOR U3868 ( .A(b[19]), .B(a[16]), .Z(n3340) );
  NANDN U3869 ( .A(n3340), .B(n18834), .Z(n3205) );
  NAND U3870 ( .A(n3206), .B(n3205), .Z(n3373) );
  XNOR U3871 ( .A(b[27]), .B(a[8]), .Z(n3343) );
  NANDN U3872 ( .A(n3343), .B(n19336), .Z(n3209) );
  NANDN U3873 ( .A(n3207), .B(n19337), .Z(n3208) );
  NAND U3874 ( .A(n3209), .B(n3208), .Z(n3370) );
  XNOR U3875 ( .A(b[5]), .B(a[30]), .Z(n3346) );
  NANDN U3876 ( .A(n3346), .B(n17310), .Z(n3212) );
  NANDN U3877 ( .A(n3210), .B(n17311), .Z(n3211) );
  AND U3878 ( .A(n3212), .B(n3211), .Z(n3371) );
  XNOR U3879 ( .A(n3370), .B(n3371), .Z(n3372) );
  XOR U3880 ( .A(n3373), .B(n3372), .Z(n3407) );
  XOR U3881 ( .A(n3406), .B(n3407), .Z(n3409) );
  XOR U3882 ( .A(n3408), .B(n3409), .Z(n3307) );
  XOR U3883 ( .A(n3306), .B(n3307), .Z(n3308) );
  XNOR U3884 ( .A(n3309), .B(n3308), .Z(n3425) );
  OR U3885 ( .A(n3214), .B(n3213), .Z(n3218) );
  NAND U3886 ( .A(n3216), .B(n3215), .Z(n3217) );
  AND U3887 ( .A(n3218), .B(n3217), .Z(n3422) );
  NANDN U3888 ( .A(n3220), .B(n3219), .Z(n3224) );
  NAND U3889 ( .A(n3222), .B(n3221), .Z(n3223) );
  NAND U3890 ( .A(n3224), .B(n3223), .Z(n3303) );
  XNOR U3891 ( .A(b[9]), .B(a[26]), .Z(n3376) );
  NANDN U3892 ( .A(n3376), .B(n17814), .Z(n3227) );
  NANDN U3893 ( .A(n3225), .B(n17815), .Z(n3226) );
  NAND U3894 ( .A(n3227), .B(n3226), .Z(n3330) );
  NAND U3895 ( .A(n3228), .B(n18513), .Z(n3230) );
  XOR U3896 ( .A(b[15]), .B(a[20]), .Z(n3379) );
  NANDN U3897 ( .A(n18512), .B(n3379), .Z(n3229) );
  AND U3898 ( .A(n3230), .B(n3229), .Z(n3328) );
  NAND U3899 ( .A(n3231), .B(n19013), .Z(n3233) );
  XNOR U3900 ( .A(b[21]), .B(a[14]), .Z(n3382) );
  NANDN U3901 ( .A(n3382), .B(n19015), .Z(n3232) );
  AND U3902 ( .A(n3233), .B(n3232), .Z(n3329) );
  XOR U3903 ( .A(n3330), .B(n3331), .Z(n3319) );
  XNOR U3904 ( .A(b[11]), .B(a[24]), .Z(n3385) );
  OR U3905 ( .A(n3385), .B(n18194), .Z(n3236) );
  NANDN U3906 ( .A(n3234), .B(n18104), .Z(n3235) );
  NAND U3907 ( .A(n3236), .B(n3235), .Z(n3317) );
  XOR U3908 ( .A(n580), .B(a[22]), .Z(n3388) );
  NANDN U3909 ( .A(n3388), .B(n18336), .Z(n3239) );
  NANDN U3910 ( .A(n3237), .B(n18337), .Z(n3238) );
  NAND U3911 ( .A(n3239), .B(n3238), .Z(n3316) );
  XOR U3912 ( .A(n3319), .B(n3318), .Z(n3313) );
  NANDN U3913 ( .A(n577), .B(a[34]), .Z(n3240) );
  XOR U3914 ( .A(n17151), .B(n3240), .Z(n3242) );
  NANDN U3915 ( .A(b[0]), .B(a[33]), .Z(n3241) );
  AND U3916 ( .A(n3242), .B(n3241), .Z(n3336) );
  NAND U3917 ( .A(n19406), .B(n3243), .Z(n3245) );
  XNOR U3918 ( .A(n584), .B(a[6]), .Z(n3391) );
  NANDN U3919 ( .A(n576), .B(n3391), .Z(n3244) );
  NAND U3920 ( .A(n3245), .B(n3244), .Z(n3334) );
  NANDN U3921 ( .A(n585), .B(a[2]), .Z(n3335) );
  XNOR U3922 ( .A(n3334), .B(n3335), .Z(n3337) );
  XNOR U3923 ( .A(n3336), .B(n3337), .Z(n3311) );
  XOR U3924 ( .A(b[23]), .B(a[12]), .Z(n3397) );
  NANDN U3925 ( .A(n19127), .B(n3397), .Z(n3248) );
  NANDN U3926 ( .A(n3246), .B(n19128), .Z(n3247) );
  NAND U3927 ( .A(n3248), .B(n3247), .Z(n3367) );
  NANDN U3928 ( .A(n3249), .B(n17553), .Z(n3251) );
  XOR U3929 ( .A(b[7]), .B(a[28]), .Z(n3400) );
  NAND U3930 ( .A(n3400), .B(n17555), .Z(n3250) );
  NAND U3931 ( .A(n3251), .B(n3250), .Z(n3364) );
  XOR U3932 ( .A(b[25]), .B(a[10]), .Z(n3403) );
  NAND U3933 ( .A(n3403), .B(n19240), .Z(n3254) );
  NAND U3934 ( .A(n3252), .B(n19242), .Z(n3253) );
  AND U3935 ( .A(n3254), .B(n3253), .Z(n3365) );
  XNOR U3936 ( .A(n3364), .B(n3365), .Z(n3366) );
  XOR U3937 ( .A(n3367), .B(n3366), .Z(n3310) );
  XNOR U3938 ( .A(n3313), .B(n3312), .Z(n3361) );
  NANDN U3939 ( .A(n3256), .B(n3255), .Z(n3260) );
  NAND U3940 ( .A(n3258), .B(n3257), .Z(n3259) );
  NAND U3941 ( .A(n3260), .B(n3259), .Z(n3358) );
  NANDN U3942 ( .A(n3262), .B(n3261), .Z(n3266) );
  NAND U3943 ( .A(n3264), .B(n3263), .Z(n3265) );
  NAND U3944 ( .A(n3266), .B(n3265), .Z(n3359) );
  XNOR U3945 ( .A(n3358), .B(n3359), .Z(n3360) );
  XNOR U3946 ( .A(n3361), .B(n3360), .Z(n3300) );
  NANDN U3947 ( .A(n3268), .B(n3267), .Z(n3272) );
  OR U3948 ( .A(n3270), .B(n3269), .Z(n3271) );
  NAND U3949 ( .A(n3272), .B(n3271), .Z(n3301) );
  XOR U3950 ( .A(n3300), .B(n3301), .Z(n3302) );
  XNOR U3951 ( .A(n3303), .B(n3302), .Z(n3423) );
  XOR U3952 ( .A(n3425), .B(n3424), .Z(n3419) );
  NANDN U3953 ( .A(n3274), .B(n3273), .Z(n3278) );
  NAND U3954 ( .A(n3276), .B(n3275), .Z(n3277) );
  NAND U3955 ( .A(n3278), .B(n3277), .Z(n3416) );
  NANDN U3956 ( .A(n3280), .B(n3279), .Z(n3284) );
  NANDN U3957 ( .A(n3282), .B(n3281), .Z(n3283) );
  AND U3958 ( .A(n3284), .B(n3283), .Z(n3417) );
  XNOR U3959 ( .A(n3416), .B(n3417), .Z(n3418) );
  XOR U3960 ( .A(n3419), .B(n3418), .Z(n3297) );
  XNOR U3961 ( .A(n3296), .B(n3297), .Z(n3290) );
  XNOR U3962 ( .A(n3291), .B(n3290), .Z(n3292) );
  XNOR U3963 ( .A(n3293), .B(n3292), .Z(n3428) );
  XNOR U3964 ( .A(n3428), .B(sreg[130]), .Z(n3430) );
  NAND U3965 ( .A(n3285), .B(sreg[129]), .Z(n3289) );
  OR U3966 ( .A(n3287), .B(n3286), .Z(n3288) );
  AND U3967 ( .A(n3289), .B(n3288), .Z(n3429) );
  XOR U3968 ( .A(n3430), .B(n3429), .Z(c[130]) );
  NANDN U3969 ( .A(n3295), .B(n3294), .Z(n3299) );
  NANDN U3970 ( .A(n3297), .B(n3296), .Z(n3298) );
  NAND U3971 ( .A(n3299), .B(n3298), .Z(n3433) );
  OR U3972 ( .A(n3301), .B(n3300), .Z(n3305) );
  NAND U3973 ( .A(n3303), .B(n3302), .Z(n3304) );
  NAND U3974 ( .A(n3305), .B(n3304), .Z(n3565) );
  XNOR U3975 ( .A(n3565), .B(n3566), .Z(n3567) );
  NANDN U3976 ( .A(n3311), .B(n3310), .Z(n3315) );
  NANDN U3977 ( .A(n3313), .B(n3312), .Z(n3314) );
  NAND U3978 ( .A(n3315), .B(n3314), .Z(n3562) );
  OR U3979 ( .A(n3317), .B(n3316), .Z(n3321) );
  NAND U3980 ( .A(n3319), .B(n3318), .Z(n3320) );
  NAND U3981 ( .A(n3321), .B(n3320), .Z(n3495) );
  OR U3982 ( .A(n3323), .B(n3322), .Z(n3327) );
  NANDN U3983 ( .A(n3325), .B(n3324), .Z(n3326) );
  NAND U3984 ( .A(n3327), .B(n3326), .Z(n3494) );
  OR U3985 ( .A(n3329), .B(n3328), .Z(n3333) );
  NANDN U3986 ( .A(n3331), .B(n3330), .Z(n3332) );
  NAND U3987 ( .A(n3333), .B(n3332), .Z(n3493) );
  XOR U3988 ( .A(n3495), .B(n3496), .Z(n3559) );
  NANDN U3989 ( .A(n3335), .B(n3334), .Z(n3339) );
  NAND U3990 ( .A(n3337), .B(n3336), .Z(n3338) );
  NAND U3991 ( .A(n3339), .B(n3338), .Z(n3508) );
  NANDN U3992 ( .A(n3340), .B(n18832), .Z(n3342) );
  XNOR U3993 ( .A(b[19]), .B(a[17]), .Z(n3451) );
  NANDN U3994 ( .A(n3451), .B(n18834), .Z(n3341) );
  NAND U3995 ( .A(n3342), .B(n3341), .Z(n3544) );
  XNOR U3996 ( .A(b[27]), .B(a[9]), .Z(n3454) );
  NANDN U3997 ( .A(n3454), .B(n19336), .Z(n3345) );
  NANDN U3998 ( .A(n3343), .B(n19337), .Z(n3344) );
  NAND U3999 ( .A(n3345), .B(n3344), .Z(n3541) );
  XOR U4000 ( .A(b[5]), .B(a[31]), .Z(n3457) );
  NAND U4001 ( .A(n3457), .B(n17310), .Z(n3348) );
  NANDN U4002 ( .A(n3346), .B(n17311), .Z(n3347) );
  AND U4003 ( .A(n3348), .B(n3347), .Z(n3542) );
  XNOR U4004 ( .A(n3541), .B(n3542), .Z(n3543) );
  XNOR U4005 ( .A(n3544), .B(n3543), .Z(n3506) );
  XOR U4006 ( .A(b[17]), .B(a[19]), .Z(n3460) );
  NAND U4007 ( .A(n3460), .B(n18673), .Z(n3351) );
  NAND U4008 ( .A(n3349), .B(n18674), .Z(n3350) );
  NAND U4009 ( .A(n3351), .B(n3350), .Z(n3478) );
  XNOR U4010 ( .A(b[31]), .B(a[5]), .Z(n3463) );
  NANDN U4011 ( .A(n3463), .B(n19472), .Z(n3354) );
  NANDN U4012 ( .A(n3352), .B(n19473), .Z(n3353) );
  NAND U4013 ( .A(n3354), .B(n3353), .Z(n3475) );
  OR U4014 ( .A(n3355), .B(n16988), .Z(n3357) );
  XNOR U4015 ( .A(b[3]), .B(a[33]), .Z(n3466) );
  NANDN U4016 ( .A(n3466), .B(n16990), .Z(n3356) );
  AND U4017 ( .A(n3357), .B(n3356), .Z(n3476) );
  XNOR U4018 ( .A(n3475), .B(n3476), .Z(n3477) );
  XOR U4019 ( .A(n3478), .B(n3477), .Z(n3505) );
  XNOR U4020 ( .A(n3506), .B(n3505), .Z(n3507) );
  XNOR U4021 ( .A(n3508), .B(n3507), .Z(n3560) );
  XNOR U4022 ( .A(n3559), .B(n3560), .Z(n3561) );
  XNOR U4023 ( .A(n3562), .B(n3561), .Z(n3574) );
  NANDN U4024 ( .A(n3359), .B(n3358), .Z(n3363) );
  NANDN U4025 ( .A(n3361), .B(n3360), .Z(n3362) );
  NAND U4026 ( .A(n3363), .B(n3362), .Z(n3556) );
  NANDN U4027 ( .A(n3365), .B(n3364), .Z(n3369) );
  NAND U4028 ( .A(n3367), .B(n3366), .Z(n3368) );
  NAND U4029 ( .A(n3369), .B(n3368), .Z(n3499) );
  NANDN U4030 ( .A(n3371), .B(n3370), .Z(n3375) );
  NAND U4031 ( .A(n3373), .B(n3372), .Z(n3374) );
  AND U4032 ( .A(n3375), .B(n3374), .Z(n3500) );
  XNOR U4033 ( .A(n3499), .B(n3500), .Z(n3501) );
  XNOR U4034 ( .A(b[9]), .B(a[27]), .Z(n3511) );
  NANDN U4035 ( .A(n3511), .B(n17814), .Z(n3378) );
  NANDN U4036 ( .A(n3376), .B(n17815), .Z(n3377) );
  NAND U4037 ( .A(n3378), .B(n3377), .Z(n3483) );
  NAND U4038 ( .A(n3379), .B(n18513), .Z(n3381) );
  XOR U4039 ( .A(b[15]), .B(a[21]), .Z(n3514) );
  NANDN U4040 ( .A(n18512), .B(n3514), .Z(n3380) );
  AND U4041 ( .A(n3381), .B(n3380), .Z(n3481) );
  NANDN U4042 ( .A(n3382), .B(n19013), .Z(n3384) );
  XOR U4043 ( .A(b[21]), .B(n5159), .Z(n3517) );
  NANDN U4044 ( .A(n3517), .B(n19015), .Z(n3383) );
  AND U4045 ( .A(n3384), .B(n3383), .Z(n3482) );
  XOR U4046 ( .A(n3483), .B(n3484), .Z(n3472) );
  XNOR U4047 ( .A(b[11]), .B(a[25]), .Z(n3520) );
  OR U4048 ( .A(n3520), .B(n18194), .Z(n3387) );
  NANDN U4049 ( .A(n3385), .B(n18104), .Z(n3386) );
  NAND U4050 ( .A(n3387), .B(n3386), .Z(n3470) );
  XOR U4051 ( .A(n580), .B(a[23]), .Z(n3523) );
  NANDN U4052 ( .A(n3523), .B(n18336), .Z(n3390) );
  NANDN U4053 ( .A(n3388), .B(n18337), .Z(n3389) );
  AND U4054 ( .A(n3390), .B(n3389), .Z(n3469) );
  XNOR U4055 ( .A(n3470), .B(n3469), .Z(n3471) );
  XOR U4056 ( .A(n3472), .B(n3471), .Z(n3489) );
  NAND U4057 ( .A(n19406), .B(n3391), .Z(n3393) );
  XNOR U4058 ( .A(n584), .B(a[7]), .Z(n3529) );
  NANDN U4059 ( .A(n576), .B(n3529), .Z(n3392) );
  NAND U4060 ( .A(n3393), .B(n3392), .Z(n3445) );
  NANDN U4061 ( .A(n585), .B(a[3]), .Z(n3446) );
  XNOR U4062 ( .A(n3445), .B(n3446), .Z(n3448) );
  NANDN U4063 ( .A(n577), .B(a[35]), .Z(n3394) );
  XOR U4064 ( .A(n17151), .B(n3394), .Z(n3396) );
  NANDN U4065 ( .A(b[0]), .B(a[34]), .Z(n3395) );
  AND U4066 ( .A(n3396), .B(n3395), .Z(n3447) );
  XOR U4067 ( .A(n3448), .B(n3447), .Z(n3487) );
  XNOR U4068 ( .A(b[23]), .B(a[13]), .Z(n3532) );
  OR U4069 ( .A(n3532), .B(n19127), .Z(n3399) );
  NAND U4070 ( .A(n3397), .B(n19128), .Z(n3398) );
  NAND U4071 ( .A(n3399), .B(n3398), .Z(n3550) );
  NAND U4072 ( .A(n3400), .B(n17553), .Z(n3402) );
  XNOR U4073 ( .A(b[7]), .B(a[29]), .Z(n3535) );
  NANDN U4074 ( .A(n3535), .B(n17555), .Z(n3401) );
  NAND U4075 ( .A(n3402), .B(n3401), .Z(n3547) );
  XNOR U4076 ( .A(b[25]), .B(a[11]), .Z(n3538) );
  NANDN U4077 ( .A(n3538), .B(n19240), .Z(n3405) );
  NAND U4078 ( .A(n3403), .B(n19242), .Z(n3404) );
  AND U4079 ( .A(n3405), .B(n3404), .Z(n3548) );
  XNOR U4080 ( .A(n3547), .B(n3548), .Z(n3549) );
  XNOR U4081 ( .A(n3550), .B(n3549), .Z(n3488) );
  XOR U4082 ( .A(n3487), .B(n3488), .Z(n3490) );
  XNOR U4083 ( .A(n3489), .B(n3490), .Z(n3502) );
  XOR U4084 ( .A(n3501), .B(n3502), .Z(n3553) );
  NANDN U4085 ( .A(n3407), .B(n3406), .Z(n3411) );
  OR U4086 ( .A(n3409), .B(n3408), .Z(n3410) );
  AND U4087 ( .A(n3411), .B(n3410), .Z(n3554) );
  XNOR U4088 ( .A(n3553), .B(n3554), .Z(n3555) );
  XOR U4089 ( .A(n3556), .B(n3555), .Z(n3572) );
  XOR U4090 ( .A(n3572), .B(n3571), .Z(n3573) );
  XNOR U4091 ( .A(n3574), .B(n3573), .Z(n3568) );
  XOR U4092 ( .A(n3567), .B(n3568), .Z(n3442) );
  NANDN U4093 ( .A(n3417), .B(n3416), .Z(n3421) );
  NANDN U4094 ( .A(n3419), .B(n3418), .Z(n3420) );
  NAND U4095 ( .A(n3421), .B(n3420), .Z(n3439) );
  OR U4096 ( .A(n3423), .B(n3422), .Z(n3427) );
  NAND U4097 ( .A(n3425), .B(n3424), .Z(n3426) );
  NAND U4098 ( .A(n3427), .B(n3426), .Z(n3440) );
  XNOR U4099 ( .A(n3439), .B(n3440), .Z(n3441) );
  XNOR U4100 ( .A(n3442), .B(n3441), .Z(n3434) );
  XNOR U4101 ( .A(n3433), .B(n3434), .Z(n3435) );
  XNOR U4102 ( .A(n3436), .B(n3435), .Z(n3577) );
  XNOR U4103 ( .A(n3577), .B(sreg[131]), .Z(n3579) );
  NAND U4104 ( .A(n3428), .B(sreg[130]), .Z(n3432) );
  OR U4105 ( .A(n3430), .B(n3429), .Z(n3431) );
  AND U4106 ( .A(n3432), .B(n3431), .Z(n3578) );
  XOR U4107 ( .A(n3579), .B(n3578), .Z(c[131]) );
  NANDN U4108 ( .A(n3434), .B(n3433), .Z(n3438) );
  NAND U4109 ( .A(n3436), .B(n3435), .Z(n3437) );
  NAND U4110 ( .A(n3438), .B(n3437), .Z(n3585) );
  NANDN U4111 ( .A(n3440), .B(n3439), .Z(n3444) );
  NAND U4112 ( .A(n3442), .B(n3441), .Z(n3443) );
  NAND U4113 ( .A(n3444), .B(n3443), .Z(n3583) );
  NANDN U4114 ( .A(n3446), .B(n3445), .Z(n3450) );
  NAND U4115 ( .A(n3448), .B(n3447), .Z(n3449) );
  NAND U4116 ( .A(n3450), .B(n3449), .Z(n3657) );
  NANDN U4117 ( .A(n3451), .B(n18832), .Z(n3453) );
  XNOR U4118 ( .A(b[19]), .B(a[18]), .Z(n3600) );
  NANDN U4119 ( .A(n3600), .B(n18834), .Z(n3452) );
  NAND U4120 ( .A(n3453), .B(n3452), .Z(n3667) );
  XNOR U4121 ( .A(b[27]), .B(a[10]), .Z(n3603) );
  NANDN U4122 ( .A(n3603), .B(n19336), .Z(n3456) );
  NANDN U4123 ( .A(n3454), .B(n19337), .Z(n3455) );
  NAND U4124 ( .A(n3456), .B(n3455), .Z(n3664) );
  XOR U4125 ( .A(b[5]), .B(a[32]), .Z(n3606) );
  NAND U4126 ( .A(n3606), .B(n17310), .Z(n3459) );
  NAND U4127 ( .A(n3457), .B(n17311), .Z(n3458) );
  AND U4128 ( .A(n3459), .B(n3458), .Z(n3665) );
  XNOR U4129 ( .A(n3664), .B(n3665), .Z(n3666) );
  XNOR U4130 ( .A(n3667), .B(n3666), .Z(n3655) );
  XOR U4131 ( .A(b[17]), .B(a[20]), .Z(n3609) );
  NAND U4132 ( .A(n3609), .B(n18673), .Z(n3462) );
  NAND U4133 ( .A(n3460), .B(n18674), .Z(n3461) );
  NAND U4134 ( .A(n3462), .B(n3461), .Z(n3627) );
  XNOR U4135 ( .A(b[31]), .B(a[6]), .Z(n3612) );
  NANDN U4136 ( .A(n3612), .B(n19472), .Z(n3465) );
  NANDN U4137 ( .A(n3463), .B(n19473), .Z(n3464) );
  NAND U4138 ( .A(n3465), .B(n3464), .Z(n3624) );
  OR U4139 ( .A(n3466), .B(n16988), .Z(n3468) );
  XNOR U4140 ( .A(b[3]), .B(a[34]), .Z(n3615) );
  NANDN U4141 ( .A(n3615), .B(n16990), .Z(n3467) );
  AND U4142 ( .A(n3468), .B(n3467), .Z(n3625) );
  XNOR U4143 ( .A(n3624), .B(n3625), .Z(n3626) );
  XOR U4144 ( .A(n3627), .B(n3626), .Z(n3654) );
  XNOR U4145 ( .A(n3655), .B(n3654), .Z(n3656) );
  XNOR U4146 ( .A(n3657), .B(n3656), .Z(n3700) );
  NANDN U4147 ( .A(n3470), .B(n3469), .Z(n3474) );
  NAND U4148 ( .A(n3472), .B(n3471), .Z(n3473) );
  NAND U4149 ( .A(n3474), .B(n3473), .Z(n3645) );
  NANDN U4150 ( .A(n3476), .B(n3475), .Z(n3480) );
  NAND U4151 ( .A(n3478), .B(n3477), .Z(n3479) );
  NAND U4152 ( .A(n3480), .B(n3479), .Z(n3643) );
  OR U4153 ( .A(n3482), .B(n3481), .Z(n3486) );
  NANDN U4154 ( .A(n3484), .B(n3483), .Z(n3485) );
  NAND U4155 ( .A(n3486), .B(n3485), .Z(n3642) );
  XNOR U4156 ( .A(n3645), .B(n3644), .Z(n3701) );
  XOR U4157 ( .A(n3700), .B(n3701), .Z(n3703) );
  NANDN U4158 ( .A(n3488), .B(n3487), .Z(n3492) );
  OR U4159 ( .A(n3490), .B(n3489), .Z(n3491) );
  NAND U4160 ( .A(n3492), .B(n3491), .Z(n3702) );
  XOR U4161 ( .A(n3703), .B(n3702), .Z(n3720) );
  OR U4162 ( .A(n3494), .B(n3493), .Z(n3498) );
  NANDN U4163 ( .A(n3496), .B(n3495), .Z(n3497) );
  NAND U4164 ( .A(n3498), .B(n3497), .Z(n3719) );
  NANDN U4165 ( .A(n3500), .B(n3499), .Z(n3504) );
  NANDN U4166 ( .A(n3502), .B(n3501), .Z(n3503) );
  NAND U4167 ( .A(n3504), .B(n3503), .Z(n3709) );
  NANDN U4168 ( .A(n3506), .B(n3505), .Z(n3510) );
  NAND U4169 ( .A(n3508), .B(n3507), .Z(n3509) );
  NAND U4170 ( .A(n3510), .B(n3509), .Z(n3706) );
  XNOR U4171 ( .A(b[9]), .B(a[28]), .Z(n3670) );
  NANDN U4172 ( .A(n3670), .B(n17814), .Z(n3513) );
  NANDN U4173 ( .A(n3511), .B(n17815), .Z(n3512) );
  NAND U4174 ( .A(n3513), .B(n3512), .Z(n3632) );
  NAND U4175 ( .A(n3514), .B(n18513), .Z(n3516) );
  XOR U4176 ( .A(b[15]), .B(a[22]), .Z(n3673) );
  NANDN U4177 ( .A(n18512), .B(n3673), .Z(n3515) );
  AND U4178 ( .A(n3516), .B(n3515), .Z(n3630) );
  NANDN U4179 ( .A(n3517), .B(n19013), .Z(n3519) );
  XNOR U4180 ( .A(b[21]), .B(a[16]), .Z(n3676) );
  NANDN U4181 ( .A(n3676), .B(n19015), .Z(n3518) );
  AND U4182 ( .A(n3519), .B(n3518), .Z(n3631) );
  XOR U4183 ( .A(n3632), .B(n3633), .Z(n3621) );
  XNOR U4184 ( .A(b[11]), .B(a[26]), .Z(n3679) );
  OR U4185 ( .A(n3679), .B(n18194), .Z(n3522) );
  NANDN U4186 ( .A(n3520), .B(n18104), .Z(n3521) );
  NAND U4187 ( .A(n3522), .B(n3521), .Z(n3619) );
  XOR U4188 ( .A(n580), .B(a[24]), .Z(n3682) );
  NANDN U4189 ( .A(n3682), .B(n18336), .Z(n3525) );
  NANDN U4190 ( .A(n3523), .B(n18337), .Z(n3524) );
  AND U4191 ( .A(n3525), .B(n3524), .Z(n3618) );
  XNOR U4192 ( .A(n3619), .B(n3618), .Z(n3620) );
  XOR U4193 ( .A(n3621), .B(n3620), .Z(n3639) );
  NANDN U4194 ( .A(n577), .B(a[36]), .Z(n3526) );
  XOR U4195 ( .A(n17151), .B(n3526), .Z(n3528) );
  NANDN U4196 ( .A(b[0]), .B(a[35]), .Z(n3527) );
  AND U4197 ( .A(n3528), .B(n3527), .Z(n3596) );
  NAND U4198 ( .A(n19406), .B(n3529), .Z(n3531) );
  XNOR U4199 ( .A(n584), .B(a[8]), .Z(n3688) );
  NANDN U4200 ( .A(n576), .B(n3688), .Z(n3530) );
  NAND U4201 ( .A(n3531), .B(n3530), .Z(n3594) );
  NANDN U4202 ( .A(n585), .B(a[4]), .Z(n3595) );
  XNOR U4203 ( .A(n3594), .B(n3595), .Z(n3597) );
  XOR U4204 ( .A(n3596), .B(n3597), .Z(n3636) );
  XOR U4205 ( .A(b[23]), .B(a[14]), .Z(n3691) );
  NANDN U4206 ( .A(n19127), .B(n3691), .Z(n3534) );
  NANDN U4207 ( .A(n3532), .B(n19128), .Z(n3533) );
  NAND U4208 ( .A(n3534), .B(n3533), .Z(n3661) );
  NANDN U4209 ( .A(n3535), .B(n17553), .Z(n3537) );
  XNOR U4210 ( .A(b[7]), .B(a[30]), .Z(n3694) );
  NANDN U4211 ( .A(n3694), .B(n17555), .Z(n3536) );
  NAND U4212 ( .A(n3537), .B(n3536), .Z(n3658) );
  XOR U4213 ( .A(b[25]), .B(a[12]), .Z(n3697) );
  NAND U4214 ( .A(n3697), .B(n19240), .Z(n3540) );
  NANDN U4215 ( .A(n3538), .B(n19242), .Z(n3539) );
  AND U4216 ( .A(n3540), .B(n3539), .Z(n3659) );
  XNOR U4217 ( .A(n3658), .B(n3659), .Z(n3660) );
  XNOR U4218 ( .A(n3661), .B(n3660), .Z(n3637) );
  XNOR U4219 ( .A(n3636), .B(n3637), .Z(n3638) );
  XNOR U4220 ( .A(n3639), .B(n3638), .Z(n3651) );
  NANDN U4221 ( .A(n3542), .B(n3541), .Z(n3546) );
  NAND U4222 ( .A(n3544), .B(n3543), .Z(n3545) );
  NAND U4223 ( .A(n3546), .B(n3545), .Z(n3649) );
  NANDN U4224 ( .A(n3548), .B(n3547), .Z(n3552) );
  NAND U4225 ( .A(n3550), .B(n3549), .Z(n3551) );
  AND U4226 ( .A(n3552), .B(n3551), .Z(n3648) );
  XNOR U4227 ( .A(n3649), .B(n3648), .Z(n3650) );
  XNOR U4228 ( .A(n3651), .B(n3650), .Z(n3707) );
  XNOR U4229 ( .A(n3706), .B(n3707), .Z(n3708) );
  XOR U4230 ( .A(n3709), .B(n3708), .Z(n3718) );
  XOR U4231 ( .A(n3719), .B(n3718), .Z(n3721) );
  NANDN U4232 ( .A(n3554), .B(n3553), .Z(n3558) );
  NAND U4233 ( .A(n3556), .B(n3555), .Z(n3557) );
  NAND U4234 ( .A(n3558), .B(n3557), .Z(n3712) );
  NANDN U4235 ( .A(n3560), .B(n3559), .Z(n3564) );
  NAND U4236 ( .A(n3562), .B(n3561), .Z(n3563) );
  NAND U4237 ( .A(n3564), .B(n3563), .Z(n3713) );
  XNOR U4238 ( .A(n3712), .B(n3713), .Z(n3714) );
  XOR U4239 ( .A(n3715), .B(n3714), .Z(n3590) );
  NANDN U4240 ( .A(n3566), .B(n3565), .Z(n3570) );
  NANDN U4241 ( .A(n3568), .B(n3567), .Z(n3569) );
  NAND U4242 ( .A(n3570), .B(n3569), .Z(n3589) );
  NANDN U4243 ( .A(n3572), .B(n3571), .Z(n3576) );
  OR U4244 ( .A(n3574), .B(n3573), .Z(n3575) );
  AND U4245 ( .A(n3576), .B(n3575), .Z(n3588) );
  XNOR U4246 ( .A(n3589), .B(n3588), .Z(n3591) );
  XOR U4247 ( .A(n3590), .B(n3591), .Z(n3582) );
  XOR U4248 ( .A(n3583), .B(n3582), .Z(n3584) );
  XNOR U4249 ( .A(n3585), .B(n3584), .Z(n3724) );
  XNOR U4250 ( .A(n3724), .B(sreg[132]), .Z(n3726) );
  NAND U4251 ( .A(n3577), .B(sreg[131]), .Z(n3581) );
  OR U4252 ( .A(n3579), .B(n3578), .Z(n3580) );
  AND U4253 ( .A(n3581), .B(n3580), .Z(n3725) );
  XOR U4254 ( .A(n3726), .B(n3725), .Z(c[132]) );
  NAND U4255 ( .A(n3583), .B(n3582), .Z(n3587) );
  NAND U4256 ( .A(n3585), .B(n3584), .Z(n3586) );
  NAND U4257 ( .A(n3587), .B(n3586), .Z(n3732) );
  NANDN U4258 ( .A(n3589), .B(n3588), .Z(n3593) );
  NAND U4259 ( .A(n3591), .B(n3590), .Z(n3592) );
  NAND U4260 ( .A(n3593), .B(n3592), .Z(n3730) );
  NANDN U4261 ( .A(n3595), .B(n3594), .Z(n3599) );
  NAND U4262 ( .A(n3597), .B(n3596), .Z(n3598) );
  NAND U4263 ( .A(n3599), .B(n3598), .Z(n3816) );
  NANDN U4264 ( .A(n3600), .B(n18832), .Z(n3602) );
  XNOR U4265 ( .A(b[19]), .B(a[19]), .Z(n3759) );
  NANDN U4266 ( .A(n3759), .B(n18834), .Z(n3601) );
  NAND U4267 ( .A(n3602), .B(n3601), .Z(n3826) );
  XOR U4268 ( .A(b[27]), .B(n4573), .Z(n3762) );
  NANDN U4269 ( .A(n3762), .B(n19336), .Z(n3605) );
  NANDN U4270 ( .A(n3603), .B(n19337), .Z(n3604) );
  NAND U4271 ( .A(n3605), .B(n3604), .Z(n3823) );
  XOR U4272 ( .A(b[5]), .B(a[33]), .Z(n3765) );
  NAND U4273 ( .A(n3765), .B(n17310), .Z(n3608) );
  NAND U4274 ( .A(n3606), .B(n17311), .Z(n3607) );
  AND U4275 ( .A(n3608), .B(n3607), .Z(n3824) );
  XNOR U4276 ( .A(n3823), .B(n3824), .Z(n3825) );
  XNOR U4277 ( .A(n3826), .B(n3825), .Z(n3814) );
  XOR U4278 ( .A(b[17]), .B(a[21]), .Z(n3768) );
  NAND U4279 ( .A(n3768), .B(n18673), .Z(n3611) );
  NAND U4280 ( .A(n3609), .B(n18674), .Z(n3610) );
  NAND U4281 ( .A(n3611), .B(n3610), .Z(n3786) );
  XNOR U4282 ( .A(b[31]), .B(a[7]), .Z(n3771) );
  NANDN U4283 ( .A(n3771), .B(n19472), .Z(n3614) );
  NANDN U4284 ( .A(n3612), .B(n19473), .Z(n3613) );
  NAND U4285 ( .A(n3614), .B(n3613), .Z(n3783) );
  OR U4286 ( .A(n3615), .B(n16988), .Z(n3617) );
  XNOR U4287 ( .A(b[3]), .B(a[35]), .Z(n3774) );
  NANDN U4288 ( .A(n3774), .B(n16990), .Z(n3616) );
  AND U4289 ( .A(n3617), .B(n3616), .Z(n3784) );
  XNOR U4290 ( .A(n3783), .B(n3784), .Z(n3785) );
  XOR U4291 ( .A(n3786), .B(n3785), .Z(n3813) );
  XNOR U4292 ( .A(n3814), .B(n3813), .Z(n3815) );
  XNOR U4293 ( .A(n3816), .B(n3815), .Z(n3859) );
  NANDN U4294 ( .A(n3619), .B(n3618), .Z(n3623) );
  NAND U4295 ( .A(n3621), .B(n3620), .Z(n3622) );
  NAND U4296 ( .A(n3623), .B(n3622), .Z(n3804) );
  NANDN U4297 ( .A(n3625), .B(n3624), .Z(n3629) );
  NAND U4298 ( .A(n3627), .B(n3626), .Z(n3628) );
  NAND U4299 ( .A(n3629), .B(n3628), .Z(n3802) );
  OR U4300 ( .A(n3631), .B(n3630), .Z(n3635) );
  NANDN U4301 ( .A(n3633), .B(n3632), .Z(n3634) );
  NAND U4302 ( .A(n3635), .B(n3634), .Z(n3801) );
  XNOR U4303 ( .A(n3804), .B(n3803), .Z(n3860) );
  XOR U4304 ( .A(n3859), .B(n3860), .Z(n3862) );
  NANDN U4305 ( .A(n3637), .B(n3636), .Z(n3641) );
  NANDN U4306 ( .A(n3639), .B(n3638), .Z(n3640) );
  NAND U4307 ( .A(n3641), .B(n3640), .Z(n3861) );
  XOR U4308 ( .A(n3862), .B(n3861), .Z(n3749) );
  OR U4309 ( .A(n3643), .B(n3642), .Z(n3647) );
  NAND U4310 ( .A(n3645), .B(n3644), .Z(n3646) );
  NAND U4311 ( .A(n3647), .B(n3646), .Z(n3748) );
  NANDN U4312 ( .A(n3649), .B(n3648), .Z(n3653) );
  NANDN U4313 ( .A(n3651), .B(n3650), .Z(n3652) );
  NAND U4314 ( .A(n3653), .B(n3652), .Z(n3867) );
  NANDN U4315 ( .A(n3659), .B(n3658), .Z(n3663) );
  NAND U4316 ( .A(n3661), .B(n3660), .Z(n3662) );
  NAND U4317 ( .A(n3663), .B(n3662), .Z(n3807) );
  NANDN U4318 ( .A(n3665), .B(n3664), .Z(n3669) );
  NAND U4319 ( .A(n3667), .B(n3666), .Z(n3668) );
  AND U4320 ( .A(n3669), .B(n3668), .Z(n3808) );
  XNOR U4321 ( .A(n3807), .B(n3808), .Z(n3809) );
  XOR U4322 ( .A(b[9]), .B(n6835), .Z(n3829) );
  NANDN U4323 ( .A(n3829), .B(n17814), .Z(n3672) );
  NANDN U4324 ( .A(n3670), .B(n17815), .Z(n3671) );
  NAND U4325 ( .A(n3672), .B(n3671), .Z(n3791) );
  NAND U4326 ( .A(n3673), .B(n18513), .Z(n3675) );
  XOR U4327 ( .A(b[15]), .B(a[23]), .Z(n3832) );
  NANDN U4328 ( .A(n18512), .B(n3832), .Z(n3674) );
  AND U4329 ( .A(n3675), .B(n3674), .Z(n3789) );
  NANDN U4330 ( .A(n3676), .B(n19013), .Z(n3678) );
  XNOR U4331 ( .A(b[21]), .B(a[17]), .Z(n3835) );
  NANDN U4332 ( .A(n3835), .B(n19015), .Z(n3677) );
  AND U4333 ( .A(n3678), .B(n3677), .Z(n3790) );
  XOR U4334 ( .A(n3791), .B(n3792), .Z(n3780) );
  XNOR U4335 ( .A(b[11]), .B(a[27]), .Z(n3838) );
  OR U4336 ( .A(n3838), .B(n18194), .Z(n3681) );
  NANDN U4337 ( .A(n3679), .B(n18104), .Z(n3680) );
  NAND U4338 ( .A(n3681), .B(n3680), .Z(n3778) );
  XOR U4339 ( .A(n580), .B(a[25]), .Z(n3841) );
  NANDN U4340 ( .A(n3841), .B(n18336), .Z(n3684) );
  NANDN U4341 ( .A(n3682), .B(n18337), .Z(n3683) );
  AND U4342 ( .A(n3684), .B(n3683), .Z(n3777) );
  XNOR U4343 ( .A(n3778), .B(n3777), .Z(n3779) );
  XOR U4344 ( .A(n3780), .B(n3779), .Z(n3797) );
  NANDN U4345 ( .A(n577), .B(a[37]), .Z(n3685) );
  XOR U4346 ( .A(n17151), .B(n3685), .Z(n3687) );
  NANDN U4347 ( .A(b[0]), .B(a[36]), .Z(n3686) );
  AND U4348 ( .A(n3687), .B(n3686), .Z(n3755) );
  NAND U4349 ( .A(n19406), .B(n3688), .Z(n3690) );
  XNOR U4350 ( .A(n584), .B(a[9]), .Z(n3844) );
  NANDN U4351 ( .A(n576), .B(n3844), .Z(n3689) );
  NAND U4352 ( .A(n3690), .B(n3689), .Z(n3753) );
  NANDN U4353 ( .A(n585), .B(a[5]), .Z(n3754) );
  XNOR U4354 ( .A(n3753), .B(n3754), .Z(n3756) );
  XOR U4355 ( .A(n3755), .B(n3756), .Z(n3795) );
  XNOR U4356 ( .A(b[23]), .B(a[15]), .Z(n3850) );
  OR U4357 ( .A(n3850), .B(n19127), .Z(n3693) );
  NAND U4358 ( .A(n3691), .B(n19128), .Z(n3692) );
  NAND U4359 ( .A(n3693), .B(n3692), .Z(n3820) );
  NANDN U4360 ( .A(n3694), .B(n17553), .Z(n3696) );
  XOR U4361 ( .A(b[7]), .B(a[31]), .Z(n3853) );
  NAND U4362 ( .A(n3853), .B(n17555), .Z(n3695) );
  NAND U4363 ( .A(n3696), .B(n3695), .Z(n3817) );
  XNOR U4364 ( .A(b[25]), .B(a[13]), .Z(n3856) );
  NANDN U4365 ( .A(n3856), .B(n19240), .Z(n3699) );
  NAND U4366 ( .A(n3697), .B(n19242), .Z(n3698) );
  AND U4367 ( .A(n3699), .B(n3698), .Z(n3818) );
  XNOR U4368 ( .A(n3817), .B(n3818), .Z(n3819) );
  XNOR U4369 ( .A(n3820), .B(n3819), .Z(n3796) );
  XOR U4370 ( .A(n3795), .B(n3796), .Z(n3798) );
  XNOR U4371 ( .A(n3797), .B(n3798), .Z(n3810) );
  XNOR U4372 ( .A(n3809), .B(n3810), .Z(n3865) );
  XNOR U4373 ( .A(n3866), .B(n3865), .Z(n3868) );
  XOR U4374 ( .A(n3867), .B(n3868), .Z(n3747) );
  XOR U4375 ( .A(n3748), .B(n3747), .Z(n3750) );
  NANDN U4376 ( .A(n3701), .B(n3700), .Z(n3705) );
  OR U4377 ( .A(n3703), .B(n3702), .Z(n3704) );
  NAND U4378 ( .A(n3705), .B(n3704), .Z(n3741) );
  NANDN U4379 ( .A(n3707), .B(n3706), .Z(n3711) );
  NAND U4380 ( .A(n3709), .B(n3708), .Z(n3710) );
  NAND U4381 ( .A(n3711), .B(n3710), .Z(n3742) );
  XNOR U4382 ( .A(n3741), .B(n3742), .Z(n3743) );
  XOR U4383 ( .A(n3744), .B(n3743), .Z(n3737) );
  NANDN U4384 ( .A(n3713), .B(n3712), .Z(n3717) );
  NAND U4385 ( .A(n3715), .B(n3714), .Z(n3716) );
  NAND U4386 ( .A(n3717), .B(n3716), .Z(n3735) );
  NANDN U4387 ( .A(n3719), .B(n3718), .Z(n3723) );
  OR U4388 ( .A(n3721), .B(n3720), .Z(n3722) );
  NAND U4389 ( .A(n3723), .B(n3722), .Z(n3736) );
  XNOR U4390 ( .A(n3735), .B(n3736), .Z(n3738) );
  XOR U4391 ( .A(n3737), .B(n3738), .Z(n3729) );
  XOR U4392 ( .A(n3730), .B(n3729), .Z(n3731) );
  XNOR U4393 ( .A(n3732), .B(n3731), .Z(n3869) );
  XNOR U4394 ( .A(n3869), .B(sreg[133]), .Z(n3871) );
  NAND U4395 ( .A(n3724), .B(sreg[132]), .Z(n3728) );
  OR U4396 ( .A(n3726), .B(n3725), .Z(n3727) );
  AND U4397 ( .A(n3728), .B(n3727), .Z(n3870) );
  XOR U4398 ( .A(n3871), .B(n3870), .Z(c[133]) );
  NAND U4399 ( .A(n3730), .B(n3729), .Z(n3734) );
  NAND U4400 ( .A(n3732), .B(n3731), .Z(n3733) );
  NAND U4401 ( .A(n3734), .B(n3733), .Z(n3877) );
  NANDN U4402 ( .A(n3736), .B(n3735), .Z(n3740) );
  NAND U4403 ( .A(n3738), .B(n3737), .Z(n3739) );
  NAND U4404 ( .A(n3740), .B(n3739), .Z(n3875) );
  NANDN U4405 ( .A(n3742), .B(n3741), .Z(n3746) );
  NAND U4406 ( .A(n3744), .B(n3743), .Z(n3745) );
  NAND U4407 ( .A(n3746), .B(n3745), .Z(n3880) );
  NANDN U4408 ( .A(n3748), .B(n3747), .Z(n3752) );
  OR U4409 ( .A(n3750), .B(n3749), .Z(n3751) );
  NAND U4410 ( .A(n3752), .B(n3751), .Z(n3881) );
  XNOR U4411 ( .A(n3880), .B(n3881), .Z(n3882) );
  NANDN U4412 ( .A(n3754), .B(n3753), .Z(n3758) );
  NAND U4413 ( .A(n3756), .B(n3755), .Z(n3757) );
  NAND U4414 ( .A(n3758), .B(n3757), .Z(n3949) );
  NANDN U4415 ( .A(n3759), .B(n18832), .Z(n3761) );
  XNOR U4416 ( .A(b[19]), .B(a[20]), .Z(n3916) );
  NANDN U4417 ( .A(n3916), .B(n18834), .Z(n3760) );
  NAND U4418 ( .A(n3761), .B(n3760), .Z(n3961) );
  XNOR U4419 ( .A(b[27]), .B(a[12]), .Z(n3919) );
  NANDN U4420 ( .A(n3919), .B(n19336), .Z(n3764) );
  NANDN U4421 ( .A(n3762), .B(n19337), .Z(n3763) );
  NAND U4422 ( .A(n3764), .B(n3763), .Z(n3958) );
  XOR U4423 ( .A(b[5]), .B(a[34]), .Z(n3922) );
  NAND U4424 ( .A(n3922), .B(n17310), .Z(n3767) );
  NAND U4425 ( .A(n3765), .B(n17311), .Z(n3766) );
  AND U4426 ( .A(n3767), .B(n3766), .Z(n3959) );
  XNOR U4427 ( .A(n3958), .B(n3959), .Z(n3960) );
  XNOR U4428 ( .A(n3961), .B(n3960), .Z(n3946) );
  XOR U4429 ( .A(b[17]), .B(a[22]), .Z(n3925) );
  NAND U4430 ( .A(n3925), .B(n18673), .Z(n3770) );
  NAND U4431 ( .A(n3768), .B(n18674), .Z(n3769) );
  NAND U4432 ( .A(n3770), .B(n3769), .Z(n3900) );
  XNOR U4433 ( .A(b[31]), .B(a[8]), .Z(n3928) );
  NANDN U4434 ( .A(n3928), .B(n19472), .Z(n3773) );
  NANDN U4435 ( .A(n3771), .B(n19473), .Z(n3772) );
  AND U4436 ( .A(n3773), .B(n3772), .Z(n3898) );
  OR U4437 ( .A(n3774), .B(n16988), .Z(n3776) );
  XNOR U4438 ( .A(b[3]), .B(a[36]), .Z(n3931) );
  NANDN U4439 ( .A(n3931), .B(n16990), .Z(n3775) );
  AND U4440 ( .A(n3776), .B(n3775), .Z(n3899) );
  XOR U4441 ( .A(n3900), .B(n3901), .Z(n3947) );
  XOR U4442 ( .A(n3946), .B(n3947), .Z(n3948) );
  XNOR U4443 ( .A(n3949), .B(n3948), .Z(n3994) );
  NANDN U4444 ( .A(n3778), .B(n3777), .Z(n3782) );
  NAND U4445 ( .A(n3780), .B(n3779), .Z(n3781) );
  NAND U4446 ( .A(n3782), .B(n3781), .Z(n3937) );
  NANDN U4447 ( .A(n3784), .B(n3783), .Z(n3788) );
  NAND U4448 ( .A(n3786), .B(n3785), .Z(n3787) );
  NAND U4449 ( .A(n3788), .B(n3787), .Z(n3935) );
  OR U4450 ( .A(n3790), .B(n3789), .Z(n3794) );
  NANDN U4451 ( .A(n3792), .B(n3791), .Z(n3793) );
  NAND U4452 ( .A(n3794), .B(n3793), .Z(n3934) );
  XNOR U4453 ( .A(n3937), .B(n3936), .Z(n3995) );
  XOR U4454 ( .A(n3994), .B(n3995), .Z(n3997) );
  NANDN U4455 ( .A(n3796), .B(n3795), .Z(n3800) );
  OR U4456 ( .A(n3798), .B(n3797), .Z(n3799) );
  NAND U4457 ( .A(n3800), .B(n3799), .Z(n3996) );
  XOR U4458 ( .A(n3997), .B(n3996), .Z(n4014) );
  OR U4459 ( .A(n3802), .B(n3801), .Z(n3806) );
  NAND U4460 ( .A(n3804), .B(n3803), .Z(n3805) );
  NAND U4461 ( .A(n3806), .B(n3805), .Z(n4013) );
  NANDN U4462 ( .A(n3808), .B(n3807), .Z(n3812) );
  NANDN U4463 ( .A(n3810), .B(n3809), .Z(n3811) );
  NAND U4464 ( .A(n3812), .B(n3811), .Z(n4002) );
  NANDN U4465 ( .A(n3818), .B(n3817), .Z(n3822) );
  NAND U4466 ( .A(n3820), .B(n3819), .Z(n3821) );
  NAND U4467 ( .A(n3822), .B(n3821), .Z(n3940) );
  NANDN U4468 ( .A(n3824), .B(n3823), .Z(n3828) );
  NAND U4469 ( .A(n3826), .B(n3825), .Z(n3827) );
  AND U4470 ( .A(n3828), .B(n3827), .Z(n3941) );
  XNOR U4471 ( .A(n3940), .B(n3941), .Z(n3942) );
  XOR U4472 ( .A(b[9]), .B(n7336), .Z(n3964) );
  NANDN U4473 ( .A(n3964), .B(n17814), .Z(n3831) );
  NANDN U4474 ( .A(n3829), .B(n17815), .Z(n3830) );
  NAND U4475 ( .A(n3831), .B(n3830), .Z(n3906) );
  NAND U4476 ( .A(n3832), .B(n18513), .Z(n3834) );
  XOR U4477 ( .A(b[15]), .B(a[24]), .Z(n3967) );
  NANDN U4478 ( .A(n18512), .B(n3967), .Z(n3833) );
  AND U4479 ( .A(n3834), .B(n3833), .Z(n3904) );
  NANDN U4480 ( .A(n3835), .B(n19013), .Z(n3837) );
  XNOR U4481 ( .A(b[21]), .B(a[18]), .Z(n3970) );
  NANDN U4482 ( .A(n3970), .B(n19015), .Z(n3836) );
  AND U4483 ( .A(n3837), .B(n3836), .Z(n3905) );
  XOR U4484 ( .A(n3906), .B(n3907), .Z(n3895) );
  XNOR U4485 ( .A(b[11]), .B(a[28]), .Z(n3973) );
  OR U4486 ( .A(n3973), .B(n18194), .Z(n3840) );
  NANDN U4487 ( .A(n3838), .B(n18104), .Z(n3839) );
  NAND U4488 ( .A(n3840), .B(n3839), .Z(n3893) );
  XOR U4489 ( .A(n580), .B(a[26]), .Z(n3976) );
  NANDN U4490 ( .A(n3976), .B(n18336), .Z(n3843) );
  NANDN U4491 ( .A(n3841), .B(n18337), .Z(n3842) );
  NAND U4492 ( .A(n3843), .B(n3842), .Z(n3892) );
  XOR U4493 ( .A(n3895), .B(n3894), .Z(n3889) );
  NAND U4494 ( .A(n19406), .B(n3844), .Z(n3846) );
  XNOR U4495 ( .A(n584), .B(a[10]), .Z(n3982) );
  NANDN U4496 ( .A(n576), .B(n3982), .Z(n3845) );
  NAND U4497 ( .A(n3846), .B(n3845), .Z(n3910) );
  NANDN U4498 ( .A(n585), .B(a[6]), .Z(n3911) );
  XNOR U4499 ( .A(n3910), .B(n3911), .Z(n3913) );
  NANDN U4500 ( .A(n577), .B(a[38]), .Z(n3847) );
  XOR U4501 ( .A(n17151), .B(n3847), .Z(n3849) );
  NANDN U4502 ( .A(b[0]), .B(a[37]), .Z(n3848) );
  AND U4503 ( .A(n3849), .B(n3848), .Z(n3912) );
  XNOR U4504 ( .A(n3913), .B(n3912), .Z(n3887) );
  XOR U4505 ( .A(b[23]), .B(a[16]), .Z(n3985) );
  NANDN U4506 ( .A(n19127), .B(n3985), .Z(n3852) );
  NANDN U4507 ( .A(n3850), .B(n19128), .Z(n3851) );
  NAND U4508 ( .A(n3852), .B(n3851), .Z(n3955) );
  NAND U4509 ( .A(n3853), .B(n17553), .Z(n3855) );
  XOR U4510 ( .A(b[7]), .B(a[32]), .Z(n3988) );
  NAND U4511 ( .A(n3988), .B(n17555), .Z(n3854) );
  NAND U4512 ( .A(n3855), .B(n3854), .Z(n3952) );
  XOR U4513 ( .A(b[25]), .B(a[14]), .Z(n3991) );
  NAND U4514 ( .A(n3991), .B(n19240), .Z(n3858) );
  NANDN U4515 ( .A(n3856), .B(n19242), .Z(n3857) );
  AND U4516 ( .A(n3858), .B(n3857), .Z(n3953) );
  XNOR U4517 ( .A(n3952), .B(n3953), .Z(n3954) );
  XOR U4518 ( .A(n3955), .B(n3954), .Z(n3886) );
  XOR U4519 ( .A(n3889), .B(n3888), .Z(n3943) );
  XNOR U4520 ( .A(n3942), .B(n3943), .Z(n4000) );
  XNOR U4521 ( .A(n4001), .B(n4000), .Z(n4003) );
  XNOR U4522 ( .A(n4002), .B(n4003), .Z(n4012) );
  XOR U4523 ( .A(n4013), .B(n4012), .Z(n4015) );
  NANDN U4524 ( .A(n3860), .B(n3859), .Z(n3864) );
  OR U4525 ( .A(n3862), .B(n3861), .Z(n3863) );
  NAND U4526 ( .A(n3864), .B(n3863), .Z(n4006) );
  XNOR U4527 ( .A(n4006), .B(n4007), .Z(n4008) );
  XOR U4528 ( .A(n4009), .B(n4008), .Z(n3883) );
  XOR U4529 ( .A(n3882), .B(n3883), .Z(n3874) );
  XOR U4530 ( .A(n3875), .B(n3874), .Z(n3876) );
  XNOR U4531 ( .A(n3877), .B(n3876), .Z(n4018) );
  XNOR U4532 ( .A(n4018), .B(sreg[134]), .Z(n4020) );
  NAND U4533 ( .A(n3869), .B(sreg[133]), .Z(n3873) );
  OR U4534 ( .A(n3871), .B(n3870), .Z(n3872) );
  AND U4535 ( .A(n3873), .B(n3872), .Z(n4019) );
  XOR U4536 ( .A(n4020), .B(n4019), .Z(c[134]) );
  NAND U4537 ( .A(n3875), .B(n3874), .Z(n3879) );
  NAND U4538 ( .A(n3877), .B(n3876), .Z(n3878) );
  NAND U4539 ( .A(n3879), .B(n3878), .Z(n4026) );
  NANDN U4540 ( .A(n3881), .B(n3880), .Z(n3885) );
  NAND U4541 ( .A(n3883), .B(n3882), .Z(n3884) );
  NAND U4542 ( .A(n3885), .B(n3884), .Z(n4024) );
  NANDN U4543 ( .A(n3887), .B(n3886), .Z(n3891) );
  NANDN U4544 ( .A(n3889), .B(n3888), .Z(n3890) );
  NAND U4545 ( .A(n3891), .B(n3890), .Z(n4144) );
  OR U4546 ( .A(n3893), .B(n3892), .Z(n3897) );
  NAND U4547 ( .A(n3895), .B(n3894), .Z(n3896) );
  NAND U4548 ( .A(n3897), .B(n3896), .Z(n4083) );
  OR U4549 ( .A(n3899), .B(n3898), .Z(n3903) );
  NANDN U4550 ( .A(n3901), .B(n3900), .Z(n3902) );
  NAND U4551 ( .A(n3903), .B(n3902), .Z(n4082) );
  OR U4552 ( .A(n3905), .B(n3904), .Z(n3909) );
  NANDN U4553 ( .A(n3907), .B(n3906), .Z(n3908) );
  NAND U4554 ( .A(n3909), .B(n3908), .Z(n4081) );
  XOR U4555 ( .A(n4083), .B(n4084), .Z(n4141) );
  NANDN U4556 ( .A(n3911), .B(n3910), .Z(n3915) );
  NAND U4557 ( .A(n3913), .B(n3912), .Z(n3914) );
  NAND U4558 ( .A(n3915), .B(n3914), .Z(n4096) );
  NANDN U4559 ( .A(n3916), .B(n18832), .Z(n3918) );
  XNOR U4560 ( .A(b[19]), .B(a[21]), .Z(n4063) );
  NANDN U4561 ( .A(n4063), .B(n18834), .Z(n3917) );
  NAND U4562 ( .A(n3918), .B(n3917), .Z(n4108) );
  XOR U4563 ( .A(b[27]), .B(n4875), .Z(n4066) );
  NANDN U4564 ( .A(n4066), .B(n19336), .Z(n3921) );
  NANDN U4565 ( .A(n3919), .B(n19337), .Z(n3920) );
  NAND U4566 ( .A(n3921), .B(n3920), .Z(n4105) );
  XOR U4567 ( .A(b[5]), .B(a[35]), .Z(n4069) );
  NAND U4568 ( .A(n4069), .B(n17310), .Z(n3924) );
  NAND U4569 ( .A(n3922), .B(n17311), .Z(n3923) );
  AND U4570 ( .A(n3924), .B(n3923), .Z(n4106) );
  XNOR U4571 ( .A(n4105), .B(n4106), .Z(n4107) );
  XNOR U4572 ( .A(n4108), .B(n4107), .Z(n4093) );
  XOR U4573 ( .A(b[17]), .B(a[23]), .Z(n4072) );
  NAND U4574 ( .A(n4072), .B(n18673), .Z(n3927) );
  NAND U4575 ( .A(n3925), .B(n18674), .Z(n3926) );
  NAND U4576 ( .A(n3927), .B(n3926), .Z(n4047) );
  XNOR U4577 ( .A(b[31]), .B(a[9]), .Z(n4075) );
  NANDN U4578 ( .A(n4075), .B(n19472), .Z(n3930) );
  NANDN U4579 ( .A(n3928), .B(n19473), .Z(n3929) );
  AND U4580 ( .A(n3930), .B(n3929), .Z(n4045) );
  OR U4581 ( .A(n3931), .B(n16988), .Z(n3933) );
  XNOR U4582 ( .A(b[3]), .B(a[37]), .Z(n4078) );
  NANDN U4583 ( .A(n4078), .B(n16990), .Z(n3932) );
  AND U4584 ( .A(n3933), .B(n3932), .Z(n4046) );
  XOR U4585 ( .A(n4047), .B(n4048), .Z(n4094) );
  XOR U4586 ( .A(n4093), .B(n4094), .Z(n4095) );
  XNOR U4587 ( .A(n4096), .B(n4095), .Z(n4142) );
  XNOR U4588 ( .A(n4141), .B(n4142), .Z(n4143) );
  XNOR U4589 ( .A(n4144), .B(n4143), .Z(n4162) );
  OR U4590 ( .A(n3935), .B(n3934), .Z(n3939) );
  NAND U4591 ( .A(n3937), .B(n3936), .Z(n3938) );
  NAND U4592 ( .A(n3939), .B(n3938), .Z(n4160) );
  NANDN U4593 ( .A(n3941), .B(n3940), .Z(n3945) );
  NANDN U4594 ( .A(n3943), .B(n3942), .Z(n3944) );
  NAND U4595 ( .A(n3945), .B(n3944), .Z(n4149) );
  OR U4596 ( .A(n3947), .B(n3946), .Z(n3951) );
  NAND U4597 ( .A(n3949), .B(n3948), .Z(n3950) );
  NAND U4598 ( .A(n3951), .B(n3950), .Z(n4148) );
  NANDN U4599 ( .A(n3953), .B(n3952), .Z(n3957) );
  NAND U4600 ( .A(n3955), .B(n3954), .Z(n3956) );
  NAND U4601 ( .A(n3957), .B(n3956), .Z(n4087) );
  NANDN U4602 ( .A(n3959), .B(n3958), .Z(n3963) );
  NAND U4603 ( .A(n3961), .B(n3960), .Z(n3962) );
  AND U4604 ( .A(n3963), .B(n3962), .Z(n4088) );
  XNOR U4605 ( .A(n4087), .B(n4088), .Z(n4089) );
  XNOR U4606 ( .A(n579), .B(a[31]), .Z(n4111) );
  NAND U4607 ( .A(n17814), .B(n4111), .Z(n3966) );
  NANDN U4608 ( .A(n3964), .B(n17815), .Z(n3965) );
  NAND U4609 ( .A(n3966), .B(n3965), .Z(n4053) );
  NAND U4610 ( .A(n3967), .B(n18513), .Z(n3969) );
  XOR U4611 ( .A(b[15]), .B(a[25]), .Z(n4114) );
  NANDN U4612 ( .A(n18512), .B(n4114), .Z(n3968) );
  AND U4613 ( .A(n3969), .B(n3968), .Z(n4051) );
  NANDN U4614 ( .A(n3970), .B(n19013), .Z(n3972) );
  XNOR U4615 ( .A(n582), .B(a[19]), .Z(n4117) );
  NAND U4616 ( .A(n4117), .B(n19015), .Z(n3971) );
  AND U4617 ( .A(n3972), .B(n3971), .Z(n4052) );
  XOR U4618 ( .A(n4053), .B(n4054), .Z(n4042) );
  XOR U4619 ( .A(b[11]), .B(n6835), .Z(n4120) );
  OR U4620 ( .A(n4120), .B(n18194), .Z(n3975) );
  NANDN U4621 ( .A(n3973), .B(n18104), .Z(n3974) );
  NAND U4622 ( .A(n3975), .B(n3974), .Z(n4040) );
  XOR U4623 ( .A(n580), .B(a[27]), .Z(n4123) );
  NANDN U4624 ( .A(n4123), .B(n18336), .Z(n3978) );
  NANDN U4625 ( .A(n3976), .B(n18337), .Z(n3977) );
  NAND U4626 ( .A(n3978), .B(n3977), .Z(n4039) );
  XOR U4627 ( .A(n4042), .B(n4041), .Z(n4036) );
  NANDN U4628 ( .A(n577), .B(a[39]), .Z(n3979) );
  XOR U4629 ( .A(n17151), .B(n3979), .Z(n3981) );
  IV U4630 ( .A(a[38]), .Z(n8490) );
  NANDN U4631 ( .A(n8490), .B(n577), .Z(n3980) );
  AND U4632 ( .A(n3981), .B(n3980), .Z(n4059) );
  NAND U4633 ( .A(n19406), .B(n3982), .Z(n3984) );
  XOR U4634 ( .A(n584), .B(n4573), .Z(n4129) );
  NANDN U4635 ( .A(n576), .B(n4129), .Z(n3983) );
  NAND U4636 ( .A(n3984), .B(n3983), .Z(n4057) );
  NANDN U4637 ( .A(n585), .B(a[7]), .Z(n4058) );
  XNOR U4638 ( .A(n4057), .B(n4058), .Z(n4060) );
  XNOR U4639 ( .A(n4059), .B(n4060), .Z(n4034) );
  XOR U4640 ( .A(b[23]), .B(a[17]), .Z(n4132) );
  NANDN U4641 ( .A(n19127), .B(n4132), .Z(n3987) );
  NAND U4642 ( .A(n3985), .B(n19128), .Z(n3986) );
  NAND U4643 ( .A(n3987), .B(n3986), .Z(n4102) );
  NAND U4644 ( .A(n3988), .B(n17553), .Z(n3990) );
  XOR U4645 ( .A(b[7]), .B(a[33]), .Z(n4135) );
  NAND U4646 ( .A(n4135), .B(n17555), .Z(n3989) );
  NAND U4647 ( .A(n3990), .B(n3989), .Z(n4099) );
  XNOR U4648 ( .A(b[25]), .B(a[15]), .Z(n4138) );
  NANDN U4649 ( .A(n4138), .B(n19240), .Z(n3993) );
  NAND U4650 ( .A(n3991), .B(n19242), .Z(n3992) );
  AND U4651 ( .A(n3993), .B(n3992), .Z(n4100) );
  XNOR U4652 ( .A(n4099), .B(n4100), .Z(n4101) );
  XOR U4653 ( .A(n4102), .B(n4101), .Z(n4033) );
  XOR U4654 ( .A(n4036), .B(n4035), .Z(n4090) );
  XNOR U4655 ( .A(n4089), .B(n4090), .Z(n4147) );
  XNOR U4656 ( .A(n4148), .B(n4147), .Z(n4150) );
  XNOR U4657 ( .A(n4149), .B(n4150), .Z(n4159) );
  XNOR U4658 ( .A(n4160), .B(n4159), .Z(n4161) );
  XOR U4659 ( .A(n4162), .B(n4161), .Z(n4156) );
  NANDN U4660 ( .A(n3995), .B(n3994), .Z(n3999) );
  OR U4661 ( .A(n3997), .B(n3996), .Z(n3998) );
  NAND U4662 ( .A(n3999), .B(n3998), .Z(n4153) );
  NAND U4663 ( .A(n4001), .B(n4000), .Z(n4005) );
  NANDN U4664 ( .A(n4003), .B(n4002), .Z(n4004) );
  NAND U4665 ( .A(n4005), .B(n4004), .Z(n4154) );
  XNOR U4666 ( .A(n4153), .B(n4154), .Z(n4155) );
  XNOR U4667 ( .A(n4156), .B(n4155), .Z(n4030) );
  NANDN U4668 ( .A(n4007), .B(n4006), .Z(n4011) );
  NAND U4669 ( .A(n4009), .B(n4008), .Z(n4010) );
  NAND U4670 ( .A(n4011), .B(n4010), .Z(n4027) );
  NANDN U4671 ( .A(n4013), .B(n4012), .Z(n4017) );
  OR U4672 ( .A(n4015), .B(n4014), .Z(n4016) );
  NAND U4673 ( .A(n4017), .B(n4016), .Z(n4028) );
  XNOR U4674 ( .A(n4027), .B(n4028), .Z(n4029) );
  XNOR U4675 ( .A(n4030), .B(n4029), .Z(n4023) );
  XOR U4676 ( .A(n4024), .B(n4023), .Z(n4025) );
  XNOR U4677 ( .A(n4026), .B(n4025), .Z(n4165) );
  XNOR U4678 ( .A(n4165), .B(sreg[135]), .Z(n4167) );
  NAND U4679 ( .A(n4018), .B(sreg[134]), .Z(n4022) );
  OR U4680 ( .A(n4020), .B(n4019), .Z(n4021) );
  AND U4681 ( .A(n4022), .B(n4021), .Z(n4166) );
  XOR U4682 ( .A(n4167), .B(n4166), .Z(c[135]) );
  NANDN U4683 ( .A(n4028), .B(n4027), .Z(n4032) );
  NANDN U4684 ( .A(n4030), .B(n4029), .Z(n4031) );
  NAND U4685 ( .A(n4032), .B(n4031), .Z(n4171) );
  NANDN U4686 ( .A(n4034), .B(n4033), .Z(n4038) );
  NANDN U4687 ( .A(n4036), .B(n4035), .Z(n4037) );
  NAND U4688 ( .A(n4038), .B(n4037), .Z(n4301) );
  OR U4689 ( .A(n4040), .B(n4039), .Z(n4044) );
  NAND U4690 ( .A(n4042), .B(n4041), .Z(n4043) );
  NAND U4691 ( .A(n4044), .B(n4043), .Z(n4240) );
  OR U4692 ( .A(n4046), .B(n4045), .Z(n4050) );
  NANDN U4693 ( .A(n4048), .B(n4047), .Z(n4049) );
  NAND U4694 ( .A(n4050), .B(n4049), .Z(n4239) );
  OR U4695 ( .A(n4052), .B(n4051), .Z(n4056) );
  NANDN U4696 ( .A(n4054), .B(n4053), .Z(n4055) );
  NAND U4697 ( .A(n4056), .B(n4055), .Z(n4238) );
  XOR U4698 ( .A(n4240), .B(n4241), .Z(n4298) );
  NANDN U4699 ( .A(n4058), .B(n4057), .Z(n4062) );
  NAND U4700 ( .A(n4060), .B(n4059), .Z(n4061) );
  NAND U4701 ( .A(n4062), .B(n4061), .Z(n4253) );
  NANDN U4702 ( .A(n4063), .B(n18832), .Z(n4065) );
  XNOR U4703 ( .A(b[19]), .B(a[22]), .Z(n4198) );
  NANDN U4704 ( .A(n4198), .B(n18834), .Z(n4064) );
  NAND U4705 ( .A(n4065), .B(n4064), .Z(n4265) );
  XNOR U4706 ( .A(b[27]), .B(a[14]), .Z(n4201) );
  NANDN U4707 ( .A(n4201), .B(n19336), .Z(n4068) );
  NANDN U4708 ( .A(n4066), .B(n19337), .Z(n4067) );
  NAND U4709 ( .A(n4068), .B(n4067), .Z(n4262) );
  XOR U4710 ( .A(b[5]), .B(a[36]), .Z(n4204) );
  NAND U4711 ( .A(n4204), .B(n17310), .Z(n4071) );
  NAND U4712 ( .A(n4069), .B(n17311), .Z(n4070) );
  AND U4713 ( .A(n4071), .B(n4070), .Z(n4263) );
  XNOR U4714 ( .A(n4262), .B(n4263), .Z(n4264) );
  XNOR U4715 ( .A(n4265), .B(n4264), .Z(n4251) );
  XOR U4716 ( .A(b[17]), .B(a[24]), .Z(n4207) );
  NAND U4717 ( .A(n4207), .B(n18673), .Z(n4074) );
  NAND U4718 ( .A(n4072), .B(n18674), .Z(n4073) );
  NAND U4719 ( .A(n4074), .B(n4073), .Z(n4225) );
  XNOR U4720 ( .A(b[31]), .B(a[10]), .Z(n4210) );
  NANDN U4721 ( .A(n4210), .B(n19472), .Z(n4077) );
  NANDN U4722 ( .A(n4075), .B(n19473), .Z(n4076) );
  NAND U4723 ( .A(n4077), .B(n4076), .Z(n4222) );
  OR U4724 ( .A(n4078), .B(n16988), .Z(n4080) );
  XOR U4725 ( .A(b[3]), .B(n8490), .Z(n4213) );
  NANDN U4726 ( .A(n4213), .B(n16990), .Z(n4079) );
  AND U4727 ( .A(n4080), .B(n4079), .Z(n4223) );
  XNOR U4728 ( .A(n4222), .B(n4223), .Z(n4224) );
  XOR U4729 ( .A(n4225), .B(n4224), .Z(n4250) );
  XNOR U4730 ( .A(n4251), .B(n4250), .Z(n4252) );
  XNOR U4731 ( .A(n4253), .B(n4252), .Z(n4299) );
  XNOR U4732 ( .A(n4298), .B(n4299), .Z(n4300) );
  XNOR U4733 ( .A(n4301), .B(n4300), .Z(n4189) );
  OR U4734 ( .A(n4082), .B(n4081), .Z(n4086) );
  NANDN U4735 ( .A(n4084), .B(n4083), .Z(n4085) );
  NAND U4736 ( .A(n4086), .B(n4085), .Z(n4187) );
  NANDN U4737 ( .A(n4088), .B(n4087), .Z(n4092) );
  NANDN U4738 ( .A(n4090), .B(n4089), .Z(n4091) );
  NAND U4739 ( .A(n4092), .B(n4091), .Z(n4306) );
  OR U4740 ( .A(n4094), .B(n4093), .Z(n4098) );
  NAND U4741 ( .A(n4096), .B(n4095), .Z(n4097) );
  NAND U4742 ( .A(n4098), .B(n4097), .Z(n4305) );
  NANDN U4743 ( .A(n4100), .B(n4099), .Z(n4104) );
  NAND U4744 ( .A(n4102), .B(n4101), .Z(n4103) );
  NAND U4745 ( .A(n4104), .B(n4103), .Z(n4244) );
  NANDN U4746 ( .A(n4106), .B(n4105), .Z(n4110) );
  NAND U4747 ( .A(n4108), .B(n4107), .Z(n4109) );
  AND U4748 ( .A(n4110), .B(n4109), .Z(n4245) );
  XNOR U4749 ( .A(n4244), .B(n4245), .Z(n4246) );
  XNOR U4750 ( .A(b[9]), .B(a[32]), .Z(n4268) );
  NANDN U4751 ( .A(n4268), .B(n17814), .Z(n4113) );
  NAND U4752 ( .A(n17815), .B(n4111), .Z(n4112) );
  NAND U4753 ( .A(n4113), .B(n4112), .Z(n4230) );
  XNOR U4754 ( .A(b[15]), .B(a[26]), .Z(n4271) );
  OR U4755 ( .A(n4271), .B(n18512), .Z(n4116) );
  NAND U4756 ( .A(n4114), .B(n18513), .Z(n4115) );
  NAND U4757 ( .A(n4116), .B(n4115), .Z(n4228) );
  XNOR U4758 ( .A(b[21]), .B(a[20]), .Z(n4274) );
  NANDN U4759 ( .A(n4274), .B(n19015), .Z(n4119) );
  NAND U4760 ( .A(n19013), .B(n4117), .Z(n4118) );
  NAND U4761 ( .A(n4119), .B(n4118), .Z(n4229) );
  XNOR U4762 ( .A(n4228), .B(n4229), .Z(n4231) );
  XOR U4763 ( .A(n4230), .B(n4231), .Z(n4219) );
  XOR U4764 ( .A(b[11]), .B(n7336), .Z(n4277) );
  OR U4765 ( .A(n4277), .B(n18194), .Z(n4122) );
  NANDN U4766 ( .A(n4120), .B(n18104), .Z(n4121) );
  NAND U4767 ( .A(n4122), .B(n4121), .Z(n4217) );
  XOR U4768 ( .A(n580), .B(a[28]), .Z(n4280) );
  NANDN U4769 ( .A(n4280), .B(n18336), .Z(n4125) );
  NANDN U4770 ( .A(n4123), .B(n18337), .Z(n4124) );
  AND U4771 ( .A(n4125), .B(n4124), .Z(n4216) );
  XNOR U4772 ( .A(n4217), .B(n4216), .Z(n4218) );
  XNOR U4773 ( .A(n4219), .B(n4218), .Z(n4235) );
  NANDN U4774 ( .A(n577), .B(a[40]), .Z(n4126) );
  XOR U4775 ( .A(n17151), .B(n4126), .Z(n4128) );
  NANDN U4776 ( .A(b[0]), .B(a[39]), .Z(n4127) );
  AND U4777 ( .A(n4128), .B(n4127), .Z(n4194) );
  NAND U4778 ( .A(n19406), .B(n4129), .Z(n4131) );
  XNOR U4779 ( .A(n584), .B(a[12]), .Z(n4283) );
  NANDN U4780 ( .A(n576), .B(n4283), .Z(n4130) );
  NAND U4781 ( .A(n4131), .B(n4130), .Z(n4192) );
  NANDN U4782 ( .A(n585), .B(a[8]), .Z(n4193) );
  XNOR U4783 ( .A(n4192), .B(n4193), .Z(n4195) );
  XNOR U4784 ( .A(n4194), .B(n4195), .Z(n4233) );
  XOR U4785 ( .A(b[23]), .B(a[18]), .Z(n4289) );
  NANDN U4786 ( .A(n19127), .B(n4289), .Z(n4134) );
  NAND U4787 ( .A(n4132), .B(n19128), .Z(n4133) );
  NAND U4788 ( .A(n4134), .B(n4133), .Z(n4259) );
  NAND U4789 ( .A(n4135), .B(n17553), .Z(n4137) );
  XOR U4790 ( .A(b[7]), .B(a[34]), .Z(n4292) );
  NAND U4791 ( .A(n4292), .B(n17555), .Z(n4136) );
  NAND U4792 ( .A(n4137), .B(n4136), .Z(n4256) );
  XOR U4793 ( .A(b[25]), .B(a[16]), .Z(n4295) );
  NAND U4794 ( .A(n4295), .B(n19240), .Z(n4140) );
  NANDN U4795 ( .A(n4138), .B(n19242), .Z(n4139) );
  AND U4796 ( .A(n4140), .B(n4139), .Z(n4257) );
  XNOR U4797 ( .A(n4256), .B(n4257), .Z(n4258) );
  XOR U4798 ( .A(n4259), .B(n4258), .Z(n4232) );
  XOR U4799 ( .A(n4235), .B(n4234), .Z(n4247) );
  XOR U4800 ( .A(n4246), .B(n4247), .Z(n4304) );
  XNOR U4801 ( .A(n4305), .B(n4304), .Z(n4307) );
  XNOR U4802 ( .A(n4306), .B(n4307), .Z(n4186) );
  XNOR U4803 ( .A(n4187), .B(n4186), .Z(n4188) );
  XOR U4804 ( .A(n4189), .B(n4188), .Z(n4183) );
  NANDN U4805 ( .A(n4142), .B(n4141), .Z(n4146) );
  NAND U4806 ( .A(n4144), .B(n4143), .Z(n4145) );
  NAND U4807 ( .A(n4146), .B(n4145), .Z(n4181) );
  NAND U4808 ( .A(n4148), .B(n4147), .Z(n4152) );
  NANDN U4809 ( .A(n4150), .B(n4149), .Z(n4151) );
  AND U4810 ( .A(n4152), .B(n4151), .Z(n4180) );
  XNOR U4811 ( .A(n4181), .B(n4180), .Z(n4182) );
  XNOR U4812 ( .A(n4183), .B(n4182), .Z(n4177) );
  NANDN U4813 ( .A(n4154), .B(n4153), .Z(n4158) );
  NAND U4814 ( .A(n4156), .B(n4155), .Z(n4157) );
  NAND U4815 ( .A(n4158), .B(n4157), .Z(n4174) );
  NANDN U4816 ( .A(n4160), .B(n4159), .Z(n4164) );
  NANDN U4817 ( .A(n4162), .B(n4161), .Z(n4163) );
  NAND U4818 ( .A(n4164), .B(n4163), .Z(n4175) );
  XNOR U4819 ( .A(n4174), .B(n4175), .Z(n4176) );
  XNOR U4820 ( .A(n4177), .B(n4176), .Z(n4170) );
  XOR U4821 ( .A(n4171), .B(n4170), .Z(n4172) );
  XNOR U4822 ( .A(n4173), .B(n4172), .Z(n4310) );
  XNOR U4823 ( .A(n4310), .B(sreg[136]), .Z(n4312) );
  NAND U4824 ( .A(n4165), .B(sreg[135]), .Z(n4169) );
  OR U4825 ( .A(n4167), .B(n4166), .Z(n4168) );
  AND U4826 ( .A(n4169), .B(n4168), .Z(n4311) );
  XOR U4827 ( .A(n4312), .B(n4311), .Z(c[136]) );
  NANDN U4828 ( .A(n4175), .B(n4174), .Z(n4179) );
  NANDN U4829 ( .A(n4177), .B(n4176), .Z(n4178) );
  NAND U4830 ( .A(n4179), .B(n4178), .Z(n4316) );
  NANDN U4831 ( .A(n4181), .B(n4180), .Z(n4185) );
  NAND U4832 ( .A(n4183), .B(n4182), .Z(n4184) );
  NAND U4833 ( .A(n4185), .B(n4184), .Z(n4321) );
  NANDN U4834 ( .A(n4187), .B(n4186), .Z(n4191) );
  NANDN U4835 ( .A(n4189), .B(n4188), .Z(n4190) );
  NAND U4836 ( .A(n4191), .B(n4190), .Z(n4322) );
  XNOR U4837 ( .A(n4321), .B(n4322), .Z(n4323) );
  NANDN U4838 ( .A(n4193), .B(n4192), .Z(n4197) );
  NAND U4839 ( .A(n4195), .B(n4194), .Z(n4196) );
  NAND U4840 ( .A(n4197), .B(n4196), .Z(n4398) );
  NANDN U4841 ( .A(n4198), .B(n18832), .Z(n4200) );
  XNOR U4842 ( .A(b[19]), .B(a[23]), .Z(n4343) );
  NANDN U4843 ( .A(n4343), .B(n18834), .Z(n4199) );
  NAND U4844 ( .A(n4200), .B(n4199), .Z(n4408) );
  XOR U4845 ( .A(b[27]), .B(n5159), .Z(n4346) );
  NANDN U4846 ( .A(n4346), .B(n19336), .Z(n4203) );
  NANDN U4847 ( .A(n4201), .B(n19337), .Z(n4202) );
  NAND U4848 ( .A(n4203), .B(n4202), .Z(n4405) );
  XOR U4849 ( .A(b[5]), .B(a[37]), .Z(n4349) );
  NAND U4850 ( .A(n4349), .B(n17310), .Z(n4206) );
  NAND U4851 ( .A(n4204), .B(n17311), .Z(n4205) );
  AND U4852 ( .A(n4206), .B(n4205), .Z(n4406) );
  XNOR U4853 ( .A(n4405), .B(n4406), .Z(n4407) );
  XNOR U4854 ( .A(n4408), .B(n4407), .Z(n4396) );
  XOR U4855 ( .A(b[17]), .B(a[25]), .Z(n4352) );
  NAND U4856 ( .A(n4352), .B(n18673), .Z(n4209) );
  NAND U4857 ( .A(n4207), .B(n18674), .Z(n4208) );
  NAND U4858 ( .A(n4209), .B(n4208), .Z(n4370) );
  XOR U4859 ( .A(b[31]), .B(n4573), .Z(n4355) );
  NANDN U4860 ( .A(n4355), .B(n19472), .Z(n4212) );
  NANDN U4861 ( .A(n4210), .B(n19473), .Z(n4211) );
  NAND U4862 ( .A(n4212), .B(n4211), .Z(n4367) );
  OR U4863 ( .A(n4213), .B(n16988), .Z(n4215) );
  XNOR U4864 ( .A(b[3]), .B(a[39]), .Z(n4358) );
  NANDN U4865 ( .A(n4358), .B(n16990), .Z(n4214) );
  AND U4866 ( .A(n4215), .B(n4214), .Z(n4368) );
  XNOR U4867 ( .A(n4367), .B(n4368), .Z(n4369) );
  XOR U4868 ( .A(n4370), .B(n4369), .Z(n4395) );
  XNOR U4869 ( .A(n4396), .B(n4395), .Z(n4397) );
  XNOR U4870 ( .A(n4398), .B(n4397), .Z(n4334) );
  NANDN U4871 ( .A(n4217), .B(n4216), .Z(n4221) );
  NAND U4872 ( .A(n4219), .B(n4218), .Z(n4220) );
  NAND U4873 ( .A(n4221), .B(n4220), .Z(n4387) );
  NANDN U4874 ( .A(n4223), .B(n4222), .Z(n4227) );
  NAND U4875 ( .A(n4225), .B(n4224), .Z(n4226) );
  NAND U4876 ( .A(n4227), .B(n4226), .Z(n4386) );
  XNOR U4877 ( .A(n4386), .B(n4385), .Z(n4388) );
  XOR U4878 ( .A(n4387), .B(n4388), .Z(n4333) );
  XOR U4879 ( .A(n4334), .B(n4333), .Z(n4335) );
  NANDN U4880 ( .A(n4233), .B(n4232), .Z(n4237) );
  NAND U4881 ( .A(n4235), .B(n4234), .Z(n4236) );
  NAND U4882 ( .A(n4237), .B(n4236), .Z(n4336) );
  XNOR U4883 ( .A(n4335), .B(n4336), .Z(n4449) );
  OR U4884 ( .A(n4239), .B(n4238), .Z(n4243) );
  NANDN U4885 ( .A(n4241), .B(n4240), .Z(n4242) );
  NAND U4886 ( .A(n4243), .B(n4242), .Z(n4448) );
  NANDN U4887 ( .A(n4245), .B(n4244), .Z(n4249) );
  NAND U4888 ( .A(n4247), .B(n4246), .Z(n4248) );
  NAND U4889 ( .A(n4249), .B(n4248), .Z(n4329) );
  NANDN U4890 ( .A(n4251), .B(n4250), .Z(n4255) );
  NAND U4891 ( .A(n4253), .B(n4252), .Z(n4254) );
  NAND U4892 ( .A(n4255), .B(n4254), .Z(n4328) );
  NANDN U4893 ( .A(n4257), .B(n4256), .Z(n4261) );
  NAND U4894 ( .A(n4259), .B(n4258), .Z(n4260) );
  NAND U4895 ( .A(n4261), .B(n4260), .Z(n4389) );
  NANDN U4896 ( .A(n4263), .B(n4262), .Z(n4267) );
  NAND U4897 ( .A(n4265), .B(n4264), .Z(n4266) );
  AND U4898 ( .A(n4267), .B(n4266), .Z(n4390) );
  XNOR U4899 ( .A(n4389), .B(n4390), .Z(n4391) );
  XNOR U4900 ( .A(b[9]), .B(a[33]), .Z(n4411) );
  NANDN U4901 ( .A(n4411), .B(n17814), .Z(n4270) );
  NANDN U4902 ( .A(n4268), .B(n17815), .Z(n4269) );
  NAND U4903 ( .A(n4270), .B(n4269), .Z(n4375) );
  NANDN U4904 ( .A(n4271), .B(n18513), .Z(n4273) );
  XOR U4905 ( .A(b[15]), .B(a[27]), .Z(n4414) );
  NANDN U4906 ( .A(n18512), .B(n4414), .Z(n4272) );
  AND U4907 ( .A(n4273), .B(n4272), .Z(n4373) );
  NANDN U4908 ( .A(n4274), .B(n19013), .Z(n4276) );
  XNOR U4909 ( .A(b[21]), .B(a[21]), .Z(n4417) );
  NANDN U4910 ( .A(n4417), .B(n19015), .Z(n4275) );
  AND U4911 ( .A(n4276), .B(n4275), .Z(n4374) );
  XOR U4912 ( .A(n4375), .B(n4376), .Z(n4364) );
  XNOR U4913 ( .A(b[11]), .B(a[31]), .Z(n4420) );
  OR U4914 ( .A(n4420), .B(n18194), .Z(n4279) );
  NANDN U4915 ( .A(n4277), .B(n18104), .Z(n4278) );
  NAND U4916 ( .A(n4279), .B(n4278), .Z(n4362) );
  XOR U4917 ( .A(n580), .B(a[29]), .Z(n4423) );
  NANDN U4918 ( .A(n4423), .B(n18336), .Z(n4282) );
  NANDN U4919 ( .A(n4280), .B(n18337), .Z(n4281) );
  AND U4920 ( .A(n4282), .B(n4281), .Z(n4361) );
  XNOR U4921 ( .A(n4362), .B(n4361), .Z(n4363) );
  XOR U4922 ( .A(n4364), .B(n4363), .Z(n4381) );
  NAND U4923 ( .A(n19406), .B(n4283), .Z(n4285) );
  XOR U4924 ( .A(n584), .B(n4875), .Z(n4429) );
  NANDN U4925 ( .A(n576), .B(n4429), .Z(n4284) );
  NAND U4926 ( .A(n4285), .B(n4284), .Z(n4337) );
  NANDN U4927 ( .A(n585), .B(a[9]), .Z(n4338) );
  XNOR U4928 ( .A(n4337), .B(n4338), .Z(n4340) );
  NANDN U4929 ( .A(n577), .B(a[41]), .Z(n4286) );
  XOR U4930 ( .A(n17151), .B(n4286), .Z(n4288) );
  NANDN U4931 ( .A(b[0]), .B(a[40]), .Z(n4287) );
  AND U4932 ( .A(n4288), .B(n4287), .Z(n4339) );
  XOR U4933 ( .A(n4340), .B(n4339), .Z(n4379) );
  XOR U4934 ( .A(b[23]), .B(a[19]), .Z(n4432) );
  NANDN U4935 ( .A(n19127), .B(n4432), .Z(n4291) );
  NAND U4936 ( .A(n4289), .B(n19128), .Z(n4290) );
  NAND U4937 ( .A(n4291), .B(n4290), .Z(n4402) );
  NAND U4938 ( .A(n4292), .B(n17553), .Z(n4294) );
  XOR U4939 ( .A(b[7]), .B(a[35]), .Z(n4435) );
  NAND U4940 ( .A(n4435), .B(n17555), .Z(n4293) );
  NAND U4941 ( .A(n4294), .B(n4293), .Z(n4399) );
  XOR U4942 ( .A(b[25]), .B(a[17]), .Z(n4438) );
  NAND U4943 ( .A(n4438), .B(n19240), .Z(n4297) );
  NAND U4944 ( .A(n4295), .B(n19242), .Z(n4296) );
  AND U4945 ( .A(n4297), .B(n4296), .Z(n4400) );
  XNOR U4946 ( .A(n4399), .B(n4400), .Z(n4401) );
  XNOR U4947 ( .A(n4402), .B(n4401), .Z(n4380) );
  XOR U4948 ( .A(n4379), .B(n4380), .Z(n4382) );
  XNOR U4949 ( .A(n4381), .B(n4382), .Z(n4392) );
  XNOR U4950 ( .A(n4391), .B(n4392), .Z(n4327) );
  XNOR U4951 ( .A(n4328), .B(n4327), .Z(n4330) );
  XNOR U4952 ( .A(n4329), .B(n4330), .Z(n4447) );
  XOR U4953 ( .A(n4448), .B(n4447), .Z(n4450) );
  NANDN U4954 ( .A(n4299), .B(n4298), .Z(n4303) );
  NAND U4955 ( .A(n4301), .B(n4300), .Z(n4302) );
  NAND U4956 ( .A(n4303), .B(n4302), .Z(n4442) );
  NAND U4957 ( .A(n4305), .B(n4304), .Z(n4309) );
  NANDN U4958 ( .A(n4307), .B(n4306), .Z(n4308) );
  AND U4959 ( .A(n4309), .B(n4308), .Z(n4441) );
  XNOR U4960 ( .A(n4442), .B(n4441), .Z(n4443) );
  XOR U4961 ( .A(n4444), .B(n4443), .Z(n4324) );
  XOR U4962 ( .A(n4323), .B(n4324), .Z(n4315) );
  XOR U4963 ( .A(n4316), .B(n4315), .Z(n4317) );
  XNOR U4964 ( .A(n4318), .B(n4317), .Z(n4453) );
  XNOR U4965 ( .A(n4453), .B(sreg[137]), .Z(n4455) );
  NAND U4966 ( .A(n4310), .B(sreg[136]), .Z(n4314) );
  OR U4967 ( .A(n4312), .B(n4311), .Z(n4313) );
  AND U4968 ( .A(n4314), .B(n4313), .Z(n4454) );
  XOR U4969 ( .A(n4455), .B(n4454), .Z(c[137]) );
  NAND U4970 ( .A(n4316), .B(n4315), .Z(n4320) );
  NAND U4971 ( .A(n4318), .B(n4317), .Z(n4319) );
  NAND U4972 ( .A(n4320), .B(n4319), .Z(n4461) );
  NANDN U4973 ( .A(n4322), .B(n4321), .Z(n4326) );
  NAND U4974 ( .A(n4324), .B(n4323), .Z(n4325) );
  NAND U4975 ( .A(n4326), .B(n4325), .Z(n4458) );
  NAND U4976 ( .A(n4328), .B(n4327), .Z(n4332) );
  NANDN U4977 ( .A(n4330), .B(n4329), .Z(n4331) );
  NAND U4978 ( .A(n4332), .B(n4331), .Z(n4470) );
  XNOR U4979 ( .A(n4470), .B(n4471), .Z(n4472) );
  NANDN U4980 ( .A(n4338), .B(n4337), .Z(n4342) );
  NAND U4981 ( .A(n4340), .B(n4339), .Z(n4341) );
  NAND U4982 ( .A(n4342), .B(n4341), .Z(n4545) );
  NANDN U4983 ( .A(n4343), .B(n18832), .Z(n4345) );
  XNOR U4984 ( .A(b[19]), .B(a[24]), .Z(n4488) );
  NANDN U4985 ( .A(n4488), .B(n18834), .Z(n4344) );
  NAND U4986 ( .A(n4345), .B(n4344), .Z(n4555) );
  XNOR U4987 ( .A(b[27]), .B(a[16]), .Z(n4491) );
  NANDN U4988 ( .A(n4491), .B(n19336), .Z(n4348) );
  NANDN U4989 ( .A(n4346), .B(n19337), .Z(n4347) );
  NAND U4990 ( .A(n4348), .B(n4347), .Z(n4552) );
  XNOR U4991 ( .A(b[5]), .B(a[38]), .Z(n4494) );
  NANDN U4992 ( .A(n4494), .B(n17310), .Z(n4351) );
  NAND U4993 ( .A(n4349), .B(n17311), .Z(n4350) );
  AND U4994 ( .A(n4351), .B(n4350), .Z(n4553) );
  XNOR U4995 ( .A(n4552), .B(n4553), .Z(n4554) );
  XNOR U4996 ( .A(n4555), .B(n4554), .Z(n4543) );
  XOR U4997 ( .A(b[17]), .B(a[26]), .Z(n4497) );
  NAND U4998 ( .A(n4497), .B(n18673), .Z(n4354) );
  NAND U4999 ( .A(n4352), .B(n18674), .Z(n4353) );
  NAND U5000 ( .A(n4354), .B(n4353), .Z(n4515) );
  XNOR U5001 ( .A(b[31]), .B(a[12]), .Z(n4500) );
  NANDN U5002 ( .A(n4500), .B(n19472), .Z(n4357) );
  NANDN U5003 ( .A(n4355), .B(n19473), .Z(n4356) );
  NAND U5004 ( .A(n4357), .B(n4356), .Z(n4512) );
  OR U5005 ( .A(n4358), .B(n16988), .Z(n4360) );
  XNOR U5006 ( .A(b[3]), .B(a[40]), .Z(n4503) );
  NANDN U5007 ( .A(n4503), .B(n16990), .Z(n4359) );
  AND U5008 ( .A(n4360), .B(n4359), .Z(n4513) );
  XNOR U5009 ( .A(n4512), .B(n4513), .Z(n4514) );
  XOR U5010 ( .A(n4515), .B(n4514), .Z(n4542) );
  XNOR U5011 ( .A(n4543), .B(n4542), .Z(n4544) );
  XNOR U5012 ( .A(n4545), .B(n4544), .Z(n4589) );
  NANDN U5013 ( .A(n4362), .B(n4361), .Z(n4366) );
  NAND U5014 ( .A(n4364), .B(n4363), .Z(n4365) );
  NAND U5015 ( .A(n4366), .B(n4365), .Z(n4533) );
  NANDN U5016 ( .A(n4368), .B(n4367), .Z(n4372) );
  NAND U5017 ( .A(n4370), .B(n4369), .Z(n4371) );
  NAND U5018 ( .A(n4372), .B(n4371), .Z(n4531) );
  OR U5019 ( .A(n4374), .B(n4373), .Z(n4378) );
  NANDN U5020 ( .A(n4376), .B(n4375), .Z(n4377) );
  NAND U5021 ( .A(n4378), .B(n4377), .Z(n4530) );
  XNOR U5022 ( .A(n4533), .B(n4532), .Z(n4590) );
  XNOR U5023 ( .A(n4589), .B(n4590), .Z(n4591) );
  NANDN U5024 ( .A(n4380), .B(n4379), .Z(n4384) );
  OR U5025 ( .A(n4382), .B(n4381), .Z(n4383) );
  AND U5026 ( .A(n4384), .B(n4383), .Z(n4592) );
  XOR U5027 ( .A(n4591), .B(n4592), .Z(n4478) );
  NANDN U5028 ( .A(n4390), .B(n4389), .Z(n4394) );
  NANDN U5029 ( .A(n4392), .B(n4391), .Z(n4393) );
  NAND U5030 ( .A(n4394), .B(n4393), .Z(n4598) );
  NANDN U5031 ( .A(n4400), .B(n4399), .Z(n4404) );
  NAND U5032 ( .A(n4402), .B(n4401), .Z(n4403) );
  NAND U5033 ( .A(n4404), .B(n4403), .Z(n4536) );
  NANDN U5034 ( .A(n4406), .B(n4405), .Z(n4410) );
  NAND U5035 ( .A(n4408), .B(n4407), .Z(n4409) );
  AND U5036 ( .A(n4410), .B(n4409), .Z(n4537) );
  XNOR U5037 ( .A(n4536), .B(n4537), .Z(n4538) );
  XNOR U5038 ( .A(b[9]), .B(a[34]), .Z(n4558) );
  NANDN U5039 ( .A(n4558), .B(n17814), .Z(n4413) );
  NANDN U5040 ( .A(n4411), .B(n17815), .Z(n4412) );
  NAND U5041 ( .A(n4413), .B(n4412), .Z(n4520) );
  NAND U5042 ( .A(n4414), .B(n18513), .Z(n4416) );
  XOR U5043 ( .A(b[15]), .B(a[28]), .Z(n4561) );
  NANDN U5044 ( .A(n18512), .B(n4561), .Z(n4415) );
  AND U5045 ( .A(n4416), .B(n4415), .Z(n4518) );
  NANDN U5046 ( .A(n4417), .B(n19013), .Z(n4419) );
  XNOR U5047 ( .A(b[21]), .B(a[22]), .Z(n4564) );
  NANDN U5048 ( .A(n4564), .B(n19015), .Z(n4418) );
  AND U5049 ( .A(n4419), .B(n4418), .Z(n4519) );
  XOR U5050 ( .A(n4520), .B(n4521), .Z(n4509) );
  XNOR U5051 ( .A(b[11]), .B(a[32]), .Z(n4567) );
  OR U5052 ( .A(n4567), .B(n18194), .Z(n4422) );
  NANDN U5053 ( .A(n4420), .B(n18104), .Z(n4421) );
  NAND U5054 ( .A(n4422), .B(n4421), .Z(n4507) );
  XOR U5055 ( .A(n580), .B(a[30]), .Z(n4570) );
  NANDN U5056 ( .A(n4570), .B(n18336), .Z(n4425) );
  NANDN U5057 ( .A(n4423), .B(n18337), .Z(n4424) );
  AND U5058 ( .A(n4425), .B(n4424), .Z(n4506) );
  XNOR U5059 ( .A(n4507), .B(n4506), .Z(n4508) );
  XOR U5060 ( .A(n4509), .B(n4508), .Z(n4526) );
  NANDN U5061 ( .A(n577), .B(a[42]), .Z(n4426) );
  XOR U5062 ( .A(n17151), .B(n4426), .Z(n4428) );
  IV U5063 ( .A(a[41]), .Z(n8930) );
  NANDN U5064 ( .A(n8930), .B(n577), .Z(n4427) );
  AND U5065 ( .A(n4428), .B(n4427), .Z(n4484) );
  NAND U5066 ( .A(n19406), .B(n4429), .Z(n4431) );
  XNOR U5067 ( .A(b[29]), .B(a[14]), .Z(n4574) );
  OR U5068 ( .A(n4574), .B(n576), .Z(n4430) );
  NAND U5069 ( .A(n4431), .B(n4430), .Z(n4482) );
  NANDN U5070 ( .A(n585), .B(a[10]), .Z(n4483) );
  XNOR U5071 ( .A(n4482), .B(n4483), .Z(n4485) );
  XOR U5072 ( .A(n4484), .B(n4485), .Z(n4524) );
  XOR U5073 ( .A(b[23]), .B(a[20]), .Z(n4580) );
  NANDN U5074 ( .A(n19127), .B(n4580), .Z(n4434) );
  NAND U5075 ( .A(n4432), .B(n19128), .Z(n4433) );
  NAND U5076 ( .A(n4434), .B(n4433), .Z(n4549) );
  NAND U5077 ( .A(n4435), .B(n17553), .Z(n4437) );
  XOR U5078 ( .A(b[7]), .B(a[36]), .Z(n4583) );
  NAND U5079 ( .A(n4583), .B(n17555), .Z(n4436) );
  NAND U5080 ( .A(n4437), .B(n4436), .Z(n4546) );
  XOR U5081 ( .A(b[25]), .B(a[18]), .Z(n4586) );
  NAND U5082 ( .A(n4586), .B(n19240), .Z(n4440) );
  NAND U5083 ( .A(n4438), .B(n19242), .Z(n4439) );
  AND U5084 ( .A(n4440), .B(n4439), .Z(n4547) );
  XNOR U5085 ( .A(n4546), .B(n4547), .Z(n4548) );
  XNOR U5086 ( .A(n4549), .B(n4548), .Z(n4525) );
  XOR U5087 ( .A(n4524), .B(n4525), .Z(n4527) );
  XNOR U5088 ( .A(n4526), .B(n4527), .Z(n4539) );
  XOR U5089 ( .A(n4538), .B(n4539), .Z(n4596) );
  XNOR U5090 ( .A(n4595), .B(n4596), .Z(n4597) );
  XNOR U5091 ( .A(n4598), .B(n4597), .Z(n4476) );
  XNOR U5092 ( .A(n4477), .B(n4476), .Z(n4479) );
  XNOR U5093 ( .A(n4478), .B(n4479), .Z(n4473) );
  XOR U5094 ( .A(n4472), .B(n4473), .Z(n4467) );
  NANDN U5095 ( .A(n4442), .B(n4441), .Z(n4446) );
  NAND U5096 ( .A(n4444), .B(n4443), .Z(n4445) );
  NAND U5097 ( .A(n4446), .B(n4445), .Z(n4464) );
  NANDN U5098 ( .A(n4448), .B(n4447), .Z(n4452) );
  OR U5099 ( .A(n4450), .B(n4449), .Z(n4451) );
  NAND U5100 ( .A(n4452), .B(n4451), .Z(n4465) );
  XNOR U5101 ( .A(n4464), .B(n4465), .Z(n4466) );
  XNOR U5102 ( .A(n4467), .B(n4466), .Z(n4459) );
  XNOR U5103 ( .A(n4458), .B(n4459), .Z(n4460) );
  XNOR U5104 ( .A(n4461), .B(n4460), .Z(n4601) );
  XNOR U5105 ( .A(n4601), .B(sreg[138]), .Z(n4603) );
  NAND U5106 ( .A(n4453), .B(sreg[137]), .Z(n4457) );
  OR U5107 ( .A(n4455), .B(n4454), .Z(n4456) );
  AND U5108 ( .A(n4457), .B(n4456), .Z(n4602) );
  XOR U5109 ( .A(n4603), .B(n4602), .Z(c[138]) );
  NANDN U5110 ( .A(n4459), .B(n4458), .Z(n4463) );
  NAND U5111 ( .A(n4461), .B(n4460), .Z(n4462) );
  NAND U5112 ( .A(n4463), .B(n4462), .Z(n4609) );
  NANDN U5113 ( .A(n4465), .B(n4464), .Z(n4469) );
  NAND U5114 ( .A(n4467), .B(n4466), .Z(n4468) );
  NAND U5115 ( .A(n4469), .B(n4468), .Z(n4607) );
  NANDN U5116 ( .A(n4471), .B(n4470), .Z(n4475) );
  NANDN U5117 ( .A(n4473), .B(n4472), .Z(n4474) );
  NAND U5118 ( .A(n4475), .B(n4474), .Z(n4613) );
  OR U5119 ( .A(n4477), .B(n4476), .Z(n4481) );
  OR U5120 ( .A(n4479), .B(n4478), .Z(n4480) );
  AND U5121 ( .A(n4481), .B(n4480), .Z(n4612) );
  XNOR U5122 ( .A(n4613), .B(n4612), .Z(n4614) );
  NANDN U5123 ( .A(n4483), .B(n4482), .Z(n4487) );
  NAND U5124 ( .A(n4485), .B(n4484), .Z(n4486) );
  NAND U5125 ( .A(n4487), .B(n4486), .Z(n4693) );
  NANDN U5126 ( .A(n4488), .B(n18832), .Z(n4490) );
  XNOR U5127 ( .A(b[19]), .B(a[25]), .Z(n4660) );
  NANDN U5128 ( .A(n4660), .B(n18834), .Z(n4489) );
  NAND U5129 ( .A(n4490), .B(n4489), .Z(n4729) );
  XNOR U5130 ( .A(b[27]), .B(a[17]), .Z(n4663) );
  NANDN U5131 ( .A(n4663), .B(n19336), .Z(n4493) );
  NANDN U5132 ( .A(n4491), .B(n19337), .Z(n4492) );
  NAND U5133 ( .A(n4493), .B(n4492), .Z(n4726) );
  XOR U5134 ( .A(b[5]), .B(a[39]), .Z(n4666) );
  NAND U5135 ( .A(n4666), .B(n17310), .Z(n4496) );
  NANDN U5136 ( .A(n4494), .B(n17311), .Z(n4495) );
  AND U5137 ( .A(n4496), .B(n4495), .Z(n4727) );
  XNOR U5138 ( .A(n4726), .B(n4727), .Z(n4728) );
  XNOR U5139 ( .A(n4729), .B(n4728), .Z(n4690) );
  XOR U5140 ( .A(b[17]), .B(a[27]), .Z(n4669) );
  NAND U5141 ( .A(n4669), .B(n18673), .Z(n4499) );
  NAND U5142 ( .A(n4497), .B(n18674), .Z(n4498) );
  NAND U5143 ( .A(n4499), .B(n4498), .Z(n4644) );
  XOR U5144 ( .A(b[31]), .B(n4875), .Z(n4672) );
  NANDN U5145 ( .A(n4672), .B(n19472), .Z(n4502) );
  NANDN U5146 ( .A(n4500), .B(n19473), .Z(n4501) );
  AND U5147 ( .A(n4502), .B(n4501), .Z(n4642) );
  OR U5148 ( .A(n4503), .B(n16988), .Z(n4505) );
  XOR U5149 ( .A(b[3]), .B(n8930), .Z(n4675) );
  NANDN U5150 ( .A(n4675), .B(n16990), .Z(n4504) );
  AND U5151 ( .A(n4505), .B(n4504), .Z(n4643) );
  XOR U5152 ( .A(n4644), .B(n4645), .Z(n4691) );
  XOR U5153 ( .A(n4690), .B(n4691), .Z(n4692) );
  XNOR U5154 ( .A(n4693), .B(n4692), .Z(n4738) );
  NANDN U5155 ( .A(n4507), .B(n4506), .Z(n4511) );
  NAND U5156 ( .A(n4509), .B(n4508), .Z(n4510) );
  NAND U5157 ( .A(n4511), .B(n4510), .Z(n4681) );
  NANDN U5158 ( .A(n4513), .B(n4512), .Z(n4517) );
  NAND U5159 ( .A(n4515), .B(n4514), .Z(n4516) );
  NAND U5160 ( .A(n4517), .B(n4516), .Z(n4679) );
  OR U5161 ( .A(n4519), .B(n4518), .Z(n4523) );
  NANDN U5162 ( .A(n4521), .B(n4520), .Z(n4522) );
  NAND U5163 ( .A(n4523), .B(n4522), .Z(n4678) );
  XNOR U5164 ( .A(n4681), .B(n4680), .Z(n4739) );
  XOR U5165 ( .A(n4738), .B(n4739), .Z(n4741) );
  NANDN U5166 ( .A(n4525), .B(n4524), .Z(n4529) );
  OR U5167 ( .A(n4527), .B(n4526), .Z(n4528) );
  NAND U5168 ( .A(n4529), .B(n4528), .Z(n4740) );
  XOR U5169 ( .A(n4741), .B(n4740), .Z(n4626) );
  OR U5170 ( .A(n4531), .B(n4530), .Z(n4535) );
  NAND U5171 ( .A(n4533), .B(n4532), .Z(n4534) );
  NAND U5172 ( .A(n4535), .B(n4534), .Z(n4625) );
  NANDN U5173 ( .A(n4537), .B(n4536), .Z(n4541) );
  NANDN U5174 ( .A(n4539), .B(n4538), .Z(n4540) );
  NAND U5175 ( .A(n4541), .B(n4540), .Z(n4746) );
  NANDN U5176 ( .A(n4547), .B(n4546), .Z(n4551) );
  NAND U5177 ( .A(n4549), .B(n4548), .Z(n4550) );
  NAND U5178 ( .A(n4551), .B(n4550), .Z(n4684) );
  NANDN U5179 ( .A(n4553), .B(n4552), .Z(n4557) );
  NAND U5180 ( .A(n4555), .B(n4554), .Z(n4556) );
  AND U5181 ( .A(n4557), .B(n4556), .Z(n4685) );
  XNOR U5182 ( .A(n4684), .B(n4685), .Z(n4686) );
  XNOR U5183 ( .A(b[9]), .B(a[35]), .Z(n4696) );
  NANDN U5184 ( .A(n4696), .B(n17814), .Z(n4560) );
  NANDN U5185 ( .A(n4558), .B(n17815), .Z(n4559) );
  NAND U5186 ( .A(n4560), .B(n4559), .Z(n4650) );
  NAND U5187 ( .A(n4561), .B(n18513), .Z(n4563) );
  XNOR U5188 ( .A(b[15]), .B(a[29]), .Z(n4699) );
  OR U5189 ( .A(n4699), .B(n18512), .Z(n4562) );
  AND U5190 ( .A(n4563), .B(n4562), .Z(n4648) );
  NANDN U5191 ( .A(n4564), .B(n19013), .Z(n4566) );
  XNOR U5192 ( .A(b[21]), .B(a[23]), .Z(n4702) );
  NANDN U5193 ( .A(n4702), .B(n19015), .Z(n4565) );
  AND U5194 ( .A(n4566), .B(n4565), .Z(n4649) );
  XOR U5195 ( .A(n4650), .B(n4651), .Z(n4639) );
  XNOR U5196 ( .A(b[11]), .B(a[33]), .Z(n4705) );
  OR U5197 ( .A(n4705), .B(n18194), .Z(n4569) );
  NANDN U5198 ( .A(n4567), .B(n18104), .Z(n4568) );
  NAND U5199 ( .A(n4569), .B(n4568), .Z(n4637) );
  XOR U5200 ( .A(n580), .B(a[31]), .Z(n4708) );
  NANDN U5201 ( .A(n4708), .B(n18336), .Z(n4572) );
  NANDN U5202 ( .A(n4570), .B(n18337), .Z(n4571) );
  NAND U5203 ( .A(n4572), .B(n4571), .Z(n4636) );
  XOR U5204 ( .A(n4639), .B(n4638), .Z(n4633) );
  ANDN U5205 ( .B(b[31]), .A(n4573), .Z(n4654) );
  NANDN U5206 ( .A(n4574), .B(n19406), .Z(n4576) );
  XNOR U5207 ( .A(n584), .B(a[15]), .Z(n4714) );
  NANDN U5208 ( .A(n576), .B(n4714), .Z(n4575) );
  NAND U5209 ( .A(n4576), .B(n4575), .Z(n4655) );
  XOR U5210 ( .A(n4654), .B(n4655), .Z(n4656) );
  NANDN U5211 ( .A(n577), .B(a[43]), .Z(n4577) );
  XOR U5212 ( .A(n17151), .B(n4577), .Z(n4579) );
  IV U5213 ( .A(a[42]), .Z(n9080) );
  NANDN U5214 ( .A(n9080), .B(n577), .Z(n4578) );
  AND U5215 ( .A(n4579), .B(n4578), .Z(n4657) );
  XNOR U5216 ( .A(n4656), .B(n4657), .Z(n4630) );
  XOR U5217 ( .A(b[23]), .B(a[21]), .Z(n4717) );
  NANDN U5218 ( .A(n19127), .B(n4717), .Z(n4582) );
  NAND U5219 ( .A(n4580), .B(n19128), .Z(n4581) );
  NAND U5220 ( .A(n4582), .B(n4581), .Z(n4735) );
  NAND U5221 ( .A(n4583), .B(n17553), .Z(n4585) );
  XOR U5222 ( .A(b[7]), .B(a[37]), .Z(n4720) );
  NAND U5223 ( .A(n4720), .B(n17555), .Z(n4584) );
  NAND U5224 ( .A(n4585), .B(n4584), .Z(n4732) );
  XOR U5225 ( .A(b[25]), .B(a[19]), .Z(n4723) );
  NAND U5226 ( .A(n4723), .B(n19240), .Z(n4588) );
  NAND U5227 ( .A(n4586), .B(n19242), .Z(n4587) );
  AND U5228 ( .A(n4588), .B(n4587), .Z(n4733) );
  XNOR U5229 ( .A(n4732), .B(n4733), .Z(n4734) );
  XNOR U5230 ( .A(n4735), .B(n4734), .Z(n4631) );
  XOR U5231 ( .A(n4633), .B(n4632), .Z(n4687) );
  XNOR U5232 ( .A(n4686), .B(n4687), .Z(n4744) );
  XNOR U5233 ( .A(n4745), .B(n4744), .Z(n4747) );
  XNOR U5234 ( .A(n4746), .B(n4747), .Z(n4624) );
  XOR U5235 ( .A(n4625), .B(n4624), .Z(n4627) );
  NANDN U5236 ( .A(n4590), .B(n4589), .Z(n4594) );
  NAND U5237 ( .A(n4592), .B(n4591), .Z(n4593) );
  NAND U5238 ( .A(n4594), .B(n4593), .Z(n4618) );
  NANDN U5239 ( .A(n4596), .B(n4595), .Z(n4600) );
  NAND U5240 ( .A(n4598), .B(n4597), .Z(n4599) );
  NAND U5241 ( .A(n4600), .B(n4599), .Z(n4619) );
  XNOR U5242 ( .A(n4618), .B(n4619), .Z(n4620) );
  XOR U5243 ( .A(n4621), .B(n4620), .Z(n4615) );
  XOR U5244 ( .A(n4614), .B(n4615), .Z(n4606) );
  XOR U5245 ( .A(n4607), .B(n4606), .Z(n4608) );
  XNOR U5246 ( .A(n4609), .B(n4608), .Z(n4750) );
  XNOR U5247 ( .A(n4750), .B(sreg[139]), .Z(n4752) );
  NAND U5248 ( .A(n4601), .B(sreg[138]), .Z(n4605) );
  OR U5249 ( .A(n4603), .B(n4602), .Z(n4604) );
  AND U5250 ( .A(n4605), .B(n4604), .Z(n4751) );
  XOR U5251 ( .A(n4752), .B(n4751), .Z(c[139]) );
  NAND U5252 ( .A(n4607), .B(n4606), .Z(n4611) );
  NAND U5253 ( .A(n4609), .B(n4608), .Z(n4610) );
  NAND U5254 ( .A(n4611), .B(n4610), .Z(n4758) );
  NANDN U5255 ( .A(n4613), .B(n4612), .Z(n4617) );
  NAND U5256 ( .A(n4615), .B(n4614), .Z(n4616) );
  NAND U5257 ( .A(n4617), .B(n4616), .Z(n4756) );
  NANDN U5258 ( .A(n4619), .B(n4618), .Z(n4623) );
  NAND U5259 ( .A(n4621), .B(n4620), .Z(n4622) );
  NAND U5260 ( .A(n4623), .B(n4622), .Z(n4761) );
  NANDN U5261 ( .A(n4625), .B(n4624), .Z(n4629) );
  OR U5262 ( .A(n4627), .B(n4626), .Z(n4628) );
  NAND U5263 ( .A(n4629), .B(n4628), .Z(n4762) );
  XNOR U5264 ( .A(n4761), .B(n4762), .Z(n4763) );
  OR U5265 ( .A(n4631), .B(n4630), .Z(n4635) );
  NANDN U5266 ( .A(n4633), .B(n4632), .Z(n4634) );
  NAND U5267 ( .A(n4635), .B(n4634), .Z(n4891) );
  OR U5268 ( .A(n4637), .B(n4636), .Z(n4641) );
  NAND U5269 ( .A(n4639), .B(n4638), .Z(n4640) );
  NAND U5270 ( .A(n4641), .B(n4640), .Z(n4829) );
  OR U5271 ( .A(n4643), .B(n4642), .Z(n4647) );
  NANDN U5272 ( .A(n4645), .B(n4644), .Z(n4646) );
  NAND U5273 ( .A(n4647), .B(n4646), .Z(n4828) );
  OR U5274 ( .A(n4649), .B(n4648), .Z(n4653) );
  NANDN U5275 ( .A(n4651), .B(n4650), .Z(n4652) );
  NAND U5276 ( .A(n4653), .B(n4652), .Z(n4827) );
  XOR U5277 ( .A(n4829), .B(n4830), .Z(n4889) );
  OR U5278 ( .A(n4655), .B(n4654), .Z(n4659) );
  NANDN U5279 ( .A(n4657), .B(n4656), .Z(n4658) );
  NAND U5280 ( .A(n4659), .B(n4658), .Z(n4842) );
  NANDN U5281 ( .A(n4660), .B(n18832), .Z(n4662) );
  XNOR U5282 ( .A(b[19]), .B(a[26]), .Z(n4809) );
  NANDN U5283 ( .A(n4809), .B(n18834), .Z(n4661) );
  NAND U5284 ( .A(n4662), .B(n4661), .Z(n4854) );
  XNOR U5285 ( .A(b[27]), .B(a[18]), .Z(n4812) );
  NANDN U5286 ( .A(n4812), .B(n19336), .Z(n4665) );
  NANDN U5287 ( .A(n4663), .B(n19337), .Z(n4664) );
  NAND U5288 ( .A(n4665), .B(n4664), .Z(n4851) );
  XOR U5289 ( .A(b[5]), .B(a[40]), .Z(n4815) );
  NAND U5290 ( .A(n4815), .B(n17310), .Z(n4668) );
  NAND U5291 ( .A(n4666), .B(n17311), .Z(n4667) );
  AND U5292 ( .A(n4668), .B(n4667), .Z(n4852) );
  XNOR U5293 ( .A(n4851), .B(n4852), .Z(n4853) );
  XNOR U5294 ( .A(n4854), .B(n4853), .Z(n4839) );
  XOR U5295 ( .A(b[17]), .B(a[28]), .Z(n4818) );
  NAND U5296 ( .A(n4818), .B(n18673), .Z(n4671) );
  NAND U5297 ( .A(n4669), .B(n18674), .Z(n4670) );
  NAND U5298 ( .A(n4671), .B(n4670), .Z(n4793) );
  XNOR U5299 ( .A(n585), .B(a[14]), .Z(n4821) );
  NAND U5300 ( .A(n4821), .B(n19472), .Z(n4674) );
  NANDN U5301 ( .A(n4672), .B(n19473), .Z(n4673) );
  AND U5302 ( .A(n4674), .B(n4673), .Z(n4791) );
  OR U5303 ( .A(n4675), .B(n16988), .Z(n4677) );
  XOR U5304 ( .A(b[3]), .B(n9080), .Z(n4824) );
  NANDN U5305 ( .A(n4824), .B(n16990), .Z(n4676) );
  AND U5306 ( .A(n4677), .B(n4676), .Z(n4792) );
  XOR U5307 ( .A(n4793), .B(n4794), .Z(n4840) );
  XOR U5308 ( .A(n4839), .B(n4840), .Z(n4841) );
  XNOR U5309 ( .A(n4842), .B(n4841), .Z(n4888) );
  XOR U5310 ( .A(n4889), .B(n4888), .Z(n4890) );
  XNOR U5311 ( .A(n4891), .B(n4890), .Z(n4776) );
  OR U5312 ( .A(n4679), .B(n4678), .Z(n4683) );
  NAND U5313 ( .A(n4681), .B(n4680), .Z(n4682) );
  NAND U5314 ( .A(n4683), .B(n4682), .Z(n4774) );
  NANDN U5315 ( .A(n4685), .B(n4684), .Z(n4689) );
  NANDN U5316 ( .A(n4687), .B(n4686), .Z(n4688) );
  NAND U5317 ( .A(n4689), .B(n4688), .Z(n4895) );
  OR U5318 ( .A(n4691), .B(n4690), .Z(n4695) );
  NAND U5319 ( .A(n4693), .B(n4692), .Z(n4694) );
  NAND U5320 ( .A(n4695), .B(n4694), .Z(n4892) );
  XNOR U5321 ( .A(n579), .B(a[36]), .Z(n4857) );
  NAND U5322 ( .A(n17814), .B(n4857), .Z(n4698) );
  NANDN U5323 ( .A(n4696), .B(n17815), .Z(n4697) );
  NAND U5324 ( .A(n4698), .B(n4697), .Z(n4799) );
  NANDN U5325 ( .A(n4699), .B(n18513), .Z(n4701) );
  XNOR U5326 ( .A(b[15]), .B(a[30]), .Z(n4860) );
  OR U5327 ( .A(n4860), .B(n18512), .Z(n4700) );
  AND U5328 ( .A(n4701), .B(n4700), .Z(n4797) );
  NANDN U5329 ( .A(n4702), .B(n19013), .Z(n4704) );
  XNOR U5330 ( .A(b[21]), .B(a[24]), .Z(n4863) );
  NANDN U5331 ( .A(n4863), .B(n19015), .Z(n4703) );
  AND U5332 ( .A(n4704), .B(n4703), .Z(n4798) );
  XOR U5333 ( .A(n4799), .B(n4800), .Z(n4788) );
  XNOR U5334 ( .A(b[11]), .B(a[34]), .Z(n4866) );
  OR U5335 ( .A(n4866), .B(n18194), .Z(n4707) );
  NANDN U5336 ( .A(n4705), .B(n18104), .Z(n4706) );
  NAND U5337 ( .A(n4707), .B(n4706), .Z(n4786) );
  XNOR U5338 ( .A(b[13]), .B(a[32]), .Z(n4869) );
  NANDN U5339 ( .A(n4869), .B(n18336), .Z(n4710) );
  NANDN U5340 ( .A(n4708), .B(n18337), .Z(n4709) );
  NAND U5341 ( .A(n4710), .B(n4709), .Z(n4785) );
  XOR U5342 ( .A(n4788), .B(n4787), .Z(n4782) );
  NANDN U5343 ( .A(n577), .B(a[44]), .Z(n4711) );
  XOR U5344 ( .A(n17151), .B(n4711), .Z(n4713) );
  NANDN U5345 ( .A(b[0]), .B(a[43]), .Z(n4712) );
  AND U5346 ( .A(n4713), .B(n4712), .Z(n4805) );
  NAND U5347 ( .A(n4714), .B(n19406), .Z(n4716) );
  XNOR U5348 ( .A(b[29]), .B(a[16]), .Z(n4876) );
  OR U5349 ( .A(n4876), .B(n576), .Z(n4715) );
  NAND U5350 ( .A(n4716), .B(n4715), .Z(n4803) );
  NANDN U5351 ( .A(n585), .B(a[12]), .Z(n4804) );
  XNOR U5352 ( .A(n4803), .B(n4804), .Z(n4806) );
  XNOR U5353 ( .A(n4805), .B(n4806), .Z(n4780) );
  XOR U5354 ( .A(b[23]), .B(a[22]), .Z(n4879) );
  NANDN U5355 ( .A(n19127), .B(n4879), .Z(n4719) );
  NAND U5356 ( .A(n4717), .B(n19128), .Z(n4718) );
  NAND U5357 ( .A(n4719), .B(n4718), .Z(n4848) );
  NAND U5358 ( .A(n4720), .B(n17553), .Z(n4722) );
  XNOR U5359 ( .A(b[7]), .B(a[38]), .Z(n4882) );
  NANDN U5360 ( .A(n4882), .B(n17555), .Z(n4721) );
  NAND U5361 ( .A(n4722), .B(n4721), .Z(n4845) );
  XOR U5362 ( .A(b[25]), .B(a[20]), .Z(n4885) );
  NAND U5363 ( .A(n4885), .B(n19240), .Z(n4725) );
  NAND U5364 ( .A(n4723), .B(n19242), .Z(n4724) );
  AND U5365 ( .A(n4725), .B(n4724), .Z(n4846) );
  XNOR U5366 ( .A(n4845), .B(n4846), .Z(n4847) );
  XOR U5367 ( .A(n4848), .B(n4847), .Z(n4779) );
  XNOR U5368 ( .A(n4782), .B(n4781), .Z(n4836) );
  NANDN U5369 ( .A(n4727), .B(n4726), .Z(n4731) );
  NAND U5370 ( .A(n4729), .B(n4728), .Z(n4730) );
  NAND U5371 ( .A(n4731), .B(n4730), .Z(n4834) );
  NANDN U5372 ( .A(n4733), .B(n4732), .Z(n4737) );
  NAND U5373 ( .A(n4735), .B(n4734), .Z(n4736) );
  AND U5374 ( .A(n4737), .B(n4736), .Z(n4833) );
  XNOR U5375 ( .A(n4834), .B(n4833), .Z(n4835) );
  XNOR U5376 ( .A(n4836), .B(n4835), .Z(n4893) );
  XNOR U5377 ( .A(n4892), .B(n4893), .Z(n4894) );
  XOR U5378 ( .A(n4895), .B(n4894), .Z(n4773) );
  XNOR U5379 ( .A(n4774), .B(n4773), .Z(n4775) );
  XOR U5380 ( .A(n4776), .B(n4775), .Z(n4770) );
  NANDN U5381 ( .A(n4739), .B(n4738), .Z(n4743) );
  OR U5382 ( .A(n4741), .B(n4740), .Z(n4742) );
  NAND U5383 ( .A(n4743), .B(n4742), .Z(n4767) );
  NAND U5384 ( .A(n4745), .B(n4744), .Z(n4749) );
  NANDN U5385 ( .A(n4747), .B(n4746), .Z(n4748) );
  NAND U5386 ( .A(n4749), .B(n4748), .Z(n4768) );
  XNOR U5387 ( .A(n4767), .B(n4768), .Z(n4769) );
  XOR U5388 ( .A(n4770), .B(n4769), .Z(n4764) );
  XOR U5389 ( .A(n4763), .B(n4764), .Z(n4755) );
  XOR U5390 ( .A(n4756), .B(n4755), .Z(n4757) );
  XNOR U5391 ( .A(n4758), .B(n4757), .Z(n4898) );
  XNOR U5392 ( .A(n4898), .B(sreg[140]), .Z(n4900) );
  NAND U5393 ( .A(n4750), .B(sreg[139]), .Z(n4754) );
  OR U5394 ( .A(n4752), .B(n4751), .Z(n4753) );
  AND U5395 ( .A(n4754), .B(n4753), .Z(n4899) );
  XOR U5396 ( .A(n4900), .B(n4899), .Z(c[140]) );
  NAND U5397 ( .A(n4756), .B(n4755), .Z(n4760) );
  NAND U5398 ( .A(n4758), .B(n4757), .Z(n4759) );
  NAND U5399 ( .A(n4760), .B(n4759), .Z(n4906) );
  NANDN U5400 ( .A(n4762), .B(n4761), .Z(n4766) );
  NAND U5401 ( .A(n4764), .B(n4763), .Z(n4765) );
  NAND U5402 ( .A(n4766), .B(n4765), .Z(n4904) );
  NANDN U5403 ( .A(n4768), .B(n4767), .Z(n4772) );
  NAND U5404 ( .A(n4770), .B(n4769), .Z(n4771) );
  NAND U5405 ( .A(n4772), .B(n4771), .Z(n4909) );
  NANDN U5406 ( .A(n4774), .B(n4773), .Z(n4778) );
  NANDN U5407 ( .A(n4776), .B(n4775), .Z(n4777) );
  NAND U5408 ( .A(n4778), .B(n4777), .Z(n4910) );
  XNOR U5409 ( .A(n4909), .B(n4910), .Z(n4911) );
  NANDN U5410 ( .A(n4780), .B(n4779), .Z(n4784) );
  NANDN U5411 ( .A(n4782), .B(n4781), .Z(n4783) );
  NAND U5412 ( .A(n4784), .B(n4783), .Z(n5020) );
  OR U5413 ( .A(n4786), .B(n4785), .Z(n4790) );
  NAND U5414 ( .A(n4788), .B(n4787), .Z(n4789) );
  NAND U5415 ( .A(n4790), .B(n4789), .Z(n4959) );
  OR U5416 ( .A(n4792), .B(n4791), .Z(n4796) );
  NANDN U5417 ( .A(n4794), .B(n4793), .Z(n4795) );
  NAND U5418 ( .A(n4796), .B(n4795), .Z(n4958) );
  OR U5419 ( .A(n4798), .B(n4797), .Z(n4802) );
  NANDN U5420 ( .A(n4800), .B(n4799), .Z(n4801) );
  NAND U5421 ( .A(n4802), .B(n4801), .Z(n4957) );
  XOR U5422 ( .A(n4959), .B(n4960), .Z(n5017) );
  NANDN U5423 ( .A(n4804), .B(n4803), .Z(n4808) );
  NAND U5424 ( .A(n4806), .B(n4805), .Z(n4807) );
  NAND U5425 ( .A(n4808), .B(n4807), .Z(n4972) );
  NANDN U5426 ( .A(n4809), .B(n18832), .Z(n4811) );
  XNOR U5427 ( .A(b[19]), .B(a[27]), .Z(n4939) );
  NANDN U5428 ( .A(n4939), .B(n18834), .Z(n4810) );
  NAND U5429 ( .A(n4811), .B(n4810), .Z(n4984) );
  XNOR U5430 ( .A(b[27]), .B(a[19]), .Z(n4942) );
  NANDN U5431 ( .A(n4942), .B(n19336), .Z(n4814) );
  NANDN U5432 ( .A(n4812), .B(n19337), .Z(n4813) );
  NAND U5433 ( .A(n4814), .B(n4813), .Z(n4981) );
  XNOR U5434 ( .A(b[5]), .B(a[41]), .Z(n4945) );
  NANDN U5435 ( .A(n4945), .B(n17310), .Z(n4817) );
  NAND U5436 ( .A(n4815), .B(n17311), .Z(n4816) );
  AND U5437 ( .A(n4817), .B(n4816), .Z(n4982) );
  XNOR U5438 ( .A(n4981), .B(n4982), .Z(n4983) );
  XNOR U5439 ( .A(n4984), .B(n4983), .Z(n4969) );
  XNOR U5440 ( .A(b[17]), .B(a[29]), .Z(n4948) );
  NANDN U5441 ( .A(n4948), .B(n18673), .Z(n4820) );
  NAND U5442 ( .A(n18674), .B(n4818), .Z(n4819) );
  NAND U5443 ( .A(n4820), .B(n4819), .Z(n4927) );
  XOR U5444 ( .A(b[31]), .B(n5159), .Z(n4951) );
  NANDN U5445 ( .A(n4951), .B(n19472), .Z(n4823) );
  NAND U5446 ( .A(n19473), .B(n4821), .Z(n4822) );
  NAND U5447 ( .A(n4823), .B(n4822), .Z(n4925) );
  OR U5448 ( .A(n4824), .B(n16988), .Z(n4826) );
  XNOR U5449 ( .A(b[3]), .B(a[43]), .Z(n4954) );
  NANDN U5450 ( .A(n4954), .B(n16990), .Z(n4825) );
  AND U5451 ( .A(n4826), .B(n4825), .Z(n4926) );
  XNOR U5452 ( .A(n4925), .B(n4926), .Z(n4928) );
  XNOR U5453 ( .A(n4927), .B(n4928), .Z(n4970) );
  XOR U5454 ( .A(n4969), .B(n4970), .Z(n4971) );
  XNOR U5455 ( .A(n4972), .B(n4971), .Z(n5018) );
  XNOR U5456 ( .A(n5017), .B(n5018), .Z(n5019) );
  XNOR U5457 ( .A(n5020), .B(n5019), .Z(n5038) );
  OR U5458 ( .A(n4828), .B(n4827), .Z(n4832) );
  NANDN U5459 ( .A(n4830), .B(n4829), .Z(n4831) );
  NAND U5460 ( .A(n4832), .B(n4831), .Z(n5036) );
  NANDN U5461 ( .A(n4834), .B(n4833), .Z(n4838) );
  NANDN U5462 ( .A(n4836), .B(n4835), .Z(n4837) );
  NAND U5463 ( .A(n4838), .B(n4837), .Z(n5026) );
  OR U5464 ( .A(n4840), .B(n4839), .Z(n4844) );
  NANDN U5465 ( .A(n4842), .B(n4841), .Z(n4843) );
  NAND U5466 ( .A(n4844), .B(n4843), .Z(n5024) );
  NANDN U5467 ( .A(n4846), .B(n4845), .Z(n4850) );
  NAND U5468 ( .A(n4848), .B(n4847), .Z(n4849) );
  NAND U5469 ( .A(n4850), .B(n4849), .Z(n4963) );
  NANDN U5470 ( .A(n4852), .B(n4851), .Z(n4856) );
  NAND U5471 ( .A(n4854), .B(n4853), .Z(n4855) );
  AND U5472 ( .A(n4856), .B(n4855), .Z(n4964) );
  XNOR U5473 ( .A(n4963), .B(n4964), .Z(n4965) );
  XNOR U5474 ( .A(b[9]), .B(a[37]), .Z(n4987) );
  NANDN U5475 ( .A(n4987), .B(n17814), .Z(n4859) );
  NAND U5476 ( .A(n17815), .B(n4857), .Z(n4858) );
  NAND U5477 ( .A(n4859), .B(n4858), .Z(n4931) );
  XNOR U5478 ( .A(b[15]), .B(a[31]), .Z(n4990) );
  OR U5479 ( .A(n4990), .B(n18512), .Z(n4862) );
  NANDN U5480 ( .A(n4860), .B(n18513), .Z(n4861) );
  NAND U5481 ( .A(n4862), .B(n4861), .Z(n4929) );
  NANDN U5482 ( .A(n4863), .B(n19013), .Z(n4865) );
  XNOR U5483 ( .A(b[21]), .B(a[25]), .Z(n4993) );
  NANDN U5484 ( .A(n4993), .B(n19015), .Z(n4864) );
  AND U5485 ( .A(n4865), .B(n4864), .Z(n4930) );
  XNOR U5486 ( .A(n4929), .B(n4930), .Z(n4932) );
  XOR U5487 ( .A(n4931), .B(n4932), .Z(n4924) );
  XNOR U5488 ( .A(b[11]), .B(a[35]), .Z(n4996) );
  OR U5489 ( .A(n4996), .B(n18194), .Z(n4868) );
  NANDN U5490 ( .A(n4866), .B(n18104), .Z(n4867) );
  NAND U5491 ( .A(n4868), .B(n4867), .Z(n4922) );
  XNOR U5492 ( .A(n580), .B(a[33]), .Z(n4999) );
  NAND U5493 ( .A(n4999), .B(n18336), .Z(n4871) );
  NANDN U5494 ( .A(n4869), .B(n18337), .Z(n4870) );
  AND U5495 ( .A(n4871), .B(n4870), .Z(n4921) );
  XNOR U5496 ( .A(n4922), .B(n4921), .Z(n4923) );
  XNOR U5497 ( .A(n4924), .B(n4923), .Z(n4917) );
  NANDN U5498 ( .A(n577), .B(a[45]), .Z(n4872) );
  XOR U5499 ( .A(n17151), .B(n4872), .Z(n4874) );
  NANDN U5500 ( .A(b[0]), .B(a[44]), .Z(n4873) );
  AND U5501 ( .A(n4874), .B(n4873), .Z(n4936) );
  ANDN U5502 ( .B(b[31]), .A(n4875), .Z(n4933) );
  NANDN U5503 ( .A(n4876), .B(n19406), .Z(n4878) );
  XNOR U5504 ( .A(n584), .B(a[17]), .Z(n5005) );
  NANDN U5505 ( .A(n576), .B(n5005), .Z(n4877) );
  NAND U5506 ( .A(n4878), .B(n4877), .Z(n4934) );
  XOR U5507 ( .A(n4933), .B(n4934), .Z(n4935) );
  XNOR U5508 ( .A(n4936), .B(n4935), .Z(n4915) );
  XOR U5509 ( .A(b[23]), .B(a[23]), .Z(n5008) );
  NANDN U5510 ( .A(n19127), .B(n5008), .Z(n4881) );
  NAND U5511 ( .A(n4879), .B(n19128), .Z(n4880) );
  NAND U5512 ( .A(n4881), .B(n4880), .Z(n4978) );
  NANDN U5513 ( .A(n4882), .B(n17553), .Z(n4884) );
  XOR U5514 ( .A(b[7]), .B(a[39]), .Z(n5011) );
  NAND U5515 ( .A(n5011), .B(n17555), .Z(n4883) );
  NAND U5516 ( .A(n4884), .B(n4883), .Z(n4975) );
  XOR U5517 ( .A(b[25]), .B(a[21]), .Z(n5014) );
  NAND U5518 ( .A(n5014), .B(n19240), .Z(n4887) );
  NAND U5519 ( .A(n4885), .B(n19242), .Z(n4886) );
  AND U5520 ( .A(n4887), .B(n4886), .Z(n4976) );
  XNOR U5521 ( .A(n4975), .B(n4976), .Z(n4977) );
  XNOR U5522 ( .A(n4978), .B(n4977), .Z(n4916) );
  XNOR U5523 ( .A(n4915), .B(n4916), .Z(n4918) );
  XOR U5524 ( .A(n4965), .B(n4966), .Z(n5023) );
  XOR U5525 ( .A(n5024), .B(n5023), .Z(n5025) );
  XNOR U5526 ( .A(n5026), .B(n5025), .Z(n5035) );
  XNOR U5527 ( .A(n5036), .B(n5035), .Z(n5037) );
  XOR U5528 ( .A(n5038), .B(n5037), .Z(n5032) );
  NANDN U5529 ( .A(n4893), .B(n4892), .Z(n4897) );
  NAND U5530 ( .A(n4895), .B(n4894), .Z(n4896) );
  AND U5531 ( .A(n4897), .B(n4896), .Z(n5029) );
  XNOR U5532 ( .A(n5030), .B(n5029), .Z(n5031) );
  XOR U5533 ( .A(n5032), .B(n5031), .Z(n4912) );
  XOR U5534 ( .A(n4911), .B(n4912), .Z(n4903) );
  XOR U5535 ( .A(n4904), .B(n4903), .Z(n4905) );
  XNOR U5536 ( .A(n4906), .B(n4905), .Z(n5041) );
  XNOR U5537 ( .A(n5041), .B(sreg[141]), .Z(n5043) );
  NAND U5538 ( .A(n4898), .B(sreg[140]), .Z(n4902) );
  OR U5539 ( .A(n4900), .B(n4899), .Z(n4901) );
  AND U5540 ( .A(n4902), .B(n4901), .Z(n5042) );
  XOR U5541 ( .A(n5043), .B(n5042), .Z(c[141]) );
  NAND U5542 ( .A(n4904), .B(n4903), .Z(n4908) );
  NAND U5543 ( .A(n4906), .B(n4905), .Z(n4907) );
  NAND U5544 ( .A(n4908), .B(n4907), .Z(n5049) );
  NANDN U5545 ( .A(n4910), .B(n4909), .Z(n4914) );
  NAND U5546 ( .A(n4912), .B(n4911), .Z(n4913) );
  NAND U5547 ( .A(n4914), .B(n4913), .Z(n5047) );
  OR U5548 ( .A(n4916), .B(n4915), .Z(n4920) );
  OR U5549 ( .A(n4918), .B(n4917), .Z(n4919) );
  NAND U5550 ( .A(n4920), .B(n4919), .Z(n5065) );
  XNOR U5551 ( .A(n5117), .B(n5116), .Z(n5119) );
  XNOR U5552 ( .A(n5118), .B(n5119), .Z(n5063) );
  OR U5553 ( .A(n4934), .B(n4933), .Z(n4938) );
  NANDN U5554 ( .A(n4936), .B(n4935), .Z(n4937) );
  NAND U5555 ( .A(n4938), .B(n4937), .Z(n5128) );
  NANDN U5556 ( .A(n4939), .B(n18832), .Z(n4941) );
  XNOR U5557 ( .A(b[19]), .B(a[28]), .Z(n5074) );
  NANDN U5558 ( .A(n5074), .B(n18834), .Z(n4940) );
  NAND U5559 ( .A(n4941), .B(n4940), .Z(n5141) );
  XNOR U5560 ( .A(b[27]), .B(a[20]), .Z(n5077) );
  NANDN U5561 ( .A(n5077), .B(n19336), .Z(n4944) );
  NANDN U5562 ( .A(n4942), .B(n19337), .Z(n4943) );
  NAND U5563 ( .A(n4944), .B(n4943), .Z(n5138) );
  XNOR U5564 ( .A(b[5]), .B(a[42]), .Z(n5080) );
  NANDN U5565 ( .A(n5080), .B(n17310), .Z(n4947) );
  NANDN U5566 ( .A(n4945), .B(n17311), .Z(n4946) );
  AND U5567 ( .A(n4947), .B(n4946), .Z(n5139) );
  XNOR U5568 ( .A(n5138), .B(n5139), .Z(n5140) );
  XNOR U5569 ( .A(n5141), .B(n5140), .Z(n5127) );
  XNOR U5570 ( .A(b[17]), .B(a[30]), .Z(n5083) );
  NANDN U5571 ( .A(n5083), .B(n18673), .Z(n4950) );
  NANDN U5572 ( .A(n4948), .B(n18674), .Z(n4949) );
  NAND U5573 ( .A(n4950), .B(n4949), .Z(n5101) );
  XNOR U5574 ( .A(b[31]), .B(a[16]), .Z(n5086) );
  NANDN U5575 ( .A(n5086), .B(n19472), .Z(n4953) );
  NANDN U5576 ( .A(n4951), .B(n19473), .Z(n4952) );
  NAND U5577 ( .A(n4953), .B(n4952), .Z(n5098) );
  OR U5578 ( .A(n4954), .B(n16988), .Z(n4956) );
  XNOR U5579 ( .A(b[3]), .B(a[44]), .Z(n5089) );
  NANDN U5580 ( .A(n5089), .B(n16990), .Z(n4955) );
  AND U5581 ( .A(n4956), .B(n4955), .Z(n5099) );
  XNOR U5582 ( .A(n5098), .B(n5099), .Z(n5100) );
  XOR U5583 ( .A(n5101), .B(n5100), .Z(n5126) );
  XOR U5584 ( .A(n5127), .B(n5126), .Z(n5129) );
  XOR U5585 ( .A(n5128), .B(n5129), .Z(n5062) );
  XNOR U5586 ( .A(n5063), .B(n5062), .Z(n5064) );
  XNOR U5587 ( .A(n5065), .B(n5064), .Z(n5184) );
  OR U5588 ( .A(n4958), .B(n4957), .Z(n4962) );
  NANDN U5589 ( .A(n4960), .B(n4959), .Z(n4961) );
  NAND U5590 ( .A(n4962), .B(n4961), .Z(n5182) );
  NANDN U5591 ( .A(n4964), .B(n4963), .Z(n4968) );
  NAND U5592 ( .A(n4966), .B(n4965), .Z(n4967) );
  NAND U5593 ( .A(n4968), .B(n4967), .Z(n5058) );
  OR U5594 ( .A(n4970), .B(n4969), .Z(n4974) );
  NAND U5595 ( .A(n4972), .B(n4971), .Z(n4973) );
  NAND U5596 ( .A(n4974), .B(n4973), .Z(n5057) );
  NANDN U5597 ( .A(n4976), .B(n4975), .Z(n4980) );
  NAND U5598 ( .A(n4978), .B(n4977), .Z(n4979) );
  NAND U5599 ( .A(n4980), .B(n4979), .Z(n5120) );
  NANDN U5600 ( .A(n4982), .B(n4981), .Z(n4986) );
  NAND U5601 ( .A(n4984), .B(n4983), .Z(n4985) );
  AND U5602 ( .A(n4986), .B(n4985), .Z(n5121) );
  XNOR U5603 ( .A(n5120), .B(n5121), .Z(n5122) );
  XOR U5604 ( .A(b[9]), .B(n8490), .Z(n5144) );
  NANDN U5605 ( .A(n5144), .B(n17814), .Z(n4989) );
  NANDN U5606 ( .A(n4987), .B(n17815), .Z(n4988) );
  NAND U5607 ( .A(n4989), .B(n4988), .Z(n5112) );
  NANDN U5608 ( .A(n4990), .B(n18513), .Z(n4992) );
  XOR U5609 ( .A(b[15]), .B(a[32]), .Z(n5147) );
  NANDN U5610 ( .A(n18512), .B(n5147), .Z(n4991) );
  AND U5611 ( .A(n4992), .B(n4991), .Z(n5110) );
  NANDN U5612 ( .A(n4993), .B(n19013), .Z(n4995) );
  XNOR U5613 ( .A(b[21]), .B(a[26]), .Z(n5150) );
  NANDN U5614 ( .A(n5150), .B(n19015), .Z(n4994) );
  AND U5615 ( .A(n4995), .B(n4994), .Z(n5111) );
  XOR U5616 ( .A(n5112), .B(n5113), .Z(n5107) );
  XNOR U5617 ( .A(b[11]), .B(a[36]), .Z(n5153) );
  OR U5618 ( .A(n5153), .B(n18194), .Z(n4998) );
  NANDN U5619 ( .A(n4996), .B(n18104), .Z(n4997) );
  NAND U5620 ( .A(n4998), .B(n4997), .Z(n5105) );
  XOR U5621 ( .A(n580), .B(a[34]), .Z(n5156) );
  NANDN U5622 ( .A(n5156), .B(n18336), .Z(n5001) );
  NAND U5623 ( .A(n18337), .B(n4999), .Z(n5000) );
  AND U5624 ( .A(n5001), .B(n5000), .Z(n5104) );
  XNOR U5625 ( .A(n5105), .B(n5104), .Z(n5106) );
  XOR U5626 ( .A(n5107), .B(n5106), .Z(n5094) );
  NANDN U5627 ( .A(n577), .B(a[46]), .Z(n5002) );
  XOR U5628 ( .A(n17151), .B(n5002), .Z(n5004) );
  NANDN U5629 ( .A(b[0]), .B(a[45]), .Z(n5003) );
  AND U5630 ( .A(n5004), .B(n5003), .Z(n5070) );
  NAND U5631 ( .A(n5005), .B(n19406), .Z(n5007) );
  XNOR U5632 ( .A(b[29]), .B(a[18]), .Z(n5160) );
  OR U5633 ( .A(n5160), .B(n576), .Z(n5006) );
  NAND U5634 ( .A(n5007), .B(n5006), .Z(n5068) );
  NANDN U5635 ( .A(n585), .B(a[14]), .Z(n5069) );
  XNOR U5636 ( .A(n5068), .B(n5069), .Z(n5071) );
  XOR U5637 ( .A(n5070), .B(n5071), .Z(n5092) );
  XOR U5638 ( .A(b[23]), .B(a[24]), .Z(n5166) );
  NANDN U5639 ( .A(n19127), .B(n5166), .Z(n5010) );
  NAND U5640 ( .A(n5008), .B(n19128), .Z(n5009) );
  NAND U5641 ( .A(n5010), .B(n5009), .Z(n5135) );
  NAND U5642 ( .A(n5011), .B(n17553), .Z(n5013) );
  XOR U5643 ( .A(b[7]), .B(a[40]), .Z(n5169) );
  NAND U5644 ( .A(n5169), .B(n17555), .Z(n5012) );
  NAND U5645 ( .A(n5013), .B(n5012), .Z(n5132) );
  XOR U5646 ( .A(b[25]), .B(a[22]), .Z(n5172) );
  NAND U5647 ( .A(n5172), .B(n19240), .Z(n5016) );
  NAND U5648 ( .A(n5014), .B(n19242), .Z(n5015) );
  AND U5649 ( .A(n5016), .B(n5015), .Z(n5133) );
  XNOR U5650 ( .A(n5132), .B(n5133), .Z(n5134) );
  XNOR U5651 ( .A(n5135), .B(n5134), .Z(n5093) );
  XOR U5652 ( .A(n5092), .B(n5093), .Z(n5095) );
  XNOR U5653 ( .A(n5094), .B(n5095), .Z(n5123) );
  XNOR U5654 ( .A(n5122), .B(n5123), .Z(n5056) );
  XNOR U5655 ( .A(n5057), .B(n5056), .Z(n5059) );
  XNOR U5656 ( .A(n5058), .B(n5059), .Z(n5181) );
  XNOR U5657 ( .A(n5182), .B(n5181), .Z(n5183) );
  XOR U5658 ( .A(n5184), .B(n5183), .Z(n5178) );
  NANDN U5659 ( .A(n5018), .B(n5017), .Z(n5022) );
  NAND U5660 ( .A(n5020), .B(n5019), .Z(n5021) );
  NAND U5661 ( .A(n5022), .B(n5021), .Z(n5176) );
  NAND U5662 ( .A(n5024), .B(n5023), .Z(n5028) );
  NANDN U5663 ( .A(n5026), .B(n5025), .Z(n5027) );
  AND U5664 ( .A(n5028), .B(n5027), .Z(n5175) );
  XNOR U5665 ( .A(n5176), .B(n5175), .Z(n5177) );
  XNOR U5666 ( .A(n5178), .B(n5177), .Z(n5053) );
  NANDN U5667 ( .A(n5030), .B(n5029), .Z(n5034) );
  NAND U5668 ( .A(n5032), .B(n5031), .Z(n5033) );
  NAND U5669 ( .A(n5034), .B(n5033), .Z(n5050) );
  NANDN U5670 ( .A(n5036), .B(n5035), .Z(n5040) );
  NANDN U5671 ( .A(n5038), .B(n5037), .Z(n5039) );
  NAND U5672 ( .A(n5040), .B(n5039), .Z(n5051) );
  XNOR U5673 ( .A(n5050), .B(n5051), .Z(n5052) );
  XNOR U5674 ( .A(n5053), .B(n5052), .Z(n5046) );
  XOR U5675 ( .A(n5047), .B(n5046), .Z(n5048) );
  XNOR U5676 ( .A(n5049), .B(n5048), .Z(n5187) );
  XNOR U5677 ( .A(n5187), .B(sreg[142]), .Z(n5189) );
  NAND U5678 ( .A(n5041), .B(sreg[141]), .Z(n5045) );
  OR U5679 ( .A(n5043), .B(n5042), .Z(n5044) );
  AND U5680 ( .A(n5045), .B(n5044), .Z(n5188) );
  XOR U5681 ( .A(n5189), .B(n5188), .Z(c[142]) );
  NANDN U5682 ( .A(n5051), .B(n5050), .Z(n5055) );
  NANDN U5683 ( .A(n5053), .B(n5052), .Z(n5054) );
  NAND U5684 ( .A(n5055), .B(n5054), .Z(n5192) );
  NAND U5685 ( .A(n5057), .B(n5056), .Z(n5061) );
  NANDN U5686 ( .A(n5059), .B(n5058), .Z(n5060) );
  NAND U5687 ( .A(n5061), .B(n5060), .Z(n5324) );
  NANDN U5688 ( .A(n5063), .B(n5062), .Z(n5067) );
  NAND U5689 ( .A(n5065), .B(n5064), .Z(n5066) );
  AND U5690 ( .A(n5067), .B(n5066), .Z(n5325) );
  XNOR U5691 ( .A(n5324), .B(n5325), .Z(n5326) );
  NANDN U5692 ( .A(n5069), .B(n5068), .Z(n5073) );
  NAND U5693 ( .A(n5071), .B(n5070), .Z(n5072) );
  NAND U5694 ( .A(n5073), .B(n5072), .Z(n5279) );
  NANDN U5695 ( .A(n5074), .B(n18832), .Z(n5076) );
  XOR U5696 ( .A(b[19]), .B(n6835), .Z(n5246) );
  NANDN U5697 ( .A(n5246), .B(n18834), .Z(n5075) );
  NAND U5698 ( .A(n5076), .B(n5075), .Z(n5291) );
  XNOR U5699 ( .A(b[27]), .B(a[21]), .Z(n5249) );
  NANDN U5700 ( .A(n5249), .B(n19336), .Z(n5079) );
  NANDN U5701 ( .A(n5077), .B(n19337), .Z(n5078) );
  NAND U5702 ( .A(n5079), .B(n5078), .Z(n5288) );
  XOR U5703 ( .A(b[5]), .B(a[43]), .Z(n5252) );
  NAND U5704 ( .A(n5252), .B(n17310), .Z(n5082) );
  NANDN U5705 ( .A(n5080), .B(n17311), .Z(n5081) );
  AND U5706 ( .A(n5082), .B(n5081), .Z(n5289) );
  XNOR U5707 ( .A(n5288), .B(n5289), .Z(n5290) );
  XNOR U5708 ( .A(n5291), .B(n5290), .Z(n5276) );
  XOR U5709 ( .A(b[17]), .B(a[31]), .Z(n5255) );
  NAND U5710 ( .A(n5255), .B(n18673), .Z(n5085) );
  NANDN U5711 ( .A(n5083), .B(n18674), .Z(n5084) );
  NAND U5712 ( .A(n5085), .B(n5084), .Z(n5230) );
  XNOR U5713 ( .A(b[31]), .B(a[17]), .Z(n5258) );
  NANDN U5714 ( .A(n5258), .B(n19472), .Z(n5088) );
  NANDN U5715 ( .A(n5086), .B(n19473), .Z(n5087) );
  AND U5716 ( .A(n5088), .B(n5087), .Z(n5228) );
  OR U5717 ( .A(n5089), .B(n16988), .Z(n5091) );
  XNOR U5718 ( .A(b[3]), .B(a[45]), .Z(n5261) );
  NANDN U5719 ( .A(n5261), .B(n16990), .Z(n5090) );
  AND U5720 ( .A(n5091), .B(n5090), .Z(n5229) );
  XOR U5721 ( .A(n5230), .B(n5231), .Z(n5277) );
  XOR U5722 ( .A(n5276), .B(n5277), .Z(n5278) );
  XNOR U5723 ( .A(n5279), .B(n5278), .Z(n5204) );
  NANDN U5724 ( .A(n5093), .B(n5092), .Z(n5097) );
  OR U5725 ( .A(n5095), .B(n5094), .Z(n5096) );
  NAND U5726 ( .A(n5097), .B(n5096), .Z(n5205) );
  XNOR U5727 ( .A(n5204), .B(n5205), .Z(n5206) );
  NANDN U5728 ( .A(n5099), .B(n5098), .Z(n5103) );
  NAND U5729 ( .A(n5101), .B(n5100), .Z(n5102) );
  NAND U5730 ( .A(n5103), .B(n5102), .Z(n5267) );
  NANDN U5731 ( .A(n5105), .B(n5104), .Z(n5109) );
  NAND U5732 ( .A(n5107), .B(n5106), .Z(n5108) );
  NAND U5733 ( .A(n5109), .B(n5108), .Z(n5264) );
  OR U5734 ( .A(n5111), .B(n5110), .Z(n5115) );
  NANDN U5735 ( .A(n5113), .B(n5112), .Z(n5114) );
  NAND U5736 ( .A(n5115), .B(n5114), .Z(n5265) );
  XNOR U5737 ( .A(n5264), .B(n5265), .Z(n5266) );
  XOR U5738 ( .A(n5267), .B(n5266), .Z(n5207) );
  XNOR U5739 ( .A(n5206), .B(n5207), .Z(n5332) );
  NANDN U5740 ( .A(n5121), .B(n5120), .Z(n5125) );
  NANDN U5741 ( .A(n5123), .B(n5122), .Z(n5124) );
  NAND U5742 ( .A(n5125), .B(n5124), .Z(n5213) );
  NANDN U5743 ( .A(n5127), .B(n5126), .Z(n5131) );
  OR U5744 ( .A(n5129), .B(n5128), .Z(n5130) );
  NAND U5745 ( .A(n5131), .B(n5130), .Z(n5211) );
  NANDN U5746 ( .A(n5133), .B(n5132), .Z(n5137) );
  NAND U5747 ( .A(n5135), .B(n5134), .Z(n5136) );
  NAND U5748 ( .A(n5137), .B(n5136), .Z(n5270) );
  NANDN U5749 ( .A(n5139), .B(n5138), .Z(n5143) );
  NAND U5750 ( .A(n5141), .B(n5140), .Z(n5142) );
  AND U5751 ( .A(n5143), .B(n5142), .Z(n5271) );
  XNOR U5752 ( .A(n5270), .B(n5271), .Z(n5272) );
  XNOR U5753 ( .A(n579), .B(a[39]), .Z(n5300) );
  NAND U5754 ( .A(n17814), .B(n5300), .Z(n5146) );
  NANDN U5755 ( .A(n5144), .B(n17815), .Z(n5145) );
  NAND U5756 ( .A(n5146), .B(n5145), .Z(n5236) );
  NAND U5757 ( .A(n5147), .B(n18513), .Z(n5149) );
  XOR U5758 ( .A(b[15]), .B(a[33]), .Z(n5297) );
  NANDN U5759 ( .A(n18512), .B(n5297), .Z(n5148) );
  AND U5760 ( .A(n5149), .B(n5148), .Z(n5234) );
  NANDN U5761 ( .A(n5150), .B(n19013), .Z(n5152) );
  XNOR U5762 ( .A(n582), .B(a[27]), .Z(n5294) );
  NAND U5763 ( .A(n5294), .B(n19015), .Z(n5151) );
  AND U5764 ( .A(n5152), .B(n5151), .Z(n5235) );
  XOR U5765 ( .A(n5236), .B(n5237), .Z(n5225) );
  XNOR U5766 ( .A(b[11]), .B(a[37]), .Z(n5303) );
  OR U5767 ( .A(n5303), .B(n18194), .Z(n5155) );
  NANDN U5768 ( .A(n5153), .B(n18104), .Z(n5154) );
  NAND U5769 ( .A(n5155), .B(n5154), .Z(n5223) );
  XOR U5770 ( .A(n580), .B(a[35]), .Z(n5306) );
  NANDN U5771 ( .A(n5306), .B(n18336), .Z(n5158) );
  NANDN U5772 ( .A(n5156), .B(n18337), .Z(n5157) );
  NAND U5773 ( .A(n5158), .B(n5157), .Z(n5222) );
  XOR U5774 ( .A(n5225), .B(n5224), .Z(n5219) );
  ANDN U5775 ( .B(b[31]), .A(n5159), .Z(n5240) );
  NANDN U5776 ( .A(n5160), .B(n19406), .Z(n5162) );
  XNOR U5777 ( .A(n584), .B(a[19]), .Z(n5312) );
  NANDN U5778 ( .A(n576), .B(n5312), .Z(n5161) );
  NAND U5779 ( .A(n5162), .B(n5161), .Z(n5241) );
  XOR U5780 ( .A(n5240), .B(n5241), .Z(n5242) );
  NANDN U5781 ( .A(n577), .B(a[47]), .Z(n5163) );
  XOR U5782 ( .A(n17151), .B(n5163), .Z(n5165) );
  NANDN U5783 ( .A(b[0]), .B(a[46]), .Z(n5164) );
  AND U5784 ( .A(n5165), .B(n5164), .Z(n5243) );
  XNOR U5785 ( .A(n5242), .B(n5243), .Z(n5216) );
  XOR U5786 ( .A(b[23]), .B(a[25]), .Z(n5315) );
  NANDN U5787 ( .A(n19127), .B(n5315), .Z(n5168) );
  NAND U5788 ( .A(n5166), .B(n19128), .Z(n5167) );
  NAND U5789 ( .A(n5168), .B(n5167), .Z(n5285) );
  NAND U5790 ( .A(n5169), .B(n17553), .Z(n5171) );
  XNOR U5791 ( .A(b[7]), .B(a[41]), .Z(n5318) );
  NANDN U5792 ( .A(n5318), .B(n17555), .Z(n5170) );
  NAND U5793 ( .A(n5171), .B(n5170), .Z(n5282) );
  XOR U5794 ( .A(b[25]), .B(a[23]), .Z(n5321) );
  NAND U5795 ( .A(n5321), .B(n19240), .Z(n5174) );
  NAND U5796 ( .A(n5172), .B(n19242), .Z(n5173) );
  AND U5797 ( .A(n5174), .B(n5173), .Z(n5283) );
  XNOR U5798 ( .A(n5282), .B(n5283), .Z(n5284) );
  XNOR U5799 ( .A(n5285), .B(n5284), .Z(n5217) );
  XOR U5800 ( .A(n5219), .B(n5218), .Z(n5273) );
  XNOR U5801 ( .A(n5272), .B(n5273), .Z(n5210) );
  XOR U5802 ( .A(n5211), .B(n5210), .Z(n5212) );
  XNOR U5803 ( .A(n5213), .B(n5212), .Z(n5330) );
  XNOR U5804 ( .A(n5331), .B(n5330), .Z(n5333) );
  XNOR U5805 ( .A(n5332), .B(n5333), .Z(n5327) );
  XOR U5806 ( .A(n5326), .B(n5327), .Z(n5201) );
  NANDN U5807 ( .A(n5176), .B(n5175), .Z(n5180) );
  NAND U5808 ( .A(n5178), .B(n5177), .Z(n5179) );
  NAND U5809 ( .A(n5180), .B(n5179), .Z(n5198) );
  NANDN U5810 ( .A(n5182), .B(n5181), .Z(n5186) );
  NANDN U5811 ( .A(n5184), .B(n5183), .Z(n5185) );
  NAND U5812 ( .A(n5186), .B(n5185), .Z(n5199) );
  XNOR U5813 ( .A(n5198), .B(n5199), .Z(n5200) );
  XNOR U5814 ( .A(n5201), .B(n5200), .Z(n5193) );
  XNOR U5815 ( .A(n5192), .B(n5193), .Z(n5194) );
  XNOR U5816 ( .A(n5195), .B(n5194), .Z(n5336) );
  XNOR U5817 ( .A(n5336), .B(sreg[143]), .Z(n5338) );
  NAND U5818 ( .A(n5187), .B(sreg[142]), .Z(n5191) );
  OR U5819 ( .A(n5189), .B(n5188), .Z(n5190) );
  AND U5820 ( .A(n5191), .B(n5190), .Z(n5337) );
  XOR U5821 ( .A(n5338), .B(n5337), .Z(c[143]) );
  NANDN U5822 ( .A(n5193), .B(n5192), .Z(n5197) );
  NAND U5823 ( .A(n5195), .B(n5194), .Z(n5196) );
  NAND U5824 ( .A(n5197), .B(n5196), .Z(n5344) );
  NANDN U5825 ( .A(n5199), .B(n5198), .Z(n5203) );
  NAND U5826 ( .A(n5201), .B(n5200), .Z(n5202) );
  NAND U5827 ( .A(n5203), .B(n5202), .Z(n5342) );
  NANDN U5828 ( .A(n5205), .B(n5204), .Z(n5209) );
  NANDN U5829 ( .A(n5207), .B(n5206), .Z(n5208) );
  NAND U5830 ( .A(n5209), .B(n5208), .Z(n5477) );
  NAND U5831 ( .A(n5211), .B(n5210), .Z(n5215) );
  NAND U5832 ( .A(n5213), .B(n5212), .Z(n5214) );
  NAND U5833 ( .A(n5215), .B(n5214), .Z(n5478) );
  XNOR U5834 ( .A(n5477), .B(n5478), .Z(n5479) );
  OR U5835 ( .A(n5217), .B(n5216), .Z(n5221) );
  NANDN U5836 ( .A(n5219), .B(n5218), .Z(n5220) );
  NAND U5837 ( .A(n5221), .B(n5220), .Z(n5462) );
  OR U5838 ( .A(n5223), .B(n5222), .Z(n5227) );
  NAND U5839 ( .A(n5225), .B(n5224), .Z(n5226) );
  NAND U5840 ( .A(n5227), .B(n5226), .Z(n5401) );
  OR U5841 ( .A(n5229), .B(n5228), .Z(n5233) );
  NANDN U5842 ( .A(n5231), .B(n5230), .Z(n5232) );
  NAND U5843 ( .A(n5233), .B(n5232), .Z(n5400) );
  OR U5844 ( .A(n5235), .B(n5234), .Z(n5239) );
  NANDN U5845 ( .A(n5237), .B(n5236), .Z(n5238) );
  NAND U5846 ( .A(n5239), .B(n5238), .Z(n5399) );
  XOR U5847 ( .A(n5401), .B(n5402), .Z(n5460) );
  OR U5848 ( .A(n5241), .B(n5240), .Z(n5245) );
  NANDN U5849 ( .A(n5243), .B(n5242), .Z(n5244) );
  NAND U5850 ( .A(n5245), .B(n5244), .Z(n5413) );
  NANDN U5851 ( .A(n5246), .B(n18832), .Z(n5248) );
  XOR U5852 ( .A(b[19]), .B(n7336), .Z(n5359) );
  NANDN U5853 ( .A(n5359), .B(n18834), .Z(n5247) );
  NAND U5854 ( .A(n5248), .B(n5247), .Z(n5426) );
  XNOR U5855 ( .A(b[27]), .B(a[22]), .Z(n5362) );
  NANDN U5856 ( .A(n5362), .B(n19336), .Z(n5251) );
  NANDN U5857 ( .A(n5249), .B(n19337), .Z(n5250) );
  NAND U5858 ( .A(n5251), .B(n5250), .Z(n5423) );
  XOR U5859 ( .A(b[5]), .B(a[44]), .Z(n5365) );
  NAND U5860 ( .A(n5365), .B(n17310), .Z(n5254) );
  NAND U5861 ( .A(n5252), .B(n17311), .Z(n5253) );
  AND U5862 ( .A(n5254), .B(n5253), .Z(n5424) );
  XNOR U5863 ( .A(n5423), .B(n5424), .Z(n5425) );
  XNOR U5864 ( .A(n5426), .B(n5425), .Z(n5412) );
  XOR U5865 ( .A(b[17]), .B(a[32]), .Z(n5368) );
  NAND U5866 ( .A(n5368), .B(n18673), .Z(n5257) );
  NAND U5867 ( .A(n5255), .B(n18674), .Z(n5256) );
  NAND U5868 ( .A(n5257), .B(n5256), .Z(n5386) );
  XNOR U5869 ( .A(b[31]), .B(a[18]), .Z(n5371) );
  NANDN U5870 ( .A(n5371), .B(n19472), .Z(n5260) );
  NANDN U5871 ( .A(n5258), .B(n19473), .Z(n5259) );
  NAND U5872 ( .A(n5260), .B(n5259), .Z(n5383) );
  OR U5873 ( .A(n5261), .B(n16988), .Z(n5263) );
  XNOR U5874 ( .A(b[3]), .B(a[46]), .Z(n5374) );
  NANDN U5875 ( .A(n5374), .B(n16990), .Z(n5262) );
  AND U5876 ( .A(n5263), .B(n5262), .Z(n5384) );
  XNOR U5877 ( .A(n5383), .B(n5384), .Z(n5385) );
  XOR U5878 ( .A(n5386), .B(n5385), .Z(n5411) );
  XOR U5879 ( .A(n5412), .B(n5411), .Z(n5414) );
  XOR U5880 ( .A(n5413), .B(n5414), .Z(n5459) );
  XOR U5881 ( .A(n5460), .B(n5459), .Z(n5461) );
  XNOR U5882 ( .A(n5462), .B(n5461), .Z(n5474) );
  NANDN U5883 ( .A(n5265), .B(n5264), .Z(n5269) );
  NANDN U5884 ( .A(n5267), .B(n5266), .Z(n5268) );
  NAND U5885 ( .A(n5269), .B(n5268), .Z(n5471) );
  NANDN U5886 ( .A(n5271), .B(n5270), .Z(n5275) );
  NANDN U5887 ( .A(n5273), .B(n5272), .Z(n5274) );
  NAND U5888 ( .A(n5275), .B(n5274), .Z(n5468) );
  OR U5889 ( .A(n5277), .B(n5276), .Z(n5281) );
  NAND U5890 ( .A(n5279), .B(n5278), .Z(n5280) );
  NAND U5891 ( .A(n5281), .B(n5280), .Z(n5466) );
  NANDN U5892 ( .A(n5283), .B(n5282), .Z(n5287) );
  NAND U5893 ( .A(n5285), .B(n5284), .Z(n5286) );
  NAND U5894 ( .A(n5287), .B(n5286), .Z(n5405) );
  NANDN U5895 ( .A(n5289), .B(n5288), .Z(n5293) );
  NAND U5896 ( .A(n5291), .B(n5290), .Z(n5292) );
  AND U5897 ( .A(n5293), .B(n5292), .Z(n5406) );
  XNOR U5898 ( .A(n5405), .B(n5406), .Z(n5407) );
  XNOR U5899 ( .A(b[21]), .B(a[28]), .Z(n5435) );
  NANDN U5900 ( .A(n5435), .B(n19015), .Z(n5296) );
  NAND U5901 ( .A(n19013), .B(n5294), .Z(n5295) );
  NAND U5902 ( .A(n5296), .B(n5295), .Z(n5395) );
  NAND U5903 ( .A(n5297), .B(n18513), .Z(n5299) );
  XOR U5904 ( .A(b[15]), .B(a[34]), .Z(n5432) );
  NANDN U5905 ( .A(n18512), .B(n5432), .Z(n5298) );
  AND U5906 ( .A(n5299), .B(n5298), .Z(n5396) );
  XNOR U5907 ( .A(n5395), .B(n5396), .Z(n5398) );
  XNOR U5908 ( .A(b[9]), .B(a[40]), .Z(n5429) );
  NANDN U5909 ( .A(n5429), .B(n17814), .Z(n5302) );
  NAND U5910 ( .A(n17815), .B(n5300), .Z(n5301) );
  NAND U5911 ( .A(n5302), .B(n5301), .Z(n5397) );
  XNOR U5912 ( .A(n5398), .B(n5397), .Z(n5391) );
  XOR U5913 ( .A(b[11]), .B(n8490), .Z(n5438) );
  OR U5914 ( .A(n5438), .B(n18194), .Z(n5305) );
  NANDN U5915 ( .A(n5303), .B(n18104), .Z(n5304) );
  NAND U5916 ( .A(n5305), .B(n5304), .Z(n5390) );
  XOR U5917 ( .A(n580), .B(a[36]), .Z(n5441) );
  NANDN U5918 ( .A(n5441), .B(n18336), .Z(n5308) );
  NANDN U5919 ( .A(n5306), .B(n18337), .Z(n5307) );
  NAND U5920 ( .A(n5308), .B(n5307), .Z(n5389) );
  XNOR U5921 ( .A(n5390), .B(n5389), .Z(n5392) );
  XNOR U5922 ( .A(n5391), .B(n5392), .Z(n5380) );
  NANDN U5923 ( .A(n577), .B(a[48]), .Z(n5309) );
  XOR U5924 ( .A(n17151), .B(n5309), .Z(n5311) );
  NANDN U5925 ( .A(b[0]), .B(a[47]), .Z(n5310) );
  AND U5926 ( .A(n5311), .B(n5310), .Z(n5355) );
  NAND U5927 ( .A(n5312), .B(n19406), .Z(n5314) );
  XNOR U5928 ( .A(n584), .B(a[20]), .Z(n5447) );
  NANDN U5929 ( .A(n576), .B(n5447), .Z(n5313) );
  NAND U5930 ( .A(n5314), .B(n5313), .Z(n5353) );
  NANDN U5931 ( .A(n585), .B(a[16]), .Z(n5354) );
  XNOR U5932 ( .A(n5353), .B(n5354), .Z(n5356) );
  XNOR U5933 ( .A(n5355), .B(n5356), .Z(n5378) );
  XOR U5934 ( .A(b[23]), .B(a[26]), .Z(n5450) );
  NANDN U5935 ( .A(n19127), .B(n5450), .Z(n5317) );
  NAND U5936 ( .A(n5315), .B(n19128), .Z(n5316) );
  NAND U5937 ( .A(n5317), .B(n5316), .Z(n5420) );
  NANDN U5938 ( .A(n5318), .B(n17553), .Z(n5320) );
  XNOR U5939 ( .A(b[7]), .B(a[42]), .Z(n5453) );
  NANDN U5940 ( .A(n5453), .B(n17555), .Z(n5319) );
  NAND U5941 ( .A(n5320), .B(n5319), .Z(n5417) );
  XOR U5942 ( .A(b[25]), .B(a[24]), .Z(n5456) );
  NAND U5943 ( .A(n5456), .B(n19240), .Z(n5323) );
  NAND U5944 ( .A(n5321), .B(n19242), .Z(n5322) );
  AND U5945 ( .A(n5323), .B(n5322), .Z(n5418) );
  XNOR U5946 ( .A(n5417), .B(n5418), .Z(n5419) );
  XOR U5947 ( .A(n5420), .B(n5419), .Z(n5377) );
  XOR U5948 ( .A(n5380), .B(n5379), .Z(n5408) );
  XNOR U5949 ( .A(n5407), .B(n5408), .Z(n5465) );
  XOR U5950 ( .A(n5466), .B(n5465), .Z(n5467) );
  XOR U5951 ( .A(n5468), .B(n5467), .Z(n5472) );
  XNOR U5952 ( .A(n5471), .B(n5472), .Z(n5473) );
  XOR U5953 ( .A(n5474), .B(n5473), .Z(n5480) );
  XOR U5954 ( .A(n5479), .B(n5480), .Z(n5349) );
  NANDN U5955 ( .A(n5325), .B(n5324), .Z(n5329) );
  NANDN U5956 ( .A(n5327), .B(n5326), .Z(n5328) );
  NAND U5957 ( .A(n5329), .B(n5328), .Z(n5348) );
  OR U5958 ( .A(n5331), .B(n5330), .Z(n5335) );
  OR U5959 ( .A(n5333), .B(n5332), .Z(n5334) );
  AND U5960 ( .A(n5335), .B(n5334), .Z(n5347) );
  XNOR U5961 ( .A(n5348), .B(n5347), .Z(n5350) );
  XOR U5962 ( .A(n5349), .B(n5350), .Z(n5341) );
  XOR U5963 ( .A(n5342), .B(n5341), .Z(n5343) );
  XNOR U5964 ( .A(n5344), .B(n5343), .Z(n5483) );
  XNOR U5965 ( .A(n5483), .B(sreg[144]), .Z(n5485) );
  NAND U5966 ( .A(n5336), .B(sreg[143]), .Z(n5340) );
  OR U5967 ( .A(n5338), .B(n5337), .Z(n5339) );
  AND U5968 ( .A(n5340), .B(n5339), .Z(n5484) );
  XOR U5969 ( .A(n5485), .B(n5484), .Z(c[144]) );
  NAND U5970 ( .A(n5342), .B(n5341), .Z(n5346) );
  NAND U5971 ( .A(n5344), .B(n5343), .Z(n5345) );
  NAND U5972 ( .A(n5346), .B(n5345), .Z(n5491) );
  NANDN U5973 ( .A(n5348), .B(n5347), .Z(n5352) );
  NAND U5974 ( .A(n5350), .B(n5349), .Z(n5351) );
  NAND U5975 ( .A(n5352), .B(n5351), .Z(n5489) );
  NANDN U5976 ( .A(n5354), .B(n5353), .Z(n5358) );
  NAND U5977 ( .A(n5356), .B(n5355), .Z(n5357) );
  NAND U5978 ( .A(n5358), .B(n5357), .Z(n5561) );
  NANDN U5979 ( .A(n5359), .B(n18832), .Z(n5361) );
  XNOR U5980 ( .A(b[19]), .B(a[31]), .Z(n5506) );
  NANDN U5981 ( .A(n5506), .B(n18834), .Z(n5360) );
  NAND U5982 ( .A(n5361), .B(n5360), .Z(n5571) );
  XNOR U5983 ( .A(b[27]), .B(a[23]), .Z(n5509) );
  NANDN U5984 ( .A(n5509), .B(n19336), .Z(n5364) );
  NANDN U5985 ( .A(n5362), .B(n19337), .Z(n5363) );
  NAND U5986 ( .A(n5364), .B(n5363), .Z(n5568) );
  XOR U5987 ( .A(b[5]), .B(a[45]), .Z(n5512) );
  NAND U5988 ( .A(n5512), .B(n17310), .Z(n5367) );
  NAND U5989 ( .A(n5365), .B(n17311), .Z(n5366) );
  AND U5990 ( .A(n5367), .B(n5366), .Z(n5569) );
  XNOR U5991 ( .A(n5568), .B(n5569), .Z(n5570) );
  XNOR U5992 ( .A(n5571), .B(n5570), .Z(n5559) );
  XOR U5993 ( .A(b[17]), .B(a[33]), .Z(n5515) );
  NAND U5994 ( .A(n5515), .B(n18673), .Z(n5370) );
  NAND U5995 ( .A(n5368), .B(n18674), .Z(n5369) );
  NAND U5996 ( .A(n5370), .B(n5369), .Z(n5533) );
  XNOR U5997 ( .A(b[31]), .B(a[19]), .Z(n5518) );
  NANDN U5998 ( .A(n5518), .B(n19472), .Z(n5373) );
  NANDN U5999 ( .A(n5371), .B(n19473), .Z(n5372) );
  NAND U6000 ( .A(n5373), .B(n5372), .Z(n5530) );
  OR U6001 ( .A(n5374), .B(n16988), .Z(n5376) );
  XNOR U6002 ( .A(b[3]), .B(a[47]), .Z(n5521) );
  NANDN U6003 ( .A(n5521), .B(n16990), .Z(n5375) );
  AND U6004 ( .A(n5376), .B(n5375), .Z(n5531) );
  XNOR U6005 ( .A(n5530), .B(n5531), .Z(n5532) );
  XOR U6006 ( .A(n5533), .B(n5532), .Z(n5558) );
  XNOR U6007 ( .A(n5559), .B(n5558), .Z(n5560) );
  XNOR U6008 ( .A(n5561), .B(n5560), .Z(n5610) );
  NANDN U6009 ( .A(n5378), .B(n5377), .Z(n5382) );
  NANDN U6010 ( .A(n5380), .B(n5379), .Z(n5381) );
  NAND U6011 ( .A(n5382), .B(n5381), .Z(n5611) );
  XNOR U6012 ( .A(n5610), .B(n5611), .Z(n5612) );
  NANDN U6013 ( .A(n5384), .B(n5383), .Z(n5388) );
  NAND U6014 ( .A(n5386), .B(n5385), .Z(n5387) );
  NAND U6015 ( .A(n5388), .B(n5387), .Z(n5551) );
  OR U6016 ( .A(n5390), .B(n5389), .Z(n5394) );
  NANDN U6017 ( .A(n5392), .B(n5391), .Z(n5393) );
  NAND U6018 ( .A(n5394), .B(n5393), .Z(n5549) );
  XNOR U6019 ( .A(n5549), .B(n5548), .Z(n5550) );
  XOR U6020 ( .A(n5551), .B(n5550), .Z(n5613) );
  XOR U6021 ( .A(n5612), .B(n5613), .Z(n5623) );
  OR U6022 ( .A(n5400), .B(n5399), .Z(n5404) );
  NANDN U6023 ( .A(n5402), .B(n5401), .Z(n5403) );
  NAND U6024 ( .A(n5404), .B(n5403), .Z(n5621) );
  NANDN U6025 ( .A(n5406), .B(n5405), .Z(n5410) );
  NANDN U6026 ( .A(n5408), .B(n5407), .Z(n5409) );
  NAND U6027 ( .A(n5410), .B(n5409), .Z(n5606) );
  NANDN U6028 ( .A(n5412), .B(n5411), .Z(n5416) );
  OR U6029 ( .A(n5414), .B(n5413), .Z(n5415) );
  NAND U6030 ( .A(n5416), .B(n5415), .Z(n5605) );
  NANDN U6031 ( .A(n5418), .B(n5417), .Z(n5422) );
  NAND U6032 ( .A(n5420), .B(n5419), .Z(n5421) );
  NAND U6033 ( .A(n5422), .B(n5421), .Z(n5552) );
  NANDN U6034 ( .A(n5424), .B(n5423), .Z(n5428) );
  NAND U6035 ( .A(n5426), .B(n5425), .Z(n5427) );
  AND U6036 ( .A(n5428), .B(n5427), .Z(n5553) );
  XNOR U6037 ( .A(n5552), .B(n5553), .Z(n5554) );
  XOR U6038 ( .A(n579), .B(n8930), .Z(n5574) );
  NAND U6039 ( .A(n17814), .B(n5574), .Z(n5431) );
  NANDN U6040 ( .A(n5429), .B(n17815), .Z(n5430) );
  NAND U6041 ( .A(n5431), .B(n5430), .Z(n5538) );
  NAND U6042 ( .A(n5432), .B(n18513), .Z(n5434) );
  XOR U6043 ( .A(b[15]), .B(a[35]), .Z(n5577) );
  NANDN U6044 ( .A(n18512), .B(n5577), .Z(n5433) );
  AND U6045 ( .A(n5434), .B(n5433), .Z(n5536) );
  NANDN U6046 ( .A(n5435), .B(n19013), .Z(n5437) );
  XOR U6047 ( .A(n582), .B(n6835), .Z(n5580) );
  NAND U6048 ( .A(n5580), .B(n19015), .Z(n5436) );
  AND U6049 ( .A(n5437), .B(n5436), .Z(n5537) );
  XOR U6050 ( .A(n5538), .B(n5539), .Z(n5527) );
  XNOR U6051 ( .A(b[11]), .B(a[39]), .Z(n5583) );
  OR U6052 ( .A(n5583), .B(n18194), .Z(n5440) );
  NANDN U6053 ( .A(n5438), .B(n18104), .Z(n5439) );
  NAND U6054 ( .A(n5440), .B(n5439), .Z(n5525) );
  XOR U6055 ( .A(n580), .B(a[37]), .Z(n5586) );
  NANDN U6056 ( .A(n5586), .B(n18336), .Z(n5443) );
  NANDN U6057 ( .A(n5441), .B(n18337), .Z(n5442) );
  AND U6058 ( .A(n5443), .B(n5442), .Z(n5524) );
  XNOR U6059 ( .A(n5525), .B(n5524), .Z(n5526) );
  XOR U6060 ( .A(n5527), .B(n5526), .Z(n5544) );
  NANDN U6061 ( .A(n577), .B(a[49]), .Z(n5444) );
  XOR U6062 ( .A(n17151), .B(n5444), .Z(n5446) );
  NANDN U6063 ( .A(b[0]), .B(a[48]), .Z(n5445) );
  AND U6064 ( .A(n5446), .B(n5445), .Z(n5502) );
  NAND U6065 ( .A(n19406), .B(n5447), .Z(n5449) );
  XNOR U6066 ( .A(n584), .B(a[21]), .Z(n5592) );
  NANDN U6067 ( .A(n576), .B(n5592), .Z(n5448) );
  NAND U6068 ( .A(n5449), .B(n5448), .Z(n5500) );
  NANDN U6069 ( .A(n585), .B(a[17]), .Z(n5501) );
  XNOR U6070 ( .A(n5500), .B(n5501), .Z(n5503) );
  XOR U6071 ( .A(n5502), .B(n5503), .Z(n5542) );
  XOR U6072 ( .A(b[23]), .B(a[27]), .Z(n5595) );
  NANDN U6073 ( .A(n19127), .B(n5595), .Z(n5452) );
  NAND U6074 ( .A(n5450), .B(n19128), .Z(n5451) );
  NAND U6075 ( .A(n5452), .B(n5451), .Z(n5565) );
  NANDN U6076 ( .A(n5453), .B(n17553), .Z(n5455) );
  XOR U6077 ( .A(b[7]), .B(a[43]), .Z(n5598) );
  NAND U6078 ( .A(n5598), .B(n17555), .Z(n5454) );
  NAND U6079 ( .A(n5455), .B(n5454), .Z(n5562) );
  XOR U6080 ( .A(b[25]), .B(a[25]), .Z(n5601) );
  NAND U6081 ( .A(n5601), .B(n19240), .Z(n5458) );
  NAND U6082 ( .A(n5456), .B(n19242), .Z(n5457) );
  AND U6083 ( .A(n5458), .B(n5457), .Z(n5563) );
  XNOR U6084 ( .A(n5562), .B(n5563), .Z(n5564) );
  XNOR U6085 ( .A(n5565), .B(n5564), .Z(n5543) );
  XOR U6086 ( .A(n5542), .B(n5543), .Z(n5545) );
  XNOR U6087 ( .A(n5544), .B(n5545), .Z(n5555) );
  XNOR U6088 ( .A(n5554), .B(n5555), .Z(n5604) );
  XNOR U6089 ( .A(n5605), .B(n5604), .Z(n5607) );
  XNOR U6090 ( .A(n5606), .B(n5607), .Z(n5620) );
  XOR U6091 ( .A(n5621), .B(n5620), .Z(n5622) );
  XNOR U6092 ( .A(n5623), .B(n5622), .Z(n5617) );
  NAND U6093 ( .A(n5460), .B(n5459), .Z(n5464) );
  NAND U6094 ( .A(n5462), .B(n5461), .Z(n5463) );
  NAND U6095 ( .A(n5464), .B(n5463), .Z(n5615) );
  NAND U6096 ( .A(n5466), .B(n5465), .Z(n5470) );
  NAND U6097 ( .A(n5468), .B(n5467), .Z(n5469) );
  AND U6098 ( .A(n5470), .B(n5469), .Z(n5614) );
  XNOR U6099 ( .A(n5615), .B(n5614), .Z(n5616) );
  XOR U6100 ( .A(n5617), .B(n5616), .Z(n5496) );
  NANDN U6101 ( .A(n5472), .B(n5471), .Z(n5476) );
  NAND U6102 ( .A(n5474), .B(n5473), .Z(n5475) );
  NAND U6103 ( .A(n5476), .B(n5475), .Z(n5494) );
  NANDN U6104 ( .A(n5478), .B(n5477), .Z(n5482) );
  NAND U6105 ( .A(n5480), .B(n5479), .Z(n5481) );
  AND U6106 ( .A(n5482), .B(n5481), .Z(n5495) );
  XNOR U6107 ( .A(n5494), .B(n5495), .Z(n5497) );
  XOR U6108 ( .A(n5496), .B(n5497), .Z(n5488) );
  XOR U6109 ( .A(n5489), .B(n5488), .Z(n5490) );
  XNOR U6110 ( .A(n5491), .B(n5490), .Z(n5626) );
  XNOR U6111 ( .A(n5626), .B(sreg[145]), .Z(n5628) );
  NAND U6112 ( .A(n5483), .B(sreg[144]), .Z(n5487) );
  OR U6113 ( .A(n5485), .B(n5484), .Z(n5486) );
  AND U6114 ( .A(n5487), .B(n5486), .Z(n5627) );
  XOR U6115 ( .A(n5628), .B(n5627), .Z(c[145]) );
  NAND U6116 ( .A(n5489), .B(n5488), .Z(n5493) );
  NAND U6117 ( .A(n5491), .B(n5490), .Z(n5492) );
  NAND U6118 ( .A(n5493), .B(n5492), .Z(n5634) );
  NANDN U6119 ( .A(n5495), .B(n5494), .Z(n5499) );
  NAND U6120 ( .A(n5497), .B(n5496), .Z(n5498) );
  NAND U6121 ( .A(n5499), .B(n5498), .Z(n5632) );
  NANDN U6122 ( .A(n5501), .B(n5500), .Z(n5505) );
  NAND U6123 ( .A(n5503), .B(n5502), .Z(n5504) );
  NAND U6124 ( .A(n5505), .B(n5504), .Z(n5702) );
  NANDN U6125 ( .A(n5506), .B(n18832), .Z(n5508) );
  XNOR U6126 ( .A(b[19]), .B(a[32]), .Z(n5647) );
  NANDN U6127 ( .A(n5647), .B(n18834), .Z(n5507) );
  NAND U6128 ( .A(n5508), .B(n5507), .Z(n5712) );
  XNOR U6129 ( .A(b[27]), .B(a[24]), .Z(n5650) );
  NANDN U6130 ( .A(n5650), .B(n19336), .Z(n5511) );
  NANDN U6131 ( .A(n5509), .B(n19337), .Z(n5510) );
  NAND U6132 ( .A(n5511), .B(n5510), .Z(n5709) );
  XOR U6133 ( .A(b[5]), .B(a[46]), .Z(n5653) );
  NAND U6134 ( .A(n5653), .B(n17310), .Z(n5514) );
  NAND U6135 ( .A(n5512), .B(n17311), .Z(n5513) );
  AND U6136 ( .A(n5514), .B(n5513), .Z(n5710) );
  XNOR U6137 ( .A(n5709), .B(n5710), .Z(n5711) );
  XNOR U6138 ( .A(n5712), .B(n5711), .Z(n5700) );
  XOR U6139 ( .A(b[17]), .B(a[34]), .Z(n5656) );
  NAND U6140 ( .A(n5656), .B(n18673), .Z(n5517) );
  NAND U6141 ( .A(n5515), .B(n18674), .Z(n5516) );
  NAND U6142 ( .A(n5517), .B(n5516), .Z(n5674) );
  XNOR U6143 ( .A(b[31]), .B(a[20]), .Z(n5659) );
  NANDN U6144 ( .A(n5659), .B(n19472), .Z(n5520) );
  NANDN U6145 ( .A(n5518), .B(n19473), .Z(n5519) );
  NAND U6146 ( .A(n5520), .B(n5519), .Z(n5671) );
  OR U6147 ( .A(n5521), .B(n16988), .Z(n5523) );
  XNOR U6148 ( .A(b[3]), .B(a[48]), .Z(n5662) );
  NANDN U6149 ( .A(n5662), .B(n16990), .Z(n5522) );
  AND U6150 ( .A(n5523), .B(n5522), .Z(n5672) );
  XNOR U6151 ( .A(n5671), .B(n5672), .Z(n5673) );
  XOR U6152 ( .A(n5674), .B(n5673), .Z(n5699) );
  XNOR U6153 ( .A(n5700), .B(n5699), .Z(n5701) );
  XNOR U6154 ( .A(n5702), .B(n5701), .Z(n5745) );
  NANDN U6155 ( .A(n5525), .B(n5524), .Z(n5529) );
  NAND U6156 ( .A(n5527), .B(n5526), .Z(n5528) );
  NAND U6157 ( .A(n5529), .B(n5528), .Z(n5690) );
  NANDN U6158 ( .A(n5531), .B(n5530), .Z(n5535) );
  NAND U6159 ( .A(n5533), .B(n5532), .Z(n5534) );
  NAND U6160 ( .A(n5535), .B(n5534), .Z(n5688) );
  OR U6161 ( .A(n5537), .B(n5536), .Z(n5541) );
  NANDN U6162 ( .A(n5539), .B(n5538), .Z(n5540) );
  NAND U6163 ( .A(n5541), .B(n5540), .Z(n5687) );
  XNOR U6164 ( .A(n5690), .B(n5689), .Z(n5746) );
  XNOR U6165 ( .A(n5745), .B(n5746), .Z(n5747) );
  NANDN U6166 ( .A(n5543), .B(n5542), .Z(n5547) );
  OR U6167 ( .A(n5545), .B(n5544), .Z(n5546) );
  AND U6168 ( .A(n5547), .B(n5546), .Z(n5748) );
  XNOR U6169 ( .A(n5747), .B(n5748), .Z(n5760) );
  NANDN U6170 ( .A(n5553), .B(n5552), .Z(n5557) );
  NANDN U6171 ( .A(n5555), .B(n5554), .Z(n5556) );
  NAND U6172 ( .A(n5557), .B(n5556), .Z(n5754) );
  NANDN U6173 ( .A(n5563), .B(n5562), .Z(n5567) );
  NAND U6174 ( .A(n5565), .B(n5564), .Z(n5566) );
  NAND U6175 ( .A(n5567), .B(n5566), .Z(n5693) );
  NANDN U6176 ( .A(n5569), .B(n5568), .Z(n5573) );
  NAND U6177 ( .A(n5571), .B(n5570), .Z(n5572) );
  AND U6178 ( .A(n5573), .B(n5572), .Z(n5694) );
  XNOR U6179 ( .A(n5693), .B(n5694), .Z(n5695) );
  XOR U6180 ( .A(b[9]), .B(n9080), .Z(n5715) );
  NANDN U6181 ( .A(n5715), .B(n17814), .Z(n5576) );
  NAND U6182 ( .A(n17815), .B(n5574), .Z(n5575) );
  NAND U6183 ( .A(n5576), .B(n5575), .Z(n5679) );
  XNOR U6184 ( .A(b[15]), .B(a[36]), .Z(n5718) );
  OR U6185 ( .A(n5718), .B(n18512), .Z(n5579) );
  NAND U6186 ( .A(n5577), .B(n18513), .Z(n5578) );
  NAND U6187 ( .A(n5579), .B(n5578), .Z(n5677) );
  XOR U6188 ( .A(b[21]), .B(n7336), .Z(n5721) );
  NANDN U6189 ( .A(n5721), .B(n19015), .Z(n5582) );
  NAND U6190 ( .A(n19013), .B(n5580), .Z(n5581) );
  NAND U6191 ( .A(n5582), .B(n5581), .Z(n5678) );
  XNOR U6192 ( .A(n5677), .B(n5678), .Z(n5680) );
  XOR U6193 ( .A(n5679), .B(n5680), .Z(n5668) );
  XNOR U6194 ( .A(b[11]), .B(a[40]), .Z(n5724) );
  OR U6195 ( .A(n5724), .B(n18194), .Z(n5585) );
  NANDN U6196 ( .A(n5583), .B(n18104), .Z(n5584) );
  NAND U6197 ( .A(n5585), .B(n5584), .Z(n5666) );
  XOR U6198 ( .A(n580), .B(a[38]), .Z(n5727) );
  NANDN U6199 ( .A(n5727), .B(n18336), .Z(n5588) );
  NANDN U6200 ( .A(n5586), .B(n18337), .Z(n5587) );
  AND U6201 ( .A(n5588), .B(n5587), .Z(n5665) );
  XNOR U6202 ( .A(n5666), .B(n5665), .Z(n5667) );
  XNOR U6203 ( .A(n5668), .B(n5667), .Z(n5684) );
  NANDN U6204 ( .A(n577), .B(a[50]), .Z(n5589) );
  XOR U6205 ( .A(n17151), .B(n5589), .Z(n5591) );
  IV U6206 ( .A(a[49]), .Z(n10083) );
  NANDN U6207 ( .A(n10083), .B(n577), .Z(n5590) );
  AND U6208 ( .A(n5591), .B(n5590), .Z(n5643) );
  NAND U6209 ( .A(n19406), .B(n5592), .Z(n5594) );
  XNOR U6210 ( .A(n584), .B(a[22]), .Z(n5733) );
  NANDN U6211 ( .A(n576), .B(n5733), .Z(n5593) );
  NAND U6212 ( .A(n5594), .B(n5593), .Z(n5641) );
  NANDN U6213 ( .A(n585), .B(a[18]), .Z(n5642) );
  XNOR U6214 ( .A(n5641), .B(n5642), .Z(n5644) );
  XNOR U6215 ( .A(n5643), .B(n5644), .Z(n5682) );
  XOR U6216 ( .A(b[23]), .B(a[28]), .Z(n5736) );
  NANDN U6217 ( .A(n19127), .B(n5736), .Z(n5597) );
  NAND U6218 ( .A(n5595), .B(n19128), .Z(n5596) );
  NAND U6219 ( .A(n5597), .B(n5596), .Z(n5706) );
  NAND U6220 ( .A(n5598), .B(n17553), .Z(n5600) );
  XOR U6221 ( .A(b[7]), .B(a[44]), .Z(n5739) );
  NAND U6222 ( .A(n5739), .B(n17555), .Z(n5599) );
  NAND U6223 ( .A(n5600), .B(n5599), .Z(n5703) );
  XOR U6224 ( .A(b[25]), .B(a[26]), .Z(n5742) );
  NAND U6225 ( .A(n5742), .B(n19240), .Z(n5603) );
  NAND U6226 ( .A(n5601), .B(n19242), .Z(n5602) );
  AND U6227 ( .A(n5603), .B(n5602), .Z(n5704) );
  XNOR U6228 ( .A(n5703), .B(n5704), .Z(n5705) );
  XOR U6229 ( .A(n5706), .B(n5705), .Z(n5681) );
  XOR U6230 ( .A(n5684), .B(n5683), .Z(n5696) );
  XOR U6231 ( .A(n5695), .B(n5696), .Z(n5751) );
  XOR U6232 ( .A(n5752), .B(n5751), .Z(n5753) );
  XOR U6233 ( .A(n5754), .B(n5753), .Z(n5758) );
  XNOR U6234 ( .A(n5757), .B(n5758), .Z(n5759) );
  XNOR U6235 ( .A(n5760), .B(n5759), .Z(n5764) );
  NAND U6236 ( .A(n5605), .B(n5604), .Z(n5609) );
  NANDN U6237 ( .A(n5607), .B(n5606), .Z(n5608) );
  NAND U6238 ( .A(n5609), .B(n5608), .Z(n5761) );
  XNOR U6239 ( .A(n5761), .B(n5762), .Z(n5763) );
  XNOR U6240 ( .A(n5764), .B(n5763), .Z(n5638) );
  NANDN U6241 ( .A(n5615), .B(n5614), .Z(n5619) );
  NAND U6242 ( .A(n5617), .B(n5616), .Z(n5618) );
  NAND U6243 ( .A(n5619), .B(n5618), .Z(n5635) );
  NANDN U6244 ( .A(n5621), .B(n5620), .Z(n5625) );
  OR U6245 ( .A(n5623), .B(n5622), .Z(n5624) );
  NAND U6246 ( .A(n5625), .B(n5624), .Z(n5636) );
  XNOR U6247 ( .A(n5635), .B(n5636), .Z(n5637) );
  XNOR U6248 ( .A(n5638), .B(n5637), .Z(n5631) );
  XOR U6249 ( .A(n5632), .B(n5631), .Z(n5633) );
  XNOR U6250 ( .A(n5634), .B(n5633), .Z(n5767) );
  XNOR U6251 ( .A(n5767), .B(sreg[146]), .Z(n5769) );
  NAND U6252 ( .A(n5626), .B(sreg[145]), .Z(n5630) );
  OR U6253 ( .A(n5628), .B(n5627), .Z(n5629) );
  AND U6254 ( .A(n5630), .B(n5629), .Z(n5768) );
  XOR U6255 ( .A(n5769), .B(n5768), .Z(c[146]) );
  NANDN U6256 ( .A(n5636), .B(n5635), .Z(n5640) );
  NANDN U6257 ( .A(n5638), .B(n5637), .Z(n5639) );
  NAND U6258 ( .A(n5640), .B(n5639), .Z(n5773) );
  NANDN U6259 ( .A(n5642), .B(n5641), .Z(n5646) );
  NAND U6260 ( .A(n5644), .B(n5643), .Z(n5645) );
  NAND U6261 ( .A(n5646), .B(n5645), .Z(n5855) );
  NANDN U6262 ( .A(n5647), .B(n18832), .Z(n5649) );
  XNOR U6263 ( .A(b[19]), .B(a[33]), .Z(n5800) );
  NANDN U6264 ( .A(n5800), .B(n18834), .Z(n5648) );
  NAND U6265 ( .A(n5649), .B(n5648), .Z(n5865) );
  XNOR U6266 ( .A(b[27]), .B(a[25]), .Z(n5803) );
  NANDN U6267 ( .A(n5803), .B(n19336), .Z(n5652) );
  NANDN U6268 ( .A(n5650), .B(n19337), .Z(n5651) );
  NAND U6269 ( .A(n5652), .B(n5651), .Z(n5862) );
  XOR U6270 ( .A(b[5]), .B(a[47]), .Z(n5806) );
  NAND U6271 ( .A(n5806), .B(n17310), .Z(n5655) );
  NAND U6272 ( .A(n5653), .B(n17311), .Z(n5654) );
  AND U6273 ( .A(n5655), .B(n5654), .Z(n5863) );
  XNOR U6274 ( .A(n5862), .B(n5863), .Z(n5864) );
  XNOR U6275 ( .A(n5865), .B(n5864), .Z(n5853) );
  XOR U6276 ( .A(b[17]), .B(a[35]), .Z(n5809) );
  NAND U6277 ( .A(n5809), .B(n18673), .Z(n5658) );
  NAND U6278 ( .A(n5656), .B(n18674), .Z(n5657) );
  NAND U6279 ( .A(n5658), .B(n5657), .Z(n5827) );
  XNOR U6280 ( .A(b[31]), .B(a[21]), .Z(n5812) );
  NANDN U6281 ( .A(n5812), .B(n19472), .Z(n5661) );
  NANDN U6282 ( .A(n5659), .B(n19473), .Z(n5660) );
  NAND U6283 ( .A(n5661), .B(n5660), .Z(n5824) );
  OR U6284 ( .A(n5662), .B(n16988), .Z(n5664) );
  XOR U6285 ( .A(b[3]), .B(n10083), .Z(n5815) );
  NANDN U6286 ( .A(n5815), .B(n16990), .Z(n5663) );
  AND U6287 ( .A(n5664), .B(n5663), .Z(n5825) );
  XNOR U6288 ( .A(n5824), .B(n5825), .Z(n5826) );
  XOR U6289 ( .A(n5827), .B(n5826), .Z(n5852) );
  XNOR U6290 ( .A(n5853), .B(n5852), .Z(n5854) );
  XNOR U6291 ( .A(n5855), .B(n5854), .Z(n5791) );
  NANDN U6292 ( .A(n5666), .B(n5665), .Z(n5670) );
  NAND U6293 ( .A(n5668), .B(n5667), .Z(n5669) );
  NAND U6294 ( .A(n5670), .B(n5669), .Z(n5844) );
  NANDN U6295 ( .A(n5672), .B(n5671), .Z(n5676) );
  NAND U6296 ( .A(n5674), .B(n5673), .Z(n5675) );
  NAND U6297 ( .A(n5676), .B(n5675), .Z(n5843) );
  XNOR U6298 ( .A(n5843), .B(n5842), .Z(n5845) );
  XOR U6299 ( .A(n5844), .B(n5845), .Z(n5790) );
  XOR U6300 ( .A(n5791), .B(n5790), .Z(n5792) );
  NANDN U6301 ( .A(n5682), .B(n5681), .Z(n5686) );
  NAND U6302 ( .A(n5684), .B(n5683), .Z(n5685) );
  NAND U6303 ( .A(n5686), .B(n5685), .Z(n5793) );
  XNOR U6304 ( .A(n5792), .B(n5793), .Z(n5906) );
  OR U6305 ( .A(n5688), .B(n5687), .Z(n5692) );
  NAND U6306 ( .A(n5690), .B(n5689), .Z(n5691) );
  NAND U6307 ( .A(n5692), .B(n5691), .Z(n5905) );
  NANDN U6308 ( .A(n5694), .B(n5693), .Z(n5698) );
  NAND U6309 ( .A(n5696), .B(n5695), .Z(n5697) );
  NAND U6310 ( .A(n5698), .B(n5697), .Z(n5786) );
  NANDN U6311 ( .A(n5704), .B(n5703), .Z(n5708) );
  NAND U6312 ( .A(n5706), .B(n5705), .Z(n5707) );
  NAND U6313 ( .A(n5708), .B(n5707), .Z(n5846) );
  NANDN U6314 ( .A(n5710), .B(n5709), .Z(n5714) );
  NAND U6315 ( .A(n5712), .B(n5711), .Z(n5713) );
  AND U6316 ( .A(n5714), .B(n5713), .Z(n5847) );
  XNOR U6317 ( .A(n5846), .B(n5847), .Z(n5848) );
  XNOR U6318 ( .A(b[9]), .B(a[43]), .Z(n5868) );
  NANDN U6319 ( .A(n5868), .B(n17814), .Z(n5717) );
  NANDN U6320 ( .A(n5715), .B(n17815), .Z(n5716) );
  NAND U6321 ( .A(n5717), .B(n5716), .Z(n5832) );
  NANDN U6322 ( .A(n5718), .B(n18513), .Z(n5720) );
  XOR U6323 ( .A(b[15]), .B(a[37]), .Z(n5871) );
  NANDN U6324 ( .A(n18512), .B(n5871), .Z(n5719) );
  AND U6325 ( .A(n5720), .B(n5719), .Z(n5830) );
  NANDN U6326 ( .A(n5721), .B(n19013), .Z(n5723) );
  XNOR U6327 ( .A(b[21]), .B(a[31]), .Z(n5874) );
  NANDN U6328 ( .A(n5874), .B(n19015), .Z(n5722) );
  AND U6329 ( .A(n5723), .B(n5722), .Z(n5831) );
  XOR U6330 ( .A(n5832), .B(n5833), .Z(n5821) );
  XOR U6331 ( .A(b[11]), .B(n8930), .Z(n5877) );
  OR U6332 ( .A(n5877), .B(n18194), .Z(n5726) );
  NANDN U6333 ( .A(n5724), .B(n18104), .Z(n5725) );
  NAND U6334 ( .A(n5726), .B(n5725), .Z(n5819) );
  XOR U6335 ( .A(n580), .B(a[39]), .Z(n5880) );
  NANDN U6336 ( .A(n5880), .B(n18336), .Z(n5729) );
  NANDN U6337 ( .A(n5727), .B(n18337), .Z(n5728) );
  AND U6338 ( .A(n5729), .B(n5728), .Z(n5818) );
  XNOR U6339 ( .A(n5819), .B(n5818), .Z(n5820) );
  XOR U6340 ( .A(n5821), .B(n5820), .Z(n5838) );
  NANDN U6341 ( .A(n577), .B(a[51]), .Z(n5730) );
  XOR U6342 ( .A(n17151), .B(n5730), .Z(n5732) );
  NANDN U6343 ( .A(b[0]), .B(a[50]), .Z(n5731) );
  AND U6344 ( .A(n5732), .B(n5731), .Z(n5796) );
  NAND U6345 ( .A(n19406), .B(n5733), .Z(n5735) );
  XNOR U6346 ( .A(n584), .B(a[23]), .Z(n5883) );
  NANDN U6347 ( .A(n576), .B(n5883), .Z(n5734) );
  NAND U6348 ( .A(n5735), .B(n5734), .Z(n5794) );
  NANDN U6349 ( .A(n585), .B(a[19]), .Z(n5795) );
  XNOR U6350 ( .A(n5794), .B(n5795), .Z(n5797) );
  XOR U6351 ( .A(n5796), .B(n5797), .Z(n5836) );
  XNOR U6352 ( .A(b[23]), .B(a[29]), .Z(n5889) );
  OR U6353 ( .A(n5889), .B(n19127), .Z(n5738) );
  NAND U6354 ( .A(n5736), .B(n19128), .Z(n5737) );
  NAND U6355 ( .A(n5738), .B(n5737), .Z(n5859) );
  NAND U6356 ( .A(n5739), .B(n17553), .Z(n5741) );
  XOR U6357 ( .A(b[7]), .B(a[45]), .Z(n5892) );
  NAND U6358 ( .A(n5892), .B(n17555), .Z(n5740) );
  NAND U6359 ( .A(n5741), .B(n5740), .Z(n5856) );
  XOR U6360 ( .A(b[25]), .B(a[27]), .Z(n5895) );
  NAND U6361 ( .A(n5895), .B(n19240), .Z(n5744) );
  NAND U6362 ( .A(n5742), .B(n19242), .Z(n5743) );
  AND U6363 ( .A(n5744), .B(n5743), .Z(n5857) );
  XNOR U6364 ( .A(n5856), .B(n5857), .Z(n5858) );
  XNOR U6365 ( .A(n5859), .B(n5858), .Z(n5837) );
  XOR U6366 ( .A(n5836), .B(n5837), .Z(n5839) );
  XNOR U6367 ( .A(n5838), .B(n5839), .Z(n5849) );
  XNOR U6368 ( .A(n5848), .B(n5849), .Z(n5784) );
  XNOR U6369 ( .A(n5785), .B(n5784), .Z(n5787) );
  XNOR U6370 ( .A(n5786), .B(n5787), .Z(n5904) );
  XOR U6371 ( .A(n5905), .B(n5904), .Z(n5907) );
  NANDN U6372 ( .A(n5746), .B(n5745), .Z(n5750) );
  NAND U6373 ( .A(n5748), .B(n5747), .Z(n5749) );
  NAND U6374 ( .A(n5750), .B(n5749), .Z(n5898) );
  NAND U6375 ( .A(n5752), .B(n5751), .Z(n5756) );
  NAND U6376 ( .A(n5754), .B(n5753), .Z(n5755) );
  NAND U6377 ( .A(n5756), .B(n5755), .Z(n5899) );
  XNOR U6378 ( .A(n5898), .B(n5899), .Z(n5900) );
  XOR U6379 ( .A(n5901), .B(n5900), .Z(n5780) );
  NANDN U6380 ( .A(n5762), .B(n5761), .Z(n5766) );
  NANDN U6381 ( .A(n5764), .B(n5763), .Z(n5765) );
  NAND U6382 ( .A(n5766), .B(n5765), .Z(n5779) );
  XNOR U6383 ( .A(n5778), .B(n5779), .Z(n5781) );
  XOR U6384 ( .A(n5780), .B(n5781), .Z(n5772) );
  XOR U6385 ( .A(n5773), .B(n5772), .Z(n5774) );
  XNOR U6386 ( .A(n5775), .B(n5774), .Z(n5910) );
  XNOR U6387 ( .A(n5910), .B(sreg[147]), .Z(n5912) );
  NAND U6388 ( .A(n5767), .B(sreg[146]), .Z(n5771) );
  OR U6389 ( .A(n5769), .B(n5768), .Z(n5770) );
  AND U6390 ( .A(n5771), .B(n5770), .Z(n5911) );
  XOR U6391 ( .A(n5912), .B(n5911), .Z(c[147]) );
  NAND U6392 ( .A(n5773), .B(n5772), .Z(n5777) );
  NAND U6393 ( .A(n5775), .B(n5774), .Z(n5776) );
  NAND U6394 ( .A(n5777), .B(n5776), .Z(n5918) );
  NANDN U6395 ( .A(n5779), .B(n5778), .Z(n5783) );
  NAND U6396 ( .A(n5781), .B(n5780), .Z(n5782) );
  NAND U6397 ( .A(n5783), .B(n5782), .Z(n5915) );
  NAND U6398 ( .A(n5785), .B(n5784), .Z(n5789) );
  NANDN U6399 ( .A(n5787), .B(n5786), .Z(n5788) );
  NAND U6400 ( .A(n5789), .B(n5788), .Z(n5927) );
  XNOR U6401 ( .A(n5927), .B(n5928), .Z(n5929) );
  NANDN U6402 ( .A(n5795), .B(n5794), .Z(n5799) );
  NAND U6403 ( .A(n5797), .B(n5796), .Z(n5798) );
  NAND U6404 ( .A(n5799), .B(n5798), .Z(n6002) );
  NANDN U6405 ( .A(n5800), .B(n18832), .Z(n5802) );
  XNOR U6406 ( .A(b[19]), .B(a[34]), .Z(n5969) );
  NANDN U6407 ( .A(n5969), .B(n18834), .Z(n5801) );
  NAND U6408 ( .A(n5802), .B(n5801), .Z(n6014) );
  XNOR U6409 ( .A(b[27]), .B(a[26]), .Z(n5972) );
  NANDN U6410 ( .A(n5972), .B(n19336), .Z(n5805) );
  NANDN U6411 ( .A(n5803), .B(n19337), .Z(n5804) );
  NAND U6412 ( .A(n5805), .B(n5804), .Z(n6011) );
  XOR U6413 ( .A(b[5]), .B(a[48]), .Z(n5975) );
  NAND U6414 ( .A(n5975), .B(n17310), .Z(n5808) );
  NAND U6415 ( .A(n5806), .B(n17311), .Z(n5807) );
  AND U6416 ( .A(n5808), .B(n5807), .Z(n6012) );
  XNOR U6417 ( .A(n6011), .B(n6012), .Z(n6013) );
  XNOR U6418 ( .A(n6014), .B(n6013), .Z(n5999) );
  XOR U6419 ( .A(b[17]), .B(a[36]), .Z(n5978) );
  NAND U6420 ( .A(n5978), .B(n18673), .Z(n5811) );
  NAND U6421 ( .A(n5809), .B(n18674), .Z(n5810) );
  NAND U6422 ( .A(n5811), .B(n5810), .Z(n5953) );
  XNOR U6423 ( .A(b[31]), .B(a[22]), .Z(n5981) );
  NANDN U6424 ( .A(n5981), .B(n19472), .Z(n5814) );
  NANDN U6425 ( .A(n5812), .B(n19473), .Z(n5813) );
  AND U6426 ( .A(n5814), .B(n5813), .Z(n5951) );
  OR U6427 ( .A(n5815), .B(n16988), .Z(n5817) );
  XNOR U6428 ( .A(b[3]), .B(a[50]), .Z(n5984) );
  NANDN U6429 ( .A(n5984), .B(n16990), .Z(n5816) );
  AND U6430 ( .A(n5817), .B(n5816), .Z(n5952) );
  XOR U6431 ( .A(n5953), .B(n5954), .Z(n6000) );
  XOR U6432 ( .A(n5999), .B(n6000), .Z(n6001) );
  XNOR U6433 ( .A(n6002), .B(n6001), .Z(n6047) );
  NANDN U6434 ( .A(n5819), .B(n5818), .Z(n5823) );
  NAND U6435 ( .A(n5821), .B(n5820), .Z(n5822) );
  NAND U6436 ( .A(n5823), .B(n5822), .Z(n5990) );
  NANDN U6437 ( .A(n5825), .B(n5824), .Z(n5829) );
  NAND U6438 ( .A(n5827), .B(n5826), .Z(n5828) );
  NAND U6439 ( .A(n5829), .B(n5828), .Z(n5988) );
  OR U6440 ( .A(n5831), .B(n5830), .Z(n5835) );
  NANDN U6441 ( .A(n5833), .B(n5832), .Z(n5834) );
  NAND U6442 ( .A(n5835), .B(n5834), .Z(n5987) );
  XNOR U6443 ( .A(n5990), .B(n5989), .Z(n6048) );
  XNOR U6444 ( .A(n6047), .B(n6048), .Z(n6049) );
  NANDN U6445 ( .A(n5837), .B(n5836), .Z(n5841) );
  OR U6446 ( .A(n5839), .B(n5838), .Z(n5840) );
  AND U6447 ( .A(n5841), .B(n5840), .Z(n6050) );
  XOR U6448 ( .A(n6049), .B(n6050), .Z(n5935) );
  NANDN U6449 ( .A(n5847), .B(n5846), .Z(n5851) );
  NANDN U6450 ( .A(n5849), .B(n5848), .Z(n5850) );
  NAND U6451 ( .A(n5851), .B(n5850), .Z(n6056) );
  NANDN U6452 ( .A(n5857), .B(n5856), .Z(n5861) );
  NAND U6453 ( .A(n5859), .B(n5858), .Z(n5860) );
  NAND U6454 ( .A(n5861), .B(n5860), .Z(n5993) );
  NANDN U6455 ( .A(n5863), .B(n5862), .Z(n5867) );
  NAND U6456 ( .A(n5865), .B(n5864), .Z(n5866) );
  AND U6457 ( .A(n5867), .B(n5866), .Z(n5994) );
  XNOR U6458 ( .A(n5993), .B(n5994), .Z(n5995) );
  XNOR U6459 ( .A(b[9]), .B(a[44]), .Z(n6017) );
  NANDN U6460 ( .A(n6017), .B(n17814), .Z(n5870) );
  NANDN U6461 ( .A(n5868), .B(n17815), .Z(n5869) );
  NAND U6462 ( .A(n5870), .B(n5869), .Z(n5959) );
  NAND U6463 ( .A(n5871), .B(n18513), .Z(n5873) );
  XNOR U6464 ( .A(b[15]), .B(a[38]), .Z(n6020) );
  OR U6465 ( .A(n6020), .B(n18512), .Z(n5872) );
  AND U6466 ( .A(n5873), .B(n5872), .Z(n5957) );
  NANDN U6467 ( .A(n5874), .B(n19013), .Z(n5876) );
  XNOR U6468 ( .A(b[21]), .B(a[32]), .Z(n6023) );
  NANDN U6469 ( .A(n6023), .B(n19015), .Z(n5875) );
  AND U6470 ( .A(n5876), .B(n5875), .Z(n5958) );
  XOR U6471 ( .A(n5959), .B(n5960), .Z(n5948) );
  XOR U6472 ( .A(b[11]), .B(n9080), .Z(n6026) );
  OR U6473 ( .A(n6026), .B(n18194), .Z(n5879) );
  NANDN U6474 ( .A(n5877), .B(n18104), .Z(n5878) );
  NAND U6475 ( .A(n5879), .B(n5878), .Z(n5946) );
  XOR U6476 ( .A(n580), .B(a[40]), .Z(n6029) );
  NANDN U6477 ( .A(n6029), .B(n18336), .Z(n5882) );
  NANDN U6478 ( .A(n5880), .B(n18337), .Z(n5881) );
  NAND U6479 ( .A(n5882), .B(n5881), .Z(n5945) );
  XOR U6480 ( .A(n5948), .B(n5947), .Z(n5942) );
  NAND U6481 ( .A(n19406), .B(n5883), .Z(n5885) );
  XNOR U6482 ( .A(n584), .B(a[24]), .Z(n6035) );
  NANDN U6483 ( .A(n576), .B(n6035), .Z(n5884) );
  NAND U6484 ( .A(n5885), .B(n5884), .Z(n5963) );
  NANDN U6485 ( .A(n585), .B(a[20]), .Z(n5964) );
  XNOR U6486 ( .A(n5963), .B(n5964), .Z(n5966) );
  NANDN U6487 ( .A(n577), .B(a[52]), .Z(n5886) );
  XOR U6488 ( .A(n17151), .B(n5886), .Z(n5888) );
  NANDN U6489 ( .A(b[0]), .B(a[51]), .Z(n5887) );
  AND U6490 ( .A(n5888), .B(n5887), .Z(n5965) );
  XNOR U6491 ( .A(n5966), .B(n5965), .Z(n5940) );
  XNOR U6492 ( .A(b[23]), .B(a[30]), .Z(n6038) );
  OR U6493 ( .A(n6038), .B(n19127), .Z(n5891) );
  NANDN U6494 ( .A(n5889), .B(n19128), .Z(n5890) );
  NAND U6495 ( .A(n5891), .B(n5890), .Z(n6008) );
  NAND U6496 ( .A(n5892), .B(n17553), .Z(n5894) );
  XOR U6497 ( .A(b[7]), .B(a[46]), .Z(n6041) );
  NAND U6498 ( .A(n6041), .B(n17555), .Z(n5893) );
  NAND U6499 ( .A(n5894), .B(n5893), .Z(n6005) );
  XOR U6500 ( .A(b[25]), .B(a[28]), .Z(n6044) );
  NAND U6501 ( .A(n6044), .B(n19240), .Z(n5897) );
  NAND U6502 ( .A(n5895), .B(n19242), .Z(n5896) );
  AND U6503 ( .A(n5897), .B(n5896), .Z(n6006) );
  XNOR U6504 ( .A(n6005), .B(n6006), .Z(n6007) );
  XOR U6505 ( .A(n6008), .B(n6007), .Z(n5939) );
  XOR U6506 ( .A(n5942), .B(n5941), .Z(n5996) );
  XNOR U6507 ( .A(n5995), .B(n5996), .Z(n6053) );
  XOR U6508 ( .A(n6054), .B(n6053), .Z(n6055) );
  XNOR U6509 ( .A(n6056), .B(n6055), .Z(n5933) );
  XNOR U6510 ( .A(n5934), .B(n5933), .Z(n5936) );
  XNOR U6511 ( .A(n5935), .B(n5936), .Z(n5930) );
  XOR U6512 ( .A(n5929), .B(n5930), .Z(n5924) );
  NANDN U6513 ( .A(n5899), .B(n5898), .Z(n5903) );
  NAND U6514 ( .A(n5901), .B(n5900), .Z(n5902) );
  NAND U6515 ( .A(n5903), .B(n5902), .Z(n5921) );
  NANDN U6516 ( .A(n5905), .B(n5904), .Z(n5909) );
  OR U6517 ( .A(n5907), .B(n5906), .Z(n5908) );
  NAND U6518 ( .A(n5909), .B(n5908), .Z(n5922) );
  XNOR U6519 ( .A(n5921), .B(n5922), .Z(n5923) );
  XNOR U6520 ( .A(n5924), .B(n5923), .Z(n5916) );
  XNOR U6521 ( .A(n5915), .B(n5916), .Z(n5917) );
  XNOR U6522 ( .A(n5918), .B(n5917), .Z(n6059) );
  XNOR U6523 ( .A(n6059), .B(sreg[148]), .Z(n6061) );
  NAND U6524 ( .A(n5910), .B(sreg[147]), .Z(n5914) );
  OR U6525 ( .A(n5912), .B(n5911), .Z(n5913) );
  AND U6526 ( .A(n5914), .B(n5913), .Z(n6060) );
  XOR U6527 ( .A(n6061), .B(n6060), .Z(c[148]) );
  NANDN U6528 ( .A(n5916), .B(n5915), .Z(n5920) );
  NAND U6529 ( .A(n5918), .B(n5917), .Z(n5919) );
  NAND U6530 ( .A(n5920), .B(n5919), .Z(n6067) );
  NANDN U6531 ( .A(n5922), .B(n5921), .Z(n5926) );
  NAND U6532 ( .A(n5924), .B(n5923), .Z(n5925) );
  NAND U6533 ( .A(n5926), .B(n5925), .Z(n6065) );
  NANDN U6534 ( .A(n5928), .B(n5927), .Z(n5932) );
  NANDN U6535 ( .A(n5930), .B(n5929), .Z(n5931) );
  NAND U6536 ( .A(n5932), .B(n5931), .Z(n6071) );
  OR U6537 ( .A(n5934), .B(n5933), .Z(n5938) );
  OR U6538 ( .A(n5936), .B(n5935), .Z(n5937) );
  AND U6539 ( .A(n5938), .B(n5937), .Z(n6070) );
  XNOR U6540 ( .A(n6071), .B(n6070), .Z(n6072) );
  NANDN U6541 ( .A(n5940), .B(n5939), .Z(n5944) );
  NANDN U6542 ( .A(n5942), .B(n5941), .Z(n5943) );
  NAND U6543 ( .A(n5944), .B(n5943), .Z(n6199) );
  OR U6544 ( .A(n5946), .B(n5945), .Z(n5950) );
  NAND U6545 ( .A(n5948), .B(n5947), .Z(n5949) );
  NAND U6546 ( .A(n5950), .B(n5949), .Z(n6138) );
  OR U6547 ( .A(n5952), .B(n5951), .Z(n5956) );
  NANDN U6548 ( .A(n5954), .B(n5953), .Z(n5955) );
  NAND U6549 ( .A(n5956), .B(n5955), .Z(n6137) );
  OR U6550 ( .A(n5958), .B(n5957), .Z(n5962) );
  NANDN U6551 ( .A(n5960), .B(n5959), .Z(n5961) );
  NAND U6552 ( .A(n5962), .B(n5961), .Z(n6136) );
  XOR U6553 ( .A(n6138), .B(n6139), .Z(n6196) );
  NANDN U6554 ( .A(n5964), .B(n5963), .Z(n5968) );
  NAND U6555 ( .A(n5966), .B(n5965), .Z(n5967) );
  NAND U6556 ( .A(n5968), .B(n5967), .Z(n6151) );
  NANDN U6557 ( .A(n5969), .B(n18832), .Z(n5971) );
  XNOR U6558 ( .A(b[19]), .B(a[35]), .Z(n6094) );
  NANDN U6559 ( .A(n6094), .B(n18834), .Z(n5970) );
  NAND U6560 ( .A(n5971), .B(n5970), .Z(n6163) );
  XNOR U6561 ( .A(b[27]), .B(a[27]), .Z(n6097) );
  NANDN U6562 ( .A(n6097), .B(n19336), .Z(n5974) );
  NANDN U6563 ( .A(n5972), .B(n19337), .Z(n5973) );
  NAND U6564 ( .A(n5974), .B(n5973), .Z(n6160) );
  XNOR U6565 ( .A(b[5]), .B(a[49]), .Z(n6100) );
  NANDN U6566 ( .A(n6100), .B(n17310), .Z(n5977) );
  NAND U6567 ( .A(n5975), .B(n17311), .Z(n5976) );
  AND U6568 ( .A(n5977), .B(n5976), .Z(n6161) );
  XNOR U6569 ( .A(n6160), .B(n6161), .Z(n6162) );
  XNOR U6570 ( .A(n6163), .B(n6162), .Z(n6149) );
  XOR U6571 ( .A(b[17]), .B(a[37]), .Z(n6103) );
  NAND U6572 ( .A(n6103), .B(n18673), .Z(n5980) );
  NAND U6573 ( .A(n5978), .B(n18674), .Z(n5979) );
  NAND U6574 ( .A(n5980), .B(n5979), .Z(n6121) );
  XNOR U6575 ( .A(b[31]), .B(a[23]), .Z(n6106) );
  NANDN U6576 ( .A(n6106), .B(n19472), .Z(n5983) );
  NANDN U6577 ( .A(n5981), .B(n19473), .Z(n5982) );
  NAND U6578 ( .A(n5983), .B(n5982), .Z(n6118) );
  OR U6579 ( .A(n5984), .B(n16988), .Z(n5986) );
  XNOR U6580 ( .A(b[3]), .B(a[51]), .Z(n6109) );
  NANDN U6581 ( .A(n6109), .B(n16990), .Z(n5985) );
  AND U6582 ( .A(n5986), .B(n5985), .Z(n6119) );
  XNOR U6583 ( .A(n6118), .B(n6119), .Z(n6120) );
  XOR U6584 ( .A(n6121), .B(n6120), .Z(n6148) );
  XNOR U6585 ( .A(n6149), .B(n6148), .Z(n6150) );
  XNOR U6586 ( .A(n6151), .B(n6150), .Z(n6197) );
  XNOR U6587 ( .A(n6196), .B(n6197), .Z(n6198) );
  XNOR U6588 ( .A(n6199), .B(n6198), .Z(n6085) );
  OR U6589 ( .A(n5988), .B(n5987), .Z(n5992) );
  NAND U6590 ( .A(n5990), .B(n5989), .Z(n5991) );
  NAND U6591 ( .A(n5992), .B(n5991), .Z(n6083) );
  NANDN U6592 ( .A(n5994), .B(n5993), .Z(n5998) );
  NANDN U6593 ( .A(n5996), .B(n5995), .Z(n5997) );
  NAND U6594 ( .A(n5998), .B(n5997), .Z(n6204) );
  OR U6595 ( .A(n6000), .B(n5999), .Z(n6004) );
  NAND U6596 ( .A(n6002), .B(n6001), .Z(n6003) );
  NAND U6597 ( .A(n6004), .B(n6003), .Z(n6203) );
  NANDN U6598 ( .A(n6006), .B(n6005), .Z(n6010) );
  NAND U6599 ( .A(n6008), .B(n6007), .Z(n6009) );
  NAND U6600 ( .A(n6010), .B(n6009), .Z(n6142) );
  NANDN U6601 ( .A(n6012), .B(n6011), .Z(n6016) );
  NAND U6602 ( .A(n6014), .B(n6013), .Z(n6015) );
  AND U6603 ( .A(n6016), .B(n6015), .Z(n6143) );
  XNOR U6604 ( .A(n6142), .B(n6143), .Z(n6144) );
  XNOR U6605 ( .A(b[9]), .B(a[45]), .Z(n6166) );
  NANDN U6606 ( .A(n6166), .B(n17814), .Z(n6019) );
  NANDN U6607 ( .A(n6017), .B(n17815), .Z(n6018) );
  NAND U6608 ( .A(n6019), .B(n6018), .Z(n6126) );
  NANDN U6609 ( .A(n6020), .B(n18513), .Z(n6022) );
  XOR U6610 ( .A(b[15]), .B(a[39]), .Z(n6169) );
  NANDN U6611 ( .A(n18512), .B(n6169), .Z(n6021) );
  AND U6612 ( .A(n6022), .B(n6021), .Z(n6124) );
  NANDN U6613 ( .A(n6023), .B(n19013), .Z(n6025) );
  XNOR U6614 ( .A(b[21]), .B(a[33]), .Z(n6172) );
  NANDN U6615 ( .A(n6172), .B(n19015), .Z(n6024) );
  AND U6616 ( .A(n6025), .B(n6024), .Z(n6125) );
  XOR U6617 ( .A(n6126), .B(n6127), .Z(n6115) );
  XNOR U6618 ( .A(b[11]), .B(a[43]), .Z(n6175) );
  OR U6619 ( .A(n6175), .B(n18194), .Z(n6028) );
  NANDN U6620 ( .A(n6026), .B(n18104), .Z(n6027) );
  NAND U6621 ( .A(n6028), .B(n6027), .Z(n6113) );
  XOR U6622 ( .A(n580), .B(a[41]), .Z(n6178) );
  NANDN U6623 ( .A(n6178), .B(n18336), .Z(n6031) );
  NANDN U6624 ( .A(n6029), .B(n18337), .Z(n6030) );
  AND U6625 ( .A(n6031), .B(n6030), .Z(n6112) );
  XNOR U6626 ( .A(n6113), .B(n6112), .Z(n6114) );
  XOR U6627 ( .A(n6115), .B(n6114), .Z(n6132) );
  NANDN U6628 ( .A(n577), .B(a[53]), .Z(n6032) );
  XOR U6629 ( .A(n17151), .B(n6032), .Z(n6034) );
  NANDN U6630 ( .A(b[0]), .B(a[52]), .Z(n6033) );
  AND U6631 ( .A(n6034), .B(n6033), .Z(n6090) );
  NAND U6632 ( .A(n19406), .B(n6035), .Z(n6037) );
  XNOR U6633 ( .A(n584), .B(a[25]), .Z(n6181) );
  NANDN U6634 ( .A(n576), .B(n6181), .Z(n6036) );
  NAND U6635 ( .A(n6037), .B(n6036), .Z(n6088) );
  NANDN U6636 ( .A(n585), .B(a[21]), .Z(n6089) );
  XNOR U6637 ( .A(n6088), .B(n6089), .Z(n6091) );
  XOR U6638 ( .A(n6090), .B(n6091), .Z(n6130) );
  XOR U6639 ( .A(b[23]), .B(a[31]), .Z(n6187) );
  NANDN U6640 ( .A(n19127), .B(n6187), .Z(n6040) );
  NANDN U6641 ( .A(n6038), .B(n19128), .Z(n6039) );
  NAND U6642 ( .A(n6040), .B(n6039), .Z(n6157) );
  NAND U6643 ( .A(n6041), .B(n17553), .Z(n6043) );
  XOR U6644 ( .A(b[7]), .B(a[47]), .Z(n6190) );
  NAND U6645 ( .A(n6190), .B(n17555), .Z(n6042) );
  NAND U6646 ( .A(n6043), .B(n6042), .Z(n6154) );
  XNOR U6647 ( .A(b[25]), .B(a[29]), .Z(n6193) );
  NANDN U6648 ( .A(n6193), .B(n19240), .Z(n6046) );
  NAND U6649 ( .A(n6044), .B(n19242), .Z(n6045) );
  AND U6650 ( .A(n6046), .B(n6045), .Z(n6155) );
  XNOR U6651 ( .A(n6154), .B(n6155), .Z(n6156) );
  XNOR U6652 ( .A(n6157), .B(n6156), .Z(n6131) );
  XOR U6653 ( .A(n6130), .B(n6131), .Z(n6133) );
  XNOR U6654 ( .A(n6132), .B(n6133), .Z(n6145) );
  XNOR U6655 ( .A(n6144), .B(n6145), .Z(n6202) );
  XNOR U6656 ( .A(n6203), .B(n6202), .Z(n6205) );
  XNOR U6657 ( .A(n6204), .B(n6205), .Z(n6082) );
  XNOR U6658 ( .A(n6083), .B(n6082), .Z(n6084) );
  XOR U6659 ( .A(n6085), .B(n6084), .Z(n6079) );
  NANDN U6660 ( .A(n6048), .B(n6047), .Z(n6052) );
  NAND U6661 ( .A(n6050), .B(n6049), .Z(n6051) );
  NAND U6662 ( .A(n6052), .B(n6051), .Z(n6076) );
  NAND U6663 ( .A(n6054), .B(n6053), .Z(n6058) );
  NAND U6664 ( .A(n6056), .B(n6055), .Z(n6057) );
  NAND U6665 ( .A(n6058), .B(n6057), .Z(n6077) );
  XNOR U6666 ( .A(n6076), .B(n6077), .Z(n6078) );
  XOR U6667 ( .A(n6079), .B(n6078), .Z(n6073) );
  XOR U6668 ( .A(n6072), .B(n6073), .Z(n6064) );
  XOR U6669 ( .A(n6065), .B(n6064), .Z(n6066) );
  XNOR U6670 ( .A(n6067), .B(n6066), .Z(n6208) );
  XNOR U6671 ( .A(n6208), .B(sreg[149]), .Z(n6210) );
  NAND U6672 ( .A(n6059), .B(sreg[148]), .Z(n6063) );
  OR U6673 ( .A(n6061), .B(n6060), .Z(n6062) );
  AND U6674 ( .A(n6063), .B(n6062), .Z(n6209) );
  XOR U6675 ( .A(n6210), .B(n6209), .Z(c[149]) );
  NAND U6676 ( .A(n6065), .B(n6064), .Z(n6069) );
  NAND U6677 ( .A(n6067), .B(n6066), .Z(n6068) );
  NAND U6678 ( .A(n6069), .B(n6068), .Z(n6216) );
  NANDN U6679 ( .A(n6071), .B(n6070), .Z(n6075) );
  NAND U6680 ( .A(n6073), .B(n6072), .Z(n6074) );
  NAND U6681 ( .A(n6075), .B(n6074), .Z(n6214) );
  NANDN U6682 ( .A(n6077), .B(n6076), .Z(n6081) );
  NAND U6683 ( .A(n6079), .B(n6078), .Z(n6080) );
  NAND U6684 ( .A(n6081), .B(n6080), .Z(n6219) );
  NANDN U6685 ( .A(n6083), .B(n6082), .Z(n6087) );
  NANDN U6686 ( .A(n6085), .B(n6084), .Z(n6086) );
  NAND U6687 ( .A(n6087), .B(n6086), .Z(n6220) );
  XNOR U6688 ( .A(n6219), .B(n6220), .Z(n6221) );
  NANDN U6689 ( .A(n6089), .B(n6088), .Z(n6093) );
  NAND U6690 ( .A(n6091), .B(n6090), .Z(n6092) );
  NAND U6691 ( .A(n6093), .B(n6092), .Z(n6288) );
  NANDN U6692 ( .A(n6094), .B(n18832), .Z(n6096) );
  XNOR U6693 ( .A(b[19]), .B(a[36]), .Z(n6255) );
  NANDN U6694 ( .A(n6255), .B(n18834), .Z(n6095) );
  NAND U6695 ( .A(n6096), .B(n6095), .Z(n6300) );
  XNOR U6696 ( .A(b[27]), .B(a[28]), .Z(n6258) );
  NANDN U6697 ( .A(n6258), .B(n19336), .Z(n6099) );
  NANDN U6698 ( .A(n6097), .B(n19337), .Z(n6098) );
  NAND U6699 ( .A(n6099), .B(n6098), .Z(n6297) );
  XOR U6700 ( .A(b[5]), .B(a[50]), .Z(n6261) );
  NAND U6701 ( .A(n6261), .B(n17310), .Z(n6102) );
  NANDN U6702 ( .A(n6100), .B(n17311), .Z(n6101) );
  AND U6703 ( .A(n6102), .B(n6101), .Z(n6298) );
  XNOR U6704 ( .A(n6297), .B(n6298), .Z(n6299) );
  XNOR U6705 ( .A(n6300), .B(n6299), .Z(n6285) );
  XNOR U6706 ( .A(b[17]), .B(a[38]), .Z(n6264) );
  NANDN U6707 ( .A(n6264), .B(n18673), .Z(n6105) );
  NAND U6708 ( .A(n6103), .B(n18674), .Z(n6104) );
  NAND U6709 ( .A(n6105), .B(n6104), .Z(n6239) );
  XNOR U6710 ( .A(b[31]), .B(a[24]), .Z(n6267) );
  NANDN U6711 ( .A(n6267), .B(n19472), .Z(n6108) );
  NANDN U6712 ( .A(n6106), .B(n19473), .Z(n6107) );
  AND U6713 ( .A(n6108), .B(n6107), .Z(n6237) );
  OR U6714 ( .A(n6109), .B(n16988), .Z(n6111) );
  XNOR U6715 ( .A(b[3]), .B(a[52]), .Z(n6270) );
  NANDN U6716 ( .A(n6270), .B(n16990), .Z(n6110) );
  AND U6717 ( .A(n6111), .B(n6110), .Z(n6238) );
  XOR U6718 ( .A(n6239), .B(n6240), .Z(n6286) );
  XOR U6719 ( .A(n6285), .B(n6286), .Z(n6287) );
  XNOR U6720 ( .A(n6288), .B(n6287), .Z(n6333) );
  NANDN U6721 ( .A(n6113), .B(n6112), .Z(n6117) );
  NAND U6722 ( .A(n6115), .B(n6114), .Z(n6116) );
  NAND U6723 ( .A(n6117), .B(n6116), .Z(n6276) );
  NANDN U6724 ( .A(n6119), .B(n6118), .Z(n6123) );
  NAND U6725 ( .A(n6121), .B(n6120), .Z(n6122) );
  NAND U6726 ( .A(n6123), .B(n6122), .Z(n6274) );
  OR U6727 ( .A(n6125), .B(n6124), .Z(n6129) );
  NANDN U6728 ( .A(n6127), .B(n6126), .Z(n6128) );
  NAND U6729 ( .A(n6129), .B(n6128), .Z(n6273) );
  XNOR U6730 ( .A(n6276), .B(n6275), .Z(n6334) );
  XOR U6731 ( .A(n6333), .B(n6334), .Z(n6336) );
  NANDN U6732 ( .A(n6131), .B(n6130), .Z(n6135) );
  OR U6733 ( .A(n6133), .B(n6132), .Z(n6134) );
  NAND U6734 ( .A(n6135), .B(n6134), .Z(n6335) );
  XOR U6735 ( .A(n6336), .B(n6335), .Z(n6353) );
  OR U6736 ( .A(n6137), .B(n6136), .Z(n6141) );
  NANDN U6737 ( .A(n6139), .B(n6138), .Z(n6140) );
  NAND U6738 ( .A(n6141), .B(n6140), .Z(n6352) );
  NANDN U6739 ( .A(n6143), .B(n6142), .Z(n6147) );
  NANDN U6740 ( .A(n6145), .B(n6144), .Z(n6146) );
  NAND U6741 ( .A(n6147), .B(n6146), .Z(n6341) );
  NANDN U6742 ( .A(n6149), .B(n6148), .Z(n6153) );
  NAND U6743 ( .A(n6151), .B(n6150), .Z(n6152) );
  NAND U6744 ( .A(n6153), .B(n6152), .Z(n6340) );
  NANDN U6745 ( .A(n6155), .B(n6154), .Z(n6159) );
  NAND U6746 ( .A(n6157), .B(n6156), .Z(n6158) );
  NAND U6747 ( .A(n6159), .B(n6158), .Z(n6279) );
  NANDN U6748 ( .A(n6161), .B(n6160), .Z(n6165) );
  NAND U6749 ( .A(n6163), .B(n6162), .Z(n6164) );
  AND U6750 ( .A(n6165), .B(n6164), .Z(n6280) );
  XNOR U6751 ( .A(n6279), .B(n6280), .Z(n6281) );
  XNOR U6752 ( .A(b[9]), .B(a[46]), .Z(n6303) );
  NANDN U6753 ( .A(n6303), .B(n17814), .Z(n6168) );
  NANDN U6754 ( .A(n6166), .B(n17815), .Z(n6167) );
  NAND U6755 ( .A(n6168), .B(n6167), .Z(n6245) );
  NAND U6756 ( .A(n6169), .B(n18513), .Z(n6171) );
  XOR U6757 ( .A(b[15]), .B(a[40]), .Z(n6306) );
  NANDN U6758 ( .A(n18512), .B(n6306), .Z(n6170) );
  AND U6759 ( .A(n6171), .B(n6170), .Z(n6243) );
  NANDN U6760 ( .A(n6172), .B(n19013), .Z(n6174) );
  XNOR U6761 ( .A(b[21]), .B(a[34]), .Z(n6309) );
  NANDN U6762 ( .A(n6309), .B(n19015), .Z(n6173) );
  AND U6763 ( .A(n6174), .B(n6173), .Z(n6244) );
  XOR U6764 ( .A(n6245), .B(n6246), .Z(n6234) );
  XNOR U6765 ( .A(b[11]), .B(a[44]), .Z(n6312) );
  OR U6766 ( .A(n6312), .B(n18194), .Z(n6177) );
  NANDN U6767 ( .A(n6175), .B(n18104), .Z(n6176) );
  NAND U6768 ( .A(n6177), .B(n6176), .Z(n6232) );
  XOR U6769 ( .A(n580), .B(a[42]), .Z(n6315) );
  NANDN U6770 ( .A(n6315), .B(n18336), .Z(n6180) );
  NANDN U6771 ( .A(n6178), .B(n18337), .Z(n6179) );
  NAND U6772 ( .A(n6180), .B(n6179), .Z(n6231) );
  XOR U6773 ( .A(n6234), .B(n6233), .Z(n6228) );
  NAND U6774 ( .A(n19406), .B(n6181), .Z(n6183) );
  XNOR U6775 ( .A(n584), .B(a[26]), .Z(n6321) );
  NANDN U6776 ( .A(n576), .B(n6321), .Z(n6182) );
  NAND U6777 ( .A(n6183), .B(n6182), .Z(n6249) );
  NANDN U6778 ( .A(n585), .B(a[22]), .Z(n6250) );
  XNOR U6779 ( .A(n6249), .B(n6250), .Z(n6252) );
  NANDN U6780 ( .A(n577), .B(a[54]), .Z(n6184) );
  XOR U6781 ( .A(n17151), .B(n6184), .Z(n6186) );
  IV U6782 ( .A(a[53]), .Z(n10660) );
  NANDN U6783 ( .A(n10660), .B(n577), .Z(n6185) );
  AND U6784 ( .A(n6186), .B(n6185), .Z(n6251) );
  XNOR U6785 ( .A(n6252), .B(n6251), .Z(n6226) );
  XOR U6786 ( .A(b[23]), .B(a[32]), .Z(n6324) );
  NANDN U6787 ( .A(n19127), .B(n6324), .Z(n6189) );
  NAND U6788 ( .A(n6187), .B(n19128), .Z(n6188) );
  NAND U6789 ( .A(n6189), .B(n6188), .Z(n6294) );
  NAND U6790 ( .A(n6190), .B(n17553), .Z(n6192) );
  XOR U6791 ( .A(b[7]), .B(a[48]), .Z(n6327) );
  NAND U6792 ( .A(n6327), .B(n17555), .Z(n6191) );
  NAND U6793 ( .A(n6192), .B(n6191), .Z(n6291) );
  XNOR U6794 ( .A(b[25]), .B(a[30]), .Z(n6330) );
  NANDN U6795 ( .A(n6330), .B(n19240), .Z(n6195) );
  NANDN U6796 ( .A(n6193), .B(n19242), .Z(n6194) );
  AND U6797 ( .A(n6195), .B(n6194), .Z(n6292) );
  XNOR U6798 ( .A(n6291), .B(n6292), .Z(n6293) );
  XOR U6799 ( .A(n6294), .B(n6293), .Z(n6225) );
  XOR U6800 ( .A(n6228), .B(n6227), .Z(n6282) );
  XNOR U6801 ( .A(n6281), .B(n6282), .Z(n6339) );
  XNOR U6802 ( .A(n6340), .B(n6339), .Z(n6342) );
  XNOR U6803 ( .A(n6341), .B(n6342), .Z(n6351) );
  XOR U6804 ( .A(n6352), .B(n6351), .Z(n6354) );
  NANDN U6805 ( .A(n6197), .B(n6196), .Z(n6201) );
  NAND U6806 ( .A(n6199), .B(n6198), .Z(n6200) );
  NAND U6807 ( .A(n6201), .B(n6200), .Z(n6346) );
  NAND U6808 ( .A(n6203), .B(n6202), .Z(n6207) );
  NANDN U6809 ( .A(n6205), .B(n6204), .Z(n6206) );
  AND U6810 ( .A(n6207), .B(n6206), .Z(n6345) );
  XNOR U6811 ( .A(n6346), .B(n6345), .Z(n6347) );
  XOR U6812 ( .A(n6348), .B(n6347), .Z(n6222) );
  XOR U6813 ( .A(n6221), .B(n6222), .Z(n6213) );
  XOR U6814 ( .A(n6214), .B(n6213), .Z(n6215) );
  XNOR U6815 ( .A(n6216), .B(n6215), .Z(n6357) );
  XNOR U6816 ( .A(n6357), .B(sreg[150]), .Z(n6359) );
  NAND U6817 ( .A(n6208), .B(sreg[149]), .Z(n6212) );
  OR U6818 ( .A(n6210), .B(n6209), .Z(n6211) );
  AND U6819 ( .A(n6212), .B(n6211), .Z(n6358) );
  XOR U6820 ( .A(n6359), .B(n6358), .Z(c[150]) );
  NAND U6821 ( .A(n6214), .B(n6213), .Z(n6218) );
  NAND U6822 ( .A(n6216), .B(n6215), .Z(n6217) );
  NAND U6823 ( .A(n6218), .B(n6217), .Z(n6365) );
  NANDN U6824 ( .A(n6220), .B(n6219), .Z(n6224) );
  NAND U6825 ( .A(n6222), .B(n6221), .Z(n6223) );
  NAND U6826 ( .A(n6224), .B(n6223), .Z(n6363) );
  NANDN U6827 ( .A(n6226), .B(n6225), .Z(n6230) );
  NANDN U6828 ( .A(n6228), .B(n6227), .Z(n6229) );
  NAND U6829 ( .A(n6230), .B(n6229), .Z(n6483) );
  OR U6830 ( .A(n6232), .B(n6231), .Z(n6236) );
  NAND U6831 ( .A(n6234), .B(n6233), .Z(n6235) );
  NAND U6832 ( .A(n6236), .B(n6235), .Z(n6422) );
  OR U6833 ( .A(n6238), .B(n6237), .Z(n6242) );
  NANDN U6834 ( .A(n6240), .B(n6239), .Z(n6241) );
  NAND U6835 ( .A(n6242), .B(n6241), .Z(n6421) );
  OR U6836 ( .A(n6244), .B(n6243), .Z(n6248) );
  NANDN U6837 ( .A(n6246), .B(n6245), .Z(n6247) );
  NAND U6838 ( .A(n6248), .B(n6247), .Z(n6420) );
  XOR U6839 ( .A(n6422), .B(n6423), .Z(n6480) );
  NANDN U6840 ( .A(n6250), .B(n6249), .Z(n6254) );
  NAND U6841 ( .A(n6252), .B(n6251), .Z(n6253) );
  NAND U6842 ( .A(n6254), .B(n6253), .Z(n6435) );
  NANDN U6843 ( .A(n6255), .B(n18832), .Z(n6257) );
  XNOR U6844 ( .A(b[19]), .B(a[37]), .Z(n6378) );
  NANDN U6845 ( .A(n6378), .B(n18834), .Z(n6256) );
  NAND U6846 ( .A(n6257), .B(n6256), .Z(n6447) );
  XOR U6847 ( .A(b[27]), .B(n6835), .Z(n6381) );
  NANDN U6848 ( .A(n6381), .B(n19336), .Z(n6260) );
  NANDN U6849 ( .A(n6258), .B(n19337), .Z(n6259) );
  NAND U6850 ( .A(n6260), .B(n6259), .Z(n6444) );
  XOR U6851 ( .A(b[5]), .B(a[51]), .Z(n6384) );
  NAND U6852 ( .A(n6384), .B(n17310), .Z(n6263) );
  NAND U6853 ( .A(n6261), .B(n17311), .Z(n6262) );
  AND U6854 ( .A(n6263), .B(n6262), .Z(n6445) );
  XNOR U6855 ( .A(n6444), .B(n6445), .Z(n6446) );
  XNOR U6856 ( .A(n6447), .B(n6446), .Z(n6433) );
  XOR U6857 ( .A(b[17]), .B(a[39]), .Z(n6387) );
  NAND U6858 ( .A(n6387), .B(n18673), .Z(n6266) );
  NANDN U6859 ( .A(n6264), .B(n18674), .Z(n6265) );
  NAND U6860 ( .A(n6266), .B(n6265), .Z(n6405) );
  XNOR U6861 ( .A(b[31]), .B(a[25]), .Z(n6390) );
  NANDN U6862 ( .A(n6390), .B(n19472), .Z(n6269) );
  NANDN U6863 ( .A(n6267), .B(n19473), .Z(n6268) );
  NAND U6864 ( .A(n6269), .B(n6268), .Z(n6402) );
  OR U6865 ( .A(n6270), .B(n16988), .Z(n6272) );
  XOR U6866 ( .A(b[3]), .B(n10660), .Z(n6393) );
  NANDN U6867 ( .A(n6393), .B(n16990), .Z(n6271) );
  AND U6868 ( .A(n6272), .B(n6271), .Z(n6403) );
  XNOR U6869 ( .A(n6402), .B(n6403), .Z(n6404) );
  XOR U6870 ( .A(n6405), .B(n6404), .Z(n6432) );
  XNOR U6871 ( .A(n6433), .B(n6432), .Z(n6434) );
  XNOR U6872 ( .A(n6435), .B(n6434), .Z(n6481) );
  XNOR U6873 ( .A(n6480), .B(n6481), .Z(n6482) );
  XNOR U6874 ( .A(n6483), .B(n6482), .Z(n6501) );
  OR U6875 ( .A(n6274), .B(n6273), .Z(n6278) );
  NAND U6876 ( .A(n6276), .B(n6275), .Z(n6277) );
  NAND U6877 ( .A(n6278), .B(n6277), .Z(n6499) );
  NANDN U6878 ( .A(n6280), .B(n6279), .Z(n6284) );
  NANDN U6879 ( .A(n6282), .B(n6281), .Z(n6283) );
  NAND U6880 ( .A(n6284), .B(n6283), .Z(n6488) );
  OR U6881 ( .A(n6286), .B(n6285), .Z(n6290) );
  NAND U6882 ( .A(n6288), .B(n6287), .Z(n6289) );
  NAND U6883 ( .A(n6290), .B(n6289), .Z(n6487) );
  NANDN U6884 ( .A(n6292), .B(n6291), .Z(n6296) );
  NAND U6885 ( .A(n6294), .B(n6293), .Z(n6295) );
  NAND U6886 ( .A(n6296), .B(n6295), .Z(n6426) );
  NANDN U6887 ( .A(n6298), .B(n6297), .Z(n6302) );
  NAND U6888 ( .A(n6300), .B(n6299), .Z(n6301) );
  AND U6889 ( .A(n6302), .B(n6301), .Z(n6427) );
  XNOR U6890 ( .A(n6426), .B(n6427), .Z(n6428) );
  XNOR U6891 ( .A(n579), .B(a[47]), .Z(n6450) );
  NAND U6892 ( .A(n17814), .B(n6450), .Z(n6305) );
  NANDN U6893 ( .A(n6303), .B(n17815), .Z(n6304) );
  NAND U6894 ( .A(n6305), .B(n6304), .Z(n6410) );
  NAND U6895 ( .A(n6306), .B(n18513), .Z(n6308) );
  XNOR U6896 ( .A(b[15]), .B(a[41]), .Z(n6453) );
  OR U6897 ( .A(n6453), .B(n18512), .Z(n6307) );
  AND U6898 ( .A(n6308), .B(n6307), .Z(n6408) );
  NANDN U6899 ( .A(n6309), .B(n19013), .Z(n6311) );
  XNOR U6900 ( .A(n582), .B(a[35]), .Z(n6456) );
  NAND U6901 ( .A(n6456), .B(n19015), .Z(n6310) );
  AND U6902 ( .A(n6311), .B(n6310), .Z(n6409) );
  XOR U6903 ( .A(n6410), .B(n6411), .Z(n6399) );
  XNOR U6904 ( .A(b[11]), .B(a[45]), .Z(n6459) );
  OR U6905 ( .A(n6459), .B(n18194), .Z(n6314) );
  NANDN U6906 ( .A(n6312), .B(n18104), .Z(n6313) );
  NAND U6907 ( .A(n6314), .B(n6313), .Z(n6397) );
  XOR U6908 ( .A(n580), .B(a[43]), .Z(n6462) );
  NANDN U6909 ( .A(n6462), .B(n18336), .Z(n6317) );
  NANDN U6910 ( .A(n6315), .B(n18337), .Z(n6316) );
  AND U6911 ( .A(n6317), .B(n6316), .Z(n6396) );
  XNOR U6912 ( .A(n6397), .B(n6396), .Z(n6398) );
  XOR U6913 ( .A(n6399), .B(n6398), .Z(n6416) );
  NANDN U6914 ( .A(n577), .B(a[55]), .Z(n6318) );
  XOR U6915 ( .A(n17151), .B(n6318), .Z(n6320) );
  NANDN U6916 ( .A(b[0]), .B(a[54]), .Z(n6319) );
  AND U6917 ( .A(n6320), .B(n6319), .Z(n6374) );
  NAND U6918 ( .A(n19406), .B(n6321), .Z(n6323) );
  XNOR U6919 ( .A(n584), .B(a[27]), .Z(n6468) );
  NANDN U6920 ( .A(n576), .B(n6468), .Z(n6322) );
  NAND U6921 ( .A(n6323), .B(n6322), .Z(n6372) );
  NANDN U6922 ( .A(n585), .B(a[23]), .Z(n6373) );
  XNOR U6923 ( .A(n6372), .B(n6373), .Z(n6375) );
  XOR U6924 ( .A(n6374), .B(n6375), .Z(n6414) );
  XOR U6925 ( .A(b[23]), .B(a[33]), .Z(n6471) );
  NANDN U6926 ( .A(n19127), .B(n6471), .Z(n6326) );
  NAND U6927 ( .A(n6324), .B(n19128), .Z(n6325) );
  NAND U6928 ( .A(n6326), .B(n6325), .Z(n6441) );
  NAND U6929 ( .A(n6327), .B(n17553), .Z(n6329) );
  XNOR U6930 ( .A(b[7]), .B(a[49]), .Z(n6474) );
  NANDN U6931 ( .A(n6474), .B(n17555), .Z(n6328) );
  NAND U6932 ( .A(n6329), .B(n6328), .Z(n6438) );
  XOR U6933 ( .A(b[25]), .B(a[31]), .Z(n6477) );
  NAND U6934 ( .A(n6477), .B(n19240), .Z(n6332) );
  NANDN U6935 ( .A(n6330), .B(n19242), .Z(n6331) );
  AND U6936 ( .A(n6332), .B(n6331), .Z(n6439) );
  XNOR U6937 ( .A(n6438), .B(n6439), .Z(n6440) );
  XNOR U6938 ( .A(n6441), .B(n6440), .Z(n6415) );
  XOR U6939 ( .A(n6414), .B(n6415), .Z(n6417) );
  XNOR U6940 ( .A(n6416), .B(n6417), .Z(n6429) );
  XNOR U6941 ( .A(n6428), .B(n6429), .Z(n6486) );
  XNOR U6942 ( .A(n6487), .B(n6486), .Z(n6489) );
  XNOR U6943 ( .A(n6488), .B(n6489), .Z(n6498) );
  XNOR U6944 ( .A(n6499), .B(n6498), .Z(n6500) );
  XOR U6945 ( .A(n6501), .B(n6500), .Z(n6495) );
  NANDN U6946 ( .A(n6334), .B(n6333), .Z(n6338) );
  OR U6947 ( .A(n6336), .B(n6335), .Z(n6337) );
  NAND U6948 ( .A(n6338), .B(n6337), .Z(n6492) );
  NAND U6949 ( .A(n6340), .B(n6339), .Z(n6344) );
  NANDN U6950 ( .A(n6342), .B(n6341), .Z(n6343) );
  NAND U6951 ( .A(n6344), .B(n6343), .Z(n6493) );
  XNOR U6952 ( .A(n6492), .B(n6493), .Z(n6494) );
  XNOR U6953 ( .A(n6495), .B(n6494), .Z(n6369) );
  NANDN U6954 ( .A(n6346), .B(n6345), .Z(n6350) );
  NAND U6955 ( .A(n6348), .B(n6347), .Z(n6349) );
  NAND U6956 ( .A(n6350), .B(n6349), .Z(n6366) );
  NANDN U6957 ( .A(n6352), .B(n6351), .Z(n6356) );
  OR U6958 ( .A(n6354), .B(n6353), .Z(n6355) );
  NAND U6959 ( .A(n6356), .B(n6355), .Z(n6367) );
  XNOR U6960 ( .A(n6366), .B(n6367), .Z(n6368) );
  XNOR U6961 ( .A(n6369), .B(n6368), .Z(n6362) );
  XOR U6962 ( .A(n6363), .B(n6362), .Z(n6364) );
  XNOR U6963 ( .A(n6365), .B(n6364), .Z(n6504) );
  XNOR U6964 ( .A(n6504), .B(sreg[151]), .Z(n6506) );
  NAND U6965 ( .A(n6357), .B(sreg[150]), .Z(n6361) );
  OR U6966 ( .A(n6359), .B(n6358), .Z(n6360) );
  AND U6967 ( .A(n6361), .B(n6360), .Z(n6505) );
  XOR U6968 ( .A(n6506), .B(n6505), .Z(c[151]) );
  NANDN U6969 ( .A(n6367), .B(n6366), .Z(n6371) );
  NANDN U6970 ( .A(n6369), .B(n6368), .Z(n6370) );
  NAND U6971 ( .A(n6371), .B(n6370), .Z(n6510) );
  NANDN U6972 ( .A(n6373), .B(n6372), .Z(n6377) );
  NAND U6973 ( .A(n6375), .B(n6374), .Z(n6376) );
  NAND U6974 ( .A(n6377), .B(n6376), .Z(n6582) );
  NANDN U6975 ( .A(n6378), .B(n18832), .Z(n6380) );
  XOR U6976 ( .A(b[19]), .B(n8490), .Z(n6527) );
  NANDN U6977 ( .A(n6527), .B(n18834), .Z(n6379) );
  NAND U6978 ( .A(n6380), .B(n6379), .Z(n6592) );
  XOR U6979 ( .A(b[27]), .B(n7336), .Z(n6530) );
  NANDN U6980 ( .A(n6530), .B(n19336), .Z(n6383) );
  NANDN U6981 ( .A(n6381), .B(n19337), .Z(n6382) );
  NAND U6982 ( .A(n6383), .B(n6382), .Z(n6589) );
  XOR U6983 ( .A(b[5]), .B(a[52]), .Z(n6533) );
  NAND U6984 ( .A(n6533), .B(n17310), .Z(n6386) );
  NAND U6985 ( .A(n6384), .B(n17311), .Z(n6385) );
  AND U6986 ( .A(n6386), .B(n6385), .Z(n6590) );
  XNOR U6987 ( .A(n6589), .B(n6590), .Z(n6591) );
  XNOR U6988 ( .A(n6592), .B(n6591), .Z(n6580) );
  XOR U6989 ( .A(b[17]), .B(a[40]), .Z(n6536) );
  NAND U6990 ( .A(n6536), .B(n18673), .Z(n6389) );
  NAND U6991 ( .A(n6387), .B(n18674), .Z(n6388) );
  NAND U6992 ( .A(n6389), .B(n6388), .Z(n6554) );
  XNOR U6993 ( .A(b[31]), .B(a[26]), .Z(n6539) );
  NANDN U6994 ( .A(n6539), .B(n19472), .Z(n6392) );
  NANDN U6995 ( .A(n6390), .B(n19473), .Z(n6391) );
  NAND U6996 ( .A(n6392), .B(n6391), .Z(n6551) );
  OR U6997 ( .A(n6393), .B(n16988), .Z(n6395) );
  XNOR U6998 ( .A(b[3]), .B(a[54]), .Z(n6542) );
  NANDN U6999 ( .A(n6542), .B(n16990), .Z(n6394) );
  AND U7000 ( .A(n6395), .B(n6394), .Z(n6552) );
  XNOR U7001 ( .A(n6551), .B(n6552), .Z(n6553) );
  XOR U7002 ( .A(n6554), .B(n6553), .Z(n6579) );
  XNOR U7003 ( .A(n6580), .B(n6579), .Z(n6581) );
  XNOR U7004 ( .A(n6582), .B(n6581), .Z(n6625) );
  NANDN U7005 ( .A(n6397), .B(n6396), .Z(n6401) );
  NAND U7006 ( .A(n6399), .B(n6398), .Z(n6400) );
  NAND U7007 ( .A(n6401), .B(n6400), .Z(n6570) );
  NANDN U7008 ( .A(n6403), .B(n6402), .Z(n6407) );
  NAND U7009 ( .A(n6405), .B(n6404), .Z(n6406) );
  NAND U7010 ( .A(n6407), .B(n6406), .Z(n6568) );
  OR U7011 ( .A(n6409), .B(n6408), .Z(n6413) );
  NANDN U7012 ( .A(n6411), .B(n6410), .Z(n6412) );
  NAND U7013 ( .A(n6413), .B(n6412), .Z(n6567) );
  XNOR U7014 ( .A(n6570), .B(n6569), .Z(n6626) );
  XOR U7015 ( .A(n6625), .B(n6626), .Z(n6628) );
  NANDN U7016 ( .A(n6415), .B(n6414), .Z(n6419) );
  OR U7017 ( .A(n6417), .B(n6416), .Z(n6418) );
  NAND U7018 ( .A(n6419), .B(n6418), .Z(n6627) );
  XOR U7019 ( .A(n6628), .B(n6627), .Z(n6645) );
  OR U7020 ( .A(n6421), .B(n6420), .Z(n6425) );
  NANDN U7021 ( .A(n6423), .B(n6422), .Z(n6424) );
  NAND U7022 ( .A(n6425), .B(n6424), .Z(n6644) );
  NANDN U7023 ( .A(n6427), .B(n6426), .Z(n6431) );
  NANDN U7024 ( .A(n6429), .B(n6428), .Z(n6430) );
  NAND U7025 ( .A(n6431), .B(n6430), .Z(n6633) );
  NANDN U7026 ( .A(n6433), .B(n6432), .Z(n6437) );
  NAND U7027 ( .A(n6435), .B(n6434), .Z(n6436) );
  NAND U7028 ( .A(n6437), .B(n6436), .Z(n6632) );
  NANDN U7029 ( .A(n6439), .B(n6438), .Z(n6443) );
  NAND U7030 ( .A(n6441), .B(n6440), .Z(n6442) );
  NAND U7031 ( .A(n6443), .B(n6442), .Z(n6573) );
  NANDN U7032 ( .A(n6445), .B(n6444), .Z(n6449) );
  NAND U7033 ( .A(n6447), .B(n6446), .Z(n6448) );
  AND U7034 ( .A(n6449), .B(n6448), .Z(n6574) );
  XNOR U7035 ( .A(n6573), .B(n6574), .Z(n6575) );
  XOR U7036 ( .A(n579), .B(a[48]), .Z(n6595) );
  NANDN U7037 ( .A(n6595), .B(n17814), .Z(n6452) );
  NAND U7038 ( .A(n17815), .B(n6450), .Z(n6451) );
  NAND U7039 ( .A(n6452), .B(n6451), .Z(n6559) );
  XNOR U7040 ( .A(b[15]), .B(a[42]), .Z(n6598) );
  OR U7041 ( .A(n6598), .B(n18512), .Z(n6455) );
  NANDN U7042 ( .A(n6453), .B(n18513), .Z(n6454) );
  NAND U7043 ( .A(n6455), .B(n6454), .Z(n6557) );
  XOR U7044 ( .A(n582), .B(a[36]), .Z(n6601) );
  NANDN U7045 ( .A(n6601), .B(n19015), .Z(n6458) );
  NAND U7046 ( .A(n19013), .B(n6456), .Z(n6457) );
  NAND U7047 ( .A(n6458), .B(n6457), .Z(n6558) );
  XNOR U7048 ( .A(n6557), .B(n6558), .Z(n6560) );
  XOR U7049 ( .A(n6559), .B(n6560), .Z(n6548) );
  XNOR U7050 ( .A(b[11]), .B(a[46]), .Z(n6604) );
  OR U7051 ( .A(n6604), .B(n18194), .Z(n6461) );
  NANDN U7052 ( .A(n6459), .B(n18104), .Z(n6460) );
  NAND U7053 ( .A(n6461), .B(n6460), .Z(n6546) );
  XOR U7054 ( .A(n580), .B(a[44]), .Z(n6607) );
  NANDN U7055 ( .A(n6607), .B(n18336), .Z(n6464) );
  NANDN U7056 ( .A(n6462), .B(n18337), .Z(n6463) );
  AND U7057 ( .A(n6464), .B(n6463), .Z(n6545) );
  XNOR U7058 ( .A(n6546), .B(n6545), .Z(n6547) );
  XNOR U7059 ( .A(n6548), .B(n6547), .Z(n6564) );
  NANDN U7060 ( .A(n577), .B(a[56]), .Z(n6465) );
  XOR U7061 ( .A(n17151), .B(n6465), .Z(n6467) );
  IV U7062 ( .A(a[55]), .Z(n10959) );
  NANDN U7063 ( .A(n10959), .B(n577), .Z(n6466) );
  AND U7064 ( .A(n6467), .B(n6466), .Z(n6523) );
  NAND U7065 ( .A(n19406), .B(n6468), .Z(n6470) );
  XNOR U7066 ( .A(n584), .B(a[28]), .Z(n6613) );
  NANDN U7067 ( .A(n576), .B(n6613), .Z(n6469) );
  NAND U7068 ( .A(n6470), .B(n6469), .Z(n6521) );
  NANDN U7069 ( .A(n585), .B(a[24]), .Z(n6522) );
  XNOR U7070 ( .A(n6521), .B(n6522), .Z(n6524) );
  XNOR U7071 ( .A(n6523), .B(n6524), .Z(n6562) );
  XOR U7072 ( .A(b[23]), .B(a[34]), .Z(n6616) );
  NANDN U7073 ( .A(n19127), .B(n6616), .Z(n6473) );
  NAND U7074 ( .A(n6471), .B(n19128), .Z(n6472) );
  NAND U7075 ( .A(n6473), .B(n6472), .Z(n6586) );
  NANDN U7076 ( .A(n6474), .B(n17553), .Z(n6476) );
  XOR U7077 ( .A(b[7]), .B(a[50]), .Z(n6619) );
  NAND U7078 ( .A(n6619), .B(n17555), .Z(n6475) );
  NAND U7079 ( .A(n6476), .B(n6475), .Z(n6583) );
  XOR U7080 ( .A(b[25]), .B(a[32]), .Z(n6622) );
  NAND U7081 ( .A(n6622), .B(n19240), .Z(n6479) );
  NAND U7082 ( .A(n6477), .B(n19242), .Z(n6478) );
  AND U7083 ( .A(n6479), .B(n6478), .Z(n6584) );
  XNOR U7084 ( .A(n6583), .B(n6584), .Z(n6585) );
  XOR U7085 ( .A(n6586), .B(n6585), .Z(n6561) );
  XOR U7086 ( .A(n6564), .B(n6563), .Z(n6576) );
  XOR U7087 ( .A(n6575), .B(n6576), .Z(n6631) );
  XNOR U7088 ( .A(n6632), .B(n6631), .Z(n6634) );
  XNOR U7089 ( .A(n6633), .B(n6634), .Z(n6643) );
  XOR U7090 ( .A(n6644), .B(n6643), .Z(n6646) );
  NANDN U7091 ( .A(n6481), .B(n6480), .Z(n6485) );
  NAND U7092 ( .A(n6483), .B(n6482), .Z(n6484) );
  NAND U7093 ( .A(n6485), .B(n6484), .Z(n6638) );
  NAND U7094 ( .A(n6487), .B(n6486), .Z(n6491) );
  NANDN U7095 ( .A(n6489), .B(n6488), .Z(n6490) );
  AND U7096 ( .A(n6491), .B(n6490), .Z(n6637) );
  XNOR U7097 ( .A(n6638), .B(n6637), .Z(n6639) );
  XOR U7098 ( .A(n6640), .B(n6639), .Z(n6517) );
  NANDN U7099 ( .A(n6493), .B(n6492), .Z(n6497) );
  NAND U7100 ( .A(n6495), .B(n6494), .Z(n6496) );
  NAND U7101 ( .A(n6497), .B(n6496), .Z(n6515) );
  NANDN U7102 ( .A(n6499), .B(n6498), .Z(n6503) );
  NANDN U7103 ( .A(n6501), .B(n6500), .Z(n6502) );
  NAND U7104 ( .A(n6503), .B(n6502), .Z(n6516) );
  XNOR U7105 ( .A(n6515), .B(n6516), .Z(n6518) );
  XOR U7106 ( .A(n6517), .B(n6518), .Z(n6509) );
  XOR U7107 ( .A(n6510), .B(n6509), .Z(n6511) );
  XNOR U7108 ( .A(n6512), .B(n6511), .Z(n6649) );
  XNOR U7109 ( .A(n6649), .B(sreg[152]), .Z(n6651) );
  NAND U7110 ( .A(n6504), .B(sreg[151]), .Z(n6508) );
  OR U7111 ( .A(n6506), .B(n6505), .Z(n6507) );
  AND U7112 ( .A(n6508), .B(n6507), .Z(n6650) );
  XOR U7113 ( .A(n6651), .B(n6650), .Z(c[152]) );
  NAND U7114 ( .A(n6510), .B(n6509), .Z(n6514) );
  NAND U7115 ( .A(n6512), .B(n6511), .Z(n6513) );
  NAND U7116 ( .A(n6514), .B(n6513), .Z(n6657) );
  NANDN U7117 ( .A(n6516), .B(n6515), .Z(n6520) );
  NAND U7118 ( .A(n6518), .B(n6517), .Z(n6519) );
  NAND U7119 ( .A(n6520), .B(n6519), .Z(n6655) );
  NANDN U7120 ( .A(n6522), .B(n6521), .Z(n6526) );
  NAND U7121 ( .A(n6524), .B(n6523), .Z(n6525) );
  NAND U7122 ( .A(n6526), .B(n6525), .Z(n6735) );
  NANDN U7123 ( .A(n6527), .B(n18832), .Z(n6529) );
  XNOR U7124 ( .A(b[19]), .B(a[39]), .Z(n6682) );
  NANDN U7125 ( .A(n6682), .B(n18834), .Z(n6528) );
  NAND U7126 ( .A(n6529), .B(n6528), .Z(n6745) );
  XNOR U7127 ( .A(b[27]), .B(a[31]), .Z(n6685) );
  NANDN U7128 ( .A(n6685), .B(n19336), .Z(n6532) );
  NANDN U7129 ( .A(n6530), .B(n19337), .Z(n6531) );
  NAND U7130 ( .A(n6532), .B(n6531), .Z(n6742) );
  XNOR U7131 ( .A(b[5]), .B(a[53]), .Z(n6688) );
  NANDN U7132 ( .A(n6688), .B(n17310), .Z(n6535) );
  NAND U7133 ( .A(n6533), .B(n17311), .Z(n6534) );
  AND U7134 ( .A(n6535), .B(n6534), .Z(n6743) );
  XNOR U7135 ( .A(n6742), .B(n6743), .Z(n6744) );
  XNOR U7136 ( .A(n6745), .B(n6744), .Z(n6733) );
  XNOR U7137 ( .A(b[17]), .B(a[41]), .Z(n6691) );
  NANDN U7138 ( .A(n6691), .B(n18673), .Z(n6538) );
  NAND U7139 ( .A(n6536), .B(n18674), .Z(n6537) );
  NAND U7140 ( .A(n6538), .B(n6537), .Z(n6709) );
  XNOR U7141 ( .A(b[31]), .B(a[27]), .Z(n6694) );
  NANDN U7142 ( .A(n6694), .B(n19472), .Z(n6541) );
  NANDN U7143 ( .A(n6539), .B(n19473), .Z(n6540) );
  NAND U7144 ( .A(n6541), .B(n6540), .Z(n6706) );
  OR U7145 ( .A(n6542), .B(n16988), .Z(n6544) );
  XOR U7146 ( .A(b[3]), .B(n10959), .Z(n6697) );
  NANDN U7147 ( .A(n6697), .B(n16990), .Z(n6543) );
  AND U7148 ( .A(n6544), .B(n6543), .Z(n6707) );
  XNOR U7149 ( .A(n6706), .B(n6707), .Z(n6708) );
  XOR U7150 ( .A(n6709), .B(n6708), .Z(n6732) );
  XNOR U7151 ( .A(n6733), .B(n6732), .Z(n6734) );
  XNOR U7152 ( .A(n6735), .B(n6734), .Z(n6673) );
  NANDN U7153 ( .A(n6546), .B(n6545), .Z(n6550) );
  NAND U7154 ( .A(n6548), .B(n6547), .Z(n6549) );
  NAND U7155 ( .A(n6550), .B(n6549), .Z(n6724) );
  NANDN U7156 ( .A(n6552), .B(n6551), .Z(n6556) );
  NAND U7157 ( .A(n6554), .B(n6553), .Z(n6555) );
  NAND U7158 ( .A(n6556), .B(n6555), .Z(n6723) );
  XNOR U7159 ( .A(n6723), .B(n6722), .Z(n6725) );
  XOR U7160 ( .A(n6724), .B(n6725), .Z(n6672) );
  XOR U7161 ( .A(n6673), .B(n6672), .Z(n6674) );
  NANDN U7162 ( .A(n6562), .B(n6561), .Z(n6566) );
  NAND U7163 ( .A(n6564), .B(n6563), .Z(n6565) );
  NAND U7164 ( .A(n6566), .B(n6565), .Z(n6675) );
  XNOR U7165 ( .A(n6674), .B(n6675), .Z(n6786) );
  OR U7166 ( .A(n6568), .B(n6567), .Z(n6572) );
  NAND U7167 ( .A(n6570), .B(n6569), .Z(n6571) );
  NAND U7168 ( .A(n6572), .B(n6571), .Z(n6785) );
  NANDN U7169 ( .A(n6574), .B(n6573), .Z(n6578) );
  NAND U7170 ( .A(n6576), .B(n6575), .Z(n6577) );
  NAND U7171 ( .A(n6578), .B(n6577), .Z(n6668) );
  NANDN U7172 ( .A(n6584), .B(n6583), .Z(n6588) );
  NAND U7173 ( .A(n6586), .B(n6585), .Z(n6587) );
  NAND U7174 ( .A(n6588), .B(n6587), .Z(n6726) );
  NANDN U7175 ( .A(n6590), .B(n6589), .Z(n6594) );
  NAND U7176 ( .A(n6592), .B(n6591), .Z(n6593) );
  AND U7177 ( .A(n6594), .B(n6593), .Z(n6727) );
  XNOR U7178 ( .A(n6726), .B(n6727), .Z(n6728) );
  XOR U7179 ( .A(b[9]), .B(n10083), .Z(n6748) );
  NANDN U7180 ( .A(n6748), .B(n17814), .Z(n6597) );
  NANDN U7181 ( .A(n6595), .B(n17815), .Z(n6596) );
  NAND U7182 ( .A(n6597), .B(n6596), .Z(n6714) );
  XNOR U7183 ( .A(b[15]), .B(a[43]), .Z(n6751) );
  OR U7184 ( .A(n6751), .B(n18512), .Z(n6600) );
  NANDN U7185 ( .A(n6598), .B(n18513), .Z(n6599) );
  NAND U7186 ( .A(n6600), .B(n6599), .Z(n6712) );
  XNOR U7187 ( .A(b[21]), .B(a[37]), .Z(n6754) );
  NANDN U7188 ( .A(n6754), .B(n19015), .Z(n6603) );
  NANDN U7189 ( .A(n6601), .B(n19013), .Z(n6602) );
  NAND U7190 ( .A(n6603), .B(n6602), .Z(n6713) );
  XNOR U7191 ( .A(n6712), .B(n6713), .Z(n6715) );
  XOR U7192 ( .A(n6714), .B(n6715), .Z(n6703) );
  XNOR U7193 ( .A(b[11]), .B(a[47]), .Z(n6757) );
  OR U7194 ( .A(n6757), .B(n18194), .Z(n6606) );
  NANDN U7195 ( .A(n6604), .B(n18104), .Z(n6605) );
  NAND U7196 ( .A(n6606), .B(n6605), .Z(n6701) );
  XOR U7197 ( .A(n580), .B(a[45]), .Z(n6760) );
  NANDN U7198 ( .A(n6760), .B(n18336), .Z(n6609) );
  NANDN U7199 ( .A(n6607), .B(n18337), .Z(n6608) );
  AND U7200 ( .A(n6609), .B(n6608), .Z(n6700) );
  XNOR U7201 ( .A(n6701), .B(n6700), .Z(n6702) );
  XNOR U7202 ( .A(n6703), .B(n6702), .Z(n6719) );
  NANDN U7203 ( .A(n577), .B(a[57]), .Z(n6610) );
  XOR U7204 ( .A(n17151), .B(n6610), .Z(n6612) );
  NANDN U7205 ( .A(b[0]), .B(a[56]), .Z(n6611) );
  AND U7206 ( .A(n6612), .B(n6611), .Z(n6678) );
  NAND U7207 ( .A(n19406), .B(n6613), .Z(n6615) );
  XOR U7208 ( .A(n584), .B(n6835), .Z(n6766) );
  NANDN U7209 ( .A(n576), .B(n6766), .Z(n6614) );
  NAND U7210 ( .A(n6615), .B(n6614), .Z(n6676) );
  NANDN U7211 ( .A(n585), .B(a[25]), .Z(n6677) );
  XNOR U7212 ( .A(n6676), .B(n6677), .Z(n6679) );
  XNOR U7213 ( .A(n6678), .B(n6679), .Z(n6717) );
  XOR U7214 ( .A(b[23]), .B(a[35]), .Z(n6769) );
  NANDN U7215 ( .A(n19127), .B(n6769), .Z(n6618) );
  NAND U7216 ( .A(n6616), .B(n19128), .Z(n6617) );
  NAND U7217 ( .A(n6618), .B(n6617), .Z(n6739) );
  NAND U7218 ( .A(n6619), .B(n17553), .Z(n6621) );
  XOR U7219 ( .A(b[7]), .B(a[51]), .Z(n6772) );
  NAND U7220 ( .A(n6772), .B(n17555), .Z(n6620) );
  NAND U7221 ( .A(n6621), .B(n6620), .Z(n6736) );
  XOR U7222 ( .A(b[25]), .B(a[33]), .Z(n6775) );
  NAND U7223 ( .A(n6775), .B(n19240), .Z(n6624) );
  NAND U7224 ( .A(n6622), .B(n19242), .Z(n6623) );
  AND U7225 ( .A(n6624), .B(n6623), .Z(n6737) );
  XNOR U7226 ( .A(n6736), .B(n6737), .Z(n6738) );
  XOR U7227 ( .A(n6739), .B(n6738), .Z(n6716) );
  XOR U7228 ( .A(n6719), .B(n6718), .Z(n6729) );
  XOR U7229 ( .A(n6728), .B(n6729), .Z(n6666) );
  XNOR U7230 ( .A(n6667), .B(n6666), .Z(n6669) );
  XNOR U7231 ( .A(n6668), .B(n6669), .Z(n6784) );
  XOR U7232 ( .A(n6785), .B(n6784), .Z(n6787) );
  NANDN U7233 ( .A(n6626), .B(n6625), .Z(n6630) );
  OR U7234 ( .A(n6628), .B(n6627), .Z(n6629) );
  NAND U7235 ( .A(n6630), .B(n6629), .Z(n6778) );
  NAND U7236 ( .A(n6632), .B(n6631), .Z(n6636) );
  NANDN U7237 ( .A(n6634), .B(n6633), .Z(n6635) );
  NAND U7238 ( .A(n6636), .B(n6635), .Z(n6779) );
  XNOR U7239 ( .A(n6778), .B(n6779), .Z(n6780) );
  XOR U7240 ( .A(n6781), .B(n6780), .Z(n6662) );
  NANDN U7241 ( .A(n6638), .B(n6637), .Z(n6642) );
  NAND U7242 ( .A(n6640), .B(n6639), .Z(n6641) );
  NAND U7243 ( .A(n6642), .B(n6641), .Z(n6660) );
  NANDN U7244 ( .A(n6644), .B(n6643), .Z(n6648) );
  OR U7245 ( .A(n6646), .B(n6645), .Z(n6647) );
  NAND U7246 ( .A(n6648), .B(n6647), .Z(n6661) );
  XNOR U7247 ( .A(n6660), .B(n6661), .Z(n6663) );
  XOR U7248 ( .A(n6662), .B(n6663), .Z(n6654) );
  XOR U7249 ( .A(n6655), .B(n6654), .Z(n6656) );
  XNOR U7250 ( .A(n6657), .B(n6656), .Z(n6790) );
  XNOR U7251 ( .A(n6790), .B(sreg[153]), .Z(n6792) );
  NAND U7252 ( .A(n6649), .B(sreg[152]), .Z(n6653) );
  OR U7253 ( .A(n6651), .B(n6650), .Z(n6652) );
  AND U7254 ( .A(n6653), .B(n6652), .Z(n6791) );
  XOR U7255 ( .A(n6792), .B(n6791), .Z(c[153]) );
  NAND U7256 ( .A(n6655), .B(n6654), .Z(n6659) );
  NAND U7257 ( .A(n6657), .B(n6656), .Z(n6658) );
  NAND U7258 ( .A(n6659), .B(n6658), .Z(n6798) );
  NANDN U7259 ( .A(n6661), .B(n6660), .Z(n6665) );
  NAND U7260 ( .A(n6663), .B(n6662), .Z(n6664) );
  NAND U7261 ( .A(n6665), .B(n6664), .Z(n6795) );
  NAND U7262 ( .A(n6667), .B(n6666), .Z(n6671) );
  NANDN U7263 ( .A(n6669), .B(n6668), .Z(n6670) );
  NAND U7264 ( .A(n6671), .B(n6670), .Z(n6922) );
  XNOR U7265 ( .A(n6922), .B(n6923), .Z(n6924) );
  NANDN U7266 ( .A(n6677), .B(n6676), .Z(n6681) );
  NAND U7267 ( .A(n6679), .B(n6678), .Z(n6680) );
  NAND U7268 ( .A(n6681), .B(n6680), .Z(n6879) );
  NANDN U7269 ( .A(n6682), .B(n18832), .Z(n6684) );
  XNOR U7270 ( .A(b[19]), .B(a[40]), .Z(n6823) );
  NANDN U7271 ( .A(n6823), .B(n18834), .Z(n6683) );
  NAND U7272 ( .A(n6684), .B(n6683), .Z(n6889) );
  XNOR U7273 ( .A(b[27]), .B(a[32]), .Z(n6826) );
  NANDN U7274 ( .A(n6826), .B(n19336), .Z(n6687) );
  NANDN U7275 ( .A(n6685), .B(n19337), .Z(n6686) );
  NAND U7276 ( .A(n6687), .B(n6686), .Z(n6886) );
  XOR U7277 ( .A(b[5]), .B(a[54]), .Z(n6829) );
  NAND U7278 ( .A(n6829), .B(n17310), .Z(n6690) );
  NANDN U7279 ( .A(n6688), .B(n17311), .Z(n6689) );
  AND U7280 ( .A(n6690), .B(n6689), .Z(n6887) );
  XNOR U7281 ( .A(n6886), .B(n6887), .Z(n6888) );
  XNOR U7282 ( .A(n6889), .B(n6888), .Z(n6877) );
  XNOR U7283 ( .A(b[17]), .B(a[42]), .Z(n6832) );
  NANDN U7284 ( .A(n6832), .B(n18673), .Z(n6693) );
  NANDN U7285 ( .A(n6691), .B(n18674), .Z(n6692) );
  NAND U7286 ( .A(n6693), .B(n6692), .Z(n6851) );
  XNOR U7287 ( .A(b[31]), .B(a[28]), .Z(n6836) );
  NANDN U7288 ( .A(n6836), .B(n19472), .Z(n6696) );
  NANDN U7289 ( .A(n6694), .B(n19473), .Z(n6695) );
  NAND U7290 ( .A(n6696), .B(n6695), .Z(n6848) );
  OR U7291 ( .A(n6697), .B(n16988), .Z(n6699) );
  XNOR U7292 ( .A(b[3]), .B(a[56]), .Z(n6839) );
  NANDN U7293 ( .A(n6839), .B(n16990), .Z(n6698) );
  AND U7294 ( .A(n6699), .B(n6698), .Z(n6849) );
  XNOR U7295 ( .A(n6848), .B(n6849), .Z(n6850) );
  XOR U7296 ( .A(n6851), .B(n6850), .Z(n6876) );
  XNOR U7297 ( .A(n6877), .B(n6876), .Z(n6878) );
  XNOR U7298 ( .A(n6879), .B(n6878), .Z(n6814) );
  NANDN U7299 ( .A(n6701), .B(n6700), .Z(n6705) );
  NAND U7300 ( .A(n6703), .B(n6702), .Z(n6704) );
  NAND U7301 ( .A(n6705), .B(n6704), .Z(n6868) );
  NANDN U7302 ( .A(n6707), .B(n6706), .Z(n6711) );
  NAND U7303 ( .A(n6709), .B(n6708), .Z(n6710) );
  NAND U7304 ( .A(n6711), .B(n6710), .Z(n6867) );
  XNOR U7305 ( .A(n6867), .B(n6866), .Z(n6869) );
  XOR U7306 ( .A(n6868), .B(n6869), .Z(n6813) );
  XOR U7307 ( .A(n6814), .B(n6813), .Z(n6815) );
  NANDN U7308 ( .A(n6717), .B(n6716), .Z(n6721) );
  NAND U7309 ( .A(n6719), .B(n6718), .Z(n6720) );
  AND U7310 ( .A(n6721), .B(n6720), .Z(n6816) );
  XOR U7311 ( .A(n6815), .B(n6816), .Z(n6930) );
  NANDN U7312 ( .A(n6727), .B(n6726), .Z(n6731) );
  NAND U7313 ( .A(n6729), .B(n6728), .Z(n6730) );
  NAND U7314 ( .A(n6731), .B(n6730), .Z(n6810) );
  NANDN U7315 ( .A(n6737), .B(n6736), .Z(n6741) );
  NAND U7316 ( .A(n6739), .B(n6738), .Z(n6740) );
  NAND U7317 ( .A(n6741), .B(n6740), .Z(n6870) );
  NANDN U7318 ( .A(n6743), .B(n6742), .Z(n6747) );
  NAND U7319 ( .A(n6745), .B(n6744), .Z(n6746) );
  AND U7320 ( .A(n6747), .B(n6746), .Z(n6871) );
  XNOR U7321 ( .A(n6870), .B(n6871), .Z(n6872) );
  XNOR U7322 ( .A(n579), .B(a[50]), .Z(n6892) );
  NAND U7323 ( .A(n17814), .B(n6892), .Z(n6750) );
  NANDN U7324 ( .A(n6748), .B(n17815), .Z(n6749) );
  NAND U7325 ( .A(n6750), .B(n6749), .Z(n6856) );
  NANDN U7326 ( .A(n6751), .B(n18513), .Z(n6753) );
  XOR U7327 ( .A(b[15]), .B(a[44]), .Z(n6895) );
  NANDN U7328 ( .A(n18512), .B(n6895), .Z(n6752) );
  AND U7329 ( .A(n6753), .B(n6752), .Z(n6854) );
  NANDN U7330 ( .A(n6754), .B(n19013), .Z(n6756) );
  XOR U7331 ( .A(n582), .B(n8490), .Z(n6898) );
  NAND U7332 ( .A(n6898), .B(n19015), .Z(n6755) );
  AND U7333 ( .A(n6756), .B(n6755), .Z(n6855) );
  XOR U7334 ( .A(n6856), .B(n6857), .Z(n6845) );
  XNOR U7335 ( .A(b[11]), .B(a[48]), .Z(n6901) );
  OR U7336 ( .A(n6901), .B(n18194), .Z(n6759) );
  NANDN U7337 ( .A(n6757), .B(n18104), .Z(n6758) );
  NAND U7338 ( .A(n6759), .B(n6758), .Z(n6843) );
  XOR U7339 ( .A(n580), .B(a[46]), .Z(n6904) );
  NANDN U7340 ( .A(n6904), .B(n18336), .Z(n6762) );
  NANDN U7341 ( .A(n6760), .B(n18337), .Z(n6761) );
  AND U7342 ( .A(n6762), .B(n6761), .Z(n6842) );
  XNOR U7343 ( .A(n6843), .B(n6842), .Z(n6844) );
  XOR U7344 ( .A(n6845), .B(n6844), .Z(n6862) );
  NANDN U7345 ( .A(n577), .B(a[58]), .Z(n6763) );
  XOR U7346 ( .A(n17151), .B(n6763), .Z(n6765) );
  NANDN U7347 ( .A(b[0]), .B(a[57]), .Z(n6764) );
  AND U7348 ( .A(n6765), .B(n6764), .Z(n6819) );
  NAND U7349 ( .A(n19406), .B(n6766), .Z(n6768) );
  XOR U7350 ( .A(n584), .B(n7336), .Z(n6907) );
  NANDN U7351 ( .A(n576), .B(n6907), .Z(n6767) );
  NAND U7352 ( .A(n6768), .B(n6767), .Z(n6817) );
  NANDN U7353 ( .A(n585), .B(a[26]), .Z(n6818) );
  XNOR U7354 ( .A(n6817), .B(n6818), .Z(n6820) );
  XOR U7355 ( .A(n6819), .B(n6820), .Z(n6860) );
  XOR U7356 ( .A(b[23]), .B(a[36]), .Z(n6913) );
  NANDN U7357 ( .A(n19127), .B(n6913), .Z(n6771) );
  NAND U7358 ( .A(n6769), .B(n19128), .Z(n6770) );
  NAND U7359 ( .A(n6771), .B(n6770), .Z(n6883) );
  NAND U7360 ( .A(n6772), .B(n17553), .Z(n6774) );
  XOR U7361 ( .A(b[7]), .B(a[52]), .Z(n6916) );
  NAND U7362 ( .A(n6916), .B(n17555), .Z(n6773) );
  NAND U7363 ( .A(n6774), .B(n6773), .Z(n6880) );
  XOR U7364 ( .A(b[25]), .B(a[34]), .Z(n6919) );
  NAND U7365 ( .A(n6919), .B(n19240), .Z(n6777) );
  NAND U7366 ( .A(n6775), .B(n19242), .Z(n6776) );
  AND U7367 ( .A(n6777), .B(n6776), .Z(n6881) );
  XNOR U7368 ( .A(n6880), .B(n6881), .Z(n6882) );
  XNOR U7369 ( .A(n6883), .B(n6882), .Z(n6861) );
  XOR U7370 ( .A(n6860), .B(n6861), .Z(n6863) );
  XNOR U7371 ( .A(n6862), .B(n6863), .Z(n6873) );
  XOR U7372 ( .A(n6872), .B(n6873), .Z(n6808) );
  XNOR U7373 ( .A(n6807), .B(n6808), .Z(n6809) );
  XNOR U7374 ( .A(n6810), .B(n6809), .Z(n6928) );
  XNOR U7375 ( .A(n6929), .B(n6928), .Z(n6931) );
  XNOR U7376 ( .A(n6930), .B(n6931), .Z(n6925) );
  XOR U7377 ( .A(n6924), .B(n6925), .Z(n6804) );
  NANDN U7378 ( .A(n6779), .B(n6778), .Z(n6783) );
  NAND U7379 ( .A(n6781), .B(n6780), .Z(n6782) );
  NAND U7380 ( .A(n6783), .B(n6782), .Z(n6801) );
  NANDN U7381 ( .A(n6785), .B(n6784), .Z(n6789) );
  OR U7382 ( .A(n6787), .B(n6786), .Z(n6788) );
  NAND U7383 ( .A(n6789), .B(n6788), .Z(n6802) );
  XNOR U7384 ( .A(n6801), .B(n6802), .Z(n6803) );
  XNOR U7385 ( .A(n6804), .B(n6803), .Z(n6796) );
  XNOR U7386 ( .A(n6795), .B(n6796), .Z(n6797) );
  XNOR U7387 ( .A(n6798), .B(n6797), .Z(n6934) );
  XNOR U7388 ( .A(n6934), .B(sreg[154]), .Z(n6936) );
  NAND U7389 ( .A(n6790), .B(sreg[153]), .Z(n6794) );
  OR U7390 ( .A(n6792), .B(n6791), .Z(n6793) );
  AND U7391 ( .A(n6794), .B(n6793), .Z(n6935) );
  XOR U7392 ( .A(n6936), .B(n6935), .Z(c[154]) );
  NANDN U7393 ( .A(n6796), .B(n6795), .Z(n6800) );
  NAND U7394 ( .A(n6798), .B(n6797), .Z(n6799) );
  NAND U7395 ( .A(n6800), .B(n6799), .Z(n6942) );
  NANDN U7396 ( .A(n6802), .B(n6801), .Z(n6806) );
  NAND U7397 ( .A(n6804), .B(n6803), .Z(n6805) );
  NAND U7398 ( .A(n6806), .B(n6805), .Z(n6939) );
  NANDN U7399 ( .A(n6808), .B(n6807), .Z(n6812) );
  NAND U7400 ( .A(n6810), .B(n6809), .Z(n6811) );
  NAND U7401 ( .A(n6812), .B(n6811), .Z(n7067) );
  XNOR U7402 ( .A(n7067), .B(n7068), .Z(n7069) );
  NANDN U7403 ( .A(n6818), .B(n6817), .Z(n6822) );
  NAND U7404 ( .A(n6820), .B(n6819), .Z(n6821) );
  NAND U7405 ( .A(n6822), .B(n6821), .Z(n7012) );
  NANDN U7406 ( .A(n6823), .B(n18832), .Z(n6825) );
  XOR U7407 ( .A(b[19]), .B(n8930), .Z(n6957) );
  NANDN U7408 ( .A(n6957), .B(n18834), .Z(n6824) );
  NAND U7409 ( .A(n6825), .B(n6824), .Z(n7022) );
  XNOR U7410 ( .A(b[27]), .B(a[33]), .Z(n6960) );
  NANDN U7411 ( .A(n6960), .B(n19336), .Z(n6828) );
  NANDN U7412 ( .A(n6826), .B(n19337), .Z(n6827) );
  NAND U7413 ( .A(n6828), .B(n6827), .Z(n7019) );
  XNOR U7414 ( .A(b[5]), .B(a[55]), .Z(n6963) );
  NANDN U7415 ( .A(n6963), .B(n17310), .Z(n6831) );
  NAND U7416 ( .A(n6829), .B(n17311), .Z(n6830) );
  AND U7417 ( .A(n6831), .B(n6830), .Z(n7020) );
  XNOR U7418 ( .A(n7019), .B(n7020), .Z(n7021) );
  XNOR U7419 ( .A(n7022), .B(n7021), .Z(n7010) );
  XOR U7420 ( .A(b[17]), .B(a[43]), .Z(n6966) );
  NAND U7421 ( .A(n6966), .B(n18673), .Z(n6834) );
  NANDN U7422 ( .A(n6832), .B(n18674), .Z(n6833) );
  NAND U7423 ( .A(n6834), .B(n6833), .Z(n6984) );
  XOR U7424 ( .A(b[31]), .B(n6835), .Z(n6969) );
  NANDN U7425 ( .A(n6969), .B(n19472), .Z(n6838) );
  NANDN U7426 ( .A(n6836), .B(n19473), .Z(n6837) );
  NAND U7427 ( .A(n6838), .B(n6837), .Z(n6981) );
  OR U7428 ( .A(n6839), .B(n16988), .Z(n6841) );
  XNOR U7429 ( .A(b[3]), .B(a[57]), .Z(n6972) );
  NANDN U7430 ( .A(n6972), .B(n16990), .Z(n6840) );
  AND U7431 ( .A(n6841), .B(n6840), .Z(n6982) );
  XNOR U7432 ( .A(n6981), .B(n6982), .Z(n6983) );
  XOR U7433 ( .A(n6984), .B(n6983), .Z(n7009) );
  XNOR U7434 ( .A(n7010), .B(n7009), .Z(n7011) );
  XNOR U7435 ( .A(n7012), .B(n7011), .Z(n7055) );
  NANDN U7436 ( .A(n6843), .B(n6842), .Z(n6847) );
  NAND U7437 ( .A(n6845), .B(n6844), .Z(n6846) );
  NAND U7438 ( .A(n6847), .B(n6846), .Z(n7000) );
  NANDN U7439 ( .A(n6849), .B(n6848), .Z(n6853) );
  NAND U7440 ( .A(n6851), .B(n6850), .Z(n6852) );
  NAND U7441 ( .A(n6853), .B(n6852), .Z(n6998) );
  OR U7442 ( .A(n6855), .B(n6854), .Z(n6859) );
  NANDN U7443 ( .A(n6857), .B(n6856), .Z(n6858) );
  NAND U7444 ( .A(n6859), .B(n6858), .Z(n6997) );
  XNOR U7445 ( .A(n7000), .B(n6999), .Z(n7056) );
  XNOR U7446 ( .A(n7055), .B(n7056), .Z(n7057) );
  NANDN U7447 ( .A(n6861), .B(n6860), .Z(n6865) );
  OR U7448 ( .A(n6863), .B(n6862), .Z(n6864) );
  AND U7449 ( .A(n6865), .B(n6864), .Z(n7058) );
  XOR U7450 ( .A(n7057), .B(n7058), .Z(n7075) );
  NANDN U7451 ( .A(n6871), .B(n6870), .Z(n6875) );
  NANDN U7452 ( .A(n6873), .B(n6872), .Z(n6874) );
  NAND U7453 ( .A(n6875), .B(n6874), .Z(n7064) );
  NANDN U7454 ( .A(n6881), .B(n6880), .Z(n6885) );
  NAND U7455 ( .A(n6883), .B(n6882), .Z(n6884) );
  NAND U7456 ( .A(n6885), .B(n6884), .Z(n7003) );
  NANDN U7457 ( .A(n6887), .B(n6886), .Z(n6891) );
  NAND U7458 ( .A(n6889), .B(n6888), .Z(n6890) );
  AND U7459 ( .A(n6891), .B(n6890), .Z(n7004) );
  XNOR U7460 ( .A(n7003), .B(n7004), .Z(n7005) );
  XOR U7461 ( .A(n579), .B(a[51]), .Z(n7025) );
  NANDN U7462 ( .A(n7025), .B(n17814), .Z(n6894) );
  NAND U7463 ( .A(n17815), .B(n6892), .Z(n6893) );
  NAND U7464 ( .A(n6894), .B(n6893), .Z(n6989) );
  XNOR U7465 ( .A(b[15]), .B(a[45]), .Z(n7028) );
  OR U7466 ( .A(n7028), .B(n18512), .Z(n6897) );
  NAND U7467 ( .A(n6895), .B(n18513), .Z(n6896) );
  NAND U7468 ( .A(n6897), .B(n6896), .Z(n6987) );
  XOR U7469 ( .A(n582), .B(a[39]), .Z(n7031) );
  NANDN U7470 ( .A(n7031), .B(n19015), .Z(n6900) );
  NAND U7471 ( .A(n19013), .B(n6898), .Z(n6899) );
  NAND U7472 ( .A(n6900), .B(n6899), .Z(n6988) );
  XNOR U7473 ( .A(n6987), .B(n6988), .Z(n6990) );
  XOR U7474 ( .A(n6989), .B(n6990), .Z(n6978) );
  XOR U7475 ( .A(b[11]), .B(n10083), .Z(n7034) );
  OR U7476 ( .A(n7034), .B(n18194), .Z(n6903) );
  NANDN U7477 ( .A(n6901), .B(n18104), .Z(n6902) );
  NAND U7478 ( .A(n6903), .B(n6902), .Z(n6976) );
  XOR U7479 ( .A(n580), .B(a[47]), .Z(n7037) );
  NANDN U7480 ( .A(n7037), .B(n18336), .Z(n6906) );
  NANDN U7481 ( .A(n6904), .B(n18337), .Z(n6905) );
  AND U7482 ( .A(n6906), .B(n6905), .Z(n6975) );
  XNOR U7483 ( .A(n6976), .B(n6975), .Z(n6977) );
  XNOR U7484 ( .A(n6978), .B(n6977), .Z(n6994) );
  NAND U7485 ( .A(n19406), .B(n6907), .Z(n6909) );
  XNOR U7486 ( .A(n584), .B(a[31]), .Z(n7043) );
  NANDN U7487 ( .A(n576), .B(n7043), .Z(n6908) );
  NAND U7488 ( .A(n6909), .B(n6908), .Z(n6951) );
  NANDN U7489 ( .A(n585), .B(a[27]), .Z(n6952) );
  XNOR U7490 ( .A(n6951), .B(n6952), .Z(n6954) );
  NANDN U7491 ( .A(n577), .B(a[59]), .Z(n6910) );
  XOR U7492 ( .A(n17151), .B(n6910), .Z(n6912) );
  NANDN U7493 ( .A(b[0]), .B(a[58]), .Z(n6911) );
  AND U7494 ( .A(n6912), .B(n6911), .Z(n6953) );
  XNOR U7495 ( .A(n6954), .B(n6953), .Z(n6992) );
  XOR U7496 ( .A(b[23]), .B(a[37]), .Z(n7046) );
  NANDN U7497 ( .A(n19127), .B(n7046), .Z(n6915) );
  NAND U7498 ( .A(n6913), .B(n19128), .Z(n6914) );
  NAND U7499 ( .A(n6915), .B(n6914), .Z(n7016) );
  NAND U7500 ( .A(n6916), .B(n17553), .Z(n6918) );
  XNOR U7501 ( .A(b[7]), .B(a[53]), .Z(n7049) );
  NANDN U7502 ( .A(n7049), .B(n17555), .Z(n6917) );
  NAND U7503 ( .A(n6918), .B(n6917), .Z(n7013) );
  XOR U7504 ( .A(b[25]), .B(a[35]), .Z(n7052) );
  NAND U7505 ( .A(n7052), .B(n19240), .Z(n6921) );
  NAND U7506 ( .A(n6919), .B(n19242), .Z(n6920) );
  AND U7507 ( .A(n6921), .B(n6920), .Z(n7014) );
  XNOR U7508 ( .A(n7013), .B(n7014), .Z(n7015) );
  XOR U7509 ( .A(n7016), .B(n7015), .Z(n6991) );
  XOR U7510 ( .A(n6994), .B(n6993), .Z(n7006) );
  XOR U7511 ( .A(n7005), .B(n7006), .Z(n7061) );
  XOR U7512 ( .A(n7062), .B(n7061), .Z(n7063) );
  XNOR U7513 ( .A(n7064), .B(n7063), .Z(n7073) );
  XNOR U7514 ( .A(n7074), .B(n7073), .Z(n7076) );
  XNOR U7515 ( .A(n7075), .B(n7076), .Z(n7070) );
  XOR U7516 ( .A(n7069), .B(n7070), .Z(n6948) );
  NANDN U7517 ( .A(n6923), .B(n6922), .Z(n6927) );
  NANDN U7518 ( .A(n6925), .B(n6924), .Z(n6926) );
  NAND U7519 ( .A(n6927), .B(n6926), .Z(n6946) );
  OR U7520 ( .A(n6929), .B(n6928), .Z(n6933) );
  OR U7521 ( .A(n6931), .B(n6930), .Z(n6932) );
  AND U7522 ( .A(n6933), .B(n6932), .Z(n6945) );
  XNOR U7523 ( .A(n6946), .B(n6945), .Z(n6947) );
  XNOR U7524 ( .A(n6948), .B(n6947), .Z(n6940) );
  XNOR U7525 ( .A(n6939), .B(n6940), .Z(n6941) );
  XNOR U7526 ( .A(n6942), .B(n6941), .Z(n7079) );
  XNOR U7527 ( .A(n7079), .B(sreg[155]), .Z(n7081) );
  NAND U7528 ( .A(n6934), .B(sreg[154]), .Z(n6938) );
  OR U7529 ( .A(n6936), .B(n6935), .Z(n6937) );
  AND U7530 ( .A(n6938), .B(n6937), .Z(n7080) );
  XOR U7531 ( .A(n7081), .B(n7080), .Z(c[155]) );
  NANDN U7532 ( .A(n6940), .B(n6939), .Z(n6944) );
  NAND U7533 ( .A(n6942), .B(n6941), .Z(n6943) );
  NAND U7534 ( .A(n6944), .B(n6943), .Z(n7087) );
  NANDN U7535 ( .A(n6946), .B(n6945), .Z(n6950) );
  NAND U7536 ( .A(n6948), .B(n6947), .Z(n6949) );
  NAND U7537 ( .A(n6950), .B(n6949), .Z(n7085) );
  NANDN U7538 ( .A(n6952), .B(n6951), .Z(n6956) );
  NAND U7539 ( .A(n6954), .B(n6953), .Z(n6955) );
  NAND U7540 ( .A(n6956), .B(n6955), .Z(n7165) );
  NANDN U7541 ( .A(n6957), .B(n18832), .Z(n6959) );
  XOR U7542 ( .A(b[19]), .B(n9080), .Z(n7112) );
  NANDN U7543 ( .A(n7112), .B(n18834), .Z(n6958) );
  NAND U7544 ( .A(n6959), .B(n6958), .Z(n7175) );
  XNOR U7545 ( .A(b[27]), .B(a[34]), .Z(n7115) );
  NANDN U7546 ( .A(n7115), .B(n19336), .Z(n6962) );
  NANDN U7547 ( .A(n6960), .B(n19337), .Z(n6961) );
  NAND U7548 ( .A(n6962), .B(n6961), .Z(n7172) );
  XOR U7549 ( .A(b[5]), .B(a[56]), .Z(n7118) );
  NAND U7550 ( .A(n7118), .B(n17310), .Z(n6965) );
  NANDN U7551 ( .A(n6963), .B(n17311), .Z(n6964) );
  AND U7552 ( .A(n6965), .B(n6964), .Z(n7173) );
  XNOR U7553 ( .A(n7172), .B(n7173), .Z(n7174) );
  XNOR U7554 ( .A(n7175), .B(n7174), .Z(n7163) );
  XOR U7555 ( .A(b[17]), .B(a[44]), .Z(n7121) );
  NAND U7556 ( .A(n7121), .B(n18673), .Z(n6968) );
  NAND U7557 ( .A(n6966), .B(n18674), .Z(n6967) );
  NAND U7558 ( .A(n6968), .B(n6967), .Z(n7139) );
  XOR U7559 ( .A(b[31]), .B(n7336), .Z(n7124) );
  NANDN U7560 ( .A(n7124), .B(n19472), .Z(n6971) );
  NANDN U7561 ( .A(n6969), .B(n19473), .Z(n6970) );
  NAND U7562 ( .A(n6971), .B(n6970), .Z(n7136) );
  OR U7563 ( .A(n6972), .B(n16988), .Z(n6974) );
  XNOR U7564 ( .A(b[3]), .B(a[58]), .Z(n7127) );
  NANDN U7565 ( .A(n7127), .B(n16990), .Z(n6973) );
  AND U7566 ( .A(n6974), .B(n6973), .Z(n7137) );
  XNOR U7567 ( .A(n7136), .B(n7137), .Z(n7138) );
  XOR U7568 ( .A(n7139), .B(n7138), .Z(n7162) );
  XNOR U7569 ( .A(n7163), .B(n7162), .Z(n7164) );
  XNOR U7570 ( .A(n7165), .B(n7164), .Z(n7103) );
  NANDN U7571 ( .A(n6976), .B(n6975), .Z(n6980) );
  NAND U7572 ( .A(n6978), .B(n6977), .Z(n6979) );
  NAND U7573 ( .A(n6980), .B(n6979), .Z(n7154) );
  NANDN U7574 ( .A(n6982), .B(n6981), .Z(n6986) );
  NAND U7575 ( .A(n6984), .B(n6983), .Z(n6985) );
  NAND U7576 ( .A(n6986), .B(n6985), .Z(n7153) );
  XNOR U7577 ( .A(n7153), .B(n7152), .Z(n7155) );
  XOR U7578 ( .A(n7154), .B(n7155), .Z(n7102) );
  XOR U7579 ( .A(n7103), .B(n7102), .Z(n7104) );
  NANDN U7580 ( .A(n6992), .B(n6991), .Z(n6996) );
  NAND U7581 ( .A(n6994), .B(n6993), .Z(n6995) );
  NAND U7582 ( .A(n6996), .B(n6995), .Z(n7105) );
  XNOR U7583 ( .A(n7104), .B(n7105), .Z(n7216) );
  OR U7584 ( .A(n6998), .B(n6997), .Z(n7002) );
  NAND U7585 ( .A(n7000), .B(n6999), .Z(n7001) );
  NAND U7586 ( .A(n7002), .B(n7001), .Z(n7215) );
  NANDN U7587 ( .A(n7004), .B(n7003), .Z(n7008) );
  NAND U7588 ( .A(n7006), .B(n7005), .Z(n7007) );
  NAND U7589 ( .A(n7008), .B(n7007), .Z(n7098) );
  NANDN U7590 ( .A(n7014), .B(n7013), .Z(n7018) );
  NAND U7591 ( .A(n7016), .B(n7015), .Z(n7017) );
  NAND U7592 ( .A(n7018), .B(n7017), .Z(n7156) );
  NANDN U7593 ( .A(n7020), .B(n7019), .Z(n7024) );
  NAND U7594 ( .A(n7022), .B(n7021), .Z(n7023) );
  AND U7595 ( .A(n7024), .B(n7023), .Z(n7157) );
  XNOR U7596 ( .A(n7156), .B(n7157), .Z(n7158) );
  XNOR U7597 ( .A(b[9]), .B(a[52]), .Z(n7178) );
  NANDN U7598 ( .A(n7178), .B(n17814), .Z(n7027) );
  NANDN U7599 ( .A(n7025), .B(n17815), .Z(n7026) );
  NAND U7600 ( .A(n7027), .B(n7026), .Z(n7144) );
  XNOR U7601 ( .A(b[15]), .B(a[46]), .Z(n7181) );
  OR U7602 ( .A(n7181), .B(n18512), .Z(n7030) );
  NANDN U7603 ( .A(n7028), .B(n18513), .Z(n7029) );
  NAND U7604 ( .A(n7030), .B(n7029), .Z(n7142) );
  XNOR U7605 ( .A(b[21]), .B(a[40]), .Z(n7184) );
  NANDN U7606 ( .A(n7184), .B(n19015), .Z(n7033) );
  NANDN U7607 ( .A(n7031), .B(n19013), .Z(n7032) );
  NAND U7608 ( .A(n7033), .B(n7032), .Z(n7143) );
  XNOR U7609 ( .A(n7142), .B(n7143), .Z(n7145) );
  XOR U7610 ( .A(n7144), .B(n7145), .Z(n7133) );
  XNOR U7611 ( .A(b[11]), .B(a[50]), .Z(n7187) );
  OR U7612 ( .A(n7187), .B(n18194), .Z(n7036) );
  NANDN U7613 ( .A(n7034), .B(n18104), .Z(n7035) );
  NAND U7614 ( .A(n7036), .B(n7035), .Z(n7131) );
  XOR U7615 ( .A(n580), .B(a[48]), .Z(n7190) );
  NANDN U7616 ( .A(n7190), .B(n18336), .Z(n7039) );
  NANDN U7617 ( .A(n7037), .B(n18337), .Z(n7038) );
  AND U7618 ( .A(n7039), .B(n7038), .Z(n7130) );
  XNOR U7619 ( .A(n7131), .B(n7130), .Z(n7132) );
  XNOR U7620 ( .A(n7133), .B(n7132), .Z(n7149) );
  NANDN U7621 ( .A(n577), .B(a[60]), .Z(n7040) );
  XOR U7622 ( .A(n17151), .B(n7040), .Z(n7042) );
  NANDN U7623 ( .A(b[0]), .B(a[59]), .Z(n7041) );
  AND U7624 ( .A(n7042), .B(n7041), .Z(n7108) );
  NAND U7625 ( .A(n19406), .B(n7043), .Z(n7045) );
  XNOR U7626 ( .A(n584), .B(a[32]), .Z(n7193) );
  NANDN U7627 ( .A(n576), .B(n7193), .Z(n7044) );
  NAND U7628 ( .A(n7045), .B(n7044), .Z(n7106) );
  NANDN U7629 ( .A(n585), .B(a[28]), .Z(n7107) );
  XNOR U7630 ( .A(n7106), .B(n7107), .Z(n7109) );
  XNOR U7631 ( .A(n7108), .B(n7109), .Z(n7147) );
  XNOR U7632 ( .A(b[23]), .B(a[38]), .Z(n7199) );
  OR U7633 ( .A(n7199), .B(n19127), .Z(n7048) );
  NAND U7634 ( .A(n7046), .B(n19128), .Z(n7047) );
  NAND U7635 ( .A(n7048), .B(n7047), .Z(n7169) );
  NANDN U7636 ( .A(n7049), .B(n17553), .Z(n7051) );
  XOR U7637 ( .A(b[7]), .B(a[54]), .Z(n7202) );
  NAND U7638 ( .A(n7202), .B(n17555), .Z(n7050) );
  NAND U7639 ( .A(n7051), .B(n7050), .Z(n7166) );
  XOR U7640 ( .A(b[25]), .B(a[36]), .Z(n7205) );
  NAND U7641 ( .A(n7205), .B(n19240), .Z(n7054) );
  NAND U7642 ( .A(n7052), .B(n19242), .Z(n7053) );
  AND U7643 ( .A(n7054), .B(n7053), .Z(n7167) );
  XNOR U7644 ( .A(n7166), .B(n7167), .Z(n7168) );
  XOR U7645 ( .A(n7169), .B(n7168), .Z(n7146) );
  XOR U7646 ( .A(n7149), .B(n7148), .Z(n7159) );
  XOR U7647 ( .A(n7158), .B(n7159), .Z(n7096) );
  XNOR U7648 ( .A(n7097), .B(n7096), .Z(n7099) );
  XNOR U7649 ( .A(n7098), .B(n7099), .Z(n7214) );
  XOR U7650 ( .A(n7215), .B(n7214), .Z(n7217) );
  NANDN U7651 ( .A(n7056), .B(n7055), .Z(n7060) );
  NAND U7652 ( .A(n7058), .B(n7057), .Z(n7059) );
  NAND U7653 ( .A(n7060), .B(n7059), .Z(n7208) );
  NAND U7654 ( .A(n7062), .B(n7061), .Z(n7066) );
  NAND U7655 ( .A(n7064), .B(n7063), .Z(n7065) );
  NAND U7656 ( .A(n7066), .B(n7065), .Z(n7209) );
  XNOR U7657 ( .A(n7208), .B(n7209), .Z(n7210) );
  XOR U7658 ( .A(n7211), .B(n7210), .Z(n7092) );
  NANDN U7659 ( .A(n7068), .B(n7067), .Z(n7072) );
  NANDN U7660 ( .A(n7070), .B(n7069), .Z(n7071) );
  NAND U7661 ( .A(n7072), .B(n7071), .Z(n7091) );
  OR U7662 ( .A(n7074), .B(n7073), .Z(n7078) );
  OR U7663 ( .A(n7076), .B(n7075), .Z(n7077) );
  AND U7664 ( .A(n7078), .B(n7077), .Z(n7090) );
  XNOR U7665 ( .A(n7091), .B(n7090), .Z(n7093) );
  XOR U7666 ( .A(n7092), .B(n7093), .Z(n7084) );
  XOR U7667 ( .A(n7085), .B(n7084), .Z(n7086) );
  XNOR U7668 ( .A(n7087), .B(n7086), .Z(n7220) );
  XNOR U7669 ( .A(n7220), .B(sreg[156]), .Z(n7222) );
  NAND U7670 ( .A(n7079), .B(sreg[155]), .Z(n7083) );
  OR U7671 ( .A(n7081), .B(n7080), .Z(n7082) );
  AND U7672 ( .A(n7083), .B(n7082), .Z(n7221) );
  XOR U7673 ( .A(n7222), .B(n7221), .Z(c[156]) );
  NAND U7674 ( .A(n7085), .B(n7084), .Z(n7089) );
  NAND U7675 ( .A(n7087), .B(n7086), .Z(n7088) );
  NAND U7676 ( .A(n7089), .B(n7088), .Z(n7228) );
  NANDN U7677 ( .A(n7091), .B(n7090), .Z(n7095) );
  NAND U7678 ( .A(n7093), .B(n7092), .Z(n7094) );
  NAND U7679 ( .A(n7095), .B(n7094), .Z(n7225) );
  NAND U7680 ( .A(n7097), .B(n7096), .Z(n7101) );
  NANDN U7681 ( .A(n7099), .B(n7098), .Z(n7100) );
  NAND U7682 ( .A(n7101), .B(n7100), .Z(n7352) );
  XNOR U7683 ( .A(n7352), .B(n7353), .Z(n7354) );
  NANDN U7684 ( .A(n7107), .B(n7106), .Z(n7111) );
  NAND U7685 ( .A(n7109), .B(n7108), .Z(n7110) );
  NAND U7686 ( .A(n7111), .B(n7110), .Z(n7308) );
  NANDN U7687 ( .A(n7112), .B(n18832), .Z(n7114) );
  XNOR U7688 ( .A(b[19]), .B(a[43]), .Z(n7253) );
  NANDN U7689 ( .A(n7253), .B(n18834), .Z(n7113) );
  NAND U7690 ( .A(n7114), .B(n7113), .Z(n7318) );
  XNOR U7691 ( .A(b[27]), .B(a[35]), .Z(n7256) );
  NANDN U7692 ( .A(n7256), .B(n19336), .Z(n7117) );
  NANDN U7693 ( .A(n7115), .B(n19337), .Z(n7116) );
  NAND U7694 ( .A(n7117), .B(n7116), .Z(n7315) );
  XOR U7695 ( .A(b[5]), .B(a[57]), .Z(n7259) );
  NAND U7696 ( .A(n7259), .B(n17310), .Z(n7120) );
  NAND U7697 ( .A(n7118), .B(n17311), .Z(n7119) );
  AND U7698 ( .A(n7120), .B(n7119), .Z(n7316) );
  XNOR U7699 ( .A(n7315), .B(n7316), .Z(n7317) );
  XNOR U7700 ( .A(n7318), .B(n7317), .Z(n7306) );
  XOR U7701 ( .A(b[17]), .B(a[45]), .Z(n7262) );
  NAND U7702 ( .A(n7262), .B(n18673), .Z(n7123) );
  NAND U7703 ( .A(n7121), .B(n18674), .Z(n7122) );
  NAND U7704 ( .A(n7123), .B(n7122), .Z(n7280) );
  XNOR U7705 ( .A(b[31]), .B(a[31]), .Z(n7265) );
  NANDN U7706 ( .A(n7265), .B(n19472), .Z(n7126) );
  NANDN U7707 ( .A(n7124), .B(n19473), .Z(n7125) );
  NAND U7708 ( .A(n7126), .B(n7125), .Z(n7277) );
  OR U7709 ( .A(n7127), .B(n16988), .Z(n7129) );
  XNOR U7710 ( .A(b[3]), .B(a[59]), .Z(n7268) );
  NANDN U7711 ( .A(n7268), .B(n16990), .Z(n7128) );
  AND U7712 ( .A(n7129), .B(n7128), .Z(n7278) );
  XNOR U7713 ( .A(n7277), .B(n7278), .Z(n7279) );
  XOR U7714 ( .A(n7280), .B(n7279), .Z(n7305) );
  XNOR U7715 ( .A(n7306), .B(n7305), .Z(n7307) );
  XNOR U7716 ( .A(n7308), .B(n7307), .Z(n7244) );
  NANDN U7717 ( .A(n7131), .B(n7130), .Z(n7135) );
  NAND U7718 ( .A(n7133), .B(n7132), .Z(n7134) );
  NAND U7719 ( .A(n7135), .B(n7134), .Z(n7297) );
  NANDN U7720 ( .A(n7137), .B(n7136), .Z(n7141) );
  NAND U7721 ( .A(n7139), .B(n7138), .Z(n7140) );
  NAND U7722 ( .A(n7141), .B(n7140), .Z(n7296) );
  XNOR U7723 ( .A(n7296), .B(n7295), .Z(n7298) );
  XOR U7724 ( .A(n7297), .B(n7298), .Z(n7243) );
  XOR U7725 ( .A(n7244), .B(n7243), .Z(n7245) );
  NANDN U7726 ( .A(n7147), .B(n7146), .Z(n7151) );
  NAND U7727 ( .A(n7149), .B(n7148), .Z(n7150) );
  AND U7728 ( .A(n7151), .B(n7150), .Z(n7246) );
  XOR U7729 ( .A(n7245), .B(n7246), .Z(n7360) );
  NANDN U7730 ( .A(n7157), .B(n7156), .Z(n7161) );
  NAND U7731 ( .A(n7159), .B(n7158), .Z(n7160) );
  NAND U7732 ( .A(n7161), .B(n7160), .Z(n7240) );
  NANDN U7733 ( .A(n7167), .B(n7166), .Z(n7171) );
  NAND U7734 ( .A(n7169), .B(n7168), .Z(n7170) );
  NAND U7735 ( .A(n7171), .B(n7170), .Z(n7299) );
  NANDN U7736 ( .A(n7173), .B(n7172), .Z(n7177) );
  NAND U7737 ( .A(n7175), .B(n7174), .Z(n7176) );
  AND U7738 ( .A(n7177), .B(n7176), .Z(n7300) );
  XNOR U7739 ( .A(n7299), .B(n7300), .Z(n7301) );
  XOR U7740 ( .A(n579), .B(n10660), .Z(n7327) );
  NAND U7741 ( .A(n17814), .B(n7327), .Z(n7180) );
  NANDN U7742 ( .A(n7178), .B(n17815), .Z(n7179) );
  NAND U7743 ( .A(n7180), .B(n7179), .Z(n7285) );
  NANDN U7744 ( .A(n7181), .B(n18513), .Z(n7183) );
  XOR U7745 ( .A(b[15]), .B(a[47]), .Z(n7324) );
  NANDN U7746 ( .A(n18512), .B(n7324), .Z(n7182) );
  AND U7747 ( .A(n7183), .B(n7182), .Z(n7283) );
  NANDN U7748 ( .A(n7184), .B(n19013), .Z(n7186) );
  XOR U7749 ( .A(n582), .B(n8930), .Z(n7321) );
  NAND U7750 ( .A(n7321), .B(n19015), .Z(n7185) );
  AND U7751 ( .A(n7186), .B(n7185), .Z(n7284) );
  XOR U7752 ( .A(n7285), .B(n7286), .Z(n7274) );
  XNOR U7753 ( .A(b[11]), .B(a[51]), .Z(n7330) );
  OR U7754 ( .A(n7330), .B(n18194), .Z(n7189) );
  NANDN U7755 ( .A(n7187), .B(n18104), .Z(n7188) );
  NAND U7756 ( .A(n7189), .B(n7188), .Z(n7272) );
  XOR U7757 ( .A(n580), .B(a[49]), .Z(n7333) );
  NANDN U7758 ( .A(n7333), .B(n18336), .Z(n7192) );
  NANDN U7759 ( .A(n7190), .B(n18337), .Z(n7191) );
  AND U7760 ( .A(n7192), .B(n7191), .Z(n7271) );
  XNOR U7761 ( .A(n7272), .B(n7271), .Z(n7273) );
  XOR U7762 ( .A(n7274), .B(n7273), .Z(n7291) );
  NAND U7763 ( .A(n19406), .B(n7193), .Z(n7195) );
  XNOR U7764 ( .A(b[29]), .B(a[33]), .Z(n7337) );
  OR U7765 ( .A(n7337), .B(n576), .Z(n7194) );
  NAND U7766 ( .A(n7195), .B(n7194), .Z(n7247) );
  NANDN U7767 ( .A(n585), .B(a[29]), .Z(n7248) );
  XNOR U7768 ( .A(n7247), .B(n7248), .Z(n7250) );
  NANDN U7769 ( .A(n577), .B(a[61]), .Z(n7196) );
  XOR U7770 ( .A(n17151), .B(n7196), .Z(n7198) );
  NANDN U7771 ( .A(b[0]), .B(a[60]), .Z(n7197) );
  AND U7772 ( .A(n7198), .B(n7197), .Z(n7249) );
  XOR U7773 ( .A(n7250), .B(n7249), .Z(n7289) );
  XOR U7774 ( .A(b[23]), .B(a[39]), .Z(n7343) );
  NANDN U7775 ( .A(n19127), .B(n7343), .Z(n7201) );
  NANDN U7776 ( .A(n7199), .B(n19128), .Z(n7200) );
  NAND U7777 ( .A(n7201), .B(n7200), .Z(n7312) );
  NAND U7778 ( .A(n7202), .B(n17553), .Z(n7204) );
  XNOR U7779 ( .A(b[7]), .B(a[55]), .Z(n7346) );
  NANDN U7780 ( .A(n7346), .B(n17555), .Z(n7203) );
  NAND U7781 ( .A(n7204), .B(n7203), .Z(n7309) );
  XOR U7782 ( .A(b[25]), .B(a[37]), .Z(n7349) );
  NAND U7783 ( .A(n7349), .B(n19240), .Z(n7207) );
  NAND U7784 ( .A(n7205), .B(n19242), .Z(n7206) );
  AND U7785 ( .A(n7207), .B(n7206), .Z(n7310) );
  XNOR U7786 ( .A(n7309), .B(n7310), .Z(n7311) );
  XNOR U7787 ( .A(n7312), .B(n7311), .Z(n7290) );
  XOR U7788 ( .A(n7289), .B(n7290), .Z(n7292) );
  XNOR U7789 ( .A(n7291), .B(n7292), .Z(n7302) );
  XOR U7790 ( .A(n7301), .B(n7302), .Z(n7238) );
  XNOR U7791 ( .A(n7237), .B(n7238), .Z(n7239) );
  XNOR U7792 ( .A(n7240), .B(n7239), .Z(n7358) );
  XNOR U7793 ( .A(n7359), .B(n7358), .Z(n7361) );
  XNOR U7794 ( .A(n7360), .B(n7361), .Z(n7355) );
  XOR U7795 ( .A(n7354), .B(n7355), .Z(n7234) );
  NANDN U7796 ( .A(n7209), .B(n7208), .Z(n7213) );
  NAND U7797 ( .A(n7211), .B(n7210), .Z(n7212) );
  NAND U7798 ( .A(n7213), .B(n7212), .Z(n7231) );
  NANDN U7799 ( .A(n7215), .B(n7214), .Z(n7219) );
  OR U7800 ( .A(n7217), .B(n7216), .Z(n7218) );
  NAND U7801 ( .A(n7219), .B(n7218), .Z(n7232) );
  XNOR U7802 ( .A(n7231), .B(n7232), .Z(n7233) );
  XNOR U7803 ( .A(n7234), .B(n7233), .Z(n7226) );
  XNOR U7804 ( .A(n7225), .B(n7226), .Z(n7227) );
  XNOR U7805 ( .A(n7228), .B(n7227), .Z(n7364) );
  XNOR U7806 ( .A(n7364), .B(sreg[157]), .Z(n7366) );
  NAND U7807 ( .A(n7220), .B(sreg[156]), .Z(n7224) );
  OR U7808 ( .A(n7222), .B(n7221), .Z(n7223) );
  AND U7809 ( .A(n7224), .B(n7223), .Z(n7365) );
  XOR U7810 ( .A(n7366), .B(n7365), .Z(c[157]) );
  NANDN U7811 ( .A(n7226), .B(n7225), .Z(n7230) );
  NAND U7812 ( .A(n7228), .B(n7227), .Z(n7229) );
  NAND U7813 ( .A(n7230), .B(n7229), .Z(n7372) );
  NANDN U7814 ( .A(n7232), .B(n7231), .Z(n7236) );
  NAND U7815 ( .A(n7234), .B(n7233), .Z(n7235) );
  NAND U7816 ( .A(n7236), .B(n7235), .Z(n7369) );
  NANDN U7817 ( .A(n7238), .B(n7237), .Z(n7242) );
  NAND U7818 ( .A(n7240), .B(n7239), .Z(n7241) );
  NAND U7819 ( .A(n7242), .B(n7241), .Z(n7381) );
  XNOR U7820 ( .A(n7381), .B(n7382), .Z(n7383) );
  NANDN U7821 ( .A(n7248), .B(n7247), .Z(n7252) );
  NAND U7822 ( .A(n7250), .B(n7249), .Z(n7251) );
  NAND U7823 ( .A(n7252), .B(n7251), .Z(n7454) );
  NANDN U7824 ( .A(n7253), .B(n18832), .Z(n7255) );
  XNOR U7825 ( .A(b[19]), .B(a[44]), .Z(n7399) );
  NANDN U7826 ( .A(n7399), .B(n18834), .Z(n7254) );
  NAND U7827 ( .A(n7255), .B(n7254), .Z(n7488) );
  XNOR U7828 ( .A(b[27]), .B(a[36]), .Z(n7402) );
  NANDN U7829 ( .A(n7402), .B(n19336), .Z(n7258) );
  NANDN U7830 ( .A(n7256), .B(n19337), .Z(n7257) );
  NAND U7831 ( .A(n7258), .B(n7257), .Z(n7485) );
  XOR U7832 ( .A(b[5]), .B(a[58]), .Z(n7405) );
  NAND U7833 ( .A(n7405), .B(n17310), .Z(n7261) );
  NAND U7834 ( .A(n7259), .B(n17311), .Z(n7260) );
  AND U7835 ( .A(n7261), .B(n7260), .Z(n7486) );
  XNOR U7836 ( .A(n7485), .B(n7486), .Z(n7487) );
  XNOR U7837 ( .A(n7488), .B(n7487), .Z(n7452) );
  XOR U7838 ( .A(b[17]), .B(a[46]), .Z(n7408) );
  NAND U7839 ( .A(n7408), .B(n18673), .Z(n7264) );
  NAND U7840 ( .A(n7262), .B(n18674), .Z(n7263) );
  NAND U7841 ( .A(n7264), .B(n7263), .Z(n7426) );
  XNOR U7842 ( .A(b[31]), .B(a[32]), .Z(n7411) );
  NANDN U7843 ( .A(n7411), .B(n19472), .Z(n7267) );
  NANDN U7844 ( .A(n7265), .B(n19473), .Z(n7266) );
  NAND U7845 ( .A(n7267), .B(n7266), .Z(n7423) );
  OR U7846 ( .A(n7268), .B(n16988), .Z(n7270) );
  XNOR U7847 ( .A(b[3]), .B(a[60]), .Z(n7414) );
  NANDN U7848 ( .A(n7414), .B(n16990), .Z(n7269) );
  AND U7849 ( .A(n7270), .B(n7269), .Z(n7424) );
  XNOR U7850 ( .A(n7423), .B(n7424), .Z(n7425) );
  XOR U7851 ( .A(n7426), .B(n7425), .Z(n7451) );
  XNOR U7852 ( .A(n7452), .B(n7451), .Z(n7453) );
  XNOR U7853 ( .A(n7454), .B(n7453), .Z(n7497) );
  NANDN U7854 ( .A(n7272), .B(n7271), .Z(n7276) );
  NAND U7855 ( .A(n7274), .B(n7273), .Z(n7275) );
  NAND U7856 ( .A(n7276), .B(n7275), .Z(n7442) );
  NANDN U7857 ( .A(n7278), .B(n7277), .Z(n7282) );
  NAND U7858 ( .A(n7280), .B(n7279), .Z(n7281) );
  NAND U7859 ( .A(n7282), .B(n7281), .Z(n7440) );
  OR U7860 ( .A(n7284), .B(n7283), .Z(n7288) );
  NANDN U7861 ( .A(n7286), .B(n7285), .Z(n7287) );
  NAND U7862 ( .A(n7288), .B(n7287), .Z(n7439) );
  XNOR U7863 ( .A(n7442), .B(n7441), .Z(n7498) );
  XNOR U7864 ( .A(n7497), .B(n7498), .Z(n7499) );
  NANDN U7865 ( .A(n7290), .B(n7289), .Z(n7294) );
  OR U7866 ( .A(n7292), .B(n7291), .Z(n7293) );
  AND U7867 ( .A(n7294), .B(n7293), .Z(n7500) );
  XOR U7868 ( .A(n7499), .B(n7500), .Z(n7389) );
  NANDN U7869 ( .A(n7300), .B(n7299), .Z(n7304) );
  NANDN U7870 ( .A(n7302), .B(n7301), .Z(n7303) );
  NAND U7871 ( .A(n7304), .B(n7303), .Z(n7506) );
  NANDN U7872 ( .A(n7310), .B(n7309), .Z(n7314) );
  NAND U7873 ( .A(n7312), .B(n7311), .Z(n7313) );
  NAND U7874 ( .A(n7314), .B(n7313), .Z(n7445) );
  NANDN U7875 ( .A(n7316), .B(n7315), .Z(n7320) );
  NAND U7876 ( .A(n7318), .B(n7317), .Z(n7319) );
  AND U7877 ( .A(n7320), .B(n7319), .Z(n7446) );
  XNOR U7878 ( .A(n7445), .B(n7446), .Z(n7447) );
  XOR U7879 ( .A(n582), .B(a[42]), .Z(n7461) );
  NANDN U7880 ( .A(n7461), .B(n19015), .Z(n7323) );
  NAND U7881 ( .A(n19013), .B(n7321), .Z(n7322) );
  NAND U7882 ( .A(n7323), .B(n7322), .Z(n7435) );
  NAND U7883 ( .A(n7324), .B(n18513), .Z(n7326) );
  XOR U7884 ( .A(b[15]), .B(a[48]), .Z(n7458) );
  NANDN U7885 ( .A(n18512), .B(n7458), .Z(n7325) );
  AND U7886 ( .A(n7326), .B(n7325), .Z(n7436) );
  XNOR U7887 ( .A(n7435), .B(n7436), .Z(n7438) );
  XOR U7888 ( .A(n579), .B(a[54]), .Z(n7455) );
  NANDN U7889 ( .A(n7455), .B(n17814), .Z(n7329) );
  NAND U7890 ( .A(n17815), .B(n7327), .Z(n7328) );
  NAND U7891 ( .A(n7329), .B(n7328), .Z(n7437) );
  XNOR U7892 ( .A(n7438), .B(n7437), .Z(n7431) );
  XNOR U7893 ( .A(b[11]), .B(a[52]), .Z(n7464) );
  OR U7894 ( .A(n7464), .B(n18194), .Z(n7332) );
  NANDN U7895 ( .A(n7330), .B(n18104), .Z(n7331) );
  NAND U7896 ( .A(n7332), .B(n7331), .Z(n7430) );
  XOR U7897 ( .A(n580), .B(a[50]), .Z(n7467) );
  NANDN U7898 ( .A(n7467), .B(n18336), .Z(n7335) );
  NANDN U7899 ( .A(n7333), .B(n18337), .Z(n7334) );
  NAND U7900 ( .A(n7335), .B(n7334), .Z(n7429) );
  XNOR U7901 ( .A(n7430), .B(n7429), .Z(n7432) );
  XNOR U7902 ( .A(n7431), .B(n7432), .Z(n7420) );
  ANDN U7903 ( .B(b[31]), .A(n7336), .Z(n7393) );
  NANDN U7904 ( .A(n7337), .B(n19406), .Z(n7339) );
  XNOR U7905 ( .A(n584), .B(a[34]), .Z(n7473) );
  NANDN U7906 ( .A(n576), .B(n7473), .Z(n7338) );
  NAND U7907 ( .A(n7339), .B(n7338), .Z(n7394) );
  XOR U7908 ( .A(n7393), .B(n7394), .Z(n7395) );
  NANDN U7909 ( .A(n577), .B(a[62]), .Z(n7340) );
  XOR U7910 ( .A(n17151), .B(n7340), .Z(n7342) );
  NANDN U7911 ( .A(b[0]), .B(a[61]), .Z(n7341) );
  AND U7912 ( .A(n7342), .B(n7341), .Z(n7396) );
  XNOR U7913 ( .A(n7395), .B(n7396), .Z(n7417) );
  XOR U7914 ( .A(b[23]), .B(a[40]), .Z(n7476) );
  NANDN U7915 ( .A(n19127), .B(n7476), .Z(n7345) );
  NAND U7916 ( .A(n7343), .B(n19128), .Z(n7344) );
  NAND U7917 ( .A(n7345), .B(n7344), .Z(n7494) );
  NANDN U7918 ( .A(n7346), .B(n17553), .Z(n7348) );
  XOR U7919 ( .A(b[7]), .B(a[56]), .Z(n7479) );
  NAND U7920 ( .A(n7479), .B(n17555), .Z(n7347) );
  NAND U7921 ( .A(n7348), .B(n7347), .Z(n7491) );
  XNOR U7922 ( .A(b[25]), .B(a[38]), .Z(n7482) );
  NANDN U7923 ( .A(n7482), .B(n19240), .Z(n7351) );
  NAND U7924 ( .A(n7349), .B(n19242), .Z(n7350) );
  AND U7925 ( .A(n7351), .B(n7350), .Z(n7492) );
  XNOR U7926 ( .A(n7491), .B(n7492), .Z(n7493) );
  XNOR U7927 ( .A(n7494), .B(n7493), .Z(n7418) );
  XOR U7928 ( .A(n7420), .B(n7419), .Z(n7448) );
  XNOR U7929 ( .A(n7447), .B(n7448), .Z(n7503) );
  XOR U7930 ( .A(n7504), .B(n7503), .Z(n7505) );
  XNOR U7931 ( .A(n7506), .B(n7505), .Z(n7387) );
  XNOR U7932 ( .A(n7388), .B(n7387), .Z(n7390) );
  XNOR U7933 ( .A(n7389), .B(n7390), .Z(n7384) );
  XOR U7934 ( .A(n7383), .B(n7384), .Z(n7378) );
  NANDN U7935 ( .A(n7353), .B(n7352), .Z(n7357) );
  NANDN U7936 ( .A(n7355), .B(n7354), .Z(n7356) );
  NAND U7937 ( .A(n7357), .B(n7356), .Z(n7376) );
  OR U7938 ( .A(n7359), .B(n7358), .Z(n7363) );
  OR U7939 ( .A(n7361), .B(n7360), .Z(n7362) );
  AND U7940 ( .A(n7363), .B(n7362), .Z(n7375) );
  XNOR U7941 ( .A(n7376), .B(n7375), .Z(n7377) );
  XNOR U7942 ( .A(n7378), .B(n7377), .Z(n7370) );
  XNOR U7943 ( .A(n7369), .B(n7370), .Z(n7371) );
  XNOR U7944 ( .A(n7372), .B(n7371), .Z(n7509) );
  XNOR U7945 ( .A(n7509), .B(sreg[158]), .Z(n7511) );
  NAND U7946 ( .A(n7364), .B(sreg[157]), .Z(n7368) );
  OR U7947 ( .A(n7366), .B(n7365), .Z(n7367) );
  AND U7948 ( .A(n7368), .B(n7367), .Z(n7510) );
  XOR U7949 ( .A(n7511), .B(n7510), .Z(c[158]) );
  NANDN U7950 ( .A(n7370), .B(n7369), .Z(n7374) );
  NAND U7951 ( .A(n7372), .B(n7371), .Z(n7373) );
  NAND U7952 ( .A(n7374), .B(n7373), .Z(n7517) );
  NANDN U7953 ( .A(n7376), .B(n7375), .Z(n7380) );
  NAND U7954 ( .A(n7378), .B(n7377), .Z(n7379) );
  NAND U7955 ( .A(n7380), .B(n7379), .Z(n7515) );
  NANDN U7956 ( .A(n7382), .B(n7381), .Z(n7386) );
  NANDN U7957 ( .A(n7384), .B(n7383), .Z(n7385) );
  NAND U7958 ( .A(n7386), .B(n7385), .Z(n7521) );
  OR U7959 ( .A(n7388), .B(n7387), .Z(n7392) );
  OR U7960 ( .A(n7390), .B(n7389), .Z(n7391) );
  AND U7961 ( .A(n7392), .B(n7391), .Z(n7520) );
  XNOR U7962 ( .A(n7521), .B(n7520), .Z(n7522) );
  OR U7963 ( .A(n7394), .B(n7393), .Z(n7398) );
  NANDN U7964 ( .A(n7396), .B(n7395), .Z(n7397) );
  NAND U7965 ( .A(n7398), .B(n7397), .Z(n7584) );
  NANDN U7966 ( .A(n7399), .B(n18832), .Z(n7401) );
  XNOR U7967 ( .A(b[19]), .B(a[45]), .Z(n7532) );
  NANDN U7968 ( .A(n7532), .B(n18834), .Z(n7400) );
  NAND U7969 ( .A(n7401), .B(n7400), .Z(n7621) );
  XNOR U7970 ( .A(b[27]), .B(a[37]), .Z(n7535) );
  NANDN U7971 ( .A(n7535), .B(n19336), .Z(n7404) );
  NANDN U7972 ( .A(n7402), .B(n19337), .Z(n7403) );
  NAND U7973 ( .A(n7404), .B(n7403), .Z(n7618) );
  XOR U7974 ( .A(b[5]), .B(a[59]), .Z(n7538) );
  NAND U7975 ( .A(n7538), .B(n17310), .Z(n7407) );
  NAND U7976 ( .A(n7405), .B(n17311), .Z(n7406) );
  AND U7977 ( .A(n7407), .B(n7406), .Z(n7619) );
  XNOR U7978 ( .A(n7618), .B(n7619), .Z(n7620) );
  XNOR U7979 ( .A(n7621), .B(n7620), .Z(n7583) );
  XOR U7980 ( .A(b[17]), .B(a[47]), .Z(n7541) );
  NAND U7981 ( .A(n7541), .B(n18673), .Z(n7410) );
  NAND U7982 ( .A(n7408), .B(n18674), .Z(n7409) );
  NAND U7983 ( .A(n7410), .B(n7409), .Z(n7559) );
  XNOR U7984 ( .A(b[31]), .B(a[33]), .Z(n7544) );
  NANDN U7985 ( .A(n7544), .B(n19472), .Z(n7413) );
  NANDN U7986 ( .A(n7411), .B(n19473), .Z(n7412) );
  NAND U7987 ( .A(n7413), .B(n7412), .Z(n7556) );
  OR U7988 ( .A(n7414), .B(n16988), .Z(n7416) );
  XNOR U7989 ( .A(b[3]), .B(a[61]), .Z(n7547) );
  NANDN U7990 ( .A(n7547), .B(n16990), .Z(n7415) );
  AND U7991 ( .A(n7416), .B(n7415), .Z(n7557) );
  XNOR U7992 ( .A(n7556), .B(n7557), .Z(n7558) );
  XOR U7993 ( .A(n7559), .B(n7558), .Z(n7582) );
  XOR U7994 ( .A(n7583), .B(n7582), .Z(n7585) );
  XNOR U7995 ( .A(n7584), .B(n7585), .Z(n7636) );
  OR U7996 ( .A(n7418), .B(n7417), .Z(n7422) );
  NANDN U7997 ( .A(n7420), .B(n7419), .Z(n7421) );
  NAND U7998 ( .A(n7422), .B(n7421), .Z(n7637) );
  XNOR U7999 ( .A(n7636), .B(n7637), .Z(n7638) );
  NANDN U8000 ( .A(n7424), .B(n7423), .Z(n7428) );
  NAND U8001 ( .A(n7426), .B(n7425), .Z(n7427) );
  NAND U8002 ( .A(n7428), .B(n7427), .Z(n7575) );
  OR U8003 ( .A(n7430), .B(n7429), .Z(n7434) );
  NANDN U8004 ( .A(n7432), .B(n7431), .Z(n7433) );
  NAND U8005 ( .A(n7434), .B(n7433), .Z(n7573) );
  XNOR U8006 ( .A(n7573), .B(n7572), .Z(n7574) );
  XOR U8007 ( .A(n7575), .B(n7574), .Z(n7639) );
  XOR U8008 ( .A(n7638), .B(n7639), .Z(n7651) );
  OR U8009 ( .A(n7440), .B(n7439), .Z(n7444) );
  NAND U8010 ( .A(n7442), .B(n7441), .Z(n7443) );
  NAND U8011 ( .A(n7444), .B(n7443), .Z(n7649) );
  NANDN U8012 ( .A(n7446), .B(n7445), .Z(n7450) );
  NANDN U8013 ( .A(n7448), .B(n7447), .Z(n7449) );
  NAND U8014 ( .A(n7450), .B(n7449), .Z(n7633) );
  XOR U8015 ( .A(n579), .B(a[55]), .Z(n7594) );
  NANDN U8016 ( .A(n7594), .B(n17814), .Z(n7457) );
  NANDN U8017 ( .A(n7455), .B(n17815), .Z(n7456) );
  NAND U8018 ( .A(n7457), .B(n7456), .Z(n7564) );
  XNOR U8019 ( .A(b[15]), .B(a[49]), .Z(n7591) );
  OR U8020 ( .A(n7591), .B(n18512), .Z(n7460) );
  NAND U8021 ( .A(n7458), .B(n18513), .Z(n7459) );
  NAND U8022 ( .A(n7460), .B(n7459), .Z(n7562) );
  XOR U8023 ( .A(n582), .B(a[43]), .Z(n7588) );
  NANDN U8024 ( .A(n7588), .B(n19015), .Z(n7463) );
  NANDN U8025 ( .A(n7461), .B(n19013), .Z(n7462) );
  NAND U8026 ( .A(n7463), .B(n7462), .Z(n7563) );
  XNOR U8027 ( .A(n7562), .B(n7563), .Z(n7565) );
  XOR U8028 ( .A(n7564), .B(n7565), .Z(n7553) );
  XOR U8029 ( .A(b[11]), .B(n10660), .Z(n7597) );
  OR U8030 ( .A(n7597), .B(n18194), .Z(n7466) );
  NANDN U8031 ( .A(n7464), .B(n18104), .Z(n7465) );
  NAND U8032 ( .A(n7466), .B(n7465), .Z(n7551) );
  XOR U8033 ( .A(n580), .B(a[51]), .Z(n7600) );
  NANDN U8034 ( .A(n7600), .B(n18336), .Z(n7469) );
  NANDN U8035 ( .A(n7467), .B(n18337), .Z(n7468) );
  AND U8036 ( .A(n7469), .B(n7468), .Z(n7550) );
  XNOR U8037 ( .A(n7551), .B(n7550), .Z(n7552) );
  XNOR U8038 ( .A(n7553), .B(n7552), .Z(n7569) );
  NANDN U8039 ( .A(n577), .B(a[63]), .Z(n7470) );
  XOR U8040 ( .A(n17151), .B(n7470), .Z(n7472) );
  NANDN U8041 ( .A(b[0]), .B(a[62]), .Z(n7471) );
  AND U8042 ( .A(n7472), .B(n7471), .Z(n7528) );
  NAND U8043 ( .A(n7473), .B(n19406), .Z(n7475) );
  XNOR U8044 ( .A(n584), .B(a[35]), .Z(n7606) );
  NANDN U8045 ( .A(n576), .B(n7606), .Z(n7474) );
  NAND U8046 ( .A(n7475), .B(n7474), .Z(n7526) );
  NANDN U8047 ( .A(n585), .B(a[31]), .Z(n7527) );
  XNOR U8048 ( .A(n7526), .B(n7527), .Z(n7529) );
  XNOR U8049 ( .A(n7528), .B(n7529), .Z(n7567) );
  XNOR U8050 ( .A(b[23]), .B(a[41]), .Z(n7609) );
  OR U8051 ( .A(n7609), .B(n19127), .Z(n7478) );
  NAND U8052 ( .A(n7476), .B(n19128), .Z(n7477) );
  NAND U8053 ( .A(n7478), .B(n7477), .Z(n7627) );
  NAND U8054 ( .A(n7479), .B(n17553), .Z(n7481) );
  XOR U8055 ( .A(b[7]), .B(a[57]), .Z(n7612) );
  NAND U8056 ( .A(n7612), .B(n17555), .Z(n7480) );
  NAND U8057 ( .A(n7481), .B(n7480), .Z(n7624) );
  XOR U8058 ( .A(b[25]), .B(a[39]), .Z(n7615) );
  NAND U8059 ( .A(n7615), .B(n19240), .Z(n7484) );
  NANDN U8060 ( .A(n7482), .B(n19242), .Z(n7483) );
  AND U8061 ( .A(n7484), .B(n7483), .Z(n7625) );
  XNOR U8062 ( .A(n7624), .B(n7625), .Z(n7626) );
  XOR U8063 ( .A(n7627), .B(n7626), .Z(n7566) );
  XOR U8064 ( .A(n7569), .B(n7568), .Z(n7579) );
  NANDN U8065 ( .A(n7486), .B(n7485), .Z(n7490) );
  NAND U8066 ( .A(n7488), .B(n7487), .Z(n7489) );
  NAND U8067 ( .A(n7490), .B(n7489), .Z(n7577) );
  NANDN U8068 ( .A(n7492), .B(n7491), .Z(n7496) );
  NAND U8069 ( .A(n7494), .B(n7493), .Z(n7495) );
  AND U8070 ( .A(n7496), .B(n7495), .Z(n7576) );
  XNOR U8071 ( .A(n7577), .B(n7576), .Z(n7578) );
  XNOR U8072 ( .A(n7579), .B(n7578), .Z(n7631) );
  XNOR U8073 ( .A(n7630), .B(n7631), .Z(n7632) );
  XOR U8074 ( .A(n7633), .B(n7632), .Z(n7648) );
  XOR U8075 ( .A(n7649), .B(n7648), .Z(n7650) );
  XNOR U8076 ( .A(n7651), .B(n7650), .Z(n7645) );
  NANDN U8077 ( .A(n7498), .B(n7497), .Z(n7502) );
  NAND U8078 ( .A(n7500), .B(n7499), .Z(n7501) );
  NAND U8079 ( .A(n7502), .B(n7501), .Z(n7642) );
  NAND U8080 ( .A(n7504), .B(n7503), .Z(n7508) );
  NAND U8081 ( .A(n7506), .B(n7505), .Z(n7507) );
  NAND U8082 ( .A(n7508), .B(n7507), .Z(n7643) );
  XNOR U8083 ( .A(n7642), .B(n7643), .Z(n7644) );
  XOR U8084 ( .A(n7645), .B(n7644), .Z(n7523) );
  XOR U8085 ( .A(n7522), .B(n7523), .Z(n7514) );
  XOR U8086 ( .A(n7515), .B(n7514), .Z(n7516) );
  XNOR U8087 ( .A(n7517), .B(n7516), .Z(n7654) );
  XNOR U8088 ( .A(n7654), .B(sreg[159]), .Z(n7656) );
  NAND U8089 ( .A(n7509), .B(sreg[158]), .Z(n7513) );
  OR U8090 ( .A(n7511), .B(n7510), .Z(n7512) );
  AND U8091 ( .A(n7513), .B(n7512), .Z(n7655) );
  XOR U8092 ( .A(n7656), .B(n7655), .Z(c[159]) );
  NAND U8093 ( .A(n7515), .B(n7514), .Z(n7519) );
  NAND U8094 ( .A(n7517), .B(n7516), .Z(n7518) );
  NAND U8095 ( .A(n7519), .B(n7518), .Z(n7662) );
  NANDN U8096 ( .A(n7521), .B(n7520), .Z(n7525) );
  NAND U8097 ( .A(n7523), .B(n7522), .Z(n7524) );
  NAND U8098 ( .A(n7525), .B(n7524), .Z(n7660) );
  NANDN U8099 ( .A(n7527), .B(n7526), .Z(n7531) );
  NAND U8100 ( .A(n7529), .B(n7528), .Z(n7530) );
  NAND U8101 ( .A(n7531), .B(n7530), .Z(n7738) );
  NANDN U8102 ( .A(n7532), .B(n18832), .Z(n7534) );
  XNOR U8103 ( .A(b[19]), .B(a[46]), .Z(n7685) );
  NANDN U8104 ( .A(n7685), .B(n18834), .Z(n7533) );
  NAND U8105 ( .A(n7534), .B(n7533), .Z(n7748) );
  XOR U8106 ( .A(b[27]), .B(n8490), .Z(n7688) );
  NANDN U8107 ( .A(n7688), .B(n19336), .Z(n7537) );
  NANDN U8108 ( .A(n7535), .B(n19337), .Z(n7536) );
  NAND U8109 ( .A(n7537), .B(n7536), .Z(n7745) );
  XOR U8110 ( .A(b[5]), .B(a[60]), .Z(n7691) );
  NAND U8111 ( .A(n7691), .B(n17310), .Z(n7540) );
  NAND U8112 ( .A(n7538), .B(n17311), .Z(n7539) );
  AND U8113 ( .A(n7540), .B(n7539), .Z(n7746) );
  XNOR U8114 ( .A(n7745), .B(n7746), .Z(n7747) );
  XNOR U8115 ( .A(n7748), .B(n7747), .Z(n7736) );
  XOR U8116 ( .A(b[17]), .B(a[48]), .Z(n7694) );
  NAND U8117 ( .A(n7694), .B(n18673), .Z(n7543) );
  NAND U8118 ( .A(n7541), .B(n18674), .Z(n7542) );
  NAND U8119 ( .A(n7543), .B(n7542), .Z(n7712) );
  XNOR U8120 ( .A(b[31]), .B(a[34]), .Z(n7697) );
  NANDN U8121 ( .A(n7697), .B(n19472), .Z(n7546) );
  NANDN U8122 ( .A(n7544), .B(n19473), .Z(n7545) );
  NAND U8123 ( .A(n7546), .B(n7545), .Z(n7709) );
  OR U8124 ( .A(n7547), .B(n16988), .Z(n7549) );
  XNOR U8125 ( .A(b[3]), .B(a[62]), .Z(n7700) );
  NANDN U8126 ( .A(n7700), .B(n16990), .Z(n7548) );
  AND U8127 ( .A(n7549), .B(n7548), .Z(n7710) );
  XNOR U8128 ( .A(n7709), .B(n7710), .Z(n7711) );
  XOR U8129 ( .A(n7712), .B(n7711), .Z(n7735) );
  XNOR U8130 ( .A(n7736), .B(n7735), .Z(n7737) );
  XNOR U8131 ( .A(n7738), .B(n7737), .Z(n7676) );
  NANDN U8132 ( .A(n7551), .B(n7550), .Z(n7555) );
  NAND U8133 ( .A(n7553), .B(n7552), .Z(n7554) );
  NAND U8134 ( .A(n7555), .B(n7554), .Z(n7727) );
  NANDN U8135 ( .A(n7557), .B(n7556), .Z(n7561) );
  NAND U8136 ( .A(n7559), .B(n7558), .Z(n7560) );
  NAND U8137 ( .A(n7561), .B(n7560), .Z(n7726) );
  XNOR U8138 ( .A(n7726), .B(n7725), .Z(n7728) );
  XOR U8139 ( .A(n7727), .B(n7728), .Z(n7675) );
  XOR U8140 ( .A(n7676), .B(n7675), .Z(n7677) );
  NANDN U8141 ( .A(n7567), .B(n7566), .Z(n7571) );
  NAND U8142 ( .A(n7569), .B(n7568), .Z(n7570) );
  AND U8143 ( .A(n7571), .B(n7570), .Z(n7678) );
  XNOR U8144 ( .A(n7677), .B(n7678), .Z(n7784) );
  NANDN U8145 ( .A(n7577), .B(n7576), .Z(n7581) );
  NANDN U8146 ( .A(n7579), .B(n7578), .Z(n7580) );
  NAND U8147 ( .A(n7581), .B(n7580), .Z(n7672) );
  NANDN U8148 ( .A(n7583), .B(n7582), .Z(n7587) );
  OR U8149 ( .A(n7585), .B(n7584), .Z(n7586) );
  NAND U8150 ( .A(n7587), .B(n7586), .Z(n7669) );
  XNOR U8151 ( .A(b[21]), .B(a[44]), .Z(n7757) );
  NANDN U8152 ( .A(n7757), .B(n19015), .Z(n7590) );
  NANDN U8153 ( .A(n7588), .B(n19013), .Z(n7589) );
  NAND U8154 ( .A(n7590), .B(n7589), .Z(n7721) );
  NANDN U8155 ( .A(n7591), .B(n18513), .Z(n7593) );
  XOR U8156 ( .A(b[15]), .B(a[50]), .Z(n7754) );
  NANDN U8157 ( .A(n18512), .B(n7754), .Z(n7592) );
  AND U8158 ( .A(n7593), .B(n7592), .Z(n7722) );
  XNOR U8159 ( .A(n7721), .B(n7722), .Z(n7724) );
  XNOR U8160 ( .A(b[9]), .B(a[56]), .Z(n7751) );
  NANDN U8161 ( .A(n7751), .B(n17814), .Z(n7596) );
  NANDN U8162 ( .A(n7594), .B(n17815), .Z(n7595) );
  NAND U8163 ( .A(n7596), .B(n7595), .Z(n7723) );
  XNOR U8164 ( .A(n7724), .B(n7723), .Z(n7717) );
  XNOR U8165 ( .A(b[11]), .B(a[54]), .Z(n7760) );
  OR U8166 ( .A(n7760), .B(n18194), .Z(n7599) );
  NANDN U8167 ( .A(n7597), .B(n18104), .Z(n7598) );
  NAND U8168 ( .A(n7599), .B(n7598), .Z(n7716) );
  XOR U8169 ( .A(n580), .B(a[52]), .Z(n7763) );
  NANDN U8170 ( .A(n7763), .B(n18336), .Z(n7602) );
  NANDN U8171 ( .A(n7600), .B(n18337), .Z(n7601) );
  NAND U8172 ( .A(n7602), .B(n7601), .Z(n7715) );
  XNOR U8173 ( .A(n7716), .B(n7715), .Z(n7718) );
  XNOR U8174 ( .A(n7717), .B(n7718), .Z(n7706) );
  NANDN U8175 ( .A(n577), .B(a[64]), .Z(n7603) );
  XOR U8176 ( .A(n17151), .B(n7603), .Z(n7605) );
  NANDN U8177 ( .A(b[0]), .B(a[63]), .Z(n7604) );
  AND U8178 ( .A(n7605), .B(n7604), .Z(n7681) );
  NAND U8179 ( .A(n19406), .B(n7606), .Z(n7608) );
  XNOR U8180 ( .A(n584), .B(a[36]), .Z(n7769) );
  NANDN U8181 ( .A(n576), .B(n7769), .Z(n7607) );
  NAND U8182 ( .A(n7608), .B(n7607), .Z(n7679) );
  NANDN U8183 ( .A(n585), .B(a[32]), .Z(n7680) );
  XNOR U8184 ( .A(n7679), .B(n7680), .Z(n7682) );
  XNOR U8185 ( .A(n7681), .B(n7682), .Z(n7704) );
  XNOR U8186 ( .A(b[23]), .B(a[42]), .Z(n7772) );
  OR U8187 ( .A(n7772), .B(n19127), .Z(n7611) );
  NANDN U8188 ( .A(n7609), .B(n19128), .Z(n7610) );
  NAND U8189 ( .A(n7611), .B(n7610), .Z(n7742) );
  NAND U8190 ( .A(n7612), .B(n17553), .Z(n7614) );
  XOR U8191 ( .A(b[7]), .B(a[58]), .Z(n7775) );
  NAND U8192 ( .A(n7775), .B(n17555), .Z(n7613) );
  NAND U8193 ( .A(n7614), .B(n7613), .Z(n7739) );
  XOR U8194 ( .A(b[25]), .B(a[40]), .Z(n7778) );
  NAND U8195 ( .A(n7778), .B(n19240), .Z(n7617) );
  NAND U8196 ( .A(n7615), .B(n19242), .Z(n7616) );
  AND U8197 ( .A(n7617), .B(n7616), .Z(n7740) );
  XNOR U8198 ( .A(n7739), .B(n7740), .Z(n7741) );
  XOR U8199 ( .A(n7742), .B(n7741), .Z(n7703) );
  XNOR U8200 ( .A(n7706), .B(n7705), .Z(n7732) );
  NANDN U8201 ( .A(n7619), .B(n7618), .Z(n7623) );
  NAND U8202 ( .A(n7621), .B(n7620), .Z(n7622) );
  NAND U8203 ( .A(n7623), .B(n7622), .Z(n7730) );
  NANDN U8204 ( .A(n7625), .B(n7624), .Z(n7629) );
  NAND U8205 ( .A(n7627), .B(n7626), .Z(n7628) );
  AND U8206 ( .A(n7629), .B(n7628), .Z(n7729) );
  XNOR U8207 ( .A(n7730), .B(n7729), .Z(n7731) );
  XNOR U8208 ( .A(n7732), .B(n7731), .Z(n7670) );
  XNOR U8209 ( .A(n7669), .B(n7670), .Z(n7671) );
  XNOR U8210 ( .A(n7672), .B(n7671), .Z(n7782) );
  XNOR U8211 ( .A(n7781), .B(n7782), .Z(n7783) );
  XNOR U8212 ( .A(n7784), .B(n7783), .Z(n7788) );
  NANDN U8213 ( .A(n7631), .B(n7630), .Z(n7635) );
  NAND U8214 ( .A(n7633), .B(n7632), .Z(n7634) );
  NAND U8215 ( .A(n7635), .B(n7634), .Z(n7785) );
  NANDN U8216 ( .A(n7637), .B(n7636), .Z(n7641) );
  NAND U8217 ( .A(n7639), .B(n7638), .Z(n7640) );
  NAND U8218 ( .A(n7641), .B(n7640), .Z(n7786) );
  XNOR U8219 ( .A(n7785), .B(n7786), .Z(n7787) );
  XNOR U8220 ( .A(n7788), .B(n7787), .Z(n7666) );
  NANDN U8221 ( .A(n7643), .B(n7642), .Z(n7647) );
  NAND U8222 ( .A(n7645), .B(n7644), .Z(n7646) );
  NAND U8223 ( .A(n7647), .B(n7646), .Z(n7663) );
  NANDN U8224 ( .A(n7649), .B(n7648), .Z(n7653) );
  OR U8225 ( .A(n7651), .B(n7650), .Z(n7652) );
  NAND U8226 ( .A(n7653), .B(n7652), .Z(n7664) );
  XNOR U8227 ( .A(n7663), .B(n7664), .Z(n7665) );
  XNOR U8228 ( .A(n7666), .B(n7665), .Z(n7659) );
  XOR U8229 ( .A(n7660), .B(n7659), .Z(n7661) );
  XNOR U8230 ( .A(n7662), .B(n7661), .Z(n7791) );
  XNOR U8231 ( .A(n7791), .B(sreg[160]), .Z(n7793) );
  NAND U8232 ( .A(n7654), .B(sreg[159]), .Z(n7658) );
  OR U8233 ( .A(n7656), .B(n7655), .Z(n7657) );
  AND U8234 ( .A(n7658), .B(n7657), .Z(n7792) );
  XOR U8235 ( .A(n7793), .B(n7792), .Z(c[160]) );
  NANDN U8236 ( .A(n7664), .B(n7663), .Z(n7668) );
  NANDN U8237 ( .A(n7666), .B(n7665), .Z(n7667) );
  NAND U8238 ( .A(n7668), .B(n7667), .Z(n7796) );
  NANDN U8239 ( .A(n7670), .B(n7669), .Z(n7674) );
  NANDN U8240 ( .A(n7672), .B(n7671), .Z(n7673) );
  NAND U8241 ( .A(n7674), .B(n7673), .Z(n7924) );
  XNOR U8242 ( .A(n7924), .B(n7925), .Z(n7926) );
  NANDN U8243 ( .A(n7680), .B(n7679), .Z(n7684) );
  NAND U8244 ( .A(n7682), .B(n7681), .Z(n7683) );
  NAND U8245 ( .A(n7684), .B(n7683), .Z(n7869) );
  NANDN U8246 ( .A(n7685), .B(n18832), .Z(n7687) );
  XNOR U8247 ( .A(b[19]), .B(a[47]), .Z(n7814) );
  NANDN U8248 ( .A(n7814), .B(n18834), .Z(n7686) );
  NAND U8249 ( .A(n7687), .B(n7686), .Z(n7903) );
  XNOR U8250 ( .A(b[27]), .B(a[39]), .Z(n7817) );
  NANDN U8251 ( .A(n7817), .B(n19336), .Z(n7690) );
  NANDN U8252 ( .A(n7688), .B(n19337), .Z(n7689) );
  NAND U8253 ( .A(n7690), .B(n7689), .Z(n7900) );
  XOR U8254 ( .A(b[5]), .B(a[61]), .Z(n7820) );
  NAND U8255 ( .A(n7820), .B(n17310), .Z(n7693) );
  NAND U8256 ( .A(n7691), .B(n17311), .Z(n7692) );
  AND U8257 ( .A(n7693), .B(n7692), .Z(n7901) );
  XNOR U8258 ( .A(n7900), .B(n7901), .Z(n7902) );
  XNOR U8259 ( .A(n7903), .B(n7902), .Z(n7867) );
  XNOR U8260 ( .A(b[17]), .B(a[49]), .Z(n7823) );
  NANDN U8261 ( .A(n7823), .B(n18673), .Z(n7696) );
  NAND U8262 ( .A(n7694), .B(n18674), .Z(n7695) );
  NAND U8263 ( .A(n7696), .B(n7695), .Z(n7841) );
  XNOR U8264 ( .A(b[31]), .B(a[35]), .Z(n7826) );
  NANDN U8265 ( .A(n7826), .B(n19472), .Z(n7699) );
  NANDN U8266 ( .A(n7697), .B(n19473), .Z(n7698) );
  NAND U8267 ( .A(n7699), .B(n7698), .Z(n7838) );
  OR U8268 ( .A(n7700), .B(n16988), .Z(n7702) );
  XNOR U8269 ( .A(b[3]), .B(a[63]), .Z(n7829) );
  NANDN U8270 ( .A(n7829), .B(n16990), .Z(n7701) );
  AND U8271 ( .A(n7702), .B(n7701), .Z(n7839) );
  XNOR U8272 ( .A(n7838), .B(n7839), .Z(n7840) );
  XOR U8273 ( .A(n7841), .B(n7840), .Z(n7866) );
  XNOR U8274 ( .A(n7867), .B(n7866), .Z(n7868) );
  XNOR U8275 ( .A(n7869), .B(n7868), .Z(n7918) );
  NANDN U8276 ( .A(n7704), .B(n7703), .Z(n7708) );
  NANDN U8277 ( .A(n7706), .B(n7705), .Z(n7707) );
  NAND U8278 ( .A(n7708), .B(n7707), .Z(n7919) );
  XNOR U8279 ( .A(n7918), .B(n7919), .Z(n7920) );
  NANDN U8280 ( .A(n7710), .B(n7709), .Z(n7714) );
  NAND U8281 ( .A(n7712), .B(n7711), .Z(n7713) );
  NAND U8282 ( .A(n7714), .B(n7713), .Z(n7859) );
  OR U8283 ( .A(n7716), .B(n7715), .Z(n7720) );
  NANDN U8284 ( .A(n7718), .B(n7717), .Z(n7719) );
  NAND U8285 ( .A(n7720), .B(n7719), .Z(n7857) );
  XNOR U8286 ( .A(n7857), .B(n7856), .Z(n7858) );
  XOR U8287 ( .A(n7859), .B(n7858), .Z(n7921) );
  XOR U8288 ( .A(n7920), .B(n7921), .Z(n7933) );
  NANDN U8289 ( .A(n7730), .B(n7729), .Z(n7734) );
  NANDN U8290 ( .A(n7732), .B(n7731), .Z(n7733) );
  NAND U8291 ( .A(n7734), .B(n7733), .Z(n7915) );
  NANDN U8292 ( .A(n7740), .B(n7739), .Z(n7744) );
  NAND U8293 ( .A(n7742), .B(n7741), .Z(n7743) );
  NAND U8294 ( .A(n7744), .B(n7743), .Z(n7860) );
  NANDN U8295 ( .A(n7746), .B(n7745), .Z(n7750) );
  NAND U8296 ( .A(n7748), .B(n7747), .Z(n7749) );
  AND U8297 ( .A(n7750), .B(n7749), .Z(n7861) );
  XNOR U8298 ( .A(n7860), .B(n7861), .Z(n7862) );
  XNOR U8299 ( .A(n579), .B(a[57]), .Z(n7870) );
  NAND U8300 ( .A(n17814), .B(n7870), .Z(n7753) );
  NANDN U8301 ( .A(n7751), .B(n17815), .Z(n7752) );
  NAND U8302 ( .A(n7753), .B(n7752), .Z(n7846) );
  NAND U8303 ( .A(n7754), .B(n18513), .Z(n7756) );
  XOR U8304 ( .A(b[15]), .B(a[51]), .Z(n7873) );
  NANDN U8305 ( .A(n18512), .B(n7873), .Z(n7755) );
  AND U8306 ( .A(n7756), .B(n7755), .Z(n7844) );
  NANDN U8307 ( .A(n7757), .B(n19013), .Z(n7759) );
  XNOR U8308 ( .A(n582), .B(a[45]), .Z(n7876) );
  NAND U8309 ( .A(n7876), .B(n19015), .Z(n7758) );
  AND U8310 ( .A(n7759), .B(n7758), .Z(n7845) );
  XOR U8311 ( .A(n7846), .B(n7847), .Z(n7835) );
  XOR U8312 ( .A(b[11]), .B(n10959), .Z(n7879) );
  OR U8313 ( .A(n7879), .B(n18194), .Z(n7762) );
  NANDN U8314 ( .A(n7760), .B(n18104), .Z(n7761) );
  NAND U8315 ( .A(n7762), .B(n7761), .Z(n7833) );
  XOR U8316 ( .A(n580), .B(a[53]), .Z(n7882) );
  NANDN U8317 ( .A(n7882), .B(n18336), .Z(n7765) );
  NANDN U8318 ( .A(n7763), .B(n18337), .Z(n7764) );
  AND U8319 ( .A(n7765), .B(n7764), .Z(n7832) );
  XNOR U8320 ( .A(n7833), .B(n7832), .Z(n7834) );
  XOR U8321 ( .A(n7835), .B(n7834), .Z(n7852) );
  ANDN U8322 ( .B(a[65]), .A(n577), .Z(n7766) );
  XNOR U8323 ( .A(n17151), .B(n7766), .Z(n7768) );
  NANDN U8324 ( .A(b[0]), .B(a[64]), .Z(n7767) );
  NAND U8325 ( .A(n7768), .B(n7767), .Z(n7811) );
  NAND U8326 ( .A(n19406), .B(n7769), .Z(n7771) );
  XNOR U8327 ( .A(n584), .B(a[37]), .Z(n7888) );
  NANDN U8328 ( .A(n576), .B(n7888), .Z(n7770) );
  NAND U8329 ( .A(n7771), .B(n7770), .Z(n7808) );
  NANDN U8330 ( .A(n585), .B(a[33]), .Z(n7809) );
  XNOR U8331 ( .A(n7808), .B(n7809), .Z(n7810) );
  XNOR U8332 ( .A(n7811), .B(n7810), .Z(n7850) );
  XOR U8333 ( .A(b[23]), .B(a[43]), .Z(n7891) );
  NANDN U8334 ( .A(n19127), .B(n7891), .Z(n7774) );
  NANDN U8335 ( .A(n7772), .B(n19128), .Z(n7773) );
  NAND U8336 ( .A(n7774), .B(n7773), .Z(n7909) );
  NAND U8337 ( .A(n7775), .B(n17553), .Z(n7777) );
  XOR U8338 ( .A(b[7]), .B(a[59]), .Z(n7894) );
  NAND U8339 ( .A(n7894), .B(n17555), .Z(n7776) );
  NAND U8340 ( .A(n7777), .B(n7776), .Z(n7906) );
  XNOR U8341 ( .A(b[25]), .B(a[41]), .Z(n7897) );
  NANDN U8342 ( .A(n7897), .B(n19240), .Z(n7780) );
  NAND U8343 ( .A(n7778), .B(n19242), .Z(n7779) );
  AND U8344 ( .A(n7780), .B(n7779), .Z(n7907) );
  XNOR U8345 ( .A(n7906), .B(n7907), .Z(n7908) );
  XNOR U8346 ( .A(n7909), .B(n7908), .Z(n7851) );
  XOR U8347 ( .A(n7850), .B(n7851), .Z(n7853) );
  XNOR U8348 ( .A(n7852), .B(n7853), .Z(n7863) );
  XNOR U8349 ( .A(n7862), .B(n7863), .Z(n7912) );
  XNOR U8350 ( .A(n7913), .B(n7912), .Z(n7914) );
  XOR U8351 ( .A(n7915), .B(n7914), .Z(n7930) );
  XNOR U8352 ( .A(n7931), .B(n7930), .Z(n7932) );
  XOR U8353 ( .A(n7933), .B(n7932), .Z(n7927) );
  XOR U8354 ( .A(n7926), .B(n7927), .Z(n7805) );
  NANDN U8355 ( .A(n7786), .B(n7785), .Z(n7790) );
  NANDN U8356 ( .A(n7788), .B(n7787), .Z(n7789) );
  NAND U8357 ( .A(n7790), .B(n7789), .Z(n7803) );
  XNOR U8358 ( .A(n7802), .B(n7803), .Z(n7804) );
  XNOR U8359 ( .A(n7805), .B(n7804), .Z(n7797) );
  XNOR U8360 ( .A(n7796), .B(n7797), .Z(n7798) );
  XNOR U8361 ( .A(n7799), .B(n7798), .Z(n7934) );
  XNOR U8362 ( .A(n7934), .B(sreg[161]), .Z(n7936) );
  NAND U8363 ( .A(n7791), .B(sreg[160]), .Z(n7795) );
  OR U8364 ( .A(n7793), .B(n7792), .Z(n7794) );
  AND U8365 ( .A(n7795), .B(n7794), .Z(n7935) );
  XOR U8366 ( .A(n7936), .B(n7935), .Z(c[161]) );
  NANDN U8367 ( .A(n7797), .B(n7796), .Z(n7801) );
  NAND U8368 ( .A(n7799), .B(n7798), .Z(n7800) );
  NAND U8369 ( .A(n7801), .B(n7800), .Z(n7942) );
  NANDN U8370 ( .A(n7803), .B(n7802), .Z(n7807) );
  NAND U8371 ( .A(n7805), .B(n7804), .Z(n7806) );
  NAND U8372 ( .A(n7807), .B(n7806), .Z(n7940) );
  NANDN U8373 ( .A(n7809), .B(n7808), .Z(n7813) );
  NANDN U8374 ( .A(n7811), .B(n7810), .Z(n7812) );
  NAND U8375 ( .A(n7813), .B(n7812), .Z(n8010) );
  NANDN U8376 ( .A(n7814), .B(n18832), .Z(n7816) );
  XNOR U8377 ( .A(b[19]), .B(a[48]), .Z(n7955) );
  NANDN U8378 ( .A(n7955), .B(n18834), .Z(n7815) );
  NAND U8379 ( .A(n7816), .B(n7815), .Z(n8020) );
  XNOR U8380 ( .A(b[27]), .B(a[40]), .Z(n7958) );
  NANDN U8381 ( .A(n7958), .B(n19336), .Z(n7819) );
  NANDN U8382 ( .A(n7817), .B(n19337), .Z(n7818) );
  NAND U8383 ( .A(n7819), .B(n7818), .Z(n8017) );
  XOR U8384 ( .A(b[5]), .B(a[62]), .Z(n7961) );
  NAND U8385 ( .A(n7961), .B(n17310), .Z(n7822) );
  NAND U8386 ( .A(n7820), .B(n17311), .Z(n7821) );
  AND U8387 ( .A(n7822), .B(n7821), .Z(n8018) );
  XNOR U8388 ( .A(n8017), .B(n8018), .Z(n8019) );
  XNOR U8389 ( .A(n8020), .B(n8019), .Z(n8008) );
  XOR U8390 ( .A(b[17]), .B(a[50]), .Z(n7964) );
  NAND U8391 ( .A(n7964), .B(n18673), .Z(n7825) );
  NANDN U8392 ( .A(n7823), .B(n18674), .Z(n7824) );
  NAND U8393 ( .A(n7825), .B(n7824), .Z(n7982) );
  XNOR U8394 ( .A(b[31]), .B(a[36]), .Z(n7967) );
  NANDN U8395 ( .A(n7967), .B(n19472), .Z(n7828) );
  NANDN U8396 ( .A(n7826), .B(n19473), .Z(n7827) );
  NAND U8397 ( .A(n7828), .B(n7827), .Z(n7979) );
  OR U8398 ( .A(n7829), .B(n16988), .Z(n7831) );
  XNOR U8399 ( .A(b[3]), .B(a[64]), .Z(n7970) );
  NANDN U8400 ( .A(n7970), .B(n16990), .Z(n7830) );
  AND U8401 ( .A(n7831), .B(n7830), .Z(n7980) );
  XNOR U8402 ( .A(n7979), .B(n7980), .Z(n7981) );
  XOR U8403 ( .A(n7982), .B(n7981), .Z(n8007) );
  XNOR U8404 ( .A(n8008), .B(n8007), .Z(n8009) );
  XNOR U8405 ( .A(n8010), .B(n8009), .Z(n8053) );
  NANDN U8406 ( .A(n7833), .B(n7832), .Z(n7837) );
  NAND U8407 ( .A(n7835), .B(n7834), .Z(n7836) );
  NAND U8408 ( .A(n7837), .B(n7836), .Z(n7998) );
  NANDN U8409 ( .A(n7839), .B(n7838), .Z(n7843) );
  NAND U8410 ( .A(n7841), .B(n7840), .Z(n7842) );
  NAND U8411 ( .A(n7843), .B(n7842), .Z(n7996) );
  OR U8412 ( .A(n7845), .B(n7844), .Z(n7849) );
  NANDN U8413 ( .A(n7847), .B(n7846), .Z(n7848) );
  NAND U8414 ( .A(n7849), .B(n7848), .Z(n7995) );
  XNOR U8415 ( .A(n7998), .B(n7997), .Z(n8054) );
  XNOR U8416 ( .A(n8053), .B(n8054), .Z(n8055) );
  NANDN U8417 ( .A(n7851), .B(n7850), .Z(n7855) );
  OR U8418 ( .A(n7853), .B(n7852), .Z(n7854) );
  AND U8419 ( .A(n7855), .B(n7854), .Z(n8056) );
  XNOR U8420 ( .A(n8055), .B(n8056), .Z(n8068) );
  NANDN U8421 ( .A(n7861), .B(n7860), .Z(n7865) );
  NANDN U8422 ( .A(n7863), .B(n7862), .Z(n7864) );
  NAND U8423 ( .A(n7865), .B(n7864), .Z(n8062) );
  XNOR U8424 ( .A(b[9]), .B(a[58]), .Z(n8023) );
  NANDN U8425 ( .A(n8023), .B(n17814), .Z(n7872) );
  NAND U8426 ( .A(n17815), .B(n7870), .Z(n7871) );
  NAND U8427 ( .A(n7872), .B(n7871), .Z(n7987) );
  XNOR U8428 ( .A(b[15]), .B(a[52]), .Z(n8026) );
  OR U8429 ( .A(n8026), .B(n18512), .Z(n7875) );
  NAND U8430 ( .A(n7873), .B(n18513), .Z(n7874) );
  NAND U8431 ( .A(n7875), .B(n7874), .Z(n7985) );
  XNOR U8432 ( .A(b[21]), .B(a[46]), .Z(n8029) );
  NANDN U8433 ( .A(n8029), .B(n19015), .Z(n7878) );
  NAND U8434 ( .A(n19013), .B(n7876), .Z(n7877) );
  NAND U8435 ( .A(n7878), .B(n7877), .Z(n7986) );
  XNOR U8436 ( .A(n7985), .B(n7986), .Z(n7988) );
  XOR U8437 ( .A(n7987), .B(n7988), .Z(n7976) );
  XNOR U8438 ( .A(b[11]), .B(a[56]), .Z(n8032) );
  OR U8439 ( .A(n8032), .B(n18194), .Z(n7881) );
  NANDN U8440 ( .A(n7879), .B(n18104), .Z(n7880) );
  NAND U8441 ( .A(n7881), .B(n7880), .Z(n7974) );
  XOR U8442 ( .A(n580), .B(a[54]), .Z(n8035) );
  NANDN U8443 ( .A(n8035), .B(n18336), .Z(n7884) );
  NANDN U8444 ( .A(n7882), .B(n18337), .Z(n7883) );
  AND U8445 ( .A(n7884), .B(n7883), .Z(n7973) );
  XNOR U8446 ( .A(n7974), .B(n7973), .Z(n7975) );
  XNOR U8447 ( .A(n7976), .B(n7975), .Z(n7992) );
  NANDN U8448 ( .A(n577), .B(a[66]), .Z(n7885) );
  XOR U8449 ( .A(n17151), .B(n7885), .Z(n7887) );
  IV U8450 ( .A(a[65]), .Z(n12055) );
  NANDN U8451 ( .A(n12055), .B(n577), .Z(n7886) );
  AND U8452 ( .A(n7887), .B(n7886), .Z(n7951) );
  NAND U8453 ( .A(n19406), .B(n7888), .Z(n7890) );
  XOR U8454 ( .A(n584), .B(n8490), .Z(n8038) );
  NANDN U8455 ( .A(n576), .B(n8038), .Z(n7889) );
  NAND U8456 ( .A(n7890), .B(n7889), .Z(n7949) );
  NANDN U8457 ( .A(n585), .B(a[34]), .Z(n7950) );
  XNOR U8458 ( .A(n7949), .B(n7950), .Z(n7952) );
  XNOR U8459 ( .A(n7951), .B(n7952), .Z(n7990) );
  XOR U8460 ( .A(b[23]), .B(a[44]), .Z(n8044) );
  NANDN U8461 ( .A(n19127), .B(n8044), .Z(n7893) );
  NAND U8462 ( .A(n7891), .B(n19128), .Z(n7892) );
  NAND U8463 ( .A(n7893), .B(n7892), .Z(n8014) );
  NAND U8464 ( .A(n7894), .B(n17553), .Z(n7896) );
  XOR U8465 ( .A(b[7]), .B(a[60]), .Z(n8047) );
  NAND U8466 ( .A(n8047), .B(n17555), .Z(n7895) );
  NAND U8467 ( .A(n7896), .B(n7895), .Z(n8011) );
  XNOR U8468 ( .A(b[25]), .B(a[42]), .Z(n8050) );
  NANDN U8469 ( .A(n8050), .B(n19240), .Z(n7899) );
  NANDN U8470 ( .A(n7897), .B(n19242), .Z(n7898) );
  AND U8471 ( .A(n7899), .B(n7898), .Z(n8012) );
  XNOR U8472 ( .A(n8011), .B(n8012), .Z(n8013) );
  XOR U8473 ( .A(n8014), .B(n8013), .Z(n7989) );
  XOR U8474 ( .A(n7992), .B(n7991), .Z(n8004) );
  NANDN U8475 ( .A(n7901), .B(n7900), .Z(n7905) );
  NAND U8476 ( .A(n7903), .B(n7902), .Z(n7904) );
  NAND U8477 ( .A(n7905), .B(n7904), .Z(n8002) );
  NANDN U8478 ( .A(n7907), .B(n7906), .Z(n7911) );
  NAND U8479 ( .A(n7909), .B(n7908), .Z(n7910) );
  AND U8480 ( .A(n7911), .B(n7910), .Z(n8001) );
  XNOR U8481 ( .A(n8002), .B(n8001), .Z(n8003) );
  XNOR U8482 ( .A(n8004), .B(n8003), .Z(n8060) );
  XNOR U8483 ( .A(n8059), .B(n8060), .Z(n8061) );
  XOR U8484 ( .A(n8062), .B(n8061), .Z(n8066) );
  XNOR U8485 ( .A(n8065), .B(n8066), .Z(n8067) );
  XNOR U8486 ( .A(n8068), .B(n8067), .Z(n8072) );
  NAND U8487 ( .A(n7913), .B(n7912), .Z(n7917) );
  OR U8488 ( .A(n7915), .B(n7914), .Z(n7916) );
  NAND U8489 ( .A(n7917), .B(n7916), .Z(n8069) );
  NANDN U8490 ( .A(n7919), .B(n7918), .Z(n7923) );
  NAND U8491 ( .A(n7921), .B(n7920), .Z(n7922) );
  NAND U8492 ( .A(n7923), .B(n7922), .Z(n8070) );
  XNOR U8493 ( .A(n8069), .B(n8070), .Z(n8071) );
  XNOR U8494 ( .A(n8072), .B(n8071), .Z(n7946) );
  NANDN U8495 ( .A(n7925), .B(n7924), .Z(n7929) );
  NANDN U8496 ( .A(n7927), .B(n7926), .Z(n7928) );
  NAND U8497 ( .A(n7929), .B(n7928), .Z(n7944) );
  XNOR U8498 ( .A(n7944), .B(n7943), .Z(n7945) );
  XNOR U8499 ( .A(n7946), .B(n7945), .Z(n7939) );
  XOR U8500 ( .A(n7940), .B(n7939), .Z(n7941) );
  XNOR U8501 ( .A(n7942), .B(n7941), .Z(n8075) );
  XNOR U8502 ( .A(n8075), .B(sreg[162]), .Z(n8077) );
  NAND U8503 ( .A(n7934), .B(sreg[161]), .Z(n7938) );
  OR U8504 ( .A(n7936), .B(n7935), .Z(n7937) );
  AND U8505 ( .A(n7938), .B(n7937), .Z(n8076) );
  XOR U8506 ( .A(n8077), .B(n8076), .Z(c[162]) );
  NANDN U8507 ( .A(n7944), .B(n7943), .Z(n7948) );
  NANDN U8508 ( .A(n7946), .B(n7945), .Z(n7947) );
  NAND U8509 ( .A(n7948), .B(n7947), .Z(n8081) );
  NANDN U8510 ( .A(n7950), .B(n7949), .Z(n7954) );
  NAND U8511 ( .A(n7952), .B(n7951), .Z(n7953) );
  NAND U8512 ( .A(n7954), .B(n7953), .Z(n8163) );
  NANDN U8513 ( .A(n7955), .B(n18832), .Z(n7957) );
  XOR U8514 ( .A(b[19]), .B(n10083), .Z(n8132) );
  NANDN U8515 ( .A(n8132), .B(n18834), .Z(n7956) );
  NAND U8516 ( .A(n7957), .B(n7956), .Z(n8175) );
  XOR U8517 ( .A(b[27]), .B(n8930), .Z(n8135) );
  NANDN U8518 ( .A(n8135), .B(n19336), .Z(n7960) );
  NANDN U8519 ( .A(n7958), .B(n19337), .Z(n7959) );
  NAND U8520 ( .A(n7960), .B(n7959), .Z(n8172) );
  XOR U8521 ( .A(b[5]), .B(a[63]), .Z(n8138) );
  NAND U8522 ( .A(n8138), .B(n17310), .Z(n7963) );
  NAND U8523 ( .A(n7961), .B(n17311), .Z(n7962) );
  AND U8524 ( .A(n7963), .B(n7962), .Z(n8173) );
  XNOR U8525 ( .A(n8172), .B(n8173), .Z(n8174) );
  XNOR U8526 ( .A(n8175), .B(n8174), .Z(n8160) );
  XOR U8527 ( .A(b[17]), .B(a[51]), .Z(n8141) );
  NAND U8528 ( .A(n8141), .B(n18673), .Z(n7966) );
  NAND U8529 ( .A(n7964), .B(n18674), .Z(n7965) );
  NAND U8530 ( .A(n7966), .B(n7965), .Z(n8116) );
  XNOR U8531 ( .A(b[31]), .B(a[37]), .Z(n8144) );
  NANDN U8532 ( .A(n8144), .B(n19472), .Z(n7969) );
  NANDN U8533 ( .A(n7967), .B(n19473), .Z(n7968) );
  AND U8534 ( .A(n7969), .B(n7968), .Z(n8114) );
  OR U8535 ( .A(n7970), .B(n16988), .Z(n7972) );
  XOR U8536 ( .A(b[3]), .B(n12055), .Z(n8147) );
  NANDN U8537 ( .A(n8147), .B(n16990), .Z(n7971) );
  AND U8538 ( .A(n7972), .B(n7971), .Z(n8115) );
  XOR U8539 ( .A(n8116), .B(n8117), .Z(n8161) );
  XOR U8540 ( .A(n8160), .B(n8161), .Z(n8162) );
  XNOR U8541 ( .A(n8163), .B(n8162), .Z(n8099) );
  NANDN U8542 ( .A(n7974), .B(n7973), .Z(n7978) );
  NAND U8543 ( .A(n7976), .B(n7975), .Z(n7977) );
  NAND U8544 ( .A(n7978), .B(n7977), .Z(n8152) );
  NANDN U8545 ( .A(n7980), .B(n7979), .Z(n7984) );
  NAND U8546 ( .A(n7982), .B(n7981), .Z(n7983) );
  NAND U8547 ( .A(n7984), .B(n7983), .Z(n8151) );
  XNOR U8548 ( .A(n8151), .B(n8150), .Z(n8153) );
  XOR U8549 ( .A(n8152), .B(n8153), .Z(n8098) );
  XOR U8550 ( .A(n8099), .B(n8098), .Z(n8100) );
  NANDN U8551 ( .A(n7990), .B(n7989), .Z(n7994) );
  NAND U8552 ( .A(n7992), .B(n7991), .Z(n7993) );
  NAND U8553 ( .A(n7994), .B(n7993), .Z(n8101) );
  XNOR U8554 ( .A(n8100), .B(n8101), .Z(n8216) );
  OR U8555 ( .A(n7996), .B(n7995), .Z(n8000) );
  NAND U8556 ( .A(n7998), .B(n7997), .Z(n7999) );
  NAND U8557 ( .A(n8000), .B(n7999), .Z(n8215) );
  NANDN U8558 ( .A(n8002), .B(n8001), .Z(n8006) );
  NANDN U8559 ( .A(n8004), .B(n8003), .Z(n8005) );
  NAND U8560 ( .A(n8006), .B(n8005), .Z(n8095) );
  NANDN U8561 ( .A(n8012), .B(n8011), .Z(n8016) );
  NAND U8562 ( .A(n8014), .B(n8013), .Z(n8015) );
  NAND U8563 ( .A(n8016), .B(n8015), .Z(n8154) );
  NANDN U8564 ( .A(n8018), .B(n8017), .Z(n8022) );
  NAND U8565 ( .A(n8020), .B(n8019), .Z(n8021) );
  AND U8566 ( .A(n8022), .B(n8021), .Z(n8155) );
  XNOR U8567 ( .A(n8154), .B(n8155), .Z(n8156) );
  XNOR U8568 ( .A(b[9]), .B(a[59]), .Z(n8178) );
  NANDN U8569 ( .A(n8178), .B(n17814), .Z(n8025) );
  NANDN U8570 ( .A(n8023), .B(n17815), .Z(n8024) );
  NAND U8571 ( .A(n8025), .B(n8024), .Z(n8122) );
  NANDN U8572 ( .A(n8026), .B(n18513), .Z(n8028) );
  XNOR U8573 ( .A(b[15]), .B(a[53]), .Z(n8181) );
  OR U8574 ( .A(n8181), .B(n18512), .Z(n8027) );
  AND U8575 ( .A(n8028), .B(n8027), .Z(n8120) );
  NANDN U8576 ( .A(n8029), .B(n19013), .Z(n8031) );
  XNOR U8577 ( .A(b[21]), .B(a[47]), .Z(n8184) );
  NANDN U8578 ( .A(n8184), .B(n19015), .Z(n8030) );
  AND U8579 ( .A(n8031), .B(n8030), .Z(n8121) );
  XOR U8580 ( .A(n8122), .B(n8123), .Z(n8111) );
  XNOR U8581 ( .A(b[11]), .B(a[57]), .Z(n8187) );
  OR U8582 ( .A(n8187), .B(n18194), .Z(n8034) );
  NANDN U8583 ( .A(n8032), .B(n18104), .Z(n8033) );
  NAND U8584 ( .A(n8034), .B(n8033), .Z(n8109) );
  XOR U8585 ( .A(n580), .B(a[55]), .Z(n8190) );
  NANDN U8586 ( .A(n8190), .B(n18336), .Z(n8037) );
  NANDN U8587 ( .A(n8035), .B(n18337), .Z(n8036) );
  NAND U8588 ( .A(n8037), .B(n8036), .Z(n8108) );
  XOR U8589 ( .A(n8111), .B(n8110), .Z(n8105) );
  NAND U8590 ( .A(n19406), .B(n8038), .Z(n8040) );
  XNOR U8591 ( .A(n584), .B(a[39]), .Z(n8196) );
  NANDN U8592 ( .A(n576), .B(n8196), .Z(n8039) );
  NAND U8593 ( .A(n8040), .B(n8039), .Z(n8126) );
  NANDN U8594 ( .A(n585), .B(a[35]), .Z(n8127) );
  XNOR U8595 ( .A(n8126), .B(n8127), .Z(n8129) );
  NANDN U8596 ( .A(n577), .B(a[67]), .Z(n8041) );
  XOR U8597 ( .A(n17151), .B(n8041), .Z(n8043) );
  NANDN U8598 ( .A(b[0]), .B(a[66]), .Z(n8042) );
  AND U8599 ( .A(n8043), .B(n8042), .Z(n8128) );
  XNOR U8600 ( .A(n8129), .B(n8128), .Z(n8103) );
  XOR U8601 ( .A(b[23]), .B(a[45]), .Z(n8199) );
  NANDN U8602 ( .A(n19127), .B(n8199), .Z(n8046) );
  NAND U8603 ( .A(n8044), .B(n19128), .Z(n8045) );
  NAND U8604 ( .A(n8046), .B(n8045), .Z(n8169) );
  NAND U8605 ( .A(n8047), .B(n17553), .Z(n8049) );
  XOR U8606 ( .A(b[7]), .B(a[61]), .Z(n8202) );
  NAND U8607 ( .A(n8202), .B(n17555), .Z(n8048) );
  NAND U8608 ( .A(n8049), .B(n8048), .Z(n8166) );
  XOR U8609 ( .A(b[25]), .B(a[43]), .Z(n8205) );
  NAND U8610 ( .A(n8205), .B(n19240), .Z(n8052) );
  NANDN U8611 ( .A(n8050), .B(n19242), .Z(n8051) );
  AND U8612 ( .A(n8052), .B(n8051), .Z(n8167) );
  XNOR U8613 ( .A(n8166), .B(n8167), .Z(n8168) );
  XOR U8614 ( .A(n8169), .B(n8168), .Z(n8102) );
  XOR U8615 ( .A(n8105), .B(n8104), .Z(n8157) );
  XNOR U8616 ( .A(n8156), .B(n8157), .Z(n8092) );
  XOR U8617 ( .A(n8093), .B(n8092), .Z(n8094) );
  XNOR U8618 ( .A(n8095), .B(n8094), .Z(n8214) );
  XOR U8619 ( .A(n8215), .B(n8214), .Z(n8217) );
  NANDN U8620 ( .A(n8054), .B(n8053), .Z(n8058) );
  NAND U8621 ( .A(n8056), .B(n8055), .Z(n8057) );
  NAND U8622 ( .A(n8058), .B(n8057), .Z(n8208) );
  NANDN U8623 ( .A(n8060), .B(n8059), .Z(n8064) );
  NAND U8624 ( .A(n8062), .B(n8061), .Z(n8063) );
  NAND U8625 ( .A(n8064), .B(n8063), .Z(n8209) );
  XNOR U8626 ( .A(n8208), .B(n8209), .Z(n8210) );
  XOR U8627 ( .A(n8211), .B(n8210), .Z(n8088) );
  NANDN U8628 ( .A(n8070), .B(n8069), .Z(n8074) );
  NANDN U8629 ( .A(n8072), .B(n8071), .Z(n8073) );
  NAND U8630 ( .A(n8074), .B(n8073), .Z(n8087) );
  XNOR U8631 ( .A(n8086), .B(n8087), .Z(n8089) );
  XOR U8632 ( .A(n8088), .B(n8089), .Z(n8080) );
  XOR U8633 ( .A(n8081), .B(n8080), .Z(n8082) );
  XNOR U8634 ( .A(n8083), .B(n8082), .Z(n8220) );
  XNOR U8635 ( .A(n8220), .B(sreg[163]), .Z(n8222) );
  NAND U8636 ( .A(n8075), .B(sreg[162]), .Z(n8079) );
  OR U8637 ( .A(n8077), .B(n8076), .Z(n8078) );
  AND U8638 ( .A(n8079), .B(n8078), .Z(n8221) );
  XOR U8639 ( .A(n8222), .B(n8221), .Z(c[163]) );
  NAND U8640 ( .A(n8081), .B(n8080), .Z(n8085) );
  NAND U8641 ( .A(n8083), .B(n8082), .Z(n8084) );
  NAND U8642 ( .A(n8085), .B(n8084), .Z(n8228) );
  NANDN U8643 ( .A(n8087), .B(n8086), .Z(n8091) );
  NAND U8644 ( .A(n8089), .B(n8088), .Z(n8090) );
  NAND U8645 ( .A(n8091), .B(n8090), .Z(n8225) );
  NAND U8646 ( .A(n8093), .B(n8092), .Z(n8097) );
  NANDN U8647 ( .A(n8095), .B(n8094), .Z(n8096) );
  NAND U8648 ( .A(n8097), .B(n8096), .Z(n8357) );
  XNOR U8649 ( .A(n8357), .B(n8358), .Z(n8359) );
  NANDN U8650 ( .A(n8103), .B(n8102), .Z(n8107) );
  NANDN U8651 ( .A(n8105), .B(n8104), .Z(n8106) );
  NAND U8652 ( .A(n8107), .B(n8106), .Z(n8348) );
  OR U8653 ( .A(n8109), .B(n8108), .Z(n8113) );
  NAND U8654 ( .A(n8111), .B(n8110), .Z(n8112) );
  NAND U8655 ( .A(n8113), .B(n8112), .Z(n8287) );
  OR U8656 ( .A(n8115), .B(n8114), .Z(n8119) );
  NANDN U8657 ( .A(n8117), .B(n8116), .Z(n8118) );
  NAND U8658 ( .A(n8119), .B(n8118), .Z(n8286) );
  OR U8659 ( .A(n8121), .B(n8120), .Z(n8125) );
  NANDN U8660 ( .A(n8123), .B(n8122), .Z(n8124) );
  NAND U8661 ( .A(n8125), .B(n8124), .Z(n8285) );
  XOR U8662 ( .A(n8287), .B(n8288), .Z(n8345) );
  NANDN U8663 ( .A(n8127), .B(n8126), .Z(n8131) );
  NAND U8664 ( .A(n8129), .B(n8128), .Z(n8130) );
  NAND U8665 ( .A(n8131), .B(n8130), .Z(n8300) );
  NANDN U8666 ( .A(n8132), .B(n18832), .Z(n8134) );
  XNOR U8667 ( .A(b[19]), .B(a[50]), .Z(n8243) );
  NANDN U8668 ( .A(n8243), .B(n18834), .Z(n8133) );
  NAND U8669 ( .A(n8134), .B(n8133), .Z(n8312) );
  XOR U8670 ( .A(b[27]), .B(n9080), .Z(n8246) );
  NANDN U8671 ( .A(n8246), .B(n19336), .Z(n8137) );
  NANDN U8672 ( .A(n8135), .B(n19337), .Z(n8136) );
  NAND U8673 ( .A(n8137), .B(n8136), .Z(n8309) );
  XOR U8674 ( .A(b[5]), .B(a[64]), .Z(n8249) );
  NAND U8675 ( .A(n8249), .B(n17310), .Z(n8140) );
  NAND U8676 ( .A(n8138), .B(n17311), .Z(n8139) );
  AND U8677 ( .A(n8140), .B(n8139), .Z(n8310) );
  XNOR U8678 ( .A(n8309), .B(n8310), .Z(n8311) );
  XNOR U8679 ( .A(n8312), .B(n8311), .Z(n8298) );
  XOR U8680 ( .A(b[17]), .B(a[52]), .Z(n8252) );
  NAND U8681 ( .A(n8252), .B(n18673), .Z(n8143) );
  NAND U8682 ( .A(n8141), .B(n18674), .Z(n8142) );
  NAND U8683 ( .A(n8143), .B(n8142), .Z(n8270) );
  XOR U8684 ( .A(b[31]), .B(n8490), .Z(n8255) );
  NANDN U8685 ( .A(n8255), .B(n19472), .Z(n8146) );
  NANDN U8686 ( .A(n8144), .B(n19473), .Z(n8145) );
  NAND U8687 ( .A(n8146), .B(n8145), .Z(n8267) );
  OR U8688 ( .A(n8147), .B(n16988), .Z(n8149) );
  XNOR U8689 ( .A(b[3]), .B(a[66]), .Z(n8258) );
  NANDN U8690 ( .A(n8258), .B(n16990), .Z(n8148) );
  AND U8691 ( .A(n8149), .B(n8148), .Z(n8268) );
  XNOR U8692 ( .A(n8267), .B(n8268), .Z(n8269) );
  XOR U8693 ( .A(n8270), .B(n8269), .Z(n8297) );
  XNOR U8694 ( .A(n8298), .B(n8297), .Z(n8299) );
  XNOR U8695 ( .A(n8300), .B(n8299), .Z(n8346) );
  XNOR U8696 ( .A(n8345), .B(n8346), .Z(n8347) );
  XNOR U8697 ( .A(n8348), .B(n8347), .Z(n8366) );
  NANDN U8698 ( .A(n8155), .B(n8154), .Z(n8159) );
  NANDN U8699 ( .A(n8157), .B(n8156), .Z(n8158) );
  NAND U8700 ( .A(n8159), .B(n8158), .Z(n8353) );
  OR U8701 ( .A(n8161), .B(n8160), .Z(n8165) );
  NAND U8702 ( .A(n8163), .B(n8162), .Z(n8164) );
  NAND U8703 ( .A(n8165), .B(n8164), .Z(n8352) );
  NANDN U8704 ( .A(n8167), .B(n8166), .Z(n8171) );
  NAND U8705 ( .A(n8169), .B(n8168), .Z(n8170) );
  NAND U8706 ( .A(n8171), .B(n8170), .Z(n8291) );
  NANDN U8707 ( .A(n8173), .B(n8172), .Z(n8177) );
  NAND U8708 ( .A(n8175), .B(n8174), .Z(n8176) );
  AND U8709 ( .A(n8177), .B(n8176), .Z(n8292) );
  XNOR U8710 ( .A(n8291), .B(n8292), .Z(n8293) );
  XNOR U8711 ( .A(n579), .B(a[60]), .Z(n8315) );
  NAND U8712 ( .A(n17814), .B(n8315), .Z(n8180) );
  NANDN U8713 ( .A(n8178), .B(n17815), .Z(n8179) );
  NAND U8714 ( .A(n8180), .B(n8179), .Z(n8275) );
  NANDN U8715 ( .A(n8181), .B(n18513), .Z(n8183) );
  XOR U8716 ( .A(b[15]), .B(a[54]), .Z(n8318) );
  NANDN U8717 ( .A(n18512), .B(n8318), .Z(n8182) );
  AND U8718 ( .A(n8183), .B(n8182), .Z(n8273) );
  NANDN U8719 ( .A(n8184), .B(n19013), .Z(n8186) );
  XNOR U8720 ( .A(n582), .B(a[48]), .Z(n8321) );
  NAND U8721 ( .A(n8321), .B(n19015), .Z(n8185) );
  AND U8722 ( .A(n8186), .B(n8185), .Z(n8274) );
  XOR U8723 ( .A(n8275), .B(n8276), .Z(n8264) );
  XNOR U8724 ( .A(b[11]), .B(a[58]), .Z(n8324) );
  OR U8725 ( .A(n8324), .B(n18194), .Z(n8189) );
  NANDN U8726 ( .A(n8187), .B(n18104), .Z(n8188) );
  NAND U8727 ( .A(n8189), .B(n8188), .Z(n8262) );
  XOR U8728 ( .A(n580), .B(a[56]), .Z(n8327) );
  NANDN U8729 ( .A(n8327), .B(n18336), .Z(n8192) );
  NANDN U8730 ( .A(n8190), .B(n18337), .Z(n8191) );
  AND U8731 ( .A(n8192), .B(n8191), .Z(n8261) );
  XNOR U8732 ( .A(n8262), .B(n8261), .Z(n8263) );
  XOR U8733 ( .A(n8264), .B(n8263), .Z(n8281) );
  NANDN U8734 ( .A(n577), .B(a[68]), .Z(n8193) );
  XOR U8735 ( .A(n17151), .B(n8193), .Z(n8195) );
  NANDN U8736 ( .A(b[0]), .B(a[67]), .Z(n8194) );
  AND U8737 ( .A(n8195), .B(n8194), .Z(n8239) );
  NAND U8738 ( .A(n19406), .B(n8196), .Z(n8198) );
  XNOR U8739 ( .A(n584), .B(a[40]), .Z(n8333) );
  NANDN U8740 ( .A(n576), .B(n8333), .Z(n8197) );
  NAND U8741 ( .A(n8198), .B(n8197), .Z(n8237) );
  NANDN U8742 ( .A(n585), .B(a[36]), .Z(n8238) );
  XNOR U8743 ( .A(n8237), .B(n8238), .Z(n8240) );
  XOR U8744 ( .A(n8239), .B(n8240), .Z(n8279) );
  XOR U8745 ( .A(b[23]), .B(a[46]), .Z(n8336) );
  NANDN U8746 ( .A(n19127), .B(n8336), .Z(n8201) );
  NAND U8747 ( .A(n8199), .B(n19128), .Z(n8200) );
  NAND U8748 ( .A(n8201), .B(n8200), .Z(n8306) );
  NAND U8749 ( .A(n8202), .B(n17553), .Z(n8204) );
  XOR U8750 ( .A(b[7]), .B(a[62]), .Z(n8339) );
  NAND U8751 ( .A(n8339), .B(n17555), .Z(n8203) );
  NAND U8752 ( .A(n8204), .B(n8203), .Z(n8303) );
  XOR U8753 ( .A(b[25]), .B(a[44]), .Z(n8342) );
  NAND U8754 ( .A(n8342), .B(n19240), .Z(n8207) );
  NAND U8755 ( .A(n8205), .B(n19242), .Z(n8206) );
  AND U8756 ( .A(n8207), .B(n8206), .Z(n8304) );
  XNOR U8757 ( .A(n8303), .B(n8304), .Z(n8305) );
  XNOR U8758 ( .A(n8306), .B(n8305), .Z(n8280) );
  XOR U8759 ( .A(n8279), .B(n8280), .Z(n8282) );
  XNOR U8760 ( .A(n8281), .B(n8282), .Z(n8294) );
  XNOR U8761 ( .A(n8293), .B(n8294), .Z(n8351) );
  XNOR U8762 ( .A(n8352), .B(n8351), .Z(n8354) );
  XNOR U8763 ( .A(n8353), .B(n8354), .Z(n8363) );
  XNOR U8764 ( .A(n8364), .B(n8363), .Z(n8365) );
  XOR U8765 ( .A(n8366), .B(n8365), .Z(n8360) );
  XOR U8766 ( .A(n8359), .B(n8360), .Z(n8234) );
  NANDN U8767 ( .A(n8209), .B(n8208), .Z(n8213) );
  NAND U8768 ( .A(n8211), .B(n8210), .Z(n8212) );
  NAND U8769 ( .A(n8213), .B(n8212), .Z(n8231) );
  NANDN U8770 ( .A(n8215), .B(n8214), .Z(n8219) );
  OR U8771 ( .A(n8217), .B(n8216), .Z(n8218) );
  NAND U8772 ( .A(n8219), .B(n8218), .Z(n8232) );
  XNOR U8773 ( .A(n8231), .B(n8232), .Z(n8233) );
  XNOR U8774 ( .A(n8234), .B(n8233), .Z(n8226) );
  XNOR U8775 ( .A(n8225), .B(n8226), .Z(n8227) );
  XNOR U8776 ( .A(n8228), .B(n8227), .Z(n8369) );
  XNOR U8777 ( .A(n8369), .B(sreg[164]), .Z(n8371) );
  NAND U8778 ( .A(n8220), .B(sreg[163]), .Z(n8224) );
  OR U8779 ( .A(n8222), .B(n8221), .Z(n8223) );
  AND U8780 ( .A(n8224), .B(n8223), .Z(n8370) );
  XOR U8781 ( .A(n8371), .B(n8370), .Z(c[164]) );
  NANDN U8782 ( .A(n8226), .B(n8225), .Z(n8230) );
  NAND U8783 ( .A(n8228), .B(n8227), .Z(n8229) );
  NAND U8784 ( .A(n8230), .B(n8229), .Z(n8377) );
  NANDN U8785 ( .A(n8232), .B(n8231), .Z(n8236) );
  NAND U8786 ( .A(n8234), .B(n8233), .Z(n8235) );
  NAND U8787 ( .A(n8236), .B(n8235), .Z(n8375) );
  NANDN U8788 ( .A(n8238), .B(n8237), .Z(n8242) );
  NAND U8789 ( .A(n8240), .B(n8239), .Z(n8241) );
  NAND U8790 ( .A(n8242), .B(n8241), .Z(n8459) );
  NANDN U8791 ( .A(n8243), .B(n18832), .Z(n8245) );
  XNOR U8792 ( .A(b[19]), .B(a[51]), .Z(n8404) );
  NANDN U8793 ( .A(n8404), .B(n18834), .Z(n8244) );
  NAND U8794 ( .A(n8245), .B(n8244), .Z(n8469) );
  XNOR U8795 ( .A(b[27]), .B(a[43]), .Z(n8407) );
  NANDN U8796 ( .A(n8407), .B(n19336), .Z(n8248) );
  NANDN U8797 ( .A(n8246), .B(n19337), .Z(n8247) );
  NAND U8798 ( .A(n8248), .B(n8247), .Z(n8466) );
  XNOR U8799 ( .A(b[5]), .B(a[65]), .Z(n8410) );
  NANDN U8800 ( .A(n8410), .B(n17310), .Z(n8251) );
  NAND U8801 ( .A(n8249), .B(n17311), .Z(n8250) );
  AND U8802 ( .A(n8251), .B(n8250), .Z(n8467) );
  XNOR U8803 ( .A(n8466), .B(n8467), .Z(n8468) );
  XNOR U8804 ( .A(n8469), .B(n8468), .Z(n8457) );
  XNOR U8805 ( .A(b[17]), .B(a[53]), .Z(n8413) );
  NANDN U8806 ( .A(n8413), .B(n18673), .Z(n8254) );
  NAND U8807 ( .A(n8252), .B(n18674), .Z(n8253) );
  NAND U8808 ( .A(n8254), .B(n8253), .Z(n8431) );
  XNOR U8809 ( .A(b[31]), .B(a[39]), .Z(n8416) );
  NANDN U8810 ( .A(n8416), .B(n19472), .Z(n8257) );
  NANDN U8811 ( .A(n8255), .B(n19473), .Z(n8256) );
  NAND U8812 ( .A(n8257), .B(n8256), .Z(n8428) );
  OR U8813 ( .A(n8258), .B(n16988), .Z(n8260) );
  XNOR U8814 ( .A(b[3]), .B(a[67]), .Z(n8419) );
  NANDN U8815 ( .A(n8419), .B(n16990), .Z(n8259) );
  AND U8816 ( .A(n8260), .B(n8259), .Z(n8429) );
  XNOR U8817 ( .A(n8428), .B(n8429), .Z(n8430) );
  XOR U8818 ( .A(n8431), .B(n8430), .Z(n8456) );
  XNOR U8819 ( .A(n8457), .B(n8456), .Z(n8458) );
  XNOR U8820 ( .A(n8459), .B(n8458), .Z(n8503) );
  NANDN U8821 ( .A(n8262), .B(n8261), .Z(n8266) );
  NAND U8822 ( .A(n8264), .B(n8263), .Z(n8265) );
  NAND U8823 ( .A(n8266), .B(n8265), .Z(n8447) );
  NANDN U8824 ( .A(n8268), .B(n8267), .Z(n8272) );
  NAND U8825 ( .A(n8270), .B(n8269), .Z(n8271) );
  NAND U8826 ( .A(n8272), .B(n8271), .Z(n8445) );
  OR U8827 ( .A(n8274), .B(n8273), .Z(n8278) );
  NANDN U8828 ( .A(n8276), .B(n8275), .Z(n8277) );
  NAND U8829 ( .A(n8278), .B(n8277), .Z(n8444) );
  XNOR U8830 ( .A(n8447), .B(n8446), .Z(n8504) );
  XOR U8831 ( .A(n8503), .B(n8504), .Z(n8506) );
  NANDN U8832 ( .A(n8280), .B(n8279), .Z(n8284) );
  OR U8833 ( .A(n8282), .B(n8281), .Z(n8283) );
  NAND U8834 ( .A(n8284), .B(n8283), .Z(n8505) );
  XOR U8835 ( .A(n8506), .B(n8505), .Z(n8394) );
  OR U8836 ( .A(n8286), .B(n8285), .Z(n8290) );
  NANDN U8837 ( .A(n8288), .B(n8287), .Z(n8289) );
  NAND U8838 ( .A(n8290), .B(n8289), .Z(n8393) );
  NANDN U8839 ( .A(n8292), .B(n8291), .Z(n8296) );
  NANDN U8840 ( .A(n8294), .B(n8293), .Z(n8295) );
  NAND U8841 ( .A(n8296), .B(n8295), .Z(n8511) );
  NANDN U8842 ( .A(n8298), .B(n8297), .Z(n8302) );
  NAND U8843 ( .A(n8300), .B(n8299), .Z(n8301) );
  NAND U8844 ( .A(n8302), .B(n8301), .Z(n8510) );
  NANDN U8845 ( .A(n8304), .B(n8303), .Z(n8308) );
  NAND U8846 ( .A(n8306), .B(n8305), .Z(n8307) );
  NAND U8847 ( .A(n8308), .B(n8307), .Z(n8450) );
  NANDN U8848 ( .A(n8310), .B(n8309), .Z(n8314) );
  NAND U8849 ( .A(n8312), .B(n8311), .Z(n8313) );
  AND U8850 ( .A(n8314), .B(n8313), .Z(n8451) );
  XNOR U8851 ( .A(n8450), .B(n8451), .Z(n8452) );
  XNOR U8852 ( .A(b[9]), .B(a[61]), .Z(n8472) );
  NANDN U8853 ( .A(n8472), .B(n17814), .Z(n8317) );
  NAND U8854 ( .A(n17815), .B(n8315), .Z(n8316) );
  NAND U8855 ( .A(n8317), .B(n8316), .Z(n8436) );
  XNOR U8856 ( .A(b[15]), .B(a[55]), .Z(n8475) );
  OR U8857 ( .A(n8475), .B(n18512), .Z(n8320) );
  NAND U8858 ( .A(n8318), .B(n18513), .Z(n8319) );
  NAND U8859 ( .A(n8320), .B(n8319), .Z(n8434) );
  XOR U8860 ( .A(b[21]), .B(n10083), .Z(n8478) );
  NANDN U8861 ( .A(n8478), .B(n19015), .Z(n8323) );
  NAND U8862 ( .A(n19013), .B(n8321), .Z(n8322) );
  NAND U8863 ( .A(n8323), .B(n8322), .Z(n8435) );
  XNOR U8864 ( .A(n8434), .B(n8435), .Z(n8437) );
  XOR U8865 ( .A(n8436), .B(n8437), .Z(n8425) );
  XNOR U8866 ( .A(b[11]), .B(a[59]), .Z(n8481) );
  OR U8867 ( .A(n8481), .B(n18194), .Z(n8326) );
  NANDN U8868 ( .A(n8324), .B(n18104), .Z(n8325) );
  NAND U8869 ( .A(n8326), .B(n8325), .Z(n8423) );
  XOR U8870 ( .A(n580), .B(a[57]), .Z(n8484) );
  NANDN U8871 ( .A(n8484), .B(n18336), .Z(n8329) );
  NANDN U8872 ( .A(n8327), .B(n18337), .Z(n8328) );
  AND U8873 ( .A(n8329), .B(n8328), .Z(n8422) );
  XNOR U8874 ( .A(n8423), .B(n8422), .Z(n8424) );
  XNOR U8875 ( .A(n8425), .B(n8424), .Z(n8441) );
  NANDN U8876 ( .A(n577), .B(a[69]), .Z(n8330) );
  XOR U8877 ( .A(n17151), .B(n8330), .Z(n8332) );
  NANDN U8878 ( .A(b[0]), .B(a[68]), .Z(n8331) );
  AND U8879 ( .A(n8332), .B(n8331), .Z(n8400) );
  NAND U8880 ( .A(n19406), .B(n8333), .Z(n8335) );
  XOR U8881 ( .A(b[29]), .B(n8930), .Z(n8491) );
  OR U8882 ( .A(n8491), .B(n576), .Z(n8334) );
  NAND U8883 ( .A(n8335), .B(n8334), .Z(n8398) );
  NANDN U8884 ( .A(n585), .B(a[37]), .Z(n8399) );
  XNOR U8885 ( .A(n8398), .B(n8399), .Z(n8401) );
  XNOR U8886 ( .A(n8400), .B(n8401), .Z(n8439) );
  XOR U8887 ( .A(b[23]), .B(a[47]), .Z(n8494) );
  NANDN U8888 ( .A(n19127), .B(n8494), .Z(n8338) );
  NAND U8889 ( .A(n8336), .B(n19128), .Z(n8337) );
  NAND U8890 ( .A(n8338), .B(n8337), .Z(n8463) );
  NAND U8891 ( .A(n8339), .B(n17553), .Z(n8341) );
  XOR U8892 ( .A(b[7]), .B(a[63]), .Z(n8497) );
  NAND U8893 ( .A(n8497), .B(n17555), .Z(n8340) );
  NAND U8894 ( .A(n8341), .B(n8340), .Z(n8460) );
  XOR U8895 ( .A(b[25]), .B(a[45]), .Z(n8500) );
  NAND U8896 ( .A(n8500), .B(n19240), .Z(n8344) );
  NAND U8897 ( .A(n8342), .B(n19242), .Z(n8343) );
  AND U8898 ( .A(n8344), .B(n8343), .Z(n8461) );
  XNOR U8899 ( .A(n8460), .B(n8461), .Z(n8462) );
  XOR U8900 ( .A(n8463), .B(n8462), .Z(n8438) );
  XOR U8901 ( .A(n8441), .B(n8440), .Z(n8453) );
  XOR U8902 ( .A(n8452), .B(n8453), .Z(n8509) );
  XNOR U8903 ( .A(n8510), .B(n8509), .Z(n8512) );
  XNOR U8904 ( .A(n8511), .B(n8512), .Z(n8392) );
  XOR U8905 ( .A(n8393), .B(n8392), .Z(n8395) );
  NANDN U8906 ( .A(n8346), .B(n8345), .Z(n8350) );
  NAND U8907 ( .A(n8348), .B(n8347), .Z(n8349) );
  NAND U8908 ( .A(n8350), .B(n8349), .Z(n8387) );
  NAND U8909 ( .A(n8352), .B(n8351), .Z(n8356) );
  NANDN U8910 ( .A(n8354), .B(n8353), .Z(n8355) );
  AND U8911 ( .A(n8356), .B(n8355), .Z(n8386) );
  XNOR U8912 ( .A(n8387), .B(n8386), .Z(n8388) );
  XOR U8913 ( .A(n8389), .B(n8388), .Z(n8382) );
  NANDN U8914 ( .A(n8358), .B(n8357), .Z(n8362) );
  NANDN U8915 ( .A(n8360), .B(n8359), .Z(n8361) );
  NAND U8916 ( .A(n8362), .B(n8361), .Z(n8381) );
  NANDN U8917 ( .A(n8364), .B(n8363), .Z(n8368) );
  NANDN U8918 ( .A(n8366), .B(n8365), .Z(n8367) );
  AND U8919 ( .A(n8368), .B(n8367), .Z(n8380) );
  XNOR U8920 ( .A(n8381), .B(n8380), .Z(n8383) );
  XOR U8921 ( .A(n8382), .B(n8383), .Z(n8374) );
  XOR U8922 ( .A(n8375), .B(n8374), .Z(n8376) );
  XNOR U8923 ( .A(n8377), .B(n8376), .Z(n8515) );
  XNOR U8924 ( .A(n8515), .B(sreg[165]), .Z(n8517) );
  NAND U8925 ( .A(n8369), .B(sreg[164]), .Z(n8373) );
  OR U8926 ( .A(n8371), .B(n8370), .Z(n8372) );
  AND U8927 ( .A(n8373), .B(n8372), .Z(n8516) );
  XOR U8928 ( .A(n8517), .B(n8516), .Z(c[165]) );
  NAND U8929 ( .A(n8375), .B(n8374), .Z(n8379) );
  NAND U8930 ( .A(n8377), .B(n8376), .Z(n8378) );
  NAND U8931 ( .A(n8379), .B(n8378), .Z(n8523) );
  NANDN U8932 ( .A(n8381), .B(n8380), .Z(n8385) );
  NAND U8933 ( .A(n8383), .B(n8382), .Z(n8384) );
  NAND U8934 ( .A(n8385), .B(n8384), .Z(n8521) );
  NANDN U8935 ( .A(n8387), .B(n8386), .Z(n8391) );
  NAND U8936 ( .A(n8389), .B(n8388), .Z(n8390) );
  NAND U8937 ( .A(n8391), .B(n8390), .Z(n8526) );
  NANDN U8938 ( .A(n8393), .B(n8392), .Z(n8397) );
  OR U8939 ( .A(n8395), .B(n8394), .Z(n8396) );
  NAND U8940 ( .A(n8397), .B(n8396), .Z(n8527) );
  XNOR U8941 ( .A(n8526), .B(n8527), .Z(n8528) );
  NANDN U8942 ( .A(n8399), .B(n8398), .Z(n8403) );
  NAND U8943 ( .A(n8401), .B(n8400), .Z(n8402) );
  NAND U8944 ( .A(n8403), .B(n8402), .Z(n8603) );
  NANDN U8945 ( .A(n8404), .B(n18832), .Z(n8406) );
  XNOR U8946 ( .A(b[19]), .B(a[52]), .Z(n8548) );
  NANDN U8947 ( .A(n8548), .B(n18834), .Z(n8405) );
  NAND U8948 ( .A(n8406), .B(n8405), .Z(n8613) );
  XNOR U8949 ( .A(b[27]), .B(a[44]), .Z(n8551) );
  NANDN U8950 ( .A(n8551), .B(n19336), .Z(n8409) );
  NANDN U8951 ( .A(n8407), .B(n19337), .Z(n8408) );
  NAND U8952 ( .A(n8409), .B(n8408), .Z(n8610) );
  XOR U8953 ( .A(b[5]), .B(a[66]), .Z(n8554) );
  NAND U8954 ( .A(n8554), .B(n17310), .Z(n8412) );
  NANDN U8955 ( .A(n8410), .B(n17311), .Z(n8411) );
  AND U8956 ( .A(n8412), .B(n8411), .Z(n8611) );
  XNOR U8957 ( .A(n8610), .B(n8611), .Z(n8612) );
  XNOR U8958 ( .A(n8613), .B(n8612), .Z(n8601) );
  XOR U8959 ( .A(b[17]), .B(a[54]), .Z(n8557) );
  NAND U8960 ( .A(n8557), .B(n18673), .Z(n8415) );
  NANDN U8961 ( .A(n8413), .B(n18674), .Z(n8414) );
  NAND U8962 ( .A(n8415), .B(n8414), .Z(n8575) );
  XNOR U8963 ( .A(b[31]), .B(a[40]), .Z(n8560) );
  NANDN U8964 ( .A(n8560), .B(n19472), .Z(n8418) );
  NANDN U8965 ( .A(n8416), .B(n19473), .Z(n8417) );
  NAND U8966 ( .A(n8418), .B(n8417), .Z(n8572) );
  OR U8967 ( .A(n8419), .B(n16988), .Z(n8421) );
  XNOR U8968 ( .A(b[3]), .B(a[68]), .Z(n8563) );
  NANDN U8969 ( .A(n8563), .B(n16990), .Z(n8420) );
  AND U8970 ( .A(n8421), .B(n8420), .Z(n8573) );
  XNOR U8971 ( .A(n8572), .B(n8573), .Z(n8574) );
  XOR U8972 ( .A(n8575), .B(n8574), .Z(n8600) );
  XNOR U8973 ( .A(n8601), .B(n8600), .Z(n8602) );
  XNOR U8974 ( .A(n8603), .B(n8602), .Z(n8539) );
  NANDN U8975 ( .A(n8423), .B(n8422), .Z(n8427) );
  NAND U8976 ( .A(n8425), .B(n8424), .Z(n8426) );
  NAND U8977 ( .A(n8427), .B(n8426), .Z(n8592) );
  NANDN U8978 ( .A(n8429), .B(n8428), .Z(n8433) );
  NAND U8979 ( .A(n8431), .B(n8430), .Z(n8432) );
  NAND U8980 ( .A(n8433), .B(n8432), .Z(n8591) );
  XNOR U8981 ( .A(n8591), .B(n8590), .Z(n8593) );
  XOR U8982 ( .A(n8592), .B(n8593), .Z(n8538) );
  XOR U8983 ( .A(n8539), .B(n8538), .Z(n8540) );
  NANDN U8984 ( .A(n8439), .B(n8438), .Z(n8443) );
  NAND U8985 ( .A(n8441), .B(n8440), .Z(n8442) );
  NAND U8986 ( .A(n8443), .B(n8442), .Z(n8541) );
  XNOR U8987 ( .A(n8540), .B(n8541), .Z(n8654) );
  OR U8988 ( .A(n8445), .B(n8444), .Z(n8449) );
  NAND U8989 ( .A(n8447), .B(n8446), .Z(n8448) );
  NAND U8990 ( .A(n8449), .B(n8448), .Z(n8653) );
  NANDN U8991 ( .A(n8451), .B(n8450), .Z(n8455) );
  NAND U8992 ( .A(n8453), .B(n8452), .Z(n8454) );
  NAND U8993 ( .A(n8455), .B(n8454), .Z(n8534) );
  NANDN U8994 ( .A(n8461), .B(n8460), .Z(n8465) );
  NAND U8995 ( .A(n8463), .B(n8462), .Z(n8464) );
  NAND U8996 ( .A(n8465), .B(n8464), .Z(n8594) );
  NANDN U8997 ( .A(n8467), .B(n8466), .Z(n8471) );
  NAND U8998 ( .A(n8469), .B(n8468), .Z(n8470) );
  AND U8999 ( .A(n8471), .B(n8470), .Z(n8595) );
  XNOR U9000 ( .A(n8594), .B(n8595), .Z(n8596) );
  XNOR U9001 ( .A(b[9]), .B(a[62]), .Z(n8616) );
  NANDN U9002 ( .A(n8616), .B(n17814), .Z(n8474) );
  NANDN U9003 ( .A(n8472), .B(n17815), .Z(n8473) );
  NAND U9004 ( .A(n8474), .B(n8473), .Z(n8580) );
  NANDN U9005 ( .A(n8475), .B(n18513), .Z(n8477) );
  XOR U9006 ( .A(b[15]), .B(a[56]), .Z(n8619) );
  NANDN U9007 ( .A(n18512), .B(n8619), .Z(n8476) );
  AND U9008 ( .A(n8477), .B(n8476), .Z(n8578) );
  NANDN U9009 ( .A(n8478), .B(n19013), .Z(n8480) );
  XNOR U9010 ( .A(b[21]), .B(a[50]), .Z(n8622) );
  NANDN U9011 ( .A(n8622), .B(n19015), .Z(n8479) );
  AND U9012 ( .A(n8480), .B(n8479), .Z(n8579) );
  XOR U9013 ( .A(n8580), .B(n8581), .Z(n8569) );
  XNOR U9014 ( .A(b[11]), .B(a[60]), .Z(n8625) );
  OR U9015 ( .A(n8625), .B(n18194), .Z(n8483) );
  NANDN U9016 ( .A(n8481), .B(n18104), .Z(n8482) );
  NAND U9017 ( .A(n8483), .B(n8482), .Z(n8567) );
  XOR U9018 ( .A(n580), .B(a[58]), .Z(n8628) );
  NANDN U9019 ( .A(n8628), .B(n18336), .Z(n8486) );
  NANDN U9020 ( .A(n8484), .B(n18337), .Z(n8485) );
  AND U9021 ( .A(n8486), .B(n8485), .Z(n8566) );
  XNOR U9022 ( .A(n8567), .B(n8566), .Z(n8568) );
  XOR U9023 ( .A(n8569), .B(n8568), .Z(n8586) );
  NANDN U9024 ( .A(n577), .B(a[70]), .Z(n8487) );
  XOR U9025 ( .A(n17151), .B(n8487), .Z(n8489) );
  NANDN U9026 ( .A(b[0]), .B(a[69]), .Z(n8488) );
  AND U9027 ( .A(n8489), .B(n8488), .Z(n8545) );
  ANDN U9028 ( .B(b[31]), .A(n8490), .Z(n8542) );
  NANDN U9029 ( .A(n8491), .B(n19406), .Z(n8493) );
  XNOR U9030 ( .A(n584), .B(a[42]), .Z(n8634) );
  NANDN U9031 ( .A(n576), .B(n8634), .Z(n8492) );
  NAND U9032 ( .A(n8493), .B(n8492), .Z(n8543) );
  XOR U9033 ( .A(n8542), .B(n8543), .Z(n8544) );
  XNOR U9034 ( .A(n8545), .B(n8544), .Z(n8584) );
  XOR U9035 ( .A(b[23]), .B(a[48]), .Z(n8637) );
  NANDN U9036 ( .A(n19127), .B(n8637), .Z(n8496) );
  NAND U9037 ( .A(n8494), .B(n19128), .Z(n8495) );
  NAND U9038 ( .A(n8496), .B(n8495), .Z(n8607) );
  NAND U9039 ( .A(n8497), .B(n17553), .Z(n8499) );
  XOR U9040 ( .A(b[7]), .B(a[64]), .Z(n8640) );
  NAND U9041 ( .A(n8640), .B(n17555), .Z(n8498) );
  NAND U9042 ( .A(n8499), .B(n8498), .Z(n8604) );
  XOR U9043 ( .A(b[25]), .B(a[46]), .Z(n8643) );
  NAND U9044 ( .A(n8643), .B(n19240), .Z(n8502) );
  NAND U9045 ( .A(n8500), .B(n19242), .Z(n8501) );
  AND U9046 ( .A(n8502), .B(n8501), .Z(n8605) );
  XNOR U9047 ( .A(n8604), .B(n8605), .Z(n8606) );
  XNOR U9048 ( .A(n8607), .B(n8606), .Z(n8585) );
  XNOR U9049 ( .A(n8584), .B(n8585), .Z(n8587) );
  XNOR U9050 ( .A(n8586), .B(n8587), .Z(n8597) );
  XNOR U9051 ( .A(n8596), .B(n8597), .Z(n8532) );
  XNOR U9052 ( .A(n8533), .B(n8532), .Z(n8535) );
  XNOR U9053 ( .A(n8534), .B(n8535), .Z(n8652) );
  XOR U9054 ( .A(n8653), .B(n8652), .Z(n8655) );
  NANDN U9055 ( .A(n8504), .B(n8503), .Z(n8508) );
  OR U9056 ( .A(n8506), .B(n8505), .Z(n8507) );
  NAND U9057 ( .A(n8508), .B(n8507), .Z(n8646) );
  NAND U9058 ( .A(n8510), .B(n8509), .Z(n8514) );
  NANDN U9059 ( .A(n8512), .B(n8511), .Z(n8513) );
  NAND U9060 ( .A(n8514), .B(n8513), .Z(n8647) );
  XNOR U9061 ( .A(n8646), .B(n8647), .Z(n8648) );
  XOR U9062 ( .A(n8649), .B(n8648), .Z(n8529) );
  XOR U9063 ( .A(n8528), .B(n8529), .Z(n8520) );
  XOR U9064 ( .A(n8521), .B(n8520), .Z(n8522) );
  XNOR U9065 ( .A(n8523), .B(n8522), .Z(n8658) );
  XNOR U9066 ( .A(n8658), .B(sreg[166]), .Z(n8660) );
  NAND U9067 ( .A(n8515), .B(sreg[165]), .Z(n8519) );
  OR U9068 ( .A(n8517), .B(n8516), .Z(n8518) );
  AND U9069 ( .A(n8519), .B(n8518), .Z(n8659) );
  XOR U9070 ( .A(n8660), .B(n8659), .Z(c[166]) );
  NAND U9071 ( .A(n8521), .B(n8520), .Z(n8525) );
  NAND U9072 ( .A(n8523), .B(n8522), .Z(n8524) );
  NAND U9073 ( .A(n8525), .B(n8524), .Z(n8666) );
  NANDN U9074 ( .A(n8527), .B(n8526), .Z(n8531) );
  NAND U9075 ( .A(n8529), .B(n8528), .Z(n8530) );
  NAND U9076 ( .A(n8531), .B(n8530), .Z(n8663) );
  NAND U9077 ( .A(n8533), .B(n8532), .Z(n8537) );
  NANDN U9078 ( .A(n8535), .B(n8534), .Z(n8536) );
  NAND U9079 ( .A(n8537), .B(n8536), .Z(n8675) );
  XNOR U9080 ( .A(n8675), .B(n8676), .Z(n8677) );
  OR U9081 ( .A(n8543), .B(n8542), .Z(n8547) );
  NANDN U9082 ( .A(n8545), .B(n8544), .Z(n8546) );
  NAND U9083 ( .A(n8547), .B(n8546), .Z(n8749) );
  NANDN U9084 ( .A(n8548), .B(n18832), .Z(n8550) );
  XOR U9085 ( .A(b[19]), .B(n10660), .Z(n8693) );
  NANDN U9086 ( .A(n8693), .B(n18834), .Z(n8549) );
  NAND U9087 ( .A(n8550), .B(n8549), .Z(n8762) );
  XNOR U9088 ( .A(b[27]), .B(a[45]), .Z(n8696) );
  NANDN U9089 ( .A(n8696), .B(n19336), .Z(n8553) );
  NANDN U9090 ( .A(n8551), .B(n19337), .Z(n8552) );
  NAND U9091 ( .A(n8553), .B(n8552), .Z(n8759) );
  XOR U9092 ( .A(b[5]), .B(a[67]), .Z(n8699) );
  NAND U9093 ( .A(n8699), .B(n17310), .Z(n8556) );
  NAND U9094 ( .A(n8554), .B(n17311), .Z(n8555) );
  AND U9095 ( .A(n8556), .B(n8555), .Z(n8760) );
  XNOR U9096 ( .A(n8759), .B(n8760), .Z(n8761) );
  XNOR U9097 ( .A(n8762), .B(n8761), .Z(n8748) );
  XNOR U9098 ( .A(b[17]), .B(a[55]), .Z(n8702) );
  NANDN U9099 ( .A(n8702), .B(n18673), .Z(n8559) );
  NAND U9100 ( .A(n8557), .B(n18674), .Z(n8558) );
  NAND U9101 ( .A(n8559), .B(n8558), .Z(n8720) );
  XOR U9102 ( .A(b[31]), .B(n8930), .Z(n8705) );
  NANDN U9103 ( .A(n8705), .B(n19472), .Z(n8562) );
  NANDN U9104 ( .A(n8560), .B(n19473), .Z(n8561) );
  NAND U9105 ( .A(n8562), .B(n8561), .Z(n8717) );
  OR U9106 ( .A(n8563), .B(n16988), .Z(n8565) );
  XNOR U9107 ( .A(b[3]), .B(a[69]), .Z(n8708) );
  NANDN U9108 ( .A(n8708), .B(n16990), .Z(n8564) );
  AND U9109 ( .A(n8565), .B(n8564), .Z(n8718) );
  XNOR U9110 ( .A(n8717), .B(n8718), .Z(n8719) );
  XOR U9111 ( .A(n8720), .B(n8719), .Z(n8747) );
  XOR U9112 ( .A(n8748), .B(n8747), .Z(n8750) );
  XNOR U9113 ( .A(n8749), .B(n8750), .Z(n8795) );
  NANDN U9114 ( .A(n8567), .B(n8566), .Z(n8571) );
  NAND U9115 ( .A(n8569), .B(n8568), .Z(n8570) );
  NAND U9116 ( .A(n8571), .B(n8570), .Z(n8738) );
  NANDN U9117 ( .A(n8573), .B(n8572), .Z(n8577) );
  NAND U9118 ( .A(n8575), .B(n8574), .Z(n8576) );
  NAND U9119 ( .A(n8577), .B(n8576), .Z(n8736) );
  OR U9120 ( .A(n8579), .B(n8578), .Z(n8583) );
  NANDN U9121 ( .A(n8581), .B(n8580), .Z(n8582) );
  NAND U9122 ( .A(n8583), .B(n8582), .Z(n8735) );
  XNOR U9123 ( .A(n8738), .B(n8737), .Z(n8796) );
  XNOR U9124 ( .A(n8795), .B(n8796), .Z(n8797) );
  OR U9125 ( .A(n8585), .B(n8584), .Z(n8589) );
  OR U9126 ( .A(n8587), .B(n8586), .Z(n8588) );
  AND U9127 ( .A(n8589), .B(n8588), .Z(n8798) );
  XOR U9128 ( .A(n8797), .B(n8798), .Z(n8683) );
  NANDN U9129 ( .A(n8595), .B(n8594), .Z(n8599) );
  NANDN U9130 ( .A(n8597), .B(n8596), .Z(n8598) );
  NAND U9131 ( .A(n8599), .B(n8598), .Z(n8804) );
  NANDN U9132 ( .A(n8605), .B(n8604), .Z(n8609) );
  NAND U9133 ( .A(n8607), .B(n8606), .Z(n8608) );
  NAND U9134 ( .A(n8609), .B(n8608), .Z(n8741) );
  NANDN U9135 ( .A(n8611), .B(n8610), .Z(n8615) );
  NAND U9136 ( .A(n8613), .B(n8612), .Z(n8614) );
  AND U9137 ( .A(n8615), .B(n8614), .Z(n8742) );
  XNOR U9138 ( .A(n8741), .B(n8742), .Z(n8743) );
  XNOR U9139 ( .A(b[9]), .B(a[63]), .Z(n8765) );
  NANDN U9140 ( .A(n8765), .B(n17814), .Z(n8618) );
  NANDN U9141 ( .A(n8616), .B(n17815), .Z(n8617) );
  NAND U9142 ( .A(n8618), .B(n8617), .Z(n8725) );
  NAND U9143 ( .A(n8619), .B(n18513), .Z(n8621) );
  XOR U9144 ( .A(b[15]), .B(a[57]), .Z(n8768) );
  NANDN U9145 ( .A(n18512), .B(n8768), .Z(n8620) );
  AND U9146 ( .A(n8621), .B(n8620), .Z(n8723) );
  NANDN U9147 ( .A(n8622), .B(n19013), .Z(n8624) );
  XNOR U9148 ( .A(b[21]), .B(a[51]), .Z(n8771) );
  NANDN U9149 ( .A(n8771), .B(n19015), .Z(n8623) );
  AND U9150 ( .A(n8624), .B(n8623), .Z(n8724) );
  XOR U9151 ( .A(n8725), .B(n8726), .Z(n8714) );
  XNOR U9152 ( .A(b[11]), .B(a[61]), .Z(n8774) );
  OR U9153 ( .A(n8774), .B(n18194), .Z(n8627) );
  NANDN U9154 ( .A(n8625), .B(n18104), .Z(n8626) );
  NAND U9155 ( .A(n8627), .B(n8626), .Z(n8712) );
  XOR U9156 ( .A(n580), .B(a[59]), .Z(n8777) );
  NANDN U9157 ( .A(n8777), .B(n18336), .Z(n8630) );
  NANDN U9158 ( .A(n8628), .B(n18337), .Z(n8629) );
  AND U9159 ( .A(n8630), .B(n8629), .Z(n8711) );
  XNOR U9160 ( .A(n8712), .B(n8711), .Z(n8713) );
  XOR U9161 ( .A(n8714), .B(n8713), .Z(n8731) );
  NANDN U9162 ( .A(n577), .B(a[71]), .Z(n8631) );
  XOR U9163 ( .A(n17151), .B(n8631), .Z(n8633) );
  NANDN U9164 ( .A(b[0]), .B(a[70]), .Z(n8632) );
  AND U9165 ( .A(n8633), .B(n8632), .Z(n8689) );
  NAND U9166 ( .A(n8634), .B(n19406), .Z(n8636) );
  XNOR U9167 ( .A(n584), .B(a[43]), .Z(n8783) );
  NANDN U9168 ( .A(n576), .B(n8783), .Z(n8635) );
  NAND U9169 ( .A(n8636), .B(n8635), .Z(n8687) );
  NANDN U9170 ( .A(n585), .B(a[39]), .Z(n8688) );
  XNOR U9171 ( .A(n8687), .B(n8688), .Z(n8690) );
  XOR U9172 ( .A(n8689), .B(n8690), .Z(n8729) );
  XNOR U9173 ( .A(b[23]), .B(a[49]), .Z(n8786) );
  OR U9174 ( .A(n8786), .B(n19127), .Z(n8639) );
  NAND U9175 ( .A(n8637), .B(n19128), .Z(n8638) );
  NAND U9176 ( .A(n8639), .B(n8638), .Z(n8756) );
  NAND U9177 ( .A(n8640), .B(n17553), .Z(n8642) );
  XNOR U9178 ( .A(b[7]), .B(a[65]), .Z(n8789) );
  NANDN U9179 ( .A(n8789), .B(n17555), .Z(n8641) );
  NAND U9180 ( .A(n8642), .B(n8641), .Z(n8753) );
  XOR U9181 ( .A(b[25]), .B(a[47]), .Z(n8792) );
  NAND U9182 ( .A(n8792), .B(n19240), .Z(n8645) );
  NAND U9183 ( .A(n8643), .B(n19242), .Z(n8644) );
  AND U9184 ( .A(n8645), .B(n8644), .Z(n8754) );
  XNOR U9185 ( .A(n8753), .B(n8754), .Z(n8755) );
  XNOR U9186 ( .A(n8756), .B(n8755), .Z(n8730) );
  XOR U9187 ( .A(n8729), .B(n8730), .Z(n8732) );
  XNOR U9188 ( .A(n8731), .B(n8732), .Z(n8744) );
  XOR U9189 ( .A(n8743), .B(n8744), .Z(n8802) );
  XNOR U9190 ( .A(n8801), .B(n8802), .Z(n8803) );
  XNOR U9191 ( .A(n8804), .B(n8803), .Z(n8681) );
  XNOR U9192 ( .A(n8682), .B(n8681), .Z(n8684) );
  XNOR U9193 ( .A(n8683), .B(n8684), .Z(n8678) );
  XOR U9194 ( .A(n8677), .B(n8678), .Z(n8672) );
  NANDN U9195 ( .A(n8647), .B(n8646), .Z(n8651) );
  NAND U9196 ( .A(n8649), .B(n8648), .Z(n8650) );
  NAND U9197 ( .A(n8651), .B(n8650), .Z(n8669) );
  NANDN U9198 ( .A(n8653), .B(n8652), .Z(n8657) );
  OR U9199 ( .A(n8655), .B(n8654), .Z(n8656) );
  NAND U9200 ( .A(n8657), .B(n8656), .Z(n8670) );
  XNOR U9201 ( .A(n8669), .B(n8670), .Z(n8671) );
  XNOR U9202 ( .A(n8672), .B(n8671), .Z(n8664) );
  XNOR U9203 ( .A(n8663), .B(n8664), .Z(n8665) );
  XNOR U9204 ( .A(n8666), .B(n8665), .Z(n8807) );
  XNOR U9205 ( .A(n8807), .B(sreg[167]), .Z(n8809) );
  NAND U9206 ( .A(n8658), .B(sreg[166]), .Z(n8662) );
  OR U9207 ( .A(n8660), .B(n8659), .Z(n8661) );
  AND U9208 ( .A(n8662), .B(n8661), .Z(n8808) );
  XOR U9209 ( .A(n8809), .B(n8808), .Z(c[167]) );
  NANDN U9210 ( .A(n8664), .B(n8663), .Z(n8668) );
  NAND U9211 ( .A(n8666), .B(n8665), .Z(n8667) );
  NAND U9212 ( .A(n8668), .B(n8667), .Z(n8815) );
  NANDN U9213 ( .A(n8670), .B(n8669), .Z(n8674) );
  NAND U9214 ( .A(n8672), .B(n8671), .Z(n8673) );
  NAND U9215 ( .A(n8674), .B(n8673), .Z(n8813) );
  NANDN U9216 ( .A(n8676), .B(n8675), .Z(n8680) );
  NANDN U9217 ( .A(n8678), .B(n8677), .Z(n8679) );
  NAND U9218 ( .A(n8680), .B(n8679), .Z(n8819) );
  OR U9219 ( .A(n8682), .B(n8681), .Z(n8686) );
  OR U9220 ( .A(n8684), .B(n8683), .Z(n8685) );
  AND U9221 ( .A(n8686), .B(n8685), .Z(n8818) );
  XNOR U9222 ( .A(n8819), .B(n8818), .Z(n8820) );
  NANDN U9223 ( .A(n8688), .B(n8687), .Z(n8692) );
  NAND U9224 ( .A(n8690), .B(n8689), .Z(n8691) );
  NAND U9225 ( .A(n8692), .B(n8691), .Z(n8899) );
  NANDN U9226 ( .A(n8693), .B(n18832), .Z(n8695) );
  XNOR U9227 ( .A(b[19]), .B(a[54]), .Z(n8842) );
  NANDN U9228 ( .A(n8842), .B(n18834), .Z(n8694) );
  NAND U9229 ( .A(n8695), .B(n8694), .Z(n8909) );
  XNOR U9230 ( .A(b[27]), .B(a[46]), .Z(n8845) );
  NANDN U9231 ( .A(n8845), .B(n19336), .Z(n8698) );
  NANDN U9232 ( .A(n8696), .B(n19337), .Z(n8697) );
  NAND U9233 ( .A(n8698), .B(n8697), .Z(n8906) );
  XOR U9234 ( .A(b[5]), .B(a[68]), .Z(n8848) );
  NAND U9235 ( .A(n8848), .B(n17310), .Z(n8701) );
  NAND U9236 ( .A(n8699), .B(n17311), .Z(n8700) );
  AND U9237 ( .A(n8701), .B(n8700), .Z(n8907) );
  XNOR U9238 ( .A(n8906), .B(n8907), .Z(n8908) );
  XNOR U9239 ( .A(n8909), .B(n8908), .Z(n8897) );
  XOR U9240 ( .A(b[17]), .B(a[56]), .Z(n8851) );
  NAND U9241 ( .A(n8851), .B(n18673), .Z(n8704) );
  NANDN U9242 ( .A(n8702), .B(n18674), .Z(n8703) );
  NAND U9243 ( .A(n8704), .B(n8703), .Z(n8869) );
  XOR U9244 ( .A(b[31]), .B(n9080), .Z(n8854) );
  NANDN U9245 ( .A(n8854), .B(n19472), .Z(n8707) );
  NANDN U9246 ( .A(n8705), .B(n19473), .Z(n8706) );
  NAND U9247 ( .A(n8707), .B(n8706), .Z(n8866) );
  OR U9248 ( .A(n8708), .B(n16988), .Z(n8710) );
  XNOR U9249 ( .A(b[3]), .B(a[70]), .Z(n8857) );
  NANDN U9250 ( .A(n8857), .B(n16990), .Z(n8709) );
  AND U9251 ( .A(n8710), .B(n8709), .Z(n8867) );
  XNOR U9252 ( .A(n8866), .B(n8867), .Z(n8868) );
  XOR U9253 ( .A(n8869), .B(n8868), .Z(n8896) );
  XNOR U9254 ( .A(n8897), .B(n8896), .Z(n8898) );
  XNOR U9255 ( .A(n8899), .B(n8898), .Z(n8943) );
  NANDN U9256 ( .A(n8712), .B(n8711), .Z(n8716) );
  NAND U9257 ( .A(n8714), .B(n8713), .Z(n8715) );
  NAND U9258 ( .A(n8716), .B(n8715), .Z(n8887) );
  NANDN U9259 ( .A(n8718), .B(n8717), .Z(n8722) );
  NAND U9260 ( .A(n8720), .B(n8719), .Z(n8721) );
  NAND U9261 ( .A(n8722), .B(n8721), .Z(n8885) );
  OR U9262 ( .A(n8724), .B(n8723), .Z(n8728) );
  NANDN U9263 ( .A(n8726), .B(n8725), .Z(n8727) );
  NAND U9264 ( .A(n8728), .B(n8727), .Z(n8884) );
  XNOR U9265 ( .A(n8887), .B(n8886), .Z(n8944) );
  XOR U9266 ( .A(n8943), .B(n8944), .Z(n8946) );
  NANDN U9267 ( .A(n8730), .B(n8729), .Z(n8734) );
  OR U9268 ( .A(n8732), .B(n8731), .Z(n8733) );
  NAND U9269 ( .A(n8734), .B(n8733), .Z(n8945) );
  XOR U9270 ( .A(n8946), .B(n8945), .Z(n8832) );
  OR U9271 ( .A(n8736), .B(n8735), .Z(n8740) );
  NAND U9272 ( .A(n8738), .B(n8737), .Z(n8739) );
  NAND U9273 ( .A(n8740), .B(n8739), .Z(n8831) );
  NANDN U9274 ( .A(n8742), .B(n8741), .Z(n8746) );
  NANDN U9275 ( .A(n8744), .B(n8743), .Z(n8745) );
  NAND U9276 ( .A(n8746), .B(n8745), .Z(n8951) );
  NANDN U9277 ( .A(n8748), .B(n8747), .Z(n8752) );
  OR U9278 ( .A(n8750), .B(n8749), .Z(n8751) );
  NAND U9279 ( .A(n8752), .B(n8751), .Z(n8950) );
  NANDN U9280 ( .A(n8754), .B(n8753), .Z(n8758) );
  NAND U9281 ( .A(n8756), .B(n8755), .Z(n8757) );
  NAND U9282 ( .A(n8758), .B(n8757), .Z(n8890) );
  NANDN U9283 ( .A(n8760), .B(n8759), .Z(n8764) );
  NAND U9284 ( .A(n8762), .B(n8761), .Z(n8763) );
  AND U9285 ( .A(n8764), .B(n8763), .Z(n8891) );
  XNOR U9286 ( .A(n8890), .B(n8891), .Z(n8892) );
  XNOR U9287 ( .A(b[9]), .B(a[64]), .Z(n8912) );
  NANDN U9288 ( .A(n8912), .B(n17814), .Z(n8767) );
  NANDN U9289 ( .A(n8765), .B(n17815), .Z(n8766) );
  NAND U9290 ( .A(n8767), .B(n8766), .Z(n8874) );
  NAND U9291 ( .A(n8768), .B(n18513), .Z(n8770) );
  XOR U9292 ( .A(b[15]), .B(a[58]), .Z(n8915) );
  NANDN U9293 ( .A(n18512), .B(n8915), .Z(n8769) );
  AND U9294 ( .A(n8770), .B(n8769), .Z(n8872) );
  NANDN U9295 ( .A(n8771), .B(n19013), .Z(n8773) );
  XNOR U9296 ( .A(b[21]), .B(a[52]), .Z(n8918) );
  NANDN U9297 ( .A(n8918), .B(n19015), .Z(n8772) );
  AND U9298 ( .A(n8773), .B(n8772), .Z(n8873) );
  XOR U9299 ( .A(n8874), .B(n8875), .Z(n8863) );
  XNOR U9300 ( .A(b[11]), .B(a[62]), .Z(n8921) );
  OR U9301 ( .A(n8921), .B(n18194), .Z(n8776) );
  NANDN U9302 ( .A(n8774), .B(n18104), .Z(n8775) );
  NAND U9303 ( .A(n8776), .B(n8775), .Z(n8861) );
  XOR U9304 ( .A(n580), .B(a[60]), .Z(n8924) );
  NANDN U9305 ( .A(n8924), .B(n18336), .Z(n8779) );
  NANDN U9306 ( .A(n8777), .B(n18337), .Z(n8778) );
  AND U9307 ( .A(n8779), .B(n8778), .Z(n8860) );
  XNOR U9308 ( .A(n8861), .B(n8860), .Z(n8862) );
  XOR U9309 ( .A(n8863), .B(n8862), .Z(n8880) );
  NANDN U9310 ( .A(n577), .B(a[72]), .Z(n8780) );
  XOR U9311 ( .A(n17151), .B(n8780), .Z(n8782) );
  NANDN U9312 ( .A(b[0]), .B(a[71]), .Z(n8781) );
  AND U9313 ( .A(n8782), .B(n8781), .Z(n8838) );
  NAND U9314 ( .A(n19406), .B(n8783), .Z(n8785) );
  XNOR U9315 ( .A(b[29]), .B(a[44]), .Z(n8931) );
  OR U9316 ( .A(n8931), .B(n576), .Z(n8784) );
  NAND U9317 ( .A(n8785), .B(n8784), .Z(n8836) );
  NANDN U9318 ( .A(n585), .B(a[40]), .Z(n8837) );
  XNOR U9319 ( .A(n8836), .B(n8837), .Z(n8839) );
  XOR U9320 ( .A(n8838), .B(n8839), .Z(n8878) );
  XOR U9321 ( .A(b[23]), .B(a[50]), .Z(n8934) );
  NANDN U9322 ( .A(n19127), .B(n8934), .Z(n8788) );
  NANDN U9323 ( .A(n8786), .B(n19128), .Z(n8787) );
  NAND U9324 ( .A(n8788), .B(n8787), .Z(n8903) );
  NANDN U9325 ( .A(n8789), .B(n17553), .Z(n8791) );
  XOR U9326 ( .A(b[7]), .B(a[66]), .Z(n8937) );
  NAND U9327 ( .A(n8937), .B(n17555), .Z(n8790) );
  NAND U9328 ( .A(n8791), .B(n8790), .Z(n8900) );
  XOR U9329 ( .A(b[25]), .B(a[48]), .Z(n8940) );
  NAND U9330 ( .A(n8940), .B(n19240), .Z(n8794) );
  NAND U9331 ( .A(n8792), .B(n19242), .Z(n8793) );
  AND U9332 ( .A(n8794), .B(n8793), .Z(n8901) );
  XNOR U9333 ( .A(n8900), .B(n8901), .Z(n8902) );
  XNOR U9334 ( .A(n8903), .B(n8902), .Z(n8879) );
  XOR U9335 ( .A(n8878), .B(n8879), .Z(n8881) );
  XNOR U9336 ( .A(n8880), .B(n8881), .Z(n8893) );
  XNOR U9337 ( .A(n8892), .B(n8893), .Z(n8949) );
  XNOR U9338 ( .A(n8950), .B(n8949), .Z(n8952) );
  XNOR U9339 ( .A(n8951), .B(n8952), .Z(n8830) );
  XOR U9340 ( .A(n8831), .B(n8830), .Z(n8833) );
  NANDN U9341 ( .A(n8796), .B(n8795), .Z(n8800) );
  NAND U9342 ( .A(n8798), .B(n8797), .Z(n8799) );
  NAND U9343 ( .A(n8800), .B(n8799), .Z(n8824) );
  NANDN U9344 ( .A(n8802), .B(n8801), .Z(n8806) );
  NAND U9345 ( .A(n8804), .B(n8803), .Z(n8805) );
  NAND U9346 ( .A(n8806), .B(n8805), .Z(n8825) );
  XNOR U9347 ( .A(n8824), .B(n8825), .Z(n8826) );
  XOR U9348 ( .A(n8827), .B(n8826), .Z(n8821) );
  XOR U9349 ( .A(n8820), .B(n8821), .Z(n8812) );
  XOR U9350 ( .A(n8813), .B(n8812), .Z(n8814) );
  XNOR U9351 ( .A(n8815), .B(n8814), .Z(n8955) );
  XNOR U9352 ( .A(n8955), .B(sreg[168]), .Z(n8957) );
  NAND U9353 ( .A(n8807), .B(sreg[167]), .Z(n8811) );
  OR U9354 ( .A(n8809), .B(n8808), .Z(n8810) );
  AND U9355 ( .A(n8811), .B(n8810), .Z(n8956) );
  XOR U9356 ( .A(n8957), .B(n8956), .Z(c[168]) );
  NAND U9357 ( .A(n8813), .B(n8812), .Z(n8817) );
  NAND U9358 ( .A(n8815), .B(n8814), .Z(n8816) );
  NAND U9359 ( .A(n8817), .B(n8816), .Z(n8963) );
  NANDN U9360 ( .A(n8819), .B(n8818), .Z(n8823) );
  NAND U9361 ( .A(n8821), .B(n8820), .Z(n8822) );
  NAND U9362 ( .A(n8823), .B(n8822), .Z(n8961) );
  NANDN U9363 ( .A(n8825), .B(n8824), .Z(n8829) );
  NAND U9364 ( .A(n8827), .B(n8826), .Z(n8828) );
  NAND U9365 ( .A(n8829), .B(n8828), .Z(n8966) );
  NANDN U9366 ( .A(n8831), .B(n8830), .Z(n8835) );
  OR U9367 ( .A(n8833), .B(n8832), .Z(n8834) );
  NAND U9368 ( .A(n8835), .B(n8834), .Z(n8967) );
  XNOR U9369 ( .A(n8966), .B(n8967), .Z(n8968) );
  NANDN U9370 ( .A(n8837), .B(n8836), .Z(n8841) );
  NAND U9371 ( .A(n8839), .B(n8838), .Z(n8840) );
  NAND U9372 ( .A(n8841), .B(n8840), .Z(n9047) );
  NANDN U9373 ( .A(n8842), .B(n18832), .Z(n8844) );
  XOR U9374 ( .A(b[19]), .B(n10959), .Z(n9014) );
  NANDN U9375 ( .A(n9014), .B(n18834), .Z(n8843) );
  NAND U9376 ( .A(n8844), .B(n8843), .Z(n9059) );
  XNOR U9377 ( .A(b[27]), .B(a[47]), .Z(n9017) );
  NANDN U9378 ( .A(n9017), .B(n19336), .Z(n8847) );
  NANDN U9379 ( .A(n8845), .B(n19337), .Z(n8846) );
  NAND U9380 ( .A(n8847), .B(n8846), .Z(n9056) );
  XOR U9381 ( .A(b[5]), .B(a[69]), .Z(n9020) );
  NAND U9382 ( .A(n9020), .B(n17310), .Z(n8850) );
  NAND U9383 ( .A(n8848), .B(n17311), .Z(n8849) );
  AND U9384 ( .A(n8850), .B(n8849), .Z(n9057) );
  XNOR U9385 ( .A(n9056), .B(n9057), .Z(n9058) );
  XNOR U9386 ( .A(n9059), .B(n9058), .Z(n9044) );
  XOR U9387 ( .A(b[17]), .B(a[57]), .Z(n9023) );
  NAND U9388 ( .A(n9023), .B(n18673), .Z(n8853) );
  NAND U9389 ( .A(n8851), .B(n18674), .Z(n8852) );
  NAND U9390 ( .A(n8853), .B(n8852), .Z(n8998) );
  XNOR U9391 ( .A(b[31]), .B(a[43]), .Z(n9026) );
  NANDN U9392 ( .A(n9026), .B(n19472), .Z(n8856) );
  NANDN U9393 ( .A(n8854), .B(n19473), .Z(n8855) );
  AND U9394 ( .A(n8856), .B(n8855), .Z(n8996) );
  OR U9395 ( .A(n8857), .B(n16988), .Z(n8859) );
  XNOR U9396 ( .A(b[3]), .B(a[71]), .Z(n9029) );
  NANDN U9397 ( .A(n9029), .B(n16990), .Z(n8858) );
  AND U9398 ( .A(n8859), .B(n8858), .Z(n8997) );
  XOR U9399 ( .A(n8998), .B(n8999), .Z(n9045) );
  XOR U9400 ( .A(n9044), .B(n9045), .Z(n9046) );
  XNOR U9401 ( .A(n9047), .B(n9046), .Z(n9093) );
  NANDN U9402 ( .A(n8861), .B(n8860), .Z(n8865) );
  NAND U9403 ( .A(n8863), .B(n8862), .Z(n8864) );
  NAND U9404 ( .A(n8865), .B(n8864), .Z(n9035) );
  NANDN U9405 ( .A(n8867), .B(n8866), .Z(n8871) );
  NAND U9406 ( .A(n8869), .B(n8868), .Z(n8870) );
  NAND U9407 ( .A(n8871), .B(n8870), .Z(n9033) );
  OR U9408 ( .A(n8873), .B(n8872), .Z(n8877) );
  NANDN U9409 ( .A(n8875), .B(n8874), .Z(n8876) );
  NAND U9410 ( .A(n8877), .B(n8876), .Z(n9032) );
  XNOR U9411 ( .A(n9035), .B(n9034), .Z(n9094) );
  XOR U9412 ( .A(n9093), .B(n9094), .Z(n9096) );
  NANDN U9413 ( .A(n8879), .B(n8878), .Z(n8883) );
  OR U9414 ( .A(n8881), .B(n8880), .Z(n8882) );
  NAND U9415 ( .A(n8883), .B(n8882), .Z(n9095) );
  XOR U9416 ( .A(n9096), .B(n9095), .Z(n8980) );
  OR U9417 ( .A(n8885), .B(n8884), .Z(n8889) );
  NAND U9418 ( .A(n8887), .B(n8886), .Z(n8888) );
  NAND U9419 ( .A(n8889), .B(n8888), .Z(n8979) );
  NANDN U9420 ( .A(n8891), .B(n8890), .Z(n8895) );
  NANDN U9421 ( .A(n8893), .B(n8892), .Z(n8894) );
  NAND U9422 ( .A(n8895), .B(n8894), .Z(n9101) );
  NANDN U9423 ( .A(n8901), .B(n8900), .Z(n8905) );
  NAND U9424 ( .A(n8903), .B(n8902), .Z(n8904) );
  NAND U9425 ( .A(n8905), .B(n8904), .Z(n9038) );
  NANDN U9426 ( .A(n8907), .B(n8906), .Z(n8911) );
  NAND U9427 ( .A(n8909), .B(n8908), .Z(n8910) );
  AND U9428 ( .A(n8911), .B(n8910), .Z(n9039) );
  XNOR U9429 ( .A(n9038), .B(n9039), .Z(n9040) );
  XOR U9430 ( .A(n579), .B(n12055), .Z(n9068) );
  NAND U9431 ( .A(n17814), .B(n9068), .Z(n8914) );
  NANDN U9432 ( .A(n8912), .B(n17815), .Z(n8913) );
  NAND U9433 ( .A(n8914), .B(n8913), .Z(n9004) );
  NAND U9434 ( .A(n8915), .B(n18513), .Z(n8917) );
  XOR U9435 ( .A(b[15]), .B(a[59]), .Z(n9065) );
  NANDN U9436 ( .A(n18512), .B(n9065), .Z(n8916) );
  AND U9437 ( .A(n8917), .B(n8916), .Z(n9002) );
  NANDN U9438 ( .A(n8918), .B(n19013), .Z(n8920) );
  XOR U9439 ( .A(n582), .B(n10660), .Z(n9062) );
  NAND U9440 ( .A(n9062), .B(n19015), .Z(n8919) );
  AND U9441 ( .A(n8920), .B(n8919), .Z(n9003) );
  XOR U9442 ( .A(n9004), .B(n9005), .Z(n8993) );
  XNOR U9443 ( .A(b[11]), .B(a[63]), .Z(n9071) );
  OR U9444 ( .A(n9071), .B(n18194), .Z(n8923) );
  NANDN U9445 ( .A(n8921), .B(n18104), .Z(n8922) );
  NAND U9446 ( .A(n8923), .B(n8922), .Z(n8991) );
  XOR U9447 ( .A(n580), .B(a[61]), .Z(n9074) );
  NANDN U9448 ( .A(n9074), .B(n18336), .Z(n8926) );
  NANDN U9449 ( .A(n8924), .B(n18337), .Z(n8925) );
  NAND U9450 ( .A(n8926), .B(n8925), .Z(n8990) );
  XOR U9451 ( .A(n8993), .B(n8992), .Z(n8987) );
  NANDN U9452 ( .A(n577), .B(a[73]), .Z(n8927) );
  XOR U9453 ( .A(n17151), .B(n8927), .Z(n8929) );
  NANDN U9454 ( .A(b[0]), .B(a[72]), .Z(n8928) );
  AND U9455 ( .A(n8929), .B(n8928), .Z(n9011) );
  ANDN U9456 ( .B(b[31]), .A(n8930), .Z(n9008) );
  NANDN U9457 ( .A(n8931), .B(n19406), .Z(n8933) );
  XNOR U9458 ( .A(b[29]), .B(a[45]), .Z(n9081) );
  OR U9459 ( .A(n9081), .B(n576), .Z(n8932) );
  NAND U9460 ( .A(n8933), .B(n8932), .Z(n9009) );
  XOR U9461 ( .A(n9008), .B(n9009), .Z(n9010) );
  XNOR U9462 ( .A(n9011), .B(n9010), .Z(n8984) );
  XOR U9463 ( .A(b[23]), .B(a[51]), .Z(n9084) );
  NANDN U9464 ( .A(n19127), .B(n9084), .Z(n8936) );
  NAND U9465 ( .A(n8934), .B(n19128), .Z(n8935) );
  NAND U9466 ( .A(n8936), .B(n8935), .Z(n9053) );
  NAND U9467 ( .A(n8937), .B(n17553), .Z(n8939) );
  XOR U9468 ( .A(b[7]), .B(a[67]), .Z(n9087) );
  NAND U9469 ( .A(n9087), .B(n17555), .Z(n8938) );
  NAND U9470 ( .A(n8939), .B(n8938), .Z(n9050) );
  XNOR U9471 ( .A(b[25]), .B(a[49]), .Z(n9090) );
  NANDN U9472 ( .A(n9090), .B(n19240), .Z(n8942) );
  NAND U9473 ( .A(n8940), .B(n19242), .Z(n8941) );
  AND U9474 ( .A(n8942), .B(n8941), .Z(n9051) );
  XNOR U9475 ( .A(n9050), .B(n9051), .Z(n9052) );
  XNOR U9476 ( .A(n9053), .B(n9052), .Z(n8985) );
  XOR U9477 ( .A(n8987), .B(n8986), .Z(n9041) );
  XNOR U9478 ( .A(n9040), .B(n9041), .Z(n9099) );
  XNOR U9479 ( .A(n9100), .B(n9099), .Z(n9102) );
  XNOR U9480 ( .A(n9101), .B(n9102), .Z(n8978) );
  XOR U9481 ( .A(n8979), .B(n8978), .Z(n8981) );
  NANDN U9482 ( .A(n8944), .B(n8943), .Z(n8948) );
  OR U9483 ( .A(n8946), .B(n8945), .Z(n8947) );
  NAND U9484 ( .A(n8948), .B(n8947), .Z(n8972) );
  NAND U9485 ( .A(n8950), .B(n8949), .Z(n8954) );
  NANDN U9486 ( .A(n8952), .B(n8951), .Z(n8953) );
  NAND U9487 ( .A(n8954), .B(n8953), .Z(n8973) );
  XNOR U9488 ( .A(n8972), .B(n8973), .Z(n8974) );
  XOR U9489 ( .A(n8975), .B(n8974), .Z(n8969) );
  XOR U9490 ( .A(n8968), .B(n8969), .Z(n8960) );
  XOR U9491 ( .A(n8961), .B(n8960), .Z(n8962) );
  XNOR U9492 ( .A(n8963), .B(n8962), .Z(n9105) );
  XNOR U9493 ( .A(n9105), .B(sreg[169]), .Z(n9107) );
  NAND U9494 ( .A(n8955), .B(sreg[168]), .Z(n8959) );
  OR U9495 ( .A(n8957), .B(n8956), .Z(n8958) );
  AND U9496 ( .A(n8959), .B(n8958), .Z(n9106) );
  XOR U9497 ( .A(n9107), .B(n9106), .Z(c[169]) );
  NAND U9498 ( .A(n8961), .B(n8960), .Z(n8965) );
  NAND U9499 ( .A(n8963), .B(n8962), .Z(n8964) );
  NAND U9500 ( .A(n8965), .B(n8964), .Z(n9113) );
  NANDN U9501 ( .A(n8967), .B(n8966), .Z(n8971) );
  NAND U9502 ( .A(n8969), .B(n8968), .Z(n8970) );
  NAND U9503 ( .A(n8971), .B(n8970), .Z(n9111) );
  NANDN U9504 ( .A(n8973), .B(n8972), .Z(n8977) );
  NAND U9505 ( .A(n8975), .B(n8974), .Z(n8976) );
  NAND U9506 ( .A(n8977), .B(n8976), .Z(n9116) );
  NANDN U9507 ( .A(n8979), .B(n8978), .Z(n8983) );
  OR U9508 ( .A(n8981), .B(n8980), .Z(n8982) );
  NAND U9509 ( .A(n8983), .B(n8982), .Z(n9117) );
  XNOR U9510 ( .A(n9116), .B(n9117), .Z(n9118) );
  OR U9511 ( .A(n8985), .B(n8984), .Z(n8989) );
  NANDN U9512 ( .A(n8987), .B(n8986), .Z(n8988) );
  NAND U9513 ( .A(n8989), .B(n8988), .Z(n9231) );
  OR U9514 ( .A(n8991), .B(n8990), .Z(n8995) );
  NAND U9515 ( .A(n8993), .B(n8992), .Z(n8994) );
  NAND U9516 ( .A(n8995), .B(n8994), .Z(n9170) );
  OR U9517 ( .A(n8997), .B(n8996), .Z(n9001) );
  NANDN U9518 ( .A(n8999), .B(n8998), .Z(n9000) );
  NAND U9519 ( .A(n9001), .B(n9000), .Z(n9169) );
  OR U9520 ( .A(n9003), .B(n9002), .Z(n9007) );
  NANDN U9521 ( .A(n9005), .B(n9004), .Z(n9006) );
  NAND U9522 ( .A(n9007), .B(n9006), .Z(n9168) );
  XOR U9523 ( .A(n9170), .B(n9171), .Z(n9229) );
  OR U9524 ( .A(n9009), .B(n9008), .Z(n9013) );
  NANDN U9525 ( .A(n9011), .B(n9010), .Z(n9012) );
  NAND U9526 ( .A(n9013), .B(n9012), .Z(n9182) );
  NANDN U9527 ( .A(n9014), .B(n18832), .Z(n9016) );
  XNOR U9528 ( .A(b[19]), .B(a[56]), .Z(n9128) );
  NANDN U9529 ( .A(n9128), .B(n18834), .Z(n9015) );
  NAND U9530 ( .A(n9016), .B(n9015), .Z(n9195) );
  XNOR U9531 ( .A(b[27]), .B(a[48]), .Z(n9131) );
  NANDN U9532 ( .A(n9131), .B(n19336), .Z(n9019) );
  NANDN U9533 ( .A(n9017), .B(n19337), .Z(n9018) );
  NAND U9534 ( .A(n9019), .B(n9018), .Z(n9192) );
  XOR U9535 ( .A(b[5]), .B(a[70]), .Z(n9134) );
  NAND U9536 ( .A(n9134), .B(n17310), .Z(n9022) );
  NAND U9537 ( .A(n9020), .B(n17311), .Z(n9021) );
  AND U9538 ( .A(n9022), .B(n9021), .Z(n9193) );
  XNOR U9539 ( .A(n9192), .B(n9193), .Z(n9194) );
  XNOR U9540 ( .A(n9195), .B(n9194), .Z(n9181) );
  XOR U9541 ( .A(b[17]), .B(a[58]), .Z(n9137) );
  NAND U9542 ( .A(n9137), .B(n18673), .Z(n9025) );
  NAND U9543 ( .A(n9023), .B(n18674), .Z(n9024) );
  NAND U9544 ( .A(n9025), .B(n9024), .Z(n9155) );
  XNOR U9545 ( .A(b[31]), .B(a[44]), .Z(n9140) );
  NANDN U9546 ( .A(n9140), .B(n19472), .Z(n9028) );
  NANDN U9547 ( .A(n9026), .B(n19473), .Z(n9027) );
  NAND U9548 ( .A(n9028), .B(n9027), .Z(n9152) );
  OR U9549 ( .A(n9029), .B(n16988), .Z(n9031) );
  XNOR U9550 ( .A(b[3]), .B(a[72]), .Z(n9143) );
  NANDN U9551 ( .A(n9143), .B(n16990), .Z(n9030) );
  AND U9552 ( .A(n9031), .B(n9030), .Z(n9153) );
  XNOR U9553 ( .A(n9152), .B(n9153), .Z(n9154) );
  XOR U9554 ( .A(n9155), .B(n9154), .Z(n9180) );
  XOR U9555 ( .A(n9181), .B(n9180), .Z(n9183) );
  XOR U9556 ( .A(n9182), .B(n9183), .Z(n9228) );
  XOR U9557 ( .A(n9229), .B(n9228), .Z(n9230) );
  XNOR U9558 ( .A(n9231), .B(n9230), .Z(n9249) );
  OR U9559 ( .A(n9033), .B(n9032), .Z(n9037) );
  NAND U9560 ( .A(n9035), .B(n9034), .Z(n9036) );
  NAND U9561 ( .A(n9037), .B(n9036), .Z(n9247) );
  NANDN U9562 ( .A(n9039), .B(n9038), .Z(n9043) );
  NANDN U9563 ( .A(n9041), .B(n9040), .Z(n9042) );
  NAND U9564 ( .A(n9043), .B(n9042), .Z(n9236) );
  OR U9565 ( .A(n9045), .B(n9044), .Z(n9049) );
  NAND U9566 ( .A(n9047), .B(n9046), .Z(n9048) );
  NAND U9567 ( .A(n9049), .B(n9048), .Z(n9235) );
  NANDN U9568 ( .A(n9051), .B(n9050), .Z(n9055) );
  NAND U9569 ( .A(n9053), .B(n9052), .Z(n9054) );
  NAND U9570 ( .A(n9055), .B(n9054), .Z(n9174) );
  NANDN U9571 ( .A(n9057), .B(n9056), .Z(n9061) );
  NAND U9572 ( .A(n9059), .B(n9058), .Z(n9060) );
  AND U9573 ( .A(n9061), .B(n9060), .Z(n9175) );
  XNOR U9574 ( .A(n9174), .B(n9175), .Z(n9176) );
  XNOR U9575 ( .A(b[21]), .B(a[54]), .Z(n9204) );
  NANDN U9576 ( .A(n9204), .B(n19015), .Z(n9064) );
  NAND U9577 ( .A(n19013), .B(n9062), .Z(n9063) );
  NAND U9578 ( .A(n9064), .B(n9063), .Z(n9164) );
  NAND U9579 ( .A(n9065), .B(n18513), .Z(n9067) );
  XOR U9580 ( .A(b[15]), .B(a[60]), .Z(n9201) );
  NANDN U9581 ( .A(n18512), .B(n9201), .Z(n9066) );
  AND U9582 ( .A(n9067), .B(n9066), .Z(n9165) );
  XNOR U9583 ( .A(n9164), .B(n9165), .Z(n9167) );
  XNOR U9584 ( .A(b[9]), .B(a[66]), .Z(n9198) );
  NANDN U9585 ( .A(n9198), .B(n17814), .Z(n9070) );
  NAND U9586 ( .A(n17815), .B(n9068), .Z(n9069) );
  NAND U9587 ( .A(n9070), .B(n9069), .Z(n9166) );
  XNOR U9588 ( .A(n9167), .B(n9166), .Z(n9160) );
  XNOR U9589 ( .A(b[11]), .B(a[64]), .Z(n9207) );
  OR U9590 ( .A(n9207), .B(n18194), .Z(n9073) );
  NANDN U9591 ( .A(n9071), .B(n18104), .Z(n9072) );
  NAND U9592 ( .A(n9073), .B(n9072), .Z(n9159) );
  XOR U9593 ( .A(n580), .B(a[62]), .Z(n9210) );
  NANDN U9594 ( .A(n9210), .B(n18336), .Z(n9076) );
  NANDN U9595 ( .A(n9074), .B(n18337), .Z(n9075) );
  NAND U9596 ( .A(n9076), .B(n9075), .Z(n9158) );
  XNOR U9597 ( .A(n9159), .B(n9158), .Z(n9161) );
  XNOR U9598 ( .A(n9160), .B(n9161), .Z(n9149) );
  NANDN U9599 ( .A(n577), .B(a[74]), .Z(n9077) );
  XOR U9600 ( .A(n17151), .B(n9077), .Z(n9079) );
  NANDN U9601 ( .A(b[0]), .B(a[73]), .Z(n9078) );
  AND U9602 ( .A(n9079), .B(n9078), .Z(n9125) );
  ANDN U9603 ( .B(b[31]), .A(n9080), .Z(n9122) );
  NANDN U9604 ( .A(n9081), .B(n19406), .Z(n9083) );
  XNOR U9605 ( .A(n584), .B(a[46]), .Z(n9213) );
  NANDN U9606 ( .A(n576), .B(n9213), .Z(n9082) );
  NAND U9607 ( .A(n9083), .B(n9082), .Z(n9123) );
  XOR U9608 ( .A(n9122), .B(n9123), .Z(n9124) );
  XNOR U9609 ( .A(n9125), .B(n9124), .Z(n9146) );
  XOR U9610 ( .A(b[23]), .B(a[52]), .Z(n9219) );
  NANDN U9611 ( .A(n19127), .B(n9219), .Z(n9086) );
  NAND U9612 ( .A(n9084), .B(n19128), .Z(n9085) );
  NAND U9613 ( .A(n9086), .B(n9085), .Z(n9189) );
  NAND U9614 ( .A(n9087), .B(n17553), .Z(n9089) );
  XOR U9615 ( .A(b[7]), .B(a[68]), .Z(n9222) );
  NAND U9616 ( .A(n9222), .B(n17555), .Z(n9088) );
  NAND U9617 ( .A(n9089), .B(n9088), .Z(n9186) );
  XOR U9618 ( .A(b[25]), .B(a[50]), .Z(n9225) );
  NAND U9619 ( .A(n9225), .B(n19240), .Z(n9092) );
  NANDN U9620 ( .A(n9090), .B(n19242), .Z(n9091) );
  AND U9621 ( .A(n9092), .B(n9091), .Z(n9187) );
  XNOR U9622 ( .A(n9186), .B(n9187), .Z(n9188) );
  XNOR U9623 ( .A(n9189), .B(n9188), .Z(n9147) );
  XOR U9624 ( .A(n9149), .B(n9148), .Z(n9177) );
  XNOR U9625 ( .A(n9176), .B(n9177), .Z(n9234) );
  XNOR U9626 ( .A(n9235), .B(n9234), .Z(n9237) );
  XNOR U9627 ( .A(n9236), .B(n9237), .Z(n9246) );
  XNOR U9628 ( .A(n9247), .B(n9246), .Z(n9248) );
  XOR U9629 ( .A(n9249), .B(n9248), .Z(n9243) );
  NANDN U9630 ( .A(n9094), .B(n9093), .Z(n9098) );
  OR U9631 ( .A(n9096), .B(n9095), .Z(n9097) );
  NAND U9632 ( .A(n9098), .B(n9097), .Z(n9240) );
  NAND U9633 ( .A(n9100), .B(n9099), .Z(n9104) );
  NANDN U9634 ( .A(n9102), .B(n9101), .Z(n9103) );
  NAND U9635 ( .A(n9104), .B(n9103), .Z(n9241) );
  XNOR U9636 ( .A(n9240), .B(n9241), .Z(n9242) );
  XOR U9637 ( .A(n9243), .B(n9242), .Z(n9119) );
  XOR U9638 ( .A(n9118), .B(n9119), .Z(n9110) );
  XOR U9639 ( .A(n9111), .B(n9110), .Z(n9112) );
  XNOR U9640 ( .A(n9113), .B(n9112), .Z(n9252) );
  XNOR U9641 ( .A(n9252), .B(sreg[170]), .Z(n9254) );
  NAND U9642 ( .A(n9105), .B(sreg[169]), .Z(n9109) );
  OR U9643 ( .A(n9107), .B(n9106), .Z(n9108) );
  AND U9644 ( .A(n9109), .B(n9108), .Z(n9253) );
  XOR U9645 ( .A(n9254), .B(n9253), .Z(c[170]) );
  NAND U9646 ( .A(n9111), .B(n9110), .Z(n9115) );
  NAND U9647 ( .A(n9113), .B(n9112), .Z(n9114) );
  NAND U9648 ( .A(n9115), .B(n9114), .Z(n9260) );
  NANDN U9649 ( .A(n9117), .B(n9116), .Z(n9121) );
  NAND U9650 ( .A(n9119), .B(n9118), .Z(n9120) );
  NAND U9651 ( .A(n9121), .B(n9120), .Z(n9258) );
  OR U9652 ( .A(n9123), .B(n9122), .Z(n9127) );
  NANDN U9653 ( .A(n9125), .B(n9124), .Z(n9126) );
  NAND U9654 ( .A(n9127), .B(n9126), .Z(n9329) );
  NANDN U9655 ( .A(n9128), .B(n18832), .Z(n9130) );
  XNOR U9656 ( .A(b[19]), .B(a[57]), .Z(n9275) );
  NANDN U9657 ( .A(n9275), .B(n18834), .Z(n9129) );
  NAND U9658 ( .A(n9130), .B(n9129), .Z(n9342) );
  XOR U9659 ( .A(b[27]), .B(n10083), .Z(n9278) );
  NANDN U9660 ( .A(n9278), .B(n19336), .Z(n9133) );
  NANDN U9661 ( .A(n9131), .B(n19337), .Z(n9132) );
  NAND U9662 ( .A(n9133), .B(n9132), .Z(n9339) );
  XOR U9663 ( .A(b[5]), .B(a[71]), .Z(n9281) );
  NAND U9664 ( .A(n9281), .B(n17310), .Z(n9136) );
  NAND U9665 ( .A(n9134), .B(n17311), .Z(n9135) );
  AND U9666 ( .A(n9136), .B(n9135), .Z(n9340) );
  XNOR U9667 ( .A(n9339), .B(n9340), .Z(n9341) );
  XNOR U9668 ( .A(n9342), .B(n9341), .Z(n9328) );
  XOR U9669 ( .A(b[17]), .B(a[59]), .Z(n9284) );
  NAND U9670 ( .A(n9284), .B(n18673), .Z(n9139) );
  NAND U9671 ( .A(n9137), .B(n18674), .Z(n9138) );
  NAND U9672 ( .A(n9139), .B(n9138), .Z(n9302) );
  XNOR U9673 ( .A(b[31]), .B(a[45]), .Z(n9287) );
  NANDN U9674 ( .A(n9287), .B(n19472), .Z(n9142) );
  NANDN U9675 ( .A(n9140), .B(n19473), .Z(n9141) );
  NAND U9676 ( .A(n9142), .B(n9141), .Z(n9299) );
  OR U9677 ( .A(n9143), .B(n16988), .Z(n9145) );
  XNOR U9678 ( .A(b[3]), .B(a[73]), .Z(n9290) );
  NANDN U9679 ( .A(n9290), .B(n16990), .Z(n9144) );
  AND U9680 ( .A(n9145), .B(n9144), .Z(n9300) );
  XNOR U9681 ( .A(n9299), .B(n9300), .Z(n9301) );
  XOR U9682 ( .A(n9302), .B(n9301), .Z(n9327) );
  XOR U9683 ( .A(n9328), .B(n9327), .Z(n9330) );
  XNOR U9684 ( .A(n9329), .B(n9330), .Z(n9381) );
  OR U9685 ( .A(n9147), .B(n9146), .Z(n9151) );
  NANDN U9686 ( .A(n9149), .B(n9148), .Z(n9150) );
  NAND U9687 ( .A(n9151), .B(n9150), .Z(n9382) );
  XNOR U9688 ( .A(n9381), .B(n9382), .Z(n9383) );
  NANDN U9689 ( .A(n9153), .B(n9152), .Z(n9157) );
  NAND U9690 ( .A(n9155), .B(n9154), .Z(n9156) );
  NAND U9691 ( .A(n9157), .B(n9156), .Z(n9320) );
  OR U9692 ( .A(n9159), .B(n9158), .Z(n9163) );
  NANDN U9693 ( .A(n9161), .B(n9160), .Z(n9162) );
  NAND U9694 ( .A(n9163), .B(n9162), .Z(n9318) );
  XNOR U9695 ( .A(n9318), .B(n9317), .Z(n9319) );
  XOR U9696 ( .A(n9320), .B(n9319), .Z(n9384) );
  XOR U9697 ( .A(n9383), .B(n9384), .Z(n9396) );
  OR U9698 ( .A(n9169), .B(n9168), .Z(n9173) );
  NANDN U9699 ( .A(n9171), .B(n9170), .Z(n9172) );
  NAND U9700 ( .A(n9173), .B(n9172), .Z(n9394) );
  NANDN U9701 ( .A(n9175), .B(n9174), .Z(n9179) );
  NANDN U9702 ( .A(n9177), .B(n9176), .Z(n9178) );
  NAND U9703 ( .A(n9179), .B(n9178), .Z(n9377) );
  NANDN U9704 ( .A(n9181), .B(n9180), .Z(n9185) );
  OR U9705 ( .A(n9183), .B(n9182), .Z(n9184) );
  NAND U9706 ( .A(n9185), .B(n9184), .Z(n9376) );
  NANDN U9707 ( .A(n9187), .B(n9186), .Z(n9191) );
  NAND U9708 ( .A(n9189), .B(n9188), .Z(n9190) );
  NAND U9709 ( .A(n9191), .B(n9190), .Z(n9321) );
  NANDN U9710 ( .A(n9193), .B(n9192), .Z(n9197) );
  NAND U9711 ( .A(n9195), .B(n9194), .Z(n9196) );
  AND U9712 ( .A(n9197), .B(n9196), .Z(n9322) );
  XNOR U9713 ( .A(n9321), .B(n9322), .Z(n9323) );
  XNOR U9714 ( .A(b[9]), .B(a[67]), .Z(n9345) );
  NANDN U9715 ( .A(n9345), .B(n17814), .Z(n9200) );
  NANDN U9716 ( .A(n9198), .B(n17815), .Z(n9199) );
  NAND U9717 ( .A(n9200), .B(n9199), .Z(n9307) );
  NAND U9718 ( .A(n9201), .B(n18513), .Z(n9203) );
  XOR U9719 ( .A(b[15]), .B(a[61]), .Z(n9348) );
  NANDN U9720 ( .A(n18512), .B(n9348), .Z(n9202) );
  AND U9721 ( .A(n9203), .B(n9202), .Z(n9305) );
  NANDN U9722 ( .A(n9204), .B(n19013), .Z(n9206) );
  XOR U9723 ( .A(b[21]), .B(n10959), .Z(n9351) );
  NANDN U9724 ( .A(n9351), .B(n19015), .Z(n9205) );
  AND U9725 ( .A(n9206), .B(n9205), .Z(n9306) );
  XOR U9726 ( .A(n9307), .B(n9308), .Z(n9296) );
  XOR U9727 ( .A(b[11]), .B(n12055), .Z(n9354) );
  OR U9728 ( .A(n9354), .B(n18194), .Z(n9209) );
  NANDN U9729 ( .A(n9207), .B(n18104), .Z(n9208) );
  NAND U9730 ( .A(n9209), .B(n9208), .Z(n9294) );
  XOR U9731 ( .A(n580), .B(a[63]), .Z(n9357) );
  NANDN U9732 ( .A(n9357), .B(n18336), .Z(n9212) );
  NANDN U9733 ( .A(n9210), .B(n18337), .Z(n9211) );
  AND U9734 ( .A(n9212), .B(n9211), .Z(n9293) );
  XNOR U9735 ( .A(n9294), .B(n9293), .Z(n9295) );
  XOR U9736 ( .A(n9296), .B(n9295), .Z(n9313) );
  NAND U9737 ( .A(n9213), .B(n19406), .Z(n9215) );
  XNOR U9738 ( .A(n584), .B(a[47]), .Z(n9363) );
  NANDN U9739 ( .A(n576), .B(n9363), .Z(n9214) );
  NAND U9740 ( .A(n9215), .B(n9214), .Z(n9269) );
  NANDN U9741 ( .A(n585), .B(a[43]), .Z(n9270) );
  XNOR U9742 ( .A(n9269), .B(n9270), .Z(n9272) );
  NANDN U9743 ( .A(n577), .B(a[75]), .Z(n9216) );
  XOR U9744 ( .A(n17151), .B(n9216), .Z(n9218) );
  NANDN U9745 ( .A(b[0]), .B(a[74]), .Z(n9217) );
  AND U9746 ( .A(n9218), .B(n9217), .Z(n9271) );
  XOR U9747 ( .A(n9272), .B(n9271), .Z(n9311) );
  XNOR U9748 ( .A(b[23]), .B(a[53]), .Z(n9366) );
  OR U9749 ( .A(n9366), .B(n19127), .Z(n9221) );
  NAND U9750 ( .A(n9219), .B(n19128), .Z(n9220) );
  NAND U9751 ( .A(n9221), .B(n9220), .Z(n9336) );
  NAND U9752 ( .A(n9222), .B(n17553), .Z(n9224) );
  XOR U9753 ( .A(b[7]), .B(a[69]), .Z(n9369) );
  NAND U9754 ( .A(n9369), .B(n17555), .Z(n9223) );
  NAND U9755 ( .A(n9224), .B(n9223), .Z(n9333) );
  XOR U9756 ( .A(b[25]), .B(a[51]), .Z(n9372) );
  NAND U9757 ( .A(n9372), .B(n19240), .Z(n9227) );
  NAND U9758 ( .A(n9225), .B(n19242), .Z(n9226) );
  AND U9759 ( .A(n9227), .B(n9226), .Z(n9334) );
  XNOR U9760 ( .A(n9333), .B(n9334), .Z(n9335) );
  XNOR U9761 ( .A(n9336), .B(n9335), .Z(n9312) );
  XOR U9762 ( .A(n9311), .B(n9312), .Z(n9314) );
  XNOR U9763 ( .A(n9313), .B(n9314), .Z(n9324) );
  XNOR U9764 ( .A(n9323), .B(n9324), .Z(n9375) );
  XNOR U9765 ( .A(n9376), .B(n9375), .Z(n9378) );
  XNOR U9766 ( .A(n9377), .B(n9378), .Z(n9393) );
  XOR U9767 ( .A(n9394), .B(n9393), .Z(n9395) );
  XNOR U9768 ( .A(n9396), .B(n9395), .Z(n9390) );
  NAND U9769 ( .A(n9229), .B(n9228), .Z(n9233) );
  NAND U9770 ( .A(n9231), .B(n9230), .Z(n9232) );
  NAND U9771 ( .A(n9233), .B(n9232), .Z(n9388) );
  NAND U9772 ( .A(n9235), .B(n9234), .Z(n9239) );
  NANDN U9773 ( .A(n9237), .B(n9236), .Z(n9238) );
  AND U9774 ( .A(n9239), .B(n9238), .Z(n9387) );
  XNOR U9775 ( .A(n9388), .B(n9387), .Z(n9389) );
  XOR U9776 ( .A(n9390), .B(n9389), .Z(n9265) );
  NANDN U9777 ( .A(n9241), .B(n9240), .Z(n9245) );
  NAND U9778 ( .A(n9243), .B(n9242), .Z(n9244) );
  NAND U9779 ( .A(n9245), .B(n9244), .Z(n9263) );
  NANDN U9780 ( .A(n9247), .B(n9246), .Z(n9251) );
  NANDN U9781 ( .A(n9249), .B(n9248), .Z(n9250) );
  NAND U9782 ( .A(n9251), .B(n9250), .Z(n9264) );
  XNOR U9783 ( .A(n9263), .B(n9264), .Z(n9266) );
  XOR U9784 ( .A(n9265), .B(n9266), .Z(n9257) );
  XOR U9785 ( .A(n9258), .B(n9257), .Z(n9259) );
  XNOR U9786 ( .A(n9260), .B(n9259), .Z(n9399) );
  XNOR U9787 ( .A(n9399), .B(sreg[171]), .Z(n9401) );
  NAND U9788 ( .A(n9252), .B(sreg[170]), .Z(n9256) );
  OR U9789 ( .A(n9254), .B(n9253), .Z(n9255) );
  AND U9790 ( .A(n9256), .B(n9255), .Z(n9400) );
  XOR U9791 ( .A(n9401), .B(n9400), .Z(c[171]) );
  NAND U9792 ( .A(n9258), .B(n9257), .Z(n9262) );
  NAND U9793 ( .A(n9260), .B(n9259), .Z(n9261) );
  NAND U9794 ( .A(n9262), .B(n9261), .Z(n9407) );
  NANDN U9795 ( .A(n9264), .B(n9263), .Z(n9268) );
  NAND U9796 ( .A(n9266), .B(n9265), .Z(n9267) );
  NAND U9797 ( .A(n9268), .B(n9267), .Z(n9405) );
  NANDN U9798 ( .A(n9270), .B(n9269), .Z(n9274) );
  NAND U9799 ( .A(n9272), .B(n9271), .Z(n9273) );
  NAND U9800 ( .A(n9274), .B(n9273), .Z(n9487) );
  NANDN U9801 ( .A(n9275), .B(n18832), .Z(n9277) );
  XNOR U9802 ( .A(b[19]), .B(a[58]), .Z(n9430) );
  NANDN U9803 ( .A(n9430), .B(n18834), .Z(n9276) );
  NAND U9804 ( .A(n9277), .B(n9276), .Z(n9497) );
  XNOR U9805 ( .A(b[27]), .B(a[50]), .Z(n9433) );
  NANDN U9806 ( .A(n9433), .B(n19336), .Z(n9280) );
  NANDN U9807 ( .A(n9278), .B(n19337), .Z(n9279) );
  NAND U9808 ( .A(n9280), .B(n9279), .Z(n9494) );
  XOR U9809 ( .A(b[5]), .B(a[72]), .Z(n9436) );
  NAND U9810 ( .A(n9436), .B(n17310), .Z(n9283) );
  NAND U9811 ( .A(n9281), .B(n17311), .Z(n9282) );
  AND U9812 ( .A(n9283), .B(n9282), .Z(n9495) );
  XNOR U9813 ( .A(n9494), .B(n9495), .Z(n9496) );
  XNOR U9814 ( .A(n9497), .B(n9496), .Z(n9485) );
  XOR U9815 ( .A(b[17]), .B(a[60]), .Z(n9439) );
  NAND U9816 ( .A(n9439), .B(n18673), .Z(n9286) );
  NAND U9817 ( .A(n9284), .B(n18674), .Z(n9285) );
  NAND U9818 ( .A(n9286), .B(n9285), .Z(n9457) );
  XNOR U9819 ( .A(b[31]), .B(a[46]), .Z(n9442) );
  NANDN U9820 ( .A(n9442), .B(n19472), .Z(n9289) );
  NANDN U9821 ( .A(n9287), .B(n19473), .Z(n9288) );
  NAND U9822 ( .A(n9289), .B(n9288), .Z(n9454) );
  OR U9823 ( .A(n9290), .B(n16988), .Z(n9292) );
  XNOR U9824 ( .A(b[3]), .B(a[74]), .Z(n9445) );
  NANDN U9825 ( .A(n9445), .B(n16990), .Z(n9291) );
  AND U9826 ( .A(n9292), .B(n9291), .Z(n9455) );
  XNOR U9827 ( .A(n9454), .B(n9455), .Z(n9456) );
  XOR U9828 ( .A(n9457), .B(n9456), .Z(n9484) );
  XNOR U9829 ( .A(n9485), .B(n9484), .Z(n9486) );
  XNOR U9830 ( .A(n9487), .B(n9486), .Z(n9530) );
  NANDN U9831 ( .A(n9294), .B(n9293), .Z(n9298) );
  NAND U9832 ( .A(n9296), .B(n9295), .Z(n9297) );
  NAND U9833 ( .A(n9298), .B(n9297), .Z(n9475) );
  NANDN U9834 ( .A(n9300), .B(n9299), .Z(n9304) );
  NAND U9835 ( .A(n9302), .B(n9301), .Z(n9303) );
  NAND U9836 ( .A(n9304), .B(n9303), .Z(n9473) );
  OR U9837 ( .A(n9306), .B(n9305), .Z(n9310) );
  NANDN U9838 ( .A(n9308), .B(n9307), .Z(n9309) );
  NAND U9839 ( .A(n9310), .B(n9309), .Z(n9472) );
  XNOR U9840 ( .A(n9475), .B(n9474), .Z(n9531) );
  XNOR U9841 ( .A(n9530), .B(n9531), .Z(n9532) );
  NANDN U9842 ( .A(n9312), .B(n9311), .Z(n9316) );
  OR U9843 ( .A(n9314), .B(n9313), .Z(n9315) );
  AND U9844 ( .A(n9316), .B(n9315), .Z(n9533) );
  XNOR U9845 ( .A(n9532), .B(n9533), .Z(n9417) );
  NANDN U9846 ( .A(n9322), .B(n9321), .Z(n9326) );
  NANDN U9847 ( .A(n9324), .B(n9323), .Z(n9325) );
  NAND U9848 ( .A(n9326), .B(n9325), .Z(n9539) );
  NANDN U9849 ( .A(n9328), .B(n9327), .Z(n9332) );
  OR U9850 ( .A(n9330), .B(n9329), .Z(n9331) );
  NAND U9851 ( .A(n9332), .B(n9331), .Z(n9536) );
  NANDN U9852 ( .A(n9334), .B(n9333), .Z(n9338) );
  NAND U9853 ( .A(n9336), .B(n9335), .Z(n9337) );
  NAND U9854 ( .A(n9338), .B(n9337), .Z(n9478) );
  NANDN U9855 ( .A(n9340), .B(n9339), .Z(n9344) );
  NAND U9856 ( .A(n9342), .B(n9341), .Z(n9343) );
  AND U9857 ( .A(n9344), .B(n9343), .Z(n9479) );
  XNOR U9858 ( .A(n9478), .B(n9479), .Z(n9480) );
  XNOR U9859 ( .A(n579), .B(a[68]), .Z(n9500) );
  NAND U9860 ( .A(n17814), .B(n9500), .Z(n9347) );
  NANDN U9861 ( .A(n9345), .B(n17815), .Z(n9346) );
  NAND U9862 ( .A(n9347), .B(n9346), .Z(n9462) );
  NAND U9863 ( .A(n9348), .B(n18513), .Z(n9350) );
  XOR U9864 ( .A(b[15]), .B(a[62]), .Z(n9503) );
  NANDN U9865 ( .A(n18512), .B(n9503), .Z(n9349) );
  AND U9866 ( .A(n9350), .B(n9349), .Z(n9460) );
  NANDN U9867 ( .A(n9351), .B(n19013), .Z(n9353) );
  XNOR U9868 ( .A(n582), .B(a[56]), .Z(n9506) );
  NAND U9869 ( .A(n9506), .B(n19015), .Z(n9352) );
  AND U9870 ( .A(n9353), .B(n9352), .Z(n9461) );
  XOR U9871 ( .A(n9462), .B(n9463), .Z(n9451) );
  XNOR U9872 ( .A(b[11]), .B(a[66]), .Z(n9509) );
  OR U9873 ( .A(n9509), .B(n18194), .Z(n9356) );
  NANDN U9874 ( .A(n9354), .B(n18104), .Z(n9355) );
  NAND U9875 ( .A(n9356), .B(n9355), .Z(n9449) );
  XOR U9876 ( .A(n580), .B(a[64]), .Z(n9512) );
  NANDN U9877 ( .A(n9512), .B(n18336), .Z(n9359) );
  NANDN U9878 ( .A(n9357), .B(n18337), .Z(n9358) );
  AND U9879 ( .A(n9359), .B(n9358), .Z(n9448) );
  XNOR U9880 ( .A(n9449), .B(n9448), .Z(n9450) );
  XOR U9881 ( .A(n9451), .B(n9450), .Z(n9468) );
  NANDN U9882 ( .A(n577), .B(a[76]), .Z(n9360) );
  XOR U9883 ( .A(n17151), .B(n9360), .Z(n9362) );
  NANDN U9884 ( .A(b[0]), .B(a[75]), .Z(n9361) );
  AND U9885 ( .A(n9362), .B(n9361), .Z(n9426) );
  NAND U9886 ( .A(n19406), .B(n9363), .Z(n9365) );
  XNOR U9887 ( .A(n584), .B(a[48]), .Z(n9518) );
  NANDN U9888 ( .A(n576), .B(n9518), .Z(n9364) );
  NAND U9889 ( .A(n9365), .B(n9364), .Z(n9424) );
  NANDN U9890 ( .A(n585), .B(a[44]), .Z(n9425) );
  XNOR U9891 ( .A(n9424), .B(n9425), .Z(n9427) );
  XOR U9892 ( .A(n9426), .B(n9427), .Z(n9466) );
  XOR U9893 ( .A(b[23]), .B(a[54]), .Z(n9521) );
  NANDN U9894 ( .A(n19127), .B(n9521), .Z(n9368) );
  NANDN U9895 ( .A(n9366), .B(n19128), .Z(n9367) );
  NAND U9896 ( .A(n9368), .B(n9367), .Z(n9491) );
  NAND U9897 ( .A(n9369), .B(n17553), .Z(n9371) );
  XOR U9898 ( .A(b[7]), .B(a[70]), .Z(n9524) );
  NAND U9899 ( .A(n9524), .B(n17555), .Z(n9370) );
  NAND U9900 ( .A(n9371), .B(n9370), .Z(n9488) );
  XOR U9901 ( .A(b[25]), .B(a[52]), .Z(n9527) );
  NAND U9902 ( .A(n9527), .B(n19240), .Z(n9374) );
  NAND U9903 ( .A(n9372), .B(n19242), .Z(n9373) );
  AND U9904 ( .A(n9374), .B(n9373), .Z(n9489) );
  XNOR U9905 ( .A(n9488), .B(n9489), .Z(n9490) );
  XNOR U9906 ( .A(n9491), .B(n9490), .Z(n9467) );
  XOR U9907 ( .A(n9466), .B(n9467), .Z(n9469) );
  XNOR U9908 ( .A(n9468), .B(n9469), .Z(n9481) );
  XOR U9909 ( .A(n9480), .B(n9481), .Z(n9537) );
  XNOR U9910 ( .A(n9536), .B(n9537), .Z(n9538) );
  XOR U9911 ( .A(n9539), .B(n9538), .Z(n9415) );
  XNOR U9912 ( .A(n9414), .B(n9415), .Z(n9416) );
  XNOR U9913 ( .A(n9417), .B(n9416), .Z(n9421) );
  NAND U9914 ( .A(n9376), .B(n9375), .Z(n9380) );
  NANDN U9915 ( .A(n9378), .B(n9377), .Z(n9379) );
  NAND U9916 ( .A(n9380), .B(n9379), .Z(n9418) );
  NANDN U9917 ( .A(n9382), .B(n9381), .Z(n9386) );
  NAND U9918 ( .A(n9384), .B(n9383), .Z(n9385) );
  NAND U9919 ( .A(n9386), .B(n9385), .Z(n9419) );
  XNOR U9920 ( .A(n9418), .B(n9419), .Z(n9420) );
  XNOR U9921 ( .A(n9421), .B(n9420), .Z(n9411) );
  NANDN U9922 ( .A(n9388), .B(n9387), .Z(n9392) );
  NAND U9923 ( .A(n9390), .B(n9389), .Z(n9391) );
  NAND U9924 ( .A(n9392), .B(n9391), .Z(n9408) );
  NANDN U9925 ( .A(n9394), .B(n9393), .Z(n9398) );
  OR U9926 ( .A(n9396), .B(n9395), .Z(n9397) );
  NAND U9927 ( .A(n9398), .B(n9397), .Z(n9409) );
  XNOR U9928 ( .A(n9408), .B(n9409), .Z(n9410) );
  XNOR U9929 ( .A(n9411), .B(n9410), .Z(n9404) );
  XOR U9930 ( .A(n9405), .B(n9404), .Z(n9406) );
  XNOR U9931 ( .A(n9407), .B(n9406), .Z(n9542) );
  XNOR U9932 ( .A(n9542), .B(sreg[172]), .Z(n9544) );
  NAND U9933 ( .A(n9399), .B(sreg[171]), .Z(n9403) );
  OR U9934 ( .A(n9401), .B(n9400), .Z(n9402) );
  AND U9935 ( .A(n9403), .B(n9402), .Z(n9543) );
  XOR U9936 ( .A(n9544), .B(n9543), .Z(c[172]) );
  NANDN U9937 ( .A(n9409), .B(n9408), .Z(n9413) );
  NANDN U9938 ( .A(n9411), .B(n9410), .Z(n9412) );
  NAND U9939 ( .A(n9413), .B(n9412), .Z(n9548) );
  NANDN U9940 ( .A(n9419), .B(n9418), .Z(n9423) );
  NANDN U9941 ( .A(n9421), .B(n9420), .Z(n9422) );
  NAND U9942 ( .A(n9423), .B(n9422), .Z(n9554) );
  XNOR U9943 ( .A(n9553), .B(n9554), .Z(n9555) );
  NANDN U9944 ( .A(n9425), .B(n9424), .Z(n9429) );
  NAND U9945 ( .A(n9427), .B(n9426), .Z(n9428) );
  NAND U9946 ( .A(n9429), .B(n9428), .Z(n9632) );
  NANDN U9947 ( .A(n9430), .B(n18832), .Z(n9432) );
  XNOR U9948 ( .A(b[19]), .B(a[59]), .Z(n9577) );
  NANDN U9949 ( .A(n9577), .B(n18834), .Z(n9431) );
  NAND U9950 ( .A(n9432), .B(n9431), .Z(n9642) );
  XNOR U9951 ( .A(b[27]), .B(a[51]), .Z(n9580) );
  NANDN U9952 ( .A(n9580), .B(n19336), .Z(n9435) );
  NANDN U9953 ( .A(n9433), .B(n19337), .Z(n9434) );
  NAND U9954 ( .A(n9435), .B(n9434), .Z(n9639) );
  XOR U9955 ( .A(b[5]), .B(a[73]), .Z(n9583) );
  NAND U9956 ( .A(n9583), .B(n17310), .Z(n9438) );
  NAND U9957 ( .A(n9436), .B(n17311), .Z(n9437) );
  AND U9958 ( .A(n9438), .B(n9437), .Z(n9640) );
  XNOR U9959 ( .A(n9639), .B(n9640), .Z(n9641) );
  XNOR U9960 ( .A(n9642), .B(n9641), .Z(n9630) );
  XOR U9961 ( .A(b[17]), .B(a[61]), .Z(n9586) );
  NAND U9962 ( .A(n9586), .B(n18673), .Z(n9441) );
  NAND U9963 ( .A(n9439), .B(n18674), .Z(n9440) );
  NAND U9964 ( .A(n9441), .B(n9440), .Z(n9604) );
  XNOR U9965 ( .A(b[31]), .B(a[47]), .Z(n9589) );
  NANDN U9966 ( .A(n9589), .B(n19472), .Z(n9444) );
  NANDN U9967 ( .A(n9442), .B(n19473), .Z(n9443) );
  NAND U9968 ( .A(n9444), .B(n9443), .Z(n9601) );
  OR U9969 ( .A(n9445), .B(n16988), .Z(n9447) );
  XNOR U9970 ( .A(b[3]), .B(a[75]), .Z(n9592) );
  NANDN U9971 ( .A(n9592), .B(n16990), .Z(n9446) );
  AND U9972 ( .A(n9447), .B(n9446), .Z(n9602) );
  XNOR U9973 ( .A(n9601), .B(n9602), .Z(n9603) );
  XOR U9974 ( .A(n9604), .B(n9603), .Z(n9629) );
  XNOR U9975 ( .A(n9630), .B(n9629), .Z(n9631) );
  XNOR U9976 ( .A(n9632), .B(n9631), .Z(n9675) );
  NANDN U9977 ( .A(n9449), .B(n9448), .Z(n9453) );
  NAND U9978 ( .A(n9451), .B(n9450), .Z(n9452) );
  NAND U9979 ( .A(n9453), .B(n9452), .Z(n9620) );
  NANDN U9980 ( .A(n9455), .B(n9454), .Z(n9459) );
  NAND U9981 ( .A(n9457), .B(n9456), .Z(n9458) );
  NAND U9982 ( .A(n9459), .B(n9458), .Z(n9618) );
  OR U9983 ( .A(n9461), .B(n9460), .Z(n9465) );
  NANDN U9984 ( .A(n9463), .B(n9462), .Z(n9464) );
  NAND U9985 ( .A(n9465), .B(n9464), .Z(n9617) );
  XNOR U9986 ( .A(n9620), .B(n9619), .Z(n9676) );
  XOR U9987 ( .A(n9675), .B(n9676), .Z(n9678) );
  NANDN U9988 ( .A(n9467), .B(n9466), .Z(n9471) );
  OR U9989 ( .A(n9469), .B(n9468), .Z(n9470) );
  NAND U9990 ( .A(n9471), .B(n9470), .Z(n9677) );
  XOR U9991 ( .A(n9678), .B(n9677), .Z(n9567) );
  OR U9992 ( .A(n9473), .B(n9472), .Z(n9477) );
  NAND U9993 ( .A(n9475), .B(n9474), .Z(n9476) );
  NAND U9994 ( .A(n9477), .B(n9476), .Z(n9566) );
  NANDN U9995 ( .A(n9479), .B(n9478), .Z(n9483) );
  NANDN U9996 ( .A(n9481), .B(n9480), .Z(n9482) );
  NAND U9997 ( .A(n9483), .B(n9482), .Z(n9683) );
  NANDN U9998 ( .A(n9489), .B(n9488), .Z(n9493) );
  NAND U9999 ( .A(n9491), .B(n9490), .Z(n9492) );
  NAND U10000 ( .A(n9493), .B(n9492), .Z(n9623) );
  NANDN U10001 ( .A(n9495), .B(n9494), .Z(n9499) );
  NAND U10002 ( .A(n9497), .B(n9496), .Z(n9498) );
  AND U10003 ( .A(n9499), .B(n9498), .Z(n9624) );
  XNOR U10004 ( .A(n9623), .B(n9624), .Z(n9625) );
  XOR U10005 ( .A(n579), .B(a[69]), .Z(n9651) );
  NANDN U10006 ( .A(n9651), .B(n17814), .Z(n9502) );
  NAND U10007 ( .A(n17815), .B(n9500), .Z(n9501) );
  NAND U10008 ( .A(n9502), .B(n9501), .Z(n9609) );
  XNOR U10009 ( .A(b[15]), .B(a[63]), .Z(n9648) );
  OR U10010 ( .A(n9648), .B(n18512), .Z(n9505) );
  NAND U10011 ( .A(n9503), .B(n18513), .Z(n9504) );
  NAND U10012 ( .A(n9505), .B(n9504), .Z(n9607) );
  XOR U10013 ( .A(n582), .B(a[57]), .Z(n9645) );
  NANDN U10014 ( .A(n9645), .B(n19015), .Z(n9508) );
  NAND U10015 ( .A(n19013), .B(n9506), .Z(n9507) );
  NAND U10016 ( .A(n9508), .B(n9507), .Z(n9608) );
  XNOR U10017 ( .A(n9607), .B(n9608), .Z(n9610) );
  XOR U10018 ( .A(n9609), .B(n9610), .Z(n9598) );
  XNOR U10019 ( .A(b[11]), .B(a[67]), .Z(n9654) );
  OR U10020 ( .A(n9654), .B(n18194), .Z(n9511) );
  NANDN U10021 ( .A(n9509), .B(n18104), .Z(n9510) );
  NAND U10022 ( .A(n9511), .B(n9510), .Z(n9596) );
  XOR U10023 ( .A(n580), .B(a[65]), .Z(n9657) );
  NANDN U10024 ( .A(n9657), .B(n18336), .Z(n9514) );
  NANDN U10025 ( .A(n9512), .B(n18337), .Z(n9513) );
  AND U10026 ( .A(n9514), .B(n9513), .Z(n9595) );
  XNOR U10027 ( .A(n9596), .B(n9595), .Z(n9597) );
  XNOR U10028 ( .A(n9598), .B(n9597), .Z(n9614) );
  NANDN U10029 ( .A(n577), .B(a[77]), .Z(n9515) );
  XOR U10030 ( .A(n17151), .B(n9515), .Z(n9517) );
  NANDN U10031 ( .A(b[0]), .B(a[76]), .Z(n9516) );
  AND U10032 ( .A(n9517), .B(n9516), .Z(n9573) );
  NAND U10033 ( .A(n19406), .B(n9518), .Z(n9520) );
  XOR U10034 ( .A(n584), .B(n10083), .Z(n9663) );
  NANDN U10035 ( .A(n576), .B(n9663), .Z(n9519) );
  NAND U10036 ( .A(n9520), .B(n9519), .Z(n9571) );
  NANDN U10037 ( .A(n585), .B(a[45]), .Z(n9572) );
  XNOR U10038 ( .A(n9571), .B(n9572), .Z(n9574) );
  XNOR U10039 ( .A(n9573), .B(n9574), .Z(n9612) );
  XNOR U10040 ( .A(b[23]), .B(a[55]), .Z(n9666) );
  OR U10041 ( .A(n9666), .B(n19127), .Z(n9523) );
  NAND U10042 ( .A(n9521), .B(n19128), .Z(n9522) );
  NAND U10043 ( .A(n9523), .B(n9522), .Z(n9636) );
  NAND U10044 ( .A(n9524), .B(n17553), .Z(n9526) );
  XOR U10045 ( .A(b[7]), .B(a[71]), .Z(n9669) );
  NAND U10046 ( .A(n9669), .B(n17555), .Z(n9525) );
  NAND U10047 ( .A(n9526), .B(n9525), .Z(n9633) );
  XNOR U10048 ( .A(b[25]), .B(a[53]), .Z(n9672) );
  NANDN U10049 ( .A(n9672), .B(n19240), .Z(n9529) );
  NAND U10050 ( .A(n9527), .B(n19242), .Z(n9528) );
  AND U10051 ( .A(n9529), .B(n9528), .Z(n9634) );
  XNOR U10052 ( .A(n9633), .B(n9634), .Z(n9635) );
  XOR U10053 ( .A(n9636), .B(n9635), .Z(n9611) );
  XOR U10054 ( .A(n9614), .B(n9613), .Z(n9626) );
  XOR U10055 ( .A(n9625), .B(n9626), .Z(n9681) );
  XNOR U10056 ( .A(n9682), .B(n9681), .Z(n9684) );
  XNOR U10057 ( .A(n9683), .B(n9684), .Z(n9565) );
  XOR U10058 ( .A(n9566), .B(n9565), .Z(n9568) );
  NANDN U10059 ( .A(n9531), .B(n9530), .Z(n9535) );
  NAND U10060 ( .A(n9533), .B(n9532), .Z(n9534) );
  NAND U10061 ( .A(n9535), .B(n9534), .Z(n9559) );
  NANDN U10062 ( .A(n9537), .B(n9536), .Z(n9541) );
  NAND U10063 ( .A(n9539), .B(n9538), .Z(n9540) );
  NAND U10064 ( .A(n9541), .B(n9540), .Z(n9560) );
  XNOR U10065 ( .A(n9559), .B(n9560), .Z(n9561) );
  XOR U10066 ( .A(n9562), .B(n9561), .Z(n9556) );
  XOR U10067 ( .A(n9555), .B(n9556), .Z(n9547) );
  XOR U10068 ( .A(n9548), .B(n9547), .Z(n9549) );
  XNOR U10069 ( .A(n9550), .B(n9549), .Z(n9687) );
  XNOR U10070 ( .A(n9687), .B(sreg[173]), .Z(n9689) );
  NAND U10071 ( .A(n9542), .B(sreg[172]), .Z(n9546) );
  OR U10072 ( .A(n9544), .B(n9543), .Z(n9545) );
  AND U10073 ( .A(n9546), .B(n9545), .Z(n9688) );
  XOR U10074 ( .A(n9689), .B(n9688), .Z(c[173]) );
  NAND U10075 ( .A(n9548), .B(n9547), .Z(n9552) );
  NAND U10076 ( .A(n9550), .B(n9549), .Z(n9551) );
  NAND U10077 ( .A(n9552), .B(n9551), .Z(n9695) );
  NANDN U10078 ( .A(n9554), .B(n9553), .Z(n9558) );
  NAND U10079 ( .A(n9556), .B(n9555), .Z(n9557) );
  NAND U10080 ( .A(n9558), .B(n9557), .Z(n9693) );
  NANDN U10081 ( .A(n9560), .B(n9559), .Z(n9564) );
  NAND U10082 ( .A(n9562), .B(n9561), .Z(n9563) );
  NAND U10083 ( .A(n9564), .B(n9563), .Z(n9698) );
  NANDN U10084 ( .A(n9566), .B(n9565), .Z(n9570) );
  OR U10085 ( .A(n9568), .B(n9567), .Z(n9569) );
  NAND U10086 ( .A(n9570), .B(n9569), .Z(n9699) );
  XNOR U10087 ( .A(n9698), .B(n9699), .Z(n9700) );
  NANDN U10088 ( .A(n9572), .B(n9571), .Z(n9576) );
  NAND U10089 ( .A(n9574), .B(n9573), .Z(n9575) );
  NAND U10090 ( .A(n9576), .B(n9575), .Z(n9773) );
  NANDN U10091 ( .A(n9577), .B(n18832), .Z(n9579) );
  XNOR U10092 ( .A(b[19]), .B(a[60]), .Z(n9720) );
  NANDN U10093 ( .A(n9720), .B(n18834), .Z(n9578) );
  NAND U10094 ( .A(n9579), .B(n9578), .Z(n9783) );
  XNOR U10095 ( .A(b[27]), .B(a[52]), .Z(n9723) );
  NANDN U10096 ( .A(n9723), .B(n19336), .Z(n9582) );
  NANDN U10097 ( .A(n9580), .B(n19337), .Z(n9581) );
  NAND U10098 ( .A(n9582), .B(n9581), .Z(n9780) );
  XOR U10099 ( .A(b[5]), .B(a[74]), .Z(n9726) );
  NAND U10100 ( .A(n9726), .B(n17310), .Z(n9585) );
  NAND U10101 ( .A(n9583), .B(n17311), .Z(n9584) );
  AND U10102 ( .A(n9585), .B(n9584), .Z(n9781) );
  XNOR U10103 ( .A(n9780), .B(n9781), .Z(n9782) );
  XNOR U10104 ( .A(n9783), .B(n9782), .Z(n9771) );
  XOR U10105 ( .A(b[17]), .B(a[62]), .Z(n9729) );
  NAND U10106 ( .A(n9729), .B(n18673), .Z(n9588) );
  NAND U10107 ( .A(n9586), .B(n18674), .Z(n9587) );
  NAND U10108 ( .A(n9588), .B(n9587), .Z(n9747) );
  XNOR U10109 ( .A(b[31]), .B(a[48]), .Z(n9732) );
  NANDN U10110 ( .A(n9732), .B(n19472), .Z(n9591) );
  NANDN U10111 ( .A(n9589), .B(n19473), .Z(n9590) );
  NAND U10112 ( .A(n9591), .B(n9590), .Z(n9744) );
  OR U10113 ( .A(n9592), .B(n16988), .Z(n9594) );
  XNOR U10114 ( .A(b[3]), .B(a[76]), .Z(n9735) );
  NANDN U10115 ( .A(n9735), .B(n16990), .Z(n9593) );
  AND U10116 ( .A(n9594), .B(n9593), .Z(n9745) );
  XNOR U10117 ( .A(n9744), .B(n9745), .Z(n9746) );
  XOR U10118 ( .A(n9747), .B(n9746), .Z(n9770) );
  XNOR U10119 ( .A(n9771), .B(n9770), .Z(n9772) );
  XNOR U10120 ( .A(n9773), .B(n9772), .Z(n9711) );
  NANDN U10121 ( .A(n9596), .B(n9595), .Z(n9600) );
  NAND U10122 ( .A(n9598), .B(n9597), .Z(n9599) );
  NAND U10123 ( .A(n9600), .B(n9599), .Z(n9762) );
  NANDN U10124 ( .A(n9602), .B(n9601), .Z(n9606) );
  NAND U10125 ( .A(n9604), .B(n9603), .Z(n9605) );
  NAND U10126 ( .A(n9606), .B(n9605), .Z(n9761) );
  XNOR U10127 ( .A(n9761), .B(n9760), .Z(n9763) );
  XOR U10128 ( .A(n9762), .B(n9763), .Z(n9710) );
  XOR U10129 ( .A(n9711), .B(n9710), .Z(n9712) );
  NANDN U10130 ( .A(n9612), .B(n9611), .Z(n9616) );
  NAND U10131 ( .A(n9614), .B(n9613), .Z(n9615) );
  NAND U10132 ( .A(n9616), .B(n9615), .Z(n9713) );
  XNOR U10133 ( .A(n9712), .B(n9713), .Z(n9824) );
  OR U10134 ( .A(n9618), .B(n9617), .Z(n9622) );
  NAND U10135 ( .A(n9620), .B(n9619), .Z(n9621) );
  NAND U10136 ( .A(n9622), .B(n9621), .Z(n9823) );
  NANDN U10137 ( .A(n9624), .B(n9623), .Z(n9628) );
  NAND U10138 ( .A(n9626), .B(n9625), .Z(n9627) );
  NAND U10139 ( .A(n9628), .B(n9627), .Z(n9706) );
  NANDN U10140 ( .A(n9634), .B(n9633), .Z(n9638) );
  NAND U10141 ( .A(n9636), .B(n9635), .Z(n9637) );
  NAND U10142 ( .A(n9638), .B(n9637), .Z(n9764) );
  NANDN U10143 ( .A(n9640), .B(n9639), .Z(n9644) );
  NAND U10144 ( .A(n9642), .B(n9641), .Z(n9643) );
  AND U10145 ( .A(n9644), .B(n9643), .Z(n9765) );
  XNOR U10146 ( .A(n9764), .B(n9765), .Z(n9766) );
  XOR U10147 ( .A(n582), .B(a[58]), .Z(n9792) );
  NANDN U10148 ( .A(n9792), .B(n19015), .Z(n9647) );
  NANDN U10149 ( .A(n9645), .B(n19013), .Z(n9646) );
  NAND U10150 ( .A(n9647), .B(n9646), .Z(n9756) );
  NANDN U10151 ( .A(n9648), .B(n18513), .Z(n9650) );
  XOR U10152 ( .A(b[15]), .B(a[64]), .Z(n9789) );
  NANDN U10153 ( .A(n18512), .B(n9789), .Z(n9649) );
  AND U10154 ( .A(n9650), .B(n9649), .Z(n9757) );
  XNOR U10155 ( .A(n9756), .B(n9757), .Z(n9759) );
  XOR U10156 ( .A(n579), .B(a[70]), .Z(n9786) );
  NANDN U10157 ( .A(n9786), .B(n17814), .Z(n9653) );
  NANDN U10158 ( .A(n9651), .B(n17815), .Z(n9652) );
  NAND U10159 ( .A(n9653), .B(n9652), .Z(n9758) );
  XNOR U10160 ( .A(n9759), .B(n9758), .Z(n9752) );
  XNOR U10161 ( .A(b[11]), .B(a[68]), .Z(n9795) );
  OR U10162 ( .A(n9795), .B(n18194), .Z(n9656) );
  NANDN U10163 ( .A(n9654), .B(n18104), .Z(n9655) );
  NAND U10164 ( .A(n9656), .B(n9655), .Z(n9751) );
  XOR U10165 ( .A(n580), .B(a[66]), .Z(n9798) );
  NANDN U10166 ( .A(n9798), .B(n18336), .Z(n9659) );
  NANDN U10167 ( .A(n9657), .B(n18337), .Z(n9658) );
  NAND U10168 ( .A(n9659), .B(n9658), .Z(n9750) );
  XNOR U10169 ( .A(n9751), .B(n9750), .Z(n9753) );
  XNOR U10170 ( .A(n9752), .B(n9753), .Z(n9741) );
  NANDN U10171 ( .A(n577), .B(a[78]), .Z(n9660) );
  XOR U10172 ( .A(n17151), .B(n9660), .Z(n9662) );
  NANDN U10173 ( .A(b[0]), .B(a[77]), .Z(n9661) );
  AND U10174 ( .A(n9662), .B(n9661), .Z(n9716) );
  NAND U10175 ( .A(n19406), .B(n9663), .Z(n9665) );
  XNOR U10176 ( .A(n584), .B(a[50]), .Z(n9804) );
  NANDN U10177 ( .A(n576), .B(n9804), .Z(n9664) );
  NAND U10178 ( .A(n9665), .B(n9664), .Z(n9714) );
  NANDN U10179 ( .A(n585), .B(a[46]), .Z(n9715) );
  XNOR U10180 ( .A(n9714), .B(n9715), .Z(n9717) );
  XNOR U10181 ( .A(n9716), .B(n9717), .Z(n9739) );
  XOR U10182 ( .A(b[23]), .B(a[56]), .Z(n9807) );
  NANDN U10183 ( .A(n19127), .B(n9807), .Z(n9668) );
  NANDN U10184 ( .A(n9666), .B(n19128), .Z(n9667) );
  NAND U10185 ( .A(n9668), .B(n9667), .Z(n9777) );
  NAND U10186 ( .A(n9669), .B(n17553), .Z(n9671) );
  XOR U10187 ( .A(b[7]), .B(a[72]), .Z(n9810) );
  NAND U10188 ( .A(n9810), .B(n17555), .Z(n9670) );
  NAND U10189 ( .A(n9671), .B(n9670), .Z(n9774) );
  XOR U10190 ( .A(b[25]), .B(a[54]), .Z(n9813) );
  NAND U10191 ( .A(n9813), .B(n19240), .Z(n9674) );
  NANDN U10192 ( .A(n9672), .B(n19242), .Z(n9673) );
  AND U10193 ( .A(n9674), .B(n9673), .Z(n9775) );
  XNOR U10194 ( .A(n9774), .B(n9775), .Z(n9776) );
  XOR U10195 ( .A(n9777), .B(n9776), .Z(n9738) );
  XOR U10196 ( .A(n9741), .B(n9740), .Z(n9767) );
  XNOR U10197 ( .A(n9766), .B(n9767), .Z(n9704) );
  XNOR U10198 ( .A(n9705), .B(n9704), .Z(n9707) );
  XNOR U10199 ( .A(n9706), .B(n9707), .Z(n9822) );
  XOR U10200 ( .A(n9823), .B(n9822), .Z(n9825) );
  NANDN U10201 ( .A(n9676), .B(n9675), .Z(n9680) );
  OR U10202 ( .A(n9678), .B(n9677), .Z(n9679) );
  NAND U10203 ( .A(n9680), .B(n9679), .Z(n9816) );
  NAND U10204 ( .A(n9682), .B(n9681), .Z(n9686) );
  NANDN U10205 ( .A(n9684), .B(n9683), .Z(n9685) );
  NAND U10206 ( .A(n9686), .B(n9685), .Z(n9817) );
  XNOR U10207 ( .A(n9816), .B(n9817), .Z(n9818) );
  XOR U10208 ( .A(n9819), .B(n9818), .Z(n9701) );
  XOR U10209 ( .A(n9700), .B(n9701), .Z(n9692) );
  XOR U10210 ( .A(n9693), .B(n9692), .Z(n9694) );
  XNOR U10211 ( .A(n9695), .B(n9694), .Z(n9828) );
  XNOR U10212 ( .A(n9828), .B(sreg[174]), .Z(n9830) );
  NAND U10213 ( .A(n9687), .B(sreg[173]), .Z(n9691) );
  OR U10214 ( .A(n9689), .B(n9688), .Z(n9690) );
  AND U10215 ( .A(n9691), .B(n9690), .Z(n9829) );
  XOR U10216 ( .A(n9830), .B(n9829), .Z(c[174]) );
  NAND U10217 ( .A(n9693), .B(n9692), .Z(n9697) );
  NAND U10218 ( .A(n9695), .B(n9694), .Z(n9696) );
  NAND U10219 ( .A(n9697), .B(n9696), .Z(n9836) );
  NANDN U10220 ( .A(n9699), .B(n9698), .Z(n9703) );
  NAND U10221 ( .A(n9701), .B(n9700), .Z(n9702) );
  NAND U10222 ( .A(n9703), .B(n9702), .Z(n9833) );
  NAND U10223 ( .A(n9705), .B(n9704), .Z(n9709) );
  NANDN U10224 ( .A(n9707), .B(n9706), .Z(n9708) );
  NAND U10225 ( .A(n9709), .B(n9708), .Z(n9959) );
  XNOR U10226 ( .A(n9959), .B(n9960), .Z(n9961) );
  NANDN U10227 ( .A(n9715), .B(n9714), .Z(n9719) );
  NAND U10228 ( .A(n9717), .B(n9716), .Z(n9718) );
  NAND U10229 ( .A(n9719), .B(n9718), .Z(n9904) );
  NANDN U10230 ( .A(n9720), .B(n18832), .Z(n9722) );
  XNOR U10231 ( .A(b[19]), .B(a[61]), .Z(n9851) );
  NANDN U10232 ( .A(n9851), .B(n18834), .Z(n9721) );
  NAND U10233 ( .A(n9722), .B(n9721), .Z(n9938) );
  XOR U10234 ( .A(b[27]), .B(n10660), .Z(n9854) );
  NANDN U10235 ( .A(n9854), .B(n19336), .Z(n9725) );
  NANDN U10236 ( .A(n9723), .B(n19337), .Z(n9724) );
  NAND U10237 ( .A(n9725), .B(n9724), .Z(n9935) );
  XOR U10238 ( .A(b[5]), .B(a[75]), .Z(n9857) );
  NAND U10239 ( .A(n9857), .B(n17310), .Z(n9728) );
  NAND U10240 ( .A(n9726), .B(n17311), .Z(n9727) );
  AND U10241 ( .A(n9728), .B(n9727), .Z(n9936) );
  XNOR U10242 ( .A(n9935), .B(n9936), .Z(n9937) );
  XNOR U10243 ( .A(n9938), .B(n9937), .Z(n9902) );
  XOR U10244 ( .A(b[17]), .B(a[63]), .Z(n9860) );
  NAND U10245 ( .A(n9860), .B(n18673), .Z(n9731) );
  NAND U10246 ( .A(n9729), .B(n18674), .Z(n9730) );
  NAND U10247 ( .A(n9731), .B(n9730), .Z(n9878) );
  XOR U10248 ( .A(b[31]), .B(n10083), .Z(n9863) );
  NANDN U10249 ( .A(n9863), .B(n19472), .Z(n9734) );
  NANDN U10250 ( .A(n9732), .B(n19473), .Z(n9733) );
  NAND U10251 ( .A(n9734), .B(n9733), .Z(n9875) );
  OR U10252 ( .A(n9735), .B(n16988), .Z(n9737) );
  XNOR U10253 ( .A(b[3]), .B(a[77]), .Z(n9866) );
  NANDN U10254 ( .A(n9866), .B(n16990), .Z(n9736) );
  AND U10255 ( .A(n9737), .B(n9736), .Z(n9876) );
  XNOR U10256 ( .A(n9875), .B(n9876), .Z(n9877) );
  XOR U10257 ( .A(n9878), .B(n9877), .Z(n9901) );
  XNOR U10258 ( .A(n9902), .B(n9901), .Z(n9903) );
  XNOR U10259 ( .A(n9904), .B(n9903), .Z(n9953) );
  NANDN U10260 ( .A(n9739), .B(n9738), .Z(n9743) );
  NANDN U10261 ( .A(n9741), .B(n9740), .Z(n9742) );
  NAND U10262 ( .A(n9743), .B(n9742), .Z(n9954) );
  XNOR U10263 ( .A(n9953), .B(n9954), .Z(n9955) );
  NANDN U10264 ( .A(n9745), .B(n9744), .Z(n9749) );
  NAND U10265 ( .A(n9747), .B(n9746), .Z(n9748) );
  NAND U10266 ( .A(n9749), .B(n9748), .Z(n9894) );
  OR U10267 ( .A(n9751), .B(n9750), .Z(n9755) );
  NANDN U10268 ( .A(n9753), .B(n9752), .Z(n9754) );
  NAND U10269 ( .A(n9755), .B(n9754), .Z(n9892) );
  XNOR U10270 ( .A(n9892), .B(n9891), .Z(n9893) );
  XOR U10271 ( .A(n9894), .B(n9893), .Z(n9956) );
  XOR U10272 ( .A(n9955), .B(n9956), .Z(n9967) );
  NANDN U10273 ( .A(n9765), .B(n9764), .Z(n9769) );
  NANDN U10274 ( .A(n9767), .B(n9766), .Z(n9768) );
  NAND U10275 ( .A(n9769), .B(n9768), .Z(n9950) );
  NANDN U10276 ( .A(n9775), .B(n9774), .Z(n9779) );
  NAND U10277 ( .A(n9777), .B(n9776), .Z(n9778) );
  NAND U10278 ( .A(n9779), .B(n9778), .Z(n9895) );
  NANDN U10279 ( .A(n9781), .B(n9780), .Z(n9785) );
  NAND U10280 ( .A(n9783), .B(n9782), .Z(n9784) );
  AND U10281 ( .A(n9785), .B(n9784), .Z(n9896) );
  XNOR U10282 ( .A(n9895), .B(n9896), .Z(n9897) );
  XOR U10283 ( .A(n579), .B(a[71]), .Z(n9911) );
  NANDN U10284 ( .A(n9911), .B(n17814), .Z(n9788) );
  NANDN U10285 ( .A(n9786), .B(n17815), .Z(n9787) );
  NAND U10286 ( .A(n9788), .B(n9787), .Z(n9883) );
  XNOR U10287 ( .A(b[15]), .B(a[65]), .Z(n9908) );
  OR U10288 ( .A(n9908), .B(n18512), .Z(n9791) );
  NAND U10289 ( .A(n9789), .B(n18513), .Z(n9790) );
  NAND U10290 ( .A(n9791), .B(n9790), .Z(n9881) );
  XOR U10291 ( .A(n582), .B(a[59]), .Z(n9905) );
  NANDN U10292 ( .A(n9905), .B(n19015), .Z(n9794) );
  NANDN U10293 ( .A(n9792), .B(n19013), .Z(n9793) );
  NAND U10294 ( .A(n9794), .B(n9793), .Z(n9882) );
  XNOR U10295 ( .A(n9881), .B(n9882), .Z(n9884) );
  XOR U10296 ( .A(n9883), .B(n9884), .Z(n9872) );
  XNOR U10297 ( .A(b[11]), .B(a[69]), .Z(n9914) );
  OR U10298 ( .A(n9914), .B(n18194), .Z(n9797) );
  NANDN U10299 ( .A(n9795), .B(n18104), .Z(n9796) );
  NAND U10300 ( .A(n9797), .B(n9796), .Z(n9870) );
  XOR U10301 ( .A(n580), .B(a[67]), .Z(n9917) );
  NANDN U10302 ( .A(n9917), .B(n18336), .Z(n9800) );
  NANDN U10303 ( .A(n9798), .B(n18337), .Z(n9799) );
  AND U10304 ( .A(n9800), .B(n9799), .Z(n9869) );
  XNOR U10305 ( .A(n9870), .B(n9869), .Z(n9871) );
  XNOR U10306 ( .A(n9872), .B(n9871), .Z(n9888) );
  NANDN U10307 ( .A(n577), .B(a[79]), .Z(n9801) );
  XOR U10308 ( .A(n17151), .B(n9801), .Z(n9803) );
  NANDN U10309 ( .A(b[0]), .B(a[78]), .Z(n9802) );
  AND U10310 ( .A(n9803), .B(n9802), .Z(n9847) );
  NAND U10311 ( .A(n19406), .B(n9804), .Z(n9806) );
  XNOR U10312 ( .A(n584), .B(a[51]), .Z(n9923) );
  NANDN U10313 ( .A(n576), .B(n9923), .Z(n9805) );
  NAND U10314 ( .A(n9806), .B(n9805), .Z(n9845) );
  NANDN U10315 ( .A(n585), .B(a[47]), .Z(n9846) );
  XNOR U10316 ( .A(n9845), .B(n9846), .Z(n9848) );
  XNOR U10317 ( .A(n9847), .B(n9848), .Z(n9886) );
  XOR U10318 ( .A(b[23]), .B(a[57]), .Z(n9926) );
  NANDN U10319 ( .A(n19127), .B(n9926), .Z(n9809) );
  NAND U10320 ( .A(n9807), .B(n19128), .Z(n9808) );
  NAND U10321 ( .A(n9809), .B(n9808), .Z(n9944) );
  NAND U10322 ( .A(n9810), .B(n17553), .Z(n9812) );
  XOR U10323 ( .A(b[7]), .B(a[73]), .Z(n9929) );
  NAND U10324 ( .A(n9929), .B(n17555), .Z(n9811) );
  NAND U10325 ( .A(n9812), .B(n9811), .Z(n9941) );
  XNOR U10326 ( .A(b[25]), .B(a[55]), .Z(n9932) );
  NANDN U10327 ( .A(n9932), .B(n19240), .Z(n9815) );
  NAND U10328 ( .A(n9813), .B(n19242), .Z(n9814) );
  AND U10329 ( .A(n9815), .B(n9814), .Z(n9942) );
  XNOR U10330 ( .A(n9941), .B(n9942), .Z(n9943) );
  XOR U10331 ( .A(n9944), .B(n9943), .Z(n9885) );
  XOR U10332 ( .A(n9888), .B(n9887), .Z(n9898) );
  XOR U10333 ( .A(n9897), .B(n9898), .Z(n9947) );
  XOR U10334 ( .A(n9948), .B(n9947), .Z(n9949) );
  XNOR U10335 ( .A(n9950), .B(n9949), .Z(n9965) );
  XNOR U10336 ( .A(n9966), .B(n9965), .Z(n9968) );
  XNOR U10337 ( .A(n9967), .B(n9968), .Z(n9962) );
  XOR U10338 ( .A(n9961), .B(n9962), .Z(n9842) );
  NANDN U10339 ( .A(n9817), .B(n9816), .Z(n9821) );
  NAND U10340 ( .A(n9819), .B(n9818), .Z(n9820) );
  NAND U10341 ( .A(n9821), .B(n9820), .Z(n9839) );
  NANDN U10342 ( .A(n9823), .B(n9822), .Z(n9827) );
  OR U10343 ( .A(n9825), .B(n9824), .Z(n9826) );
  NAND U10344 ( .A(n9827), .B(n9826), .Z(n9840) );
  XNOR U10345 ( .A(n9839), .B(n9840), .Z(n9841) );
  XNOR U10346 ( .A(n9842), .B(n9841), .Z(n9834) );
  XNOR U10347 ( .A(n9833), .B(n9834), .Z(n9835) );
  XNOR U10348 ( .A(n9836), .B(n9835), .Z(n9971) );
  XNOR U10349 ( .A(n9971), .B(sreg[175]), .Z(n9973) );
  NAND U10350 ( .A(n9828), .B(sreg[174]), .Z(n9832) );
  OR U10351 ( .A(n9830), .B(n9829), .Z(n9831) );
  AND U10352 ( .A(n9832), .B(n9831), .Z(n9972) );
  XOR U10353 ( .A(n9973), .B(n9972), .Z(c[175]) );
  NANDN U10354 ( .A(n9834), .B(n9833), .Z(n9838) );
  NAND U10355 ( .A(n9836), .B(n9835), .Z(n9837) );
  NAND U10356 ( .A(n9838), .B(n9837), .Z(n9979) );
  NANDN U10357 ( .A(n9840), .B(n9839), .Z(n9844) );
  NAND U10358 ( .A(n9842), .B(n9841), .Z(n9843) );
  NAND U10359 ( .A(n9844), .B(n9843), .Z(n9977) );
  NANDN U10360 ( .A(n9846), .B(n9845), .Z(n9850) );
  NAND U10361 ( .A(n9848), .B(n9847), .Z(n9849) );
  NAND U10362 ( .A(n9850), .B(n9849), .Z(n10055) );
  NANDN U10363 ( .A(n9851), .B(n18832), .Z(n9853) );
  XNOR U10364 ( .A(b[19]), .B(a[62]), .Z(n10002) );
  NANDN U10365 ( .A(n10002), .B(n18834), .Z(n9852) );
  NAND U10366 ( .A(n9853), .B(n9852), .Z(n10065) );
  XNOR U10367 ( .A(b[27]), .B(a[54]), .Z(n10005) );
  NANDN U10368 ( .A(n10005), .B(n19336), .Z(n9856) );
  NANDN U10369 ( .A(n9854), .B(n19337), .Z(n9855) );
  NAND U10370 ( .A(n9856), .B(n9855), .Z(n10062) );
  XOR U10371 ( .A(b[5]), .B(a[76]), .Z(n10008) );
  NAND U10372 ( .A(n10008), .B(n17310), .Z(n9859) );
  NAND U10373 ( .A(n9857), .B(n17311), .Z(n9858) );
  AND U10374 ( .A(n9859), .B(n9858), .Z(n10063) );
  XNOR U10375 ( .A(n10062), .B(n10063), .Z(n10064) );
  XNOR U10376 ( .A(n10065), .B(n10064), .Z(n10053) );
  XOR U10377 ( .A(b[17]), .B(a[64]), .Z(n10011) );
  NAND U10378 ( .A(n10011), .B(n18673), .Z(n9862) );
  NAND U10379 ( .A(n9860), .B(n18674), .Z(n9861) );
  NAND U10380 ( .A(n9862), .B(n9861), .Z(n10029) );
  XNOR U10381 ( .A(b[31]), .B(a[50]), .Z(n10014) );
  NANDN U10382 ( .A(n10014), .B(n19472), .Z(n9865) );
  NANDN U10383 ( .A(n9863), .B(n19473), .Z(n9864) );
  NAND U10384 ( .A(n9865), .B(n9864), .Z(n10026) );
  OR U10385 ( .A(n9866), .B(n16988), .Z(n9868) );
  XNOR U10386 ( .A(b[3]), .B(a[78]), .Z(n10017) );
  NANDN U10387 ( .A(n10017), .B(n16990), .Z(n9867) );
  AND U10388 ( .A(n9868), .B(n9867), .Z(n10027) );
  XNOR U10389 ( .A(n10026), .B(n10027), .Z(n10028) );
  XOR U10390 ( .A(n10029), .B(n10028), .Z(n10052) );
  XNOR U10391 ( .A(n10053), .B(n10052), .Z(n10054) );
  XNOR U10392 ( .A(n10055), .B(n10054), .Z(n9993) );
  NANDN U10393 ( .A(n9870), .B(n9869), .Z(n9874) );
  NAND U10394 ( .A(n9872), .B(n9871), .Z(n9873) );
  NAND U10395 ( .A(n9874), .B(n9873), .Z(n10044) );
  NANDN U10396 ( .A(n9876), .B(n9875), .Z(n9880) );
  NAND U10397 ( .A(n9878), .B(n9877), .Z(n9879) );
  NAND U10398 ( .A(n9880), .B(n9879), .Z(n10043) );
  XNOR U10399 ( .A(n10043), .B(n10042), .Z(n10045) );
  XOR U10400 ( .A(n10044), .B(n10045), .Z(n9992) );
  XOR U10401 ( .A(n9993), .B(n9992), .Z(n9994) );
  NANDN U10402 ( .A(n9886), .B(n9885), .Z(n9890) );
  NAND U10403 ( .A(n9888), .B(n9887), .Z(n9889) );
  AND U10404 ( .A(n9890), .B(n9889), .Z(n9995) );
  XNOR U10405 ( .A(n9994), .B(n9995), .Z(n10102) );
  NANDN U10406 ( .A(n9896), .B(n9895), .Z(n9900) );
  NAND U10407 ( .A(n9898), .B(n9897), .Z(n9899) );
  NAND U10408 ( .A(n9900), .B(n9899), .Z(n9989) );
  XNOR U10409 ( .A(b[21]), .B(a[60]), .Z(n10074) );
  NANDN U10410 ( .A(n10074), .B(n19015), .Z(n9907) );
  NANDN U10411 ( .A(n9905), .B(n19013), .Z(n9906) );
  NAND U10412 ( .A(n9907), .B(n9906), .Z(n10038) );
  NANDN U10413 ( .A(n9908), .B(n18513), .Z(n9910) );
  XOR U10414 ( .A(b[15]), .B(a[66]), .Z(n10071) );
  NANDN U10415 ( .A(n18512), .B(n10071), .Z(n9909) );
  AND U10416 ( .A(n9910), .B(n9909), .Z(n10039) );
  XNOR U10417 ( .A(n10038), .B(n10039), .Z(n10041) );
  XNOR U10418 ( .A(b[9]), .B(a[72]), .Z(n10068) );
  NANDN U10419 ( .A(n10068), .B(n17814), .Z(n9913) );
  NANDN U10420 ( .A(n9911), .B(n17815), .Z(n9912) );
  NAND U10421 ( .A(n9913), .B(n9912), .Z(n10040) );
  XNOR U10422 ( .A(n10041), .B(n10040), .Z(n10034) );
  XNOR U10423 ( .A(b[11]), .B(a[70]), .Z(n10077) );
  OR U10424 ( .A(n10077), .B(n18194), .Z(n9916) );
  NANDN U10425 ( .A(n9914), .B(n18104), .Z(n9915) );
  NAND U10426 ( .A(n9916), .B(n9915), .Z(n10033) );
  XOR U10427 ( .A(n580), .B(a[68]), .Z(n10080) );
  NANDN U10428 ( .A(n10080), .B(n18336), .Z(n9919) );
  NANDN U10429 ( .A(n9917), .B(n18337), .Z(n9918) );
  NAND U10430 ( .A(n9919), .B(n9918), .Z(n10032) );
  XNOR U10431 ( .A(n10033), .B(n10032), .Z(n10035) );
  XNOR U10432 ( .A(n10034), .B(n10035), .Z(n10023) );
  NANDN U10433 ( .A(n577), .B(a[80]), .Z(n9920) );
  XOR U10434 ( .A(n17151), .B(n9920), .Z(n9922) );
  NANDN U10435 ( .A(b[0]), .B(a[79]), .Z(n9921) );
  AND U10436 ( .A(n9922), .B(n9921), .Z(n9998) );
  NAND U10437 ( .A(n19406), .B(n9923), .Z(n9925) );
  XNOR U10438 ( .A(b[29]), .B(a[52]), .Z(n10084) );
  OR U10439 ( .A(n10084), .B(n576), .Z(n9924) );
  NAND U10440 ( .A(n9925), .B(n9924), .Z(n9996) );
  NANDN U10441 ( .A(n585), .B(a[48]), .Z(n9997) );
  XNOR U10442 ( .A(n9996), .B(n9997), .Z(n9999) );
  XNOR U10443 ( .A(n9998), .B(n9999), .Z(n10021) );
  XOR U10444 ( .A(b[23]), .B(a[58]), .Z(n10090) );
  NANDN U10445 ( .A(n19127), .B(n10090), .Z(n9928) );
  NAND U10446 ( .A(n9926), .B(n19128), .Z(n9927) );
  NAND U10447 ( .A(n9928), .B(n9927), .Z(n10059) );
  NAND U10448 ( .A(n9929), .B(n17553), .Z(n9931) );
  XOR U10449 ( .A(b[7]), .B(a[74]), .Z(n10093) );
  NAND U10450 ( .A(n10093), .B(n17555), .Z(n9930) );
  NAND U10451 ( .A(n9931), .B(n9930), .Z(n10056) );
  XOR U10452 ( .A(b[25]), .B(a[56]), .Z(n10096) );
  NAND U10453 ( .A(n10096), .B(n19240), .Z(n9934) );
  NANDN U10454 ( .A(n9932), .B(n19242), .Z(n9933) );
  AND U10455 ( .A(n9934), .B(n9933), .Z(n10057) );
  XNOR U10456 ( .A(n10056), .B(n10057), .Z(n10058) );
  XOR U10457 ( .A(n10059), .B(n10058), .Z(n10020) );
  XNOR U10458 ( .A(n10023), .B(n10022), .Z(n10049) );
  NANDN U10459 ( .A(n9936), .B(n9935), .Z(n9940) );
  NAND U10460 ( .A(n9938), .B(n9937), .Z(n9939) );
  NAND U10461 ( .A(n9940), .B(n9939), .Z(n10047) );
  NANDN U10462 ( .A(n9942), .B(n9941), .Z(n9946) );
  NAND U10463 ( .A(n9944), .B(n9943), .Z(n9945) );
  AND U10464 ( .A(n9946), .B(n9945), .Z(n10046) );
  XNOR U10465 ( .A(n10047), .B(n10046), .Z(n10048) );
  XNOR U10466 ( .A(n10049), .B(n10048), .Z(n9987) );
  XNOR U10467 ( .A(n9986), .B(n9987), .Z(n9988) );
  XOR U10468 ( .A(n9989), .B(n9988), .Z(n10100) );
  XNOR U10469 ( .A(n10099), .B(n10100), .Z(n10101) );
  XNOR U10470 ( .A(n10102), .B(n10101), .Z(n10106) );
  NAND U10471 ( .A(n9948), .B(n9947), .Z(n9952) );
  NAND U10472 ( .A(n9950), .B(n9949), .Z(n9951) );
  NAND U10473 ( .A(n9952), .B(n9951), .Z(n10103) );
  NANDN U10474 ( .A(n9954), .B(n9953), .Z(n9958) );
  NAND U10475 ( .A(n9956), .B(n9955), .Z(n9957) );
  NAND U10476 ( .A(n9958), .B(n9957), .Z(n10104) );
  XNOR U10477 ( .A(n10103), .B(n10104), .Z(n10105) );
  XNOR U10478 ( .A(n10106), .B(n10105), .Z(n9983) );
  NANDN U10479 ( .A(n9960), .B(n9959), .Z(n9964) );
  NANDN U10480 ( .A(n9962), .B(n9961), .Z(n9963) );
  NAND U10481 ( .A(n9964), .B(n9963), .Z(n9981) );
  OR U10482 ( .A(n9966), .B(n9965), .Z(n9970) );
  OR U10483 ( .A(n9968), .B(n9967), .Z(n9969) );
  AND U10484 ( .A(n9970), .B(n9969), .Z(n9980) );
  XNOR U10485 ( .A(n9981), .B(n9980), .Z(n9982) );
  XNOR U10486 ( .A(n9983), .B(n9982), .Z(n9976) );
  XOR U10487 ( .A(n9977), .B(n9976), .Z(n9978) );
  XNOR U10488 ( .A(n9979), .B(n9978), .Z(n10109) );
  XNOR U10489 ( .A(n10109), .B(sreg[176]), .Z(n10111) );
  NAND U10490 ( .A(n9971), .B(sreg[175]), .Z(n9975) );
  OR U10491 ( .A(n9973), .B(n9972), .Z(n9974) );
  AND U10492 ( .A(n9975), .B(n9974), .Z(n10110) );
  XOR U10493 ( .A(n10111), .B(n10110), .Z(c[176]) );
  NANDN U10494 ( .A(n9981), .B(n9980), .Z(n9985) );
  NANDN U10495 ( .A(n9983), .B(n9982), .Z(n9984) );
  NAND U10496 ( .A(n9985), .B(n9984), .Z(n10114) );
  NANDN U10497 ( .A(n9987), .B(n9986), .Z(n9991) );
  NAND U10498 ( .A(n9989), .B(n9988), .Z(n9990) );
  NAND U10499 ( .A(n9991), .B(n9990), .Z(n10244) );
  XNOR U10500 ( .A(n10244), .B(n10245), .Z(n10246) );
  NANDN U10501 ( .A(n9997), .B(n9996), .Z(n10001) );
  NAND U10502 ( .A(n9999), .B(n9998), .Z(n10000) );
  NAND U10503 ( .A(n10001), .B(n10000), .Z(n10187) );
  NANDN U10504 ( .A(n10002), .B(n18832), .Z(n10004) );
  XNOR U10505 ( .A(b[19]), .B(a[63]), .Z(n10156) );
  NANDN U10506 ( .A(n10156), .B(n18834), .Z(n10003) );
  NAND U10507 ( .A(n10004), .B(n10003), .Z(n10199) );
  XOR U10508 ( .A(b[27]), .B(n10959), .Z(n10159) );
  NANDN U10509 ( .A(n10159), .B(n19336), .Z(n10007) );
  NANDN U10510 ( .A(n10005), .B(n19337), .Z(n10006) );
  NAND U10511 ( .A(n10007), .B(n10006), .Z(n10196) );
  XOR U10512 ( .A(b[5]), .B(a[77]), .Z(n10162) );
  NAND U10513 ( .A(n10162), .B(n17310), .Z(n10010) );
  NAND U10514 ( .A(n10008), .B(n17311), .Z(n10009) );
  AND U10515 ( .A(n10010), .B(n10009), .Z(n10197) );
  XNOR U10516 ( .A(n10196), .B(n10197), .Z(n10198) );
  XNOR U10517 ( .A(n10199), .B(n10198), .Z(n10184) );
  XNOR U10518 ( .A(b[17]), .B(a[65]), .Z(n10165) );
  NANDN U10519 ( .A(n10165), .B(n18673), .Z(n10013) );
  NAND U10520 ( .A(n10011), .B(n18674), .Z(n10012) );
  NAND U10521 ( .A(n10013), .B(n10012), .Z(n10140) );
  XNOR U10522 ( .A(b[31]), .B(a[51]), .Z(n10168) );
  NANDN U10523 ( .A(n10168), .B(n19472), .Z(n10016) );
  NANDN U10524 ( .A(n10014), .B(n19473), .Z(n10015) );
  AND U10525 ( .A(n10016), .B(n10015), .Z(n10138) );
  OR U10526 ( .A(n10017), .B(n16988), .Z(n10019) );
  XNOR U10527 ( .A(b[3]), .B(a[79]), .Z(n10171) );
  NANDN U10528 ( .A(n10171), .B(n16990), .Z(n10018) );
  AND U10529 ( .A(n10019), .B(n10018), .Z(n10139) );
  XOR U10530 ( .A(n10140), .B(n10141), .Z(n10185) );
  XOR U10531 ( .A(n10184), .B(n10185), .Z(n10186) );
  XNOR U10532 ( .A(n10187), .B(n10186), .Z(n10238) );
  NANDN U10533 ( .A(n10021), .B(n10020), .Z(n10025) );
  NANDN U10534 ( .A(n10023), .B(n10022), .Z(n10024) );
  NAND U10535 ( .A(n10025), .B(n10024), .Z(n10239) );
  XNOR U10536 ( .A(n10238), .B(n10239), .Z(n10240) );
  NANDN U10537 ( .A(n10027), .B(n10026), .Z(n10031) );
  NAND U10538 ( .A(n10029), .B(n10028), .Z(n10030) );
  NAND U10539 ( .A(n10031), .B(n10030), .Z(n10177) );
  OR U10540 ( .A(n10033), .B(n10032), .Z(n10037) );
  NANDN U10541 ( .A(n10035), .B(n10034), .Z(n10036) );
  NAND U10542 ( .A(n10037), .B(n10036), .Z(n10175) );
  XNOR U10543 ( .A(n10175), .B(n10174), .Z(n10176) );
  XOR U10544 ( .A(n10177), .B(n10176), .Z(n10241) );
  XOR U10545 ( .A(n10240), .B(n10241), .Z(n10253) );
  NANDN U10546 ( .A(n10047), .B(n10046), .Z(n10051) );
  NANDN U10547 ( .A(n10049), .B(n10048), .Z(n10050) );
  NAND U10548 ( .A(n10051), .B(n10050), .Z(n10235) );
  NANDN U10549 ( .A(n10057), .B(n10056), .Z(n10061) );
  NAND U10550 ( .A(n10059), .B(n10058), .Z(n10060) );
  NAND U10551 ( .A(n10061), .B(n10060), .Z(n10178) );
  NANDN U10552 ( .A(n10063), .B(n10062), .Z(n10067) );
  NAND U10553 ( .A(n10065), .B(n10064), .Z(n10066) );
  AND U10554 ( .A(n10067), .B(n10066), .Z(n10179) );
  XNOR U10555 ( .A(n10178), .B(n10179), .Z(n10180) );
  XNOR U10556 ( .A(b[9]), .B(a[73]), .Z(n10202) );
  NANDN U10557 ( .A(n10202), .B(n17814), .Z(n10070) );
  NANDN U10558 ( .A(n10068), .B(n17815), .Z(n10069) );
  NAND U10559 ( .A(n10070), .B(n10069), .Z(n10146) );
  NAND U10560 ( .A(n10071), .B(n18513), .Z(n10073) );
  XOR U10561 ( .A(b[15]), .B(a[67]), .Z(n10205) );
  NANDN U10562 ( .A(n18512), .B(n10205), .Z(n10072) );
  AND U10563 ( .A(n10073), .B(n10072), .Z(n10144) );
  NANDN U10564 ( .A(n10074), .B(n19013), .Z(n10076) );
  XNOR U10565 ( .A(b[21]), .B(a[61]), .Z(n10208) );
  NANDN U10566 ( .A(n10208), .B(n19015), .Z(n10075) );
  AND U10567 ( .A(n10076), .B(n10075), .Z(n10145) );
  XOR U10568 ( .A(n10146), .B(n10147), .Z(n10135) );
  XNOR U10569 ( .A(b[11]), .B(a[71]), .Z(n10211) );
  OR U10570 ( .A(n10211), .B(n18194), .Z(n10079) );
  NANDN U10571 ( .A(n10077), .B(n18104), .Z(n10078) );
  NAND U10572 ( .A(n10079), .B(n10078), .Z(n10133) );
  XOR U10573 ( .A(n580), .B(a[69]), .Z(n10214) );
  NANDN U10574 ( .A(n10214), .B(n18336), .Z(n10082) );
  NANDN U10575 ( .A(n10080), .B(n18337), .Z(n10081) );
  NAND U10576 ( .A(n10082), .B(n10081), .Z(n10132) );
  XOR U10577 ( .A(n10135), .B(n10134), .Z(n10129) );
  ANDN U10578 ( .B(b[31]), .A(n10083), .Z(n10150) );
  NANDN U10579 ( .A(n10084), .B(n19406), .Z(n10086) );
  XNOR U10580 ( .A(n584), .B(a[53]), .Z(n10220) );
  NANDN U10581 ( .A(n576), .B(n10220), .Z(n10085) );
  NAND U10582 ( .A(n10086), .B(n10085), .Z(n10151) );
  XOR U10583 ( .A(n10150), .B(n10151), .Z(n10152) );
  NANDN U10584 ( .A(n577), .B(a[81]), .Z(n10087) );
  XOR U10585 ( .A(n17151), .B(n10087), .Z(n10089) );
  IV U10586 ( .A(a[80]), .Z(n14551) );
  NANDN U10587 ( .A(n14551), .B(n577), .Z(n10088) );
  AND U10588 ( .A(n10089), .B(n10088), .Z(n10153) );
  XNOR U10589 ( .A(n10152), .B(n10153), .Z(n10126) );
  XOR U10590 ( .A(b[23]), .B(a[59]), .Z(n10223) );
  NANDN U10591 ( .A(n19127), .B(n10223), .Z(n10092) );
  NAND U10592 ( .A(n10090), .B(n19128), .Z(n10091) );
  NAND U10593 ( .A(n10092), .B(n10091), .Z(n10193) );
  NAND U10594 ( .A(n10093), .B(n17553), .Z(n10095) );
  XOR U10595 ( .A(b[7]), .B(a[75]), .Z(n10226) );
  NAND U10596 ( .A(n10226), .B(n17555), .Z(n10094) );
  NAND U10597 ( .A(n10095), .B(n10094), .Z(n10190) );
  XOR U10598 ( .A(b[25]), .B(a[57]), .Z(n10229) );
  NAND U10599 ( .A(n10229), .B(n19240), .Z(n10098) );
  NAND U10600 ( .A(n10096), .B(n19242), .Z(n10097) );
  AND U10601 ( .A(n10098), .B(n10097), .Z(n10191) );
  XNOR U10602 ( .A(n10190), .B(n10191), .Z(n10192) );
  XNOR U10603 ( .A(n10193), .B(n10192), .Z(n10127) );
  XOR U10604 ( .A(n10129), .B(n10128), .Z(n10181) );
  XNOR U10605 ( .A(n10180), .B(n10181), .Z(n10232) );
  XNOR U10606 ( .A(n10233), .B(n10232), .Z(n10234) );
  XOR U10607 ( .A(n10235), .B(n10234), .Z(n10250) );
  XNOR U10608 ( .A(n10251), .B(n10250), .Z(n10252) );
  XOR U10609 ( .A(n10253), .B(n10252), .Z(n10247) );
  XOR U10610 ( .A(n10246), .B(n10247), .Z(n10123) );
  NANDN U10611 ( .A(n10104), .B(n10103), .Z(n10108) );
  NANDN U10612 ( .A(n10106), .B(n10105), .Z(n10107) );
  NAND U10613 ( .A(n10108), .B(n10107), .Z(n10121) );
  XNOR U10614 ( .A(n10120), .B(n10121), .Z(n10122) );
  XNOR U10615 ( .A(n10123), .B(n10122), .Z(n10115) );
  XNOR U10616 ( .A(n10114), .B(n10115), .Z(n10116) );
  XNOR U10617 ( .A(n10117), .B(n10116), .Z(n10254) );
  XNOR U10618 ( .A(n10254), .B(sreg[177]), .Z(n10256) );
  NAND U10619 ( .A(n10109), .B(sreg[176]), .Z(n10113) );
  OR U10620 ( .A(n10111), .B(n10110), .Z(n10112) );
  AND U10621 ( .A(n10113), .B(n10112), .Z(n10255) );
  XOR U10622 ( .A(n10256), .B(n10255), .Z(c[177]) );
  NANDN U10623 ( .A(n10115), .B(n10114), .Z(n10119) );
  NAND U10624 ( .A(n10117), .B(n10116), .Z(n10118) );
  NAND U10625 ( .A(n10119), .B(n10118), .Z(n10262) );
  NANDN U10626 ( .A(n10121), .B(n10120), .Z(n10125) );
  NAND U10627 ( .A(n10123), .B(n10122), .Z(n10124) );
  NAND U10628 ( .A(n10125), .B(n10124), .Z(n10260) );
  OR U10629 ( .A(n10127), .B(n10126), .Z(n10131) );
  NANDN U10630 ( .A(n10129), .B(n10128), .Z(n10130) );
  NAND U10631 ( .A(n10131), .B(n10130), .Z(n10380) );
  OR U10632 ( .A(n10133), .B(n10132), .Z(n10137) );
  NAND U10633 ( .A(n10135), .B(n10134), .Z(n10136) );
  NAND U10634 ( .A(n10137), .B(n10136), .Z(n10319) );
  OR U10635 ( .A(n10139), .B(n10138), .Z(n10143) );
  NANDN U10636 ( .A(n10141), .B(n10140), .Z(n10142) );
  NAND U10637 ( .A(n10143), .B(n10142), .Z(n10318) );
  OR U10638 ( .A(n10145), .B(n10144), .Z(n10149) );
  NANDN U10639 ( .A(n10147), .B(n10146), .Z(n10148) );
  NAND U10640 ( .A(n10149), .B(n10148), .Z(n10317) );
  XOR U10641 ( .A(n10319), .B(n10320), .Z(n10378) );
  OR U10642 ( .A(n10151), .B(n10150), .Z(n10155) );
  NANDN U10643 ( .A(n10153), .B(n10152), .Z(n10154) );
  NAND U10644 ( .A(n10155), .B(n10154), .Z(n10331) );
  NANDN U10645 ( .A(n10156), .B(n18832), .Z(n10158) );
  XNOR U10646 ( .A(b[19]), .B(a[64]), .Z(n10275) );
  NANDN U10647 ( .A(n10275), .B(n18834), .Z(n10157) );
  NAND U10648 ( .A(n10158), .B(n10157), .Z(n10344) );
  XNOR U10649 ( .A(b[27]), .B(a[56]), .Z(n10278) );
  NANDN U10650 ( .A(n10278), .B(n19336), .Z(n10161) );
  NANDN U10651 ( .A(n10159), .B(n19337), .Z(n10160) );
  NAND U10652 ( .A(n10161), .B(n10160), .Z(n10341) );
  XOR U10653 ( .A(b[5]), .B(a[78]), .Z(n10281) );
  NAND U10654 ( .A(n10281), .B(n17310), .Z(n10164) );
  NAND U10655 ( .A(n10162), .B(n17311), .Z(n10163) );
  AND U10656 ( .A(n10164), .B(n10163), .Z(n10342) );
  XNOR U10657 ( .A(n10341), .B(n10342), .Z(n10343) );
  XNOR U10658 ( .A(n10344), .B(n10343), .Z(n10330) );
  XOR U10659 ( .A(b[17]), .B(a[66]), .Z(n10284) );
  NAND U10660 ( .A(n10284), .B(n18673), .Z(n10167) );
  NANDN U10661 ( .A(n10165), .B(n18674), .Z(n10166) );
  NAND U10662 ( .A(n10167), .B(n10166), .Z(n10302) );
  XNOR U10663 ( .A(b[31]), .B(a[52]), .Z(n10287) );
  NANDN U10664 ( .A(n10287), .B(n19472), .Z(n10170) );
  NANDN U10665 ( .A(n10168), .B(n19473), .Z(n10169) );
  NAND U10666 ( .A(n10170), .B(n10169), .Z(n10299) );
  OR U10667 ( .A(n10171), .B(n16988), .Z(n10173) );
  XOR U10668 ( .A(b[3]), .B(n14551), .Z(n10290) );
  NANDN U10669 ( .A(n10290), .B(n16990), .Z(n10172) );
  AND U10670 ( .A(n10173), .B(n10172), .Z(n10300) );
  XNOR U10671 ( .A(n10299), .B(n10300), .Z(n10301) );
  XOR U10672 ( .A(n10302), .B(n10301), .Z(n10329) );
  XOR U10673 ( .A(n10330), .B(n10329), .Z(n10332) );
  XOR U10674 ( .A(n10331), .B(n10332), .Z(n10377) );
  XOR U10675 ( .A(n10378), .B(n10377), .Z(n10379) );
  XOR U10676 ( .A(n10380), .B(n10379), .Z(n10392) );
  NANDN U10677 ( .A(n10179), .B(n10178), .Z(n10183) );
  NANDN U10678 ( .A(n10181), .B(n10180), .Z(n10182) );
  NAND U10679 ( .A(n10183), .B(n10182), .Z(n10385) );
  OR U10680 ( .A(n10185), .B(n10184), .Z(n10189) );
  NAND U10681 ( .A(n10187), .B(n10186), .Z(n10188) );
  NAND U10682 ( .A(n10189), .B(n10188), .Z(n10384) );
  NANDN U10683 ( .A(n10191), .B(n10190), .Z(n10195) );
  NAND U10684 ( .A(n10193), .B(n10192), .Z(n10194) );
  NAND U10685 ( .A(n10195), .B(n10194), .Z(n10323) );
  NANDN U10686 ( .A(n10197), .B(n10196), .Z(n10201) );
  NAND U10687 ( .A(n10199), .B(n10198), .Z(n10200) );
  AND U10688 ( .A(n10201), .B(n10200), .Z(n10324) );
  XNOR U10689 ( .A(n10323), .B(n10324), .Z(n10325) );
  XNOR U10690 ( .A(b[9]), .B(a[74]), .Z(n10347) );
  NANDN U10691 ( .A(n10347), .B(n17814), .Z(n10204) );
  NANDN U10692 ( .A(n10202), .B(n17815), .Z(n10203) );
  NAND U10693 ( .A(n10204), .B(n10203), .Z(n10307) );
  NAND U10694 ( .A(n10205), .B(n18513), .Z(n10207) );
  XOR U10695 ( .A(b[15]), .B(a[68]), .Z(n10350) );
  NANDN U10696 ( .A(n18512), .B(n10350), .Z(n10206) );
  AND U10697 ( .A(n10207), .B(n10206), .Z(n10305) );
  NANDN U10698 ( .A(n10208), .B(n19013), .Z(n10210) );
  XNOR U10699 ( .A(b[21]), .B(a[62]), .Z(n10353) );
  NANDN U10700 ( .A(n10353), .B(n19015), .Z(n10209) );
  AND U10701 ( .A(n10210), .B(n10209), .Z(n10306) );
  XOR U10702 ( .A(n10307), .B(n10308), .Z(n10296) );
  XNOR U10703 ( .A(b[11]), .B(a[72]), .Z(n10356) );
  OR U10704 ( .A(n10356), .B(n18194), .Z(n10213) );
  NANDN U10705 ( .A(n10211), .B(n18104), .Z(n10212) );
  NAND U10706 ( .A(n10213), .B(n10212), .Z(n10294) );
  XOR U10707 ( .A(n580), .B(a[70]), .Z(n10359) );
  NANDN U10708 ( .A(n10359), .B(n18336), .Z(n10216) );
  NANDN U10709 ( .A(n10214), .B(n18337), .Z(n10215) );
  AND U10710 ( .A(n10216), .B(n10215), .Z(n10293) );
  XNOR U10711 ( .A(n10294), .B(n10293), .Z(n10295) );
  XOR U10712 ( .A(n10296), .B(n10295), .Z(n10313) );
  NANDN U10713 ( .A(n577), .B(a[82]), .Z(n10217) );
  XOR U10714 ( .A(n17151), .B(n10217), .Z(n10219) );
  NANDN U10715 ( .A(b[0]), .B(a[81]), .Z(n10218) );
  AND U10716 ( .A(n10219), .B(n10218), .Z(n10271) );
  NAND U10717 ( .A(n10220), .B(n19406), .Z(n10222) );
  XNOR U10718 ( .A(n584), .B(a[54]), .Z(n10365) );
  NANDN U10719 ( .A(n576), .B(n10365), .Z(n10221) );
  NAND U10720 ( .A(n10222), .B(n10221), .Z(n10269) );
  NANDN U10721 ( .A(n585), .B(a[50]), .Z(n10270) );
  XNOR U10722 ( .A(n10269), .B(n10270), .Z(n10272) );
  XOR U10723 ( .A(n10271), .B(n10272), .Z(n10311) );
  XOR U10724 ( .A(b[23]), .B(a[60]), .Z(n10368) );
  NANDN U10725 ( .A(n19127), .B(n10368), .Z(n10225) );
  NAND U10726 ( .A(n10223), .B(n19128), .Z(n10224) );
  NAND U10727 ( .A(n10225), .B(n10224), .Z(n10338) );
  NAND U10728 ( .A(n10226), .B(n17553), .Z(n10228) );
  XOR U10729 ( .A(b[7]), .B(a[76]), .Z(n10371) );
  NAND U10730 ( .A(n10371), .B(n17555), .Z(n10227) );
  NAND U10731 ( .A(n10228), .B(n10227), .Z(n10335) );
  XOR U10732 ( .A(b[25]), .B(a[58]), .Z(n10374) );
  NAND U10733 ( .A(n10374), .B(n19240), .Z(n10231) );
  NAND U10734 ( .A(n10229), .B(n19242), .Z(n10230) );
  AND U10735 ( .A(n10231), .B(n10230), .Z(n10336) );
  XNOR U10736 ( .A(n10335), .B(n10336), .Z(n10337) );
  XNOR U10737 ( .A(n10338), .B(n10337), .Z(n10312) );
  XOR U10738 ( .A(n10311), .B(n10312), .Z(n10314) );
  XNOR U10739 ( .A(n10313), .B(n10314), .Z(n10326) );
  XNOR U10740 ( .A(n10325), .B(n10326), .Z(n10383) );
  XNOR U10741 ( .A(n10384), .B(n10383), .Z(n10386) );
  XNOR U10742 ( .A(n10385), .B(n10386), .Z(n10390) );
  XOR U10743 ( .A(n10389), .B(n10390), .Z(n10391) );
  XOR U10744 ( .A(n10392), .B(n10391), .Z(n10398) );
  NAND U10745 ( .A(n10233), .B(n10232), .Z(n10237) );
  OR U10746 ( .A(n10235), .B(n10234), .Z(n10236) );
  NAND U10747 ( .A(n10237), .B(n10236), .Z(n10395) );
  NANDN U10748 ( .A(n10239), .B(n10238), .Z(n10243) );
  NAND U10749 ( .A(n10241), .B(n10240), .Z(n10242) );
  NAND U10750 ( .A(n10243), .B(n10242), .Z(n10396) );
  XNOR U10751 ( .A(n10395), .B(n10396), .Z(n10397) );
  XNOR U10752 ( .A(n10398), .B(n10397), .Z(n10266) );
  NANDN U10753 ( .A(n10245), .B(n10244), .Z(n10249) );
  NANDN U10754 ( .A(n10247), .B(n10246), .Z(n10248) );
  NAND U10755 ( .A(n10249), .B(n10248), .Z(n10264) );
  XNOR U10756 ( .A(n10264), .B(n10263), .Z(n10265) );
  XNOR U10757 ( .A(n10266), .B(n10265), .Z(n10259) );
  XOR U10758 ( .A(n10260), .B(n10259), .Z(n10261) );
  XNOR U10759 ( .A(n10262), .B(n10261), .Z(n10401) );
  XNOR U10760 ( .A(n10401), .B(sreg[178]), .Z(n10403) );
  NAND U10761 ( .A(n10254), .B(sreg[177]), .Z(n10258) );
  OR U10762 ( .A(n10256), .B(n10255), .Z(n10257) );
  AND U10763 ( .A(n10258), .B(n10257), .Z(n10402) );
  XOR U10764 ( .A(n10403), .B(n10402), .Z(c[178]) );
  NANDN U10765 ( .A(n10264), .B(n10263), .Z(n10268) );
  NANDN U10766 ( .A(n10266), .B(n10265), .Z(n10267) );
  NAND U10767 ( .A(n10268), .B(n10267), .Z(n10407) );
  NANDN U10768 ( .A(n10270), .B(n10269), .Z(n10274) );
  NAND U10769 ( .A(n10272), .B(n10271), .Z(n10273) );
  NAND U10770 ( .A(n10274), .B(n10273), .Z(n10493) );
  NANDN U10771 ( .A(n10275), .B(n18832), .Z(n10277) );
  XOR U10772 ( .A(b[19]), .B(n12055), .Z(n10460) );
  NANDN U10773 ( .A(n10460), .B(n18834), .Z(n10276) );
  NAND U10774 ( .A(n10277), .B(n10276), .Z(n10505) );
  XNOR U10775 ( .A(b[27]), .B(a[57]), .Z(n10463) );
  NANDN U10776 ( .A(n10463), .B(n19336), .Z(n10280) );
  NANDN U10777 ( .A(n10278), .B(n19337), .Z(n10279) );
  NAND U10778 ( .A(n10280), .B(n10279), .Z(n10502) );
  XOR U10779 ( .A(b[5]), .B(a[79]), .Z(n10466) );
  NAND U10780 ( .A(n10466), .B(n17310), .Z(n10283) );
  NAND U10781 ( .A(n10281), .B(n17311), .Z(n10282) );
  AND U10782 ( .A(n10283), .B(n10282), .Z(n10503) );
  XNOR U10783 ( .A(n10502), .B(n10503), .Z(n10504) );
  XNOR U10784 ( .A(n10505), .B(n10504), .Z(n10490) );
  XOR U10785 ( .A(b[17]), .B(a[67]), .Z(n10469) );
  NAND U10786 ( .A(n10469), .B(n18673), .Z(n10286) );
  NAND U10787 ( .A(n10284), .B(n18674), .Z(n10285) );
  NAND U10788 ( .A(n10286), .B(n10285), .Z(n10444) );
  XOR U10789 ( .A(b[31]), .B(n10660), .Z(n10472) );
  NANDN U10790 ( .A(n10472), .B(n19472), .Z(n10289) );
  NANDN U10791 ( .A(n10287), .B(n19473), .Z(n10288) );
  AND U10792 ( .A(n10289), .B(n10288), .Z(n10442) );
  OR U10793 ( .A(n10290), .B(n16988), .Z(n10292) );
  XNOR U10794 ( .A(b[3]), .B(a[81]), .Z(n10475) );
  NANDN U10795 ( .A(n10475), .B(n16990), .Z(n10291) );
  AND U10796 ( .A(n10292), .B(n10291), .Z(n10443) );
  XOR U10797 ( .A(n10444), .B(n10445), .Z(n10491) );
  XOR U10798 ( .A(n10490), .B(n10491), .Z(n10492) );
  XNOR U10799 ( .A(n10493), .B(n10492), .Z(n10538) );
  NANDN U10800 ( .A(n10294), .B(n10293), .Z(n10298) );
  NAND U10801 ( .A(n10296), .B(n10295), .Z(n10297) );
  NAND U10802 ( .A(n10298), .B(n10297), .Z(n10481) );
  NANDN U10803 ( .A(n10300), .B(n10299), .Z(n10304) );
  NAND U10804 ( .A(n10302), .B(n10301), .Z(n10303) );
  NAND U10805 ( .A(n10304), .B(n10303), .Z(n10479) );
  OR U10806 ( .A(n10306), .B(n10305), .Z(n10310) );
  NANDN U10807 ( .A(n10308), .B(n10307), .Z(n10309) );
  NAND U10808 ( .A(n10310), .B(n10309), .Z(n10478) );
  XNOR U10809 ( .A(n10481), .B(n10480), .Z(n10539) );
  XOR U10810 ( .A(n10538), .B(n10539), .Z(n10541) );
  NANDN U10811 ( .A(n10312), .B(n10311), .Z(n10316) );
  OR U10812 ( .A(n10314), .B(n10313), .Z(n10315) );
  NAND U10813 ( .A(n10316), .B(n10315), .Z(n10540) );
  XOR U10814 ( .A(n10541), .B(n10540), .Z(n10426) );
  OR U10815 ( .A(n10318), .B(n10317), .Z(n10322) );
  NANDN U10816 ( .A(n10320), .B(n10319), .Z(n10321) );
  NAND U10817 ( .A(n10322), .B(n10321), .Z(n10425) );
  NANDN U10818 ( .A(n10324), .B(n10323), .Z(n10328) );
  NANDN U10819 ( .A(n10326), .B(n10325), .Z(n10327) );
  NAND U10820 ( .A(n10328), .B(n10327), .Z(n10546) );
  NANDN U10821 ( .A(n10330), .B(n10329), .Z(n10334) );
  OR U10822 ( .A(n10332), .B(n10331), .Z(n10333) );
  NAND U10823 ( .A(n10334), .B(n10333), .Z(n10545) );
  NANDN U10824 ( .A(n10336), .B(n10335), .Z(n10340) );
  NAND U10825 ( .A(n10338), .B(n10337), .Z(n10339) );
  NAND U10826 ( .A(n10340), .B(n10339), .Z(n10484) );
  NANDN U10827 ( .A(n10342), .B(n10341), .Z(n10346) );
  NAND U10828 ( .A(n10344), .B(n10343), .Z(n10345) );
  AND U10829 ( .A(n10346), .B(n10345), .Z(n10485) );
  XNOR U10830 ( .A(n10484), .B(n10485), .Z(n10486) );
  XNOR U10831 ( .A(b[9]), .B(a[75]), .Z(n10508) );
  NANDN U10832 ( .A(n10508), .B(n17814), .Z(n10349) );
  NANDN U10833 ( .A(n10347), .B(n17815), .Z(n10348) );
  NAND U10834 ( .A(n10349), .B(n10348), .Z(n10450) );
  NAND U10835 ( .A(n10350), .B(n18513), .Z(n10352) );
  XOR U10836 ( .A(b[15]), .B(a[69]), .Z(n10511) );
  NANDN U10837 ( .A(n18512), .B(n10511), .Z(n10351) );
  AND U10838 ( .A(n10352), .B(n10351), .Z(n10448) );
  NANDN U10839 ( .A(n10353), .B(n19013), .Z(n10355) );
  XNOR U10840 ( .A(b[21]), .B(a[63]), .Z(n10514) );
  NANDN U10841 ( .A(n10514), .B(n19015), .Z(n10354) );
  AND U10842 ( .A(n10355), .B(n10354), .Z(n10449) );
  XOR U10843 ( .A(n10450), .B(n10451), .Z(n10439) );
  XNOR U10844 ( .A(b[11]), .B(a[73]), .Z(n10517) );
  OR U10845 ( .A(n10517), .B(n18194), .Z(n10358) );
  NANDN U10846 ( .A(n10356), .B(n18104), .Z(n10357) );
  NAND U10847 ( .A(n10358), .B(n10357), .Z(n10437) );
  XOR U10848 ( .A(n580), .B(a[71]), .Z(n10520) );
  NANDN U10849 ( .A(n10520), .B(n18336), .Z(n10361) );
  NANDN U10850 ( .A(n10359), .B(n18337), .Z(n10360) );
  NAND U10851 ( .A(n10361), .B(n10360), .Z(n10436) );
  XOR U10852 ( .A(n10439), .B(n10438), .Z(n10433) );
  NANDN U10853 ( .A(n577), .B(a[83]), .Z(n10362) );
  XOR U10854 ( .A(n17151), .B(n10362), .Z(n10364) );
  NANDN U10855 ( .A(b[0]), .B(a[82]), .Z(n10363) );
  AND U10856 ( .A(n10364), .B(n10363), .Z(n10456) );
  NAND U10857 ( .A(n19406), .B(n10365), .Z(n10367) );
  XOR U10858 ( .A(n584), .B(n10959), .Z(n10526) );
  NANDN U10859 ( .A(n576), .B(n10526), .Z(n10366) );
  NAND U10860 ( .A(n10367), .B(n10366), .Z(n10454) );
  NANDN U10861 ( .A(n585), .B(a[51]), .Z(n10455) );
  XNOR U10862 ( .A(n10454), .B(n10455), .Z(n10457) );
  XNOR U10863 ( .A(n10456), .B(n10457), .Z(n10431) );
  XOR U10864 ( .A(b[23]), .B(a[61]), .Z(n10529) );
  NANDN U10865 ( .A(n19127), .B(n10529), .Z(n10370) );
  NAND U10866 ( .A(n10368), .B(n19128), .Z(n10369) );
  NAND U10867 ( .A(n10370), .B(n10369), .Z(n10499) );
  NAND U10868 ( .A(n10371), .B(n17553), .Z(n10373) );
  XOR U10869 ( .A(b[7]), .B(a[77]), .Z(n10532) );
  NAND U10870 ( .A(n10532), .B(n17555), .Z(n10372) );
  NAND U10871 ( .A(n10373), .B(n10372), .Z(n10496) );
  XOR U10872 ( .A(b[25]), .B(a[59]), .Z(n10535) );
  NAND U10873 ( .A(n10535), .B(n19240), .Z(n10376) );
  NAND U10874 ( .A(n10374), .B(n19242), .Z(n10375) );
  AND U10875 ( .A(n10376), .B(n10375), .Z(n10497) );
  XNOR U10876 ( .A(n10496), .B(n10497), .Z(n10498) );
  XOR U10877 ( .A(n10499), .B(n10498), .Z(n10430) );
  XOR U10878 ( .A(n10433), .B(n10432), .Z(n10487) );
  XNOR U10879 ( .A(n10486), .B(n10487), .Z(n10544) );
  XNOR U10880 ( .A(n10545), .B(n10544), .Z(n10547) );
  XNOR U10881 ( .A(n10546), .B(n10547), .Z(n10424) );
  XOR U10882 ( .A(n10425), .B(n10424), .Z(n10427) );
  NAND U10883 ( .A(n10378), .B(n10377), .Z(n10382) );
  NAND U10884 ( .A(n10380), .B(n10379), .Z(n10381) );
  NAND U10885 ( .A(n10382), .B(n10381), .Z(n10419) );
  NAND U10886 ( .A(n10384), .B(n10383), .Z(n10388) );
  NANDN U10887 ( .A(n10386), .B(n10385), .Z(n10387) );
  AND U10888 ( .A(n10388), .B(n10387), .Z(n10418) );
  XNOR U10889 ( .A(n10419), .B(n10418), .Z(n10420) );
  XOR U10890 ( .A(n10421), .B(n10420), .Z(n10414) );
  NANDN U10891 ( .A(n10390), .B(n10389), .Z(n10394) );
  OR U10892 ( .A(n10392), .B(n10391), .Z(n10393) );
  NAND U10893 ( .A(n10394), .B(n10393), .Z(n10412) );
  NANDN U10894 ( .A(n10396), .B(n10395), .Z(n10400) );
  NANDN U10895 ( .A(n10398), .B(n10397), .Z(n10399) );
  NAND U10896 ( .A(n10400), .B(n10399), .Z(n10413) );
  XNOR U10897 ( .A(n10412), .B(n10413), .Z(n10415) );
  XOR U10898 ( .A(n10414), .B(n10415), .Z(n10406) );
  XOR U10899 ( .A(n10407), .B(n10406), .Z(n10408) );
  XNOR U10900 ( .A(n10409), .B(n10408), .Z(n10550) );
  XNOR U10901 ( .A(n10550), .B(sreg[179]), .Z(n10552) );
  NAND U10902 ( .A(n10401), .B(sreg[178]), .Z(n10405) );
  OR U10903 ( .A(n10403), .B(n10402), .Z(n10404) );
  AND U10904 ( .A(n10405), .B(n10404), .Z(n10551) );
  XOR U10905 ( .A(n10552), .B(n10551), .Z(c[179]) );
  NAND U10906 ( .A(n10407), .B(n10406), .Z(n10411) );
  NAND U10907 ( .A(n10409), .B(n10408), .Z(n10410) );
  NAND U10908 ( .A(n10411), .B(n10410), .Z(n10558) );
  NANDN U10909 ( .A(n10413), .B(n10412), .Z(n10417) );
  NAND U10910 ( .A(n10415), .B(n10414), .Z(n10416) );
  NAND U10911 ( .A(n10417), .B(n10416), .Z(n10556) );
  NANDN U10912 ( .A(n10419), .B(n10418), .Z(n10423) );
  NAND U10913 ( .A(n10421), .B(n10420), .Z(n10422) );
  NAND U10914 ( .A(n10423), .B(n10422), .Z(n10561) );
  NANDN U10915 ( .A(n10425), .B(n10424), .Z(n10429) );
  OR U10916 ( .A(n10427), .B(n10426), .Z(n10428) );
  NAND U10917 ( .A(n10429), .B(n10428), .Z(n10562) );
  XNOR U10918 ( .A(n10561), .B(n10562), .Z(n10563) );
  NANDN U10919 ( .A(n10431), .B(n10430), .Z(n10435) );
  NANDN U10920 ( .A(n10433), .B(n10432), .Z(n10434) );
  NAND U10921 ( .A(n10435), .B(n10434), .Z(n10679) );
  OR U10922 ( .A(n10437), .B(n10436), .Z(n10441) );
  NAND U10923 ( .A(n10439), .B(n10438), .Z(n10440) );
  NAND U10924 ( .A(n10441), .B(n10440), .Z(n10617) );
  OR U10925 ( .A(n10443), .B(n10442), .Z(n10447) );
  NANDN U10926 ( .A(n10445), .B(n10444), .Z(n10446) );
  NAND U10927 ( .A(n10447), .B(n10446), .Z(n10616) );
  OR U10928 ( .A(n10449), .B(n10448), .Z(n10453) );
  NANDN U10929 ( .A(n10451), .B(n10450), .Z(n10452) );
  NAND U10930 ( .A(n10453), .B(n10452), .Z(n10615) );
  XOR U10931 ( .A(n10617), .B(n10618), .Z(n10676) );
  NANDN U10932 ( .A(n10455), .B(n10454), .Z(n10459) );
  NAND U10933 ( .A(n10457), .B(n10456), .Z(n10458) );
  NAND U10934 ( .A(n10459), .B(n10458), .Z(n10630) );
  NANDN U10935 ( .A(n10460), .B(n18832), .Z(n10462) );
  XNOR U10936 ( .A(b[19]), .B(a[66]), .Z(n10573) );
  NANDN U10937 ( .A(n10573), .B(n18834), .Z(n10461) );
  NAND U10938 ( .A(n10462), .B(n10461), .Z(n10642) );
  XNOR U10939 ( .A(b[27]), .B(a[58]), .Z(n10576) );
  NANDN U10940 ( .A(n10576), .B(n19336), .Z(n10465) );
  NANDN U10941 ( .A(n10463), .B(n19337), .Z(n10464) );
  NAND U10942 ( .A(n10465), .B(n10464), .Z(n10639) );
  XNOR U10943 ( .A(b[5]), .B(a[80]), .Z(n10579) );
  NANDN U10944 ( .A(n10579), .B(n17310), .Z(n10468) );
  NAND U10945 ( .A(n10466), .B(n17311), .Z(n10467) );
  AND U10946 ( .A(n10468), .B(n10467), .Z(n10640) );
  XNOR U10947 ( .A(n10639), .B(n10640), .Z(n10641) );
  XNOR U10948 ( .A(n10642), .B(n10641), .Z(n10628) );
  XOR U10949 ( .A(b[17]), .B(a[68]), .Z(n10582) );
  NAND U10950 ( .A(n10582), .B(n18673), .Z(n10471) );
  NAND U10951 ( .A(n10469), .B(n18674), .Z(n10470) );
  NAND U10952 ( .A(n10471), .B(n10470), .Z(n10600) );
  XNOR U10953 ( .A(b[31]), .B(a[54]), .Z(n10585) );
  NANDN U10954 ( .A(n10585), .B(n19472), .Z(n10474) );
  NANDN U10955 ( .A(n10472), .B(n19473), .Z(n10473) );
  NAND U10956 ( .A(n10474), .B(n10473), .Z(n10597) );
  OR U10957 ( .A(n10475), .B(n16988), .Z(n10477) );
  XNOR U10958 ( .A(b[3]), .B(a[82]), .Z(n10588) );
  NANDN U10959 ( .A(n10588), .B(n16990), .Z(n10476) );
  AND U10960 ( .A(n10477), .B(n10476), .Z(n10598) );
  XNOR U10961 ( .A(n10597), .B(n10598), .Z(n10599) );
  XOR U10962 ( .A(n10600), .B(n10599), .Z(n10627) );
  XNOR U10963 ( .A(n10628), .B(n10627), .Z(n10629) );
  XNOR U10964 ( .A(n10630), .B(n10629), .Z(n10677) );
  XNOR U10965 ( .A(n10676), .B(n10677), .Z(n10678) );
  XNOR U10966 ( .A(n10679), .B(n10678), .Z(n10697) );
  OR U10967 ( .A(n10479), .B(n10478), .Z(n10483) );
  NAND U10968 ( .A(n10481), .B(n10480), .Z(n10482) );
  NAND U10969 ( .A(n10483), .B(n10482), .Z(n10695) );
  NANDN U10970 ( .A(n10485), .B(n10484), .Z(n10489) );
  NANDN U10971 ( .A(n10487), .B(n10486), .Z(n10488) );
  NAND U10972 ( .A(n10489), .B(n10488), .Z(n10684) );
  OR U10973 ( .A(n10491), .B(n10490), .Z(n10495) );
  NAND U10974 ( .A(n10493), .B(n10492), .Z(n10494) );
  NAND U10975 ( .A(n10495), .B(n10494), .Z(n10683) );
  NANDN U10976 ( .A(n10497), .B(n10496), .Z(n10501) );
  NAND U10977 ( .A(n10499), .B(n10498), .Z(n10500) );
  NAND U10978 ( .A(n10501), .B(n10500), .Z(n10621) );
  NANDN U10979 ( .A(n10503), .B(n10502), .Z(n10507) );
  NAND U10980 ( .A(n10505), .B(n10504), .Z(n10506) );
  AND U10981 ( .A(n10507), .B(n10506), .Z(n10622) );
  XNOR U10982 ( .A(n10621), .B(n10622), .Z(n10623) );
  XNOR U10983 ( .A(b[9]), .B(a[76]), .Z(n10645) );
  NANDN U10984 ( .A(n10645), .B(n17814), .Z(n10510) );
  NANDN U10985 ( .A(n10508), .B(n17815), .Z(n10509) );
  NAND U10986 ( .A(n10510), .B(n10509), .Z(n10605) );
  NAND U10987 ( .A(n10511), .B(n18513), .Z(n10513) );
  XOR U10988 ( .A(b[15]), .B(a[70]), .Z(n10648) );
  NANDN U10989 ( .A(n18512), .B(n10648), .Z(n10512) );
  AND U10990 ( .A(n10513), .B(n10512), .Z(n10603) );
  NANDN U10991 ( .A(n10514), .B(n19013), .Z(n10516) );
  XNOR U10992 ( .A(b[21]), .B(a[64]), .Z(n10651) );
  NANDN U10993 ( .A(n10651), .B(n19015), .Z(n10515) );
  AND U10994 ( .A(n10516), .B(n10515), .Z(n10604) );
  XOR U10995 ( .A(n10605), .B(n10606), .Z(n10594) );
  XNOR U10996 ( .A(b[11]), .B(a[74]), .Z(n10654) );
  OR U10997 ( .A(n10654), .B(n18194), .Z(n10519) );
  NANDN U10998 ( .A(n10517), .B(n18104), .Z(n10518) );
  NAND U10999 ( .A(n10519), .B(n10518), .Z(n10592) );
  XOR U11000 ( .A(n580), .B(a[72]), .Z(n10657) );
  NANDN U11001 ( .A(n10657), .B(n18336), .Z(n10522) );
  NANDN U11002 ( .A(n10520), .B(n18337), .Z(n10521) );
  AND U11003 ( .A(n10522), .B(n10521), .Z(n10591) );
  XNOR U11004 ( .A(n10592), .B(n10591), .Z(n10593) );
  XOR U11005 ( .A(n10594), .B(n10593), .Z(n10611) );
  NANDN U11006 ( .A(n577), .B(a[84]), .Z(n10523) );
  XOR U11007 ( .A(n17151), .B(n10523), .Z(n10525) );
  NANDN U11008 ( .A(b[0]), .B(a[83]), .Z(n10524) );
  AND U11009 ( .A(n10525), .B(n10524), .Z(n10569) );
  NAND U11010 ( .A(n19406), .B(n10526), .Z(n10528) );
  XNOR U11011 ( .A(b[29]), .B(a[56]), .Z(n10661) );
  OR U11012 ( .A(n10661), .B(n576), .Z(n10527) );
  NAND U11013 ( .A(n10528), .B(n10527), .Z(n10567) );
  NANDN U11014 ( .A(n585), .B(a[52]), .Z(n10568) );
  XNOR U11015 ( .A(n10567), .B(n10568), .Z(n10570) );
  XOR U11016 ( .A(n10569), .B(n10570), .Z(n10609) );
  XOR U11017 ( .A(b[23]), .B(a[62]), .Z(n10667) );
  NANDN U11018 ( .A(n19127), .B(n10667), .Z(n10531) );
  NAND U11019 ( .A(n10529), .B(n19128), .Z(n10530) );
  NAND U11020 ( .A(n10531), .B(n10530), .Z(n10636) );
  NAND U11021 ( .A(n10532), .B(n17553), .Z(n10534) );
  XOR U11022 ( .A(b[7]), .B(a[78]), .Z(n10670) );
  NAND U11023 ( .A(n10670), .B(n17555), .Z(n10533) );
  NAND U11024 ( .A(n10534), .B(n10533), .Z(n10633) );
  XOR U11025 ( .A(b[25]), .B(a[60]), .Z(n10673) );
  NAND U11026 ( .A(n10673), .B(n19240), .Z(n10537) );
  NAND U11027 ( .A(n10535), .B(n19242), .Z(n10536) );
  AND U11028 ( .A(n10537), .B(n10536), .Z(n10634) );
  XNOR U11029 ( .A(n10633), .B(n10634), .Z(n10635) );
  XNOR U11030 ( .A(n10636), .B(n10635), .Z(n10610) );
  XOR U11031 ( .A(n10609), .B(n10610), .Z(n10612) );
  XNOR U11032 ( .A(n10611), .B(n10612), .Z(n10624) );
  XNOR U11033 ( .A(n10623), .B(n10624), .Z(n10682) );
  XNOR U11034 ( .A(n10683), .B(n10682), .Z(n10685) );
  XNOR U11035 ( .A(n10684), .B(n10685), .Z(n10694) );
  XNOR U11036 ( .A(n10695), .B(n10694), .Z(n10696) );
  XOR U11037 ( .A(n10697), .B(n10696), .Z(n10691) );
  NANDN U11038 ( .A(n10539), .B(n10538), .Z(n10543) );
  OR U11039 ( .A(n10541), .B(n10540), .Z(n10542) );
  NAND U11040 ( .A(n10543), .B(n10542), .Z(n10688) );
  NAND U11041 ( .A(n10545), .B(n10544), .Z(n10549) );
  NANDN U11042 ( .A(n10547), .B(n10546), .Z(n10548) );
  NAND U11043 ( .A(n10549), .B(n10548), .Z(n10689) );
  XNOR U11044 ( .A(n10688), .B(n10689), .Z(n10690) );
  XOR U11045 ( .A(n10691), .B(n10690), .Z(n10564) );
  XOR U11046 ( .A(n10563), .B(n10564), .Z(n10555) );
  XOR U11047 ( .A(n10556), .B(n10555), .Z(n10557) );
  XNOR U11048 ( .A(n10558), .B(n10557), .Z(n10700) );
  XNOR U11049 ( .A(n10700), .B(sreg[180]), .Z(n10702) );
  NAND U11050 ( .A(n10550), .B(sreg[179]), .Z(n10554) );
  OR U11051 ( .A(n10552), .B(n10551), .Z(n10553) );
  AND U11052 ( .A(n10554), .B(n10553), .Z(n10701) );
  XOR U11053 ( .A(n10702), .B(n10701), .Z(c[180]) );
  NAND U11054 ( .A(n10556), .B(n10555), .Z(n10560) );
  NAND U11055 ( .A(n10558), .B(n10557), .Z(n10559) );
  NAND U11056 ( .A(n10560), .B(n10559), .Z(n10708) );
  NANDN U11057 ( .A(n10562), .B(n10561), .Z(n10566) );
  NAND U11058 ( .A(n10564), .B(n10563), .Z(n10565) );
  NAND U11059 ( .A(n10566), .B(n10565), .Z(n10706) );
  NANDN U11060 ( .A(n10568), .B(n10567), .Z(n10572) );
  NAND U11061 ( .A(n10570), .B(n10569), .Z(n10571) );
  NAND U11062 ( .A(n10572), .B(n10571), .Z(n10792) );
  NANDN U11063 ( .A(n10573), .B(n18832), .Z(n10575) );
  XNOR U11064 ( .A(b[19]), .B(a[67]), .Z(n10759) );
  NANDN U11065 ( .A(n10759), .B(n18834), .Z(n10574) );
  NAND U11066 ( .A(n10575), .B(n10574), .Z(n10804) );
  XNOR U11067 ( .A(b[27]), .B(a[59]), .Z(n10762) );
  NANDN U11068 ( .A(n10762), .B(n19336), .Z(n10578) );
  NANDN U11069 ( .A(n10576), .B(n19337), .Z(n10577) );
  NAND U11070 ( .A(n10578), .B(n10577), .Z(n10801) );
  XOR U11071 ( .A(b[5]), .B(a[81]), .Z(n10765) );
  NAND U11072 ( .A(n10765), .B(n17310), .Z(n10581) );
  NANDN U11073 ( .A(n10579), .B(n17311), .Z(n10580) );
  AND U11074 ( .A(n10581), .B(n10580), .Z(n10802) );
  XNOR U11075 ( .A(n10801), .B(n10802), .Z(n10803) );
  XNOR U11076 ( .A(n10804), .B(n10803), .Z(n10789) );
  XOR U11077 ( .A(b[17]), .B(a[69]), .Z(n10768) );
  NAND U11078 ( .A(n10768), .B(n18673), .Z(n10584) );
  NAND U11079 ( .A(n10582), .B(n18674), .Z(n10583) );
  NAND U11080 ( .A(n10584), .B(n10583), .Z(n10743) );
  XOR U11081 ( .A(b[31]), .B(n10959), .Z(n10771) );
  NANDN U11082 ( .A(n10771), .B(n19472), .Z(n10587) );
  NANDN U11083 ( .A(n10585), .B(n19473), .Z(n10586) );
  AND U11084 ( .A(n10587), .B(n10586), .Z(n10741) );
  OR U11085 ( .A(n10588), .B(n16988), .Z(n10590) );
  XNOR U11086 ( .A(b[3]), .B(a[83]), .Z(n10774) );
  NANDN U11087 ( .A(n10774), .B(n16990), .Z(n10589) );
  AND U11088 ( .A(n10590), .B(n10589), .Z(n10742) );
  XOR U11089 ( .A(n10743), .B(n10744), .Z(n10790) );
  XOR U11090 ( .A(n10789), .B(n10790), .Z(n10791) );
  XNOR U11091 ( .A(n10792), .B(n10791), .Z(n10837) );
  NANDN U11092 ( .A(n10592), .B(n10591), .Z(n10596) );
  NAND U11093 ( .A(n10594), .B(n10593), .Z(n10595) );
  NAND U11094 ( .A(n10596), .B(n10595), .Z(n10780) );
  NANDN U11095 ( .A(n10598), .B(n10597), .Z(n10602) );
  NAND U11096 ( .A(n10600), .B(n10599), .Z(n10601) );
  NAND U11097 ( .A(n10602), .B(n10601), .Z(n10778) );
  OR U11098 ( .A(n10604), .B(n10603), .Z(n10608) );
  NANDN U11099 ( .A(n10606), .B(n10605), .Z(n10607) );
  NAND U11100 ( .A(n10608), .B(n10607), .Z(n10777) );
  XNOR U11101 ( .A(n10780), .B(n10779), .Z(n10838) );
  XOR U11102 ( .A(n10837), .B(n10838), .Z(n10840) );
  NANDN U11103 ( .A(n10610), .B(n10609), .Z(n10614) );
  OR U11104 ( .A(n10612), .B(n10611), .Z(n10613) );
  NAND U11105 ( .A(n10614), .B(n10613), .Z(n10839) );
  XOR U11106 ( .A(n10840), .B(n10839), .Z(n10725) );
  OR U11107 ( .A(n10616), .B(n10615), .Z(n10620) );
  NANDN U11108 ( .A(n10618), .B(n10617), .Z(n10619) );
  NAND U11109 ( .A(n10620), .B(n10619), .Z(n10724) );
  NANDN U11110 ( .A(n10622), .B(n10621), .Z(n10626) );
  NANDN U11111 ( .A(n10624), .B(n10623), .Z(n10625) );
  NAND U11112 ( .A(n10626), .B(n10625), .Z(n10845) );
  NANDN U11113 ( .A(n10628), .B(n10627), .Z(n10632) );
  NAND U11114 ( .A(n10630), .B(n10629), .Z(n10631) );
  NAND U11115 ( .A(n10632), .B(n10631), .Z(n10844) );
  NANDN U11116 ( .A(n10634), .B(n10633), .Z(n10638) );
  NAND U11117 ( .A(n10636), .B(n10635), .Z(n10637) );
  NAND U11118 ( .A(n10638), .B(n10637), .Z(n10783) );
  NANDN U11119 ( .A(n10640), .B(n10639), .Z(n10644) );
  NAND U11120 ( .A(n10642), .B(n10641), .Z(n10643) );
  AND U11121 ( .A(n10644), .B(n10643), .Z(n10784) );
  XNOR U11122 ( .A(n10783), .B(n10784), .Z(n10785) );
  XNOR U11123 ( .A(b[9]), .B(a[77]), .Z(n10807) );
  NANDN U11124 ( .A(n10807), .B(n17814), .Z(n10647) );
  NANDN U11125 ( .A(n10645), .B(n17815), .Z(n10646) );
  NAND U11126 ( .A(n10647), .B(n10646), .Z(n10749) );
  NAND U11127 ( .A(n10648), .B(n18513), .Z(n10650) );
  XOR U11128 ( .A(b[15]), .B(a[71]), .Z(n10810) );
  NANDN U11129 ( .A(n18512), .B(n10810), .Z(n10649) );
  AND U11130 ( .A(n10650), .B(n10649), .Z(n10747) );
  NANDN U11131 ( .A(n10651), .B(n19013), .Z(n10653) );
  XOR U11132 ( .A(b[21]), .B(n12055), .Z(n10813) );
  NANDN U11133 ( .A(n10813), .B(n19015), .Z(n10652) );
  AND U11134 ( .A(n10653), .B(n10652), .Z(n10748) );
  XOR U11135 ( .A(n10749), .B(n10750), .Z(n10738) );
  XNOR U11136 ( .A(b[11]), .B(a[75]), .Z(n10816) );
  OR U11137 ( .A(n10816), .B(n18194), .Z(n10656) );
  NANDN U11138 ( .A(n10654), .B(n18104), .Z(n10655) );
  NAND U11139 ( .A(n10656), .B(n10655), .Z(n10736) );
  XOR U11140 ( .A(n580), .B(a[73]), .Z(n10819) );
  NANDN U11141 ( .A(n10819), .B(n18336), .Z(n10659) );
  NANDN U11142 ( .A(n10657), .B(n18337), .Z(n10658) );
  NAND U11143 ( .A(n10659), .B(n10658), .Z(n10735) );
  XOR U11144 ( .A(n10738), .B(n10737), .Z(n10732) );
  ANDN U11145 ( .B(b[31]), .A(n10660), .Z(n10753) );
  NANDN U11146 ( .A(n10661), .B(n19406), .Z(n10663) );
  XNOR U11147 ( .A(n584), .B(a[57]), .Z(n10825) );
  NANDN U11148 ( .A(n576), .B(n10825), .Z(n10662) );
  NAND U11149 ( .A(n10663), .B(n10662), .Z(n10754) );
  XOR U11150 ( .A(n10753), .B(n10754), .Z(n10755) );
  NANDN U11151 ( .A(n577), .B(a[85]), .Z(n10664) );
  XOR U11152 ( .A(n17151), .B(n10664), .Z(n10666) );
  IV U11153 ( .A(a[84]), .Z(n15134) );
  NANDN U11154 ( .A(n15134), .B(n577), .Z(n10665) );
  AND U11155 ( .A(n10666), .B(n10665), .Z(n10756) );
  XNOR U11156 ( .A(n10755), .B(n10756), .Z(n10729) );
  XOR U11157 ( .A(b[23]), .B(a[63]), .Z(n10828) );
  NANDN U11158 ( .A(n19127), .B(n10828), .Z(n10669) );
  NAND U11159 ( .A(n10667), .B(n19128), .Z(n10668) );
  NAND U11160 ( .A(n10669), .B(n10668), .Z(n10798) );
  NAND U11161 ( .A(n10670), .B(n17553), .Z(n10672) );
  XOR U11162 ( .A(b[7]), .B(a[79]), .Z(n10831) );
  NAND U11163 ( .A(n10831), .B(n17555), .Z(n10671) );
  NAND U11164 ( .A(n10672), .B(n10671), .Z(n10795) );
  XOR U11165 ( .A(b[25]), .B(a[61]), .Z(n10834) );
  NAND U11166 ( .A(n10834), .B(n19240), .Z(n10675) );
  NAND U11167 ( .A(n10673), .B(n19242), .Z(n10674) );
  AND U11168 ( .A(n10675), .B(n10674), .Z(n10796) );
  XNOR U11169 ( .A(n10795), .B(n10796), .Z(n10797) );
  XNOR U11170 ( .A(n10798), .B(n10797), .Z(n10730) );
  XOR U11171 ( .A(n10732), .B(n10731), .Z(n10786) );
  XNOR U11172 ( .A(n10785), .B(n10786), .Z(n10843) );
  XNOR U11173 ( .A(n10844), .B(n10843), .Z(n10846) );
  XNOR U11174 ( .A(n10845), .B(n10846), .Z(n10723) );
  XOR U11175 ( .A(n10724), .B(n10723), .Z(n10726) );
  NANDN U11176 ( .A(n10677), .B(n10676), .Z(n10681) );
  NAND U11177 ( .A(n10679), .B(n10678), .Z(n10680) );
  NAND U11178 ( .A(n10681), .B(n10680), .Z(n10718) );
  NAND U11179 ( .A(n10683), .B(n10682), .Z(n10687) );
  NANDN U11180 ( .A(n10685), .B(n10684), .Z(n10686) );
  AND U11181 ( .A(n10687), .B(n10686), .Z(n10717) );
  XNOR U11182 ( .A(n10718), .B(n10717), .Z(n10719) );
  XOR U11183 ( .A(n10720), .B(n10719), .Z(n10713) );
  NANDN U11184 ( .A(n10689), .B(n10688), .Z(n10693) );
  NAND U11185 ( .A(n10691), .B(n10690), .Z(n10692) );
  NAND U11186 ( .A(n10693), .B(n10692), .Z(n10711) );
  NANDN U11187 ( .A(n10695), .B(n10694), .Z(n10699) );
  NANDN U11188 ( .A(n10697), .B(n10696), .Z(n10698) );
  NAND U11189 ( .A(n10699), .B(n10698), .Z(n10712) );
  XNOR U11190 ( .A(n10711), .B(n10712), .Z(n10714) );
  XOR U11191 ( .A(n10713), .B(n10714), .Z(n10705) );
  XOR U11192 ( .A(n10706), .B(n10705), .Z(n10707) );
  XNOR U11193 ( .A(n10708), .B(n10707), .Z(n10849) );
  XNOR U11194 ( .A(n10849), .B(sreg[181]), .Z(n10851) );
  NAND U11195 ( .A(n10700), .B(sreg[180]), .Z(n10704) );
  OR U11196 ( .A(n10702), .B(n10701), .Z(n10703) );
  AND U11197 ( .A(n10704), .B(n10703), .Z(n10850) );
  XOR U11198 ( .A(n10851), .B(n10850), .Z(c[181]) );
  NAND U11199 ( .A(n10706), .B(n10705), .Z(n10710) );
  NAND U11200 ( .A(n10708), .B(n10707), .Z(n10709) );
  NAND U11201 ( .A(n10710), .B(n10709), .Z(n10857) );
  NANDN U11202 ( .A(n10712), .B(n10711), .Z(n10716) );
  NAND U11203 ( .A(n10714), .B(n10713), .Z(n10715) );
  NAND U11204 ( .A(n10716), .B(n10715), .Z(n10855) );
  NANDN U11205 ( .A(n10718), .B(n10717), .Z(n10722) );
  NAND U11206 ( .A(n10720), .B(n10719), .Z(n10721) );
  NAND U11207 ( .A(n10722), .B(n10721), .Z(n10860) );
  NANDN U11208 ( .A(n10724), .B(n10723), .Z(n10728) );
  OR U11209 ( .A(n10726), .B(n10725), .Z(n10727) );
  NAND U11210 ( .A(n10728), .B(n10727), .Z(n10861) );
  XNOR U11211 ( .A(n10860), .B(n10861), .Z(n10862) );
  OR U11212 ( .A(n10730), .B(n10729), .Z(n10734) );
  NANDN U11213 ( .A(n10732), .B(n10731), .Z(n10733) );
  NAND U11214 ( .A(n10734), .B(n10733), .Z(n10978) );
  OR U11215 ( .A(n10736), .B(n10735), .Z(n10740) );
  NAND U11216 ( .A(n10738), .B(n10737), .Z(n10739) );
  NAND U11217 ( .A(n10740), .B(n10739), .Z(n10916) );
  OR U11218 ( .A(n10742), .B(n10741), .Z(n10746) );
  NANDN U11219 ( .A(n10744), .B(n10743), .Z(n10745) );
  NAND U11220 ( .A(n10746), .B(n10745), .Z(n10915) );
  OR U11221 ( .A(n10748), .B(n10747), .Z(n10752) );
  NANDN U11222 ( .A(n10750), .B(n10749), .Z(n10751) );
  NAND U11223 ( .A(n10752), .B(n10751), .Z(n10914) );
  XOR U11224 ( .A(n10916), .B(n10917), .Z(n10976) );
  OR U11225 ( .A(n10754), .B(n10753), .Z(n10758) );
  NANDN U11226 ( .A(n10756), .B(n10755), .Z(n10757) );
  NAND U11227 ( .A(n10758), .B(n10757), .Z(n10929) );
  NANDN U11228 ( .A(n10759), .B(n18832), .Z(n10761) );
  XNOR U11229 ( .A(b[19]), .B(a[68]), .Z(n10896) );
  NANDN U11230 ( .A(n10896), .B(n18834), .Z(n10760) );
  NAND U11231 ( .A(n10761), .B(n10760), .Z(n10941) );
  XNOR U11232 ( .A(b[27]), .B(a[60]), .Z(n10899) );
  NANDN U11233 ( .A(n10899), .B(n19336), .Z(n10764) );
  NANDN U11234 ( .A(n10762), .B(n19337), .Z(n10763) );
  NAND U11235 ( .A(n10764), .B(n10763), .Z(n10938) );
  XOR U11236 ( .A(b[5]), .B(a[82]), .Z(n10902) );
  NAND U11237 ( .A(n10902), .B(n17310), .Z(n10767) );
  NAND U11238 ( .A(n10765), .B(n17311), .Z(n10766) );
  AND U11239 ( .A(n10767), .B(n10766), .Z(n10939) );
  XNOR U11240 ( .A(n10938), .B(n10939), .Z(n10940) );
  XNOR U11241 ( .A(n10941), .B(n10940), .Z(n10926) );
  XOR U11242 ( .A(b[17]), .B(a[70]), .Z(n10905) );
  NAND U11243 ( .A(n10905), .B(n18673), .Z(n10770) );
  NAND U11244 ( .A(n10768), .B(n18674), .Z(n10769) );
  NAND U11245 ( .A(n10770), .B(n10769), .Z(n10880) );
  XNOR U11246 ( .A(b[31]), .B(a[56]), .Z(n10908) );
  NANDN U11247 ( .A(n10908), .B(n19472), .Z(n10773) );
  NANDN U11248 ( .A(n10771), .B(n19473), .Z(n10772) );
  AND U11249 ( .A(n10773), .B(n10772), .Z(n10878) );
  OR U11250 ( .A(n10774), .B(n16988), .Z(n10776) );
  XOR U11251 ( .A(b[3]), .B(n15134), .Z(n10911) );
  NANDN U11252 ( .A(n10911), .B(n16990), .Z(n10775) );
  AND U11253 ( .A(n10776), .B(n10775), .Z(n10879) );
  XOR U11254 ( .A(n10880), .B(n10881), .Z(n10927) );
  XOR U11255 ( .A(n10926), .B(n10927), .Z(n10928) );
  XNOR U11256 ( .A(n10929), .B(n10928), .Z(n10975) );
  XOR U11257 ( .A(n10976), .B(n10975), .Z(n10977) );
  XNOR U11258 ( .A(n10978), .B(n10977), .Z(n10994) );
  OR U11259 ( .A(n10778), .B(n10777), .Z(n10782) );
  NAND U11260 ( .A(n10780), .B(n10779), .Z(n10781) );
  NAND U11261 ( .A(n10782), .B(n10781), .Z(n10992) );
  NANDN U11262 ( .A(n10784), .B(n10783), .Z(n10788) );
  NANDN U11263 ( .A(n10786), .B(n10785), .Z(n10787) );
  NAND U11264 ( .A(n10788), .B(n10787), .Z(n10981) );
  OR U11265 ( .A(n10790), .B(n10789), .Z(n10794) );
  NAND U11266 ( .A(n10792), .B(n10791), .Z(n10793) );
  NAND U11267 ( .A(n10794), .B(n10793), .Z(n10980) );
  NANDN U11268 ( .A(n10796), .B(n10795), .Z(n10800) );
  NAND U11269 ( .A(n10798), .B(n10797), .Z(n10799) );
  NAND U11270 ( .A(n10800), .B(n10799), .Z(n10920) );
  NANDN U11271 ( .A(n10802), .B(n10801), .Z(n10806) );
  NAND U11272 ( .A(n10804), .B(n10803), .Z(n10805) );
  AND U11273 ( .A(n10806), .B(n10805), .Z(n10921) );
  XNOR U11274 ( .A(n10920), .B(n10921), .Z(n10922) );
  XNOR U11275 ( .A(b[9]), .B(a[78]), .Z(n10944) );
  NANDN U11276 ( .A(n10944), .B(n17814), .Z(n10809) );
  NANDN U11277 ( .A(n10807), .B(n17815), .Z(n10808) );
  NAND U11278 ( .A(n10809), .B(n10808), .Z(n10886) );
  NAND U11279 ( .A(n10810), .B(n18513), .Z(n10812) );
  XOR U11280 ( .A(b[15]), .B(a[72]), .Z(n10947) );
  NANDN U11281 ( .A(n18512), .B(n10947), .Z(n10811) );
  AND U11282 ( .A(n10812), .B(n10811), .Z(n10884) );
  NANDN U11283 ( .A(n10813), .B(n19013), .Z(n10815) );
  XNOR U11284 ( .A(b[21]), .B(a[66]), .Z(n10950) );
  NANDN U11285 ( .A(n10950), .B(n19015), .Z(n10814) );
  AND U11286 ( .A(n10815), .B(n10814), .Z(n10885) );
  XOR U11287 ( .A(n10886), .B(n10887), .Z(n10875) );
  XNOR U11288 ( .A(b[11]), .B(a[76]), .Z(n10953) );
  OR U11289 ( .A(n10953), .B(n18194), .Z(n10818) );
  NANDN U11290 ( .A(n10816), .B(n18104), .Z(n10817) );
  NAND U11291 ( .A(n10818), .B(n10817), .Z(n10873) );
  XOR U11292 ( .A(n580), .B(a[74]), .Z(n10956) );
  NANDN U11293 ( .A(n10956), .B(n18336), .Z(n10821) );
  NANDN U11294 ( .A(n10819), .B(n18337), .Z(n10820) );
  NAND U11295 ( .A(n10821), .B(n10820), .Z(n10872) );
  XOR U11296 ( .A(n10875), .B(n10874), .Z(n10869) );
  NANDN U11297 ( .A(n577), .B(a[86]), .Z(n10822) );
  XOR U11298 ( .A(n17151), .B(n10822), .Z(n10824) );
  NANDN U11299 ( .A(b[0]), .B(a[85]), .Z(n10823) );
  AND U11300 ( .A(n10824), .B(n10823), .Z(n10892) );
  NAND U11301 ( .A(n10825), .B(n19406), .Z(n10827) );
  XNOR U11302 ( .A(b[29]), .B(a[58]), .Z(n10960) );
  OR U11303 ( .A(n10960), .B(n576), .Z(n10826) );
  NAND U11304 ( .A(n10827), .B(n10826), .Z(n10890) );
  NANDN U11305 ( .A(n585), .B(a[54]), .Z(n10891) );
  XNOR U11306 ( .A(n10890), .B(n10891), .Z(n10893) );
  XNOR U11307 ( .A(n10892), .B(n10893), .Z(n10867) );
  XOR U11308 ( .A(b[23]), .B(a[64]), .Z(n10966) );
  NANDN U11309 ( .A(n19127), .B(n10966), .Z(n10830) );
  NAND U11310 ( .A(n10828), .B(n19128), .Z(n10829) );
  NAND U11311 ( .A(n10830), .B(n10829), .Z(n10935) );
  NAND U11312 ( .A(n10831), .B(n17553), .Z(n10833) );
  XNOR U11313 ( .A(b[7]), .B(a[80]), .Z(n10969) );
  NANDN U11314 ( .A(n10969), .B(n17555), .Z(n10832) );
  NAND U11315 ( .A(n10833), .B(n10832), .Z(n10932) );
  XOR U11316 ( .A(b[25]), .B(a[62]), .Z(n10972) );
  NAND U11317 ( .A(n10972), .B(n19240), .Z(n10836) );
  NAND U11318 ( .A(n10834), .B(n19242), .Z(n10835) );
  AND U11319 ( .A(n10836), .B(n10835), .Z(n10933) );
  XNOR U11320 ( .A(n10932), .B(n10933), .Z(n10934) );
  XOR U11321 ( .A(n10935), .B(n10934), .Z(n10866) );
  XOR U11322 ( .A(n10869), .B(n10868), .Z(n10923) );
  XNOR U11323 ( .A(n10922), .B(n10923), .Z(n10979) );
  XNOR U11324 ( .A(n10980), .B(n10979), .Z(n10982) );
  XNOR U11325 ( .A(n10981), .B(n10982), .Z(n10991) );
  XNOR U11326 ( .A(n10992), .B(n10991), .Z(n10993) );
  XOR U11327 ( .A(n10994), .B(n10993), .Z(n10988) );
  NANDN U11328 ( .A(n10838), .B(n10837), .Z(n10842) );
  OR U11329 ( .A(n10840), .B(n10839), .Z(n10841) );
  NAND U11330 ( .A(n10842), .B(n10841), .Z(n10985) );
  NAND U11331 ( .A(n10844), .B(n10843), .Z(n10848) );
  NANDN U11332 ( .A(n10846), .B(n10845), .Z(n10847) );
  NAND U11333 ( .A(n10848), .B(n10847), .Z(n10986) );
  XNOR U11334 ( .A(n10985), .B(n10986), .Z(n10987) );
  XOR U11335 ( .A(n10988), .B(n10987), .Z(n10863) );
  XOR U11336 ( .A(n10862), .B(n10863), .Z(n10854) );
  XOR U11337 ( .A(n10855), .B(n10854), .Z(n10856) );
  XNOR U11338 ( .A(n10857), .B(n10856), .Z(n10997) );
  XNOR U11339 ( .A(n10997), .B(sreg[182]), .Z(n10999) );
  NAND U11340 ( .A(n10849), .B(sreg[181]), .Z(n10853) );
  OR U11341 ( .A(n10851), .B(n10850), .Z(n10852) );
  AND U11342 ( .A(n10853), .B(n10852), .Z(n10998) );
  XOR U11343 ( .A(n10999), .B(n10998), .Z(c[182]) );
  NAND U11344 ( .A(n10855), .B(n10854), .Z(n10859) );
  NAND U11345 ( .A(n10857), .B(n10856), .Z(n10858) );
  NAND U11346 ( .A(n10859), .B(n10858), .Z(n11005) );
  NANDN U11347 ( .A(n10861), .B(n10860), .Z(n10865) );
  NAND U11348 ( .A(n10863), .B(n10862), .Z(n10864) );
  NAND U11349 ( .A(n10865), .B(n10864), .Z(n11003) );
  NANDN U11350 ( .A(n10867), .B(n10866), .Z(n10871) );
  NANDN U11351 ( .A(n10869), .B(n10868), .Z(n10870) );
  NAND U11352 ( .A(n10871), .B(n10870), .Z(n11123) );
  OR U11353 ( .A(n10873), .B(n10872), .Z(n10877) );
  NAND U11354 ( .A(n10875), .B(n10874), .Z(n10876) );
  NAND U11355 ( .A(n10877), .B(n10876), .Z(n11062) );
  OR U11356 ( .A(n10879), .B(n10878), .Z(n10883) );
  NANDN U11357 ( .A(n10881), .B(n10880), .Z(n10882) );
  NAND U11358 ( .A(n10883), .B(n10882), .Z(n11061) );
  OR U11359 ( .A(n10885), .B(n10884), .Z(n10889) );
  NANDN U11360 ( .A(n10887), .B(n10886), .Z(n10888) );
  NAND U11361 ( .A(n10889), .B(n10888), .Z(n11060) );
  XOR U11362 ( .A(n11062), .B(n11063), .Z(n11120) );
  NANDN U11363 ( .A(n10891), .B(n10890), .Z(n10895) );
  NAND U11364 ( .A(n10893), .B(n10892), .Z(n10894) );
  NAND U11365 ( .A(n10895), .B(n10894), .Z(n11075) );
  NANDN U11366 ( .A(n10896), .B(n18832), .Z(n10898) );
  XNOR U11367 ( .A(b[19]), .B(a[69]), .Z(n11042) );
  NANDN U11368 ( .A(n11042), .B(n18834), .Z(n10897) );
  NAND U11369 ( .A(n10898), .B(n10897), .Z(n11111) );
  XNOR U11370 ( .A(b[27]), .B(a[61]), .Z(n11045) );
  NANDN U11371 ( .A(n11045), .B(n19336), .Z(n10901) );
  NANDN U11372 ( .A(n10899), .B(n19337), .Z(n10900) );
  NAND U11373 ( .A(n10901), .B(n10900), .Z(n11108) );
  XOR U11374 ( .A(b[5]), .B(a[83]), .Z(n11048) );
  NAND U11375 ( .A(n11048), .B(n17310), .Z(n10904) );
  NAND U11376 ( .A(n10902), .B(n17311), .Z(n10903) );
  AND U11377 ( .A(n10904), .B(n10903), .Z(n11109) );
  XNOR U11378 ( .A(n11108), .B(n11109), .Z(n11110) );
  XNOR U11379 ( .A(n11111), .B(n11110), .Z(n11072) );
  XOR U11380 ( .A(b[17]), .B(a[71]), .Z(n11051) );
  NAND U11381 ( .A(n11051), .B(n18673), .Z(n10907) );
  NAND U11382 ( .A(n10905), .B(n18674), .Z(n10906) );
  NAND U11383 ( .A(n10907), .B(n10906), .Z(n11026) );
  XNOR U11384 ( .A(b[31]), .B(a[57]), .Z(n11054) );
  NANDN U11385 ( .A(n11054), .B(n19472), .Z(n10910) );
  NANDN U11386 ( .A(n10908), .B(n19473), .Z(n10909) );
  AND U11387 ( .A(n10910), .B(n10909), .Z(n11024) );
  OR U11388 ( .A(n10911), .B(n16988), .Z(n10913) );
  XNOR U11389 ( .A(b[3]), .B(a[85]), .Z(n11057) );
  NANDN U11390 ( .A(n11057), .B(n16990), .Z(n10912) );
  AND U11391 ( .A(n10913), .B(n10912), .Z(n11025) );
  XOR U11392 ( .A(n11026), .B(n11027), .Z(n11073) );
  XOR U11393 ( .A(n11072), .B(n11073), .Z(n11074) );
  XNOR U11394 ( .A(n11075), .B(n11074), .Z(n11121) );
  XNOR U11395 ( .A(n11120), .B(n11121), .Z(n11122) );
  XNOR U11396 ( .A(n11123), .B(n11122), .Z(n11141) );
  OR U11397 ( .A(n10915), .B(n10914), .Z(n10919) );
  NANDN U11398 ( .A(n10917), .B(n10916), .Z(n10918) );
  NAND U11399 ( .A(n10919), .B(n10918), .Z(n11139) );
  NANDN U11400 ( .A(n10921), .B(n10920), .Z(n10925) );
  NANDN U11401 ( .A(n10923), .B(n10922), .Z(n10924) );
  NAND U11402 ( .A(n10925), .B(n10924), .Z(n11128) );
  OR U11403 ( .A(n10927), .B(n10926), .Z(n10931) );
  NANDN U11404 ( .A(n10929), .B(n10928), .Z(n10930) );
  NAND U11405 ( .A(n10931), .B(n10930), .Z(n11127) );
  NANDN U11406 ( .A(n10933), .B(n10932), .Z(n10937) );
  NAND U11407 ( .A(n10935), .B(n10934), .Z(n10936) );
  NAND U11408 ( .A(n10937), .B(n10936), .Z(n11066) );
  NANDN U11409 ( .A(n10939), .B(n10938), .Z(n10943) );
  NAND U11410 ( .A(n10941), .B(n10940), .Z(n10942) );
  AND U11411 ( .A(n10943), .B(n10942), .Z(n11067) );
  XNOR U11412 ( .A(n11066), .B(n11067), .Z(n11068) );
  XNOR U11413 ( .A(n579), .B(a[79]), .Z(n11078) );
  NAND U11414 ( .A(n17814), .B(n11078), .Z(n10946) );
  NANDN U11415 ( .A(n10944), .B(n17815), .Z(n10945) );
  NAND U11416 ( .A(n10946), .B(n10945), .Z(n11032) );
  NAND U11417 ( .A(n10947), .B(n18513), .Z(n10949) );
  XOR U11418 ( .A(b[15]), .B(a[73]), .Z(n11081) );
  NANDN U11419 ( .A(n18512), .B(n11081), .Z(n10948) );
  AND U11420 ( .A(n10949), .B(n10948), .Z(n11030) );
  NANDN U11421 ( .A(n10950), .B(n19013), .Z(n10952) );
  XNOR U11422 ( .A(n582), .B(a[67]), .Z(n11084) );
  NAND U11423 ( .A(n11084), .B(n19015), .Z(n10951) );
  AND U11424 ( .A(n10952), .B(n10951), .Z(n11031) );
  XOR U11425 ( .A(n11032), .B(n11033), .Z(n11021) );
  XNOR U11426 ( .A(b[11]), .B(a[77]), .Z(n11087) );
  OR U11427 ( .A(n11087), .B(n18194), .Z(n10955) );
  NANDN U11428 ( .A(n10953), .B(n18104), .Z(n10954) );
  NAND U11429 ( .A(n10955), .B(n10954), .Z(n11019) );
  XOR U11430 ( .A(n580), .B(a[75]), .Z(n11090) );
  NANDN U11431 ( .A(n11090), .B(n18336), .Z(n10958) );
  NANDN U11432 ( .A(n10956), .B(n18337), .Z(n10957) );
  NAND U11433 ( .A(n10958), .B(n10957), .Z(n11018) );
  XOR U11434 ( .A(n11021), .B(n11020), .Z(n11015) );
  ANDN U11435 ( .B(b[31]), .A(n10959), .Z(n11036) );
  NANDN U11436 ( .A(n10960), .B(n19406), .Z(n10962) );
  XNOR U11437 ( .A(n584), .B(a[59]), .Z(n11096) );
  NANDN U11438 ( .A(n576), .B(n11096), .Z(n10961) );
  NAND U11439 ( .A(n10962), .B(n10961), .Z(n11037) );
  XOR U11440 ( .A(n11036), .B(n11037), .Z(n11038) );
  NANDN U11441 ( .A(n577), .B(a[87]), .Z(n10963) );
  XOR U11442 ( .A(n17151), .B(n10963), .Z(n10965) );
  IV U11443 ( .A(a[86]), .Z(n15429) );
  NANDN U11444 ( .A(n15429), .B(n577), .Z(n10964) );
  AND U11445 ( .A(n10965), .B(n10964), .Z(n11039) );
  XNOR U11446 ( .A(n11038), .B(n11039), .Z(n11012) );
  XNOR U11447 ( .A(b[23]), .B(a[65]), .Z(n11099) );
  OR U11448 ( .A(n11099), .B(n19127), .Z(n10968) );
  NAND U11449 ( .A(n10966), .B(n19128), .Z(n10967) );
  NAND U11450 ( .A(n10968), .B(n10967), .Z(n11117) );
  NANDN U11451 ( .A(n10969), .B(n17553), .Z(n10971) );
  XOR U11452 ( .A(b[7]), .B(a[81]), .Z(n11102) );
  NAND U11453 ( .A(n11102), .B(n17555), .Z(n10970) );
  NAND U11454 ( .A(n10971), .B(n10970), .Z(n11114) );
  XOR U11455 ( .A(b[25]), .B(a[63]), .Z(n11105) );
  NAND U11456 ( .A(n11105), .B(n19240), .Z(n10974) );
  NAND U11457 ( .A(n10972), .B(n19242), .Z(n10973) );
  AND U11458 ( .A(n10974), .B(n10973), .Z(n11115) );
  XNOR U11459 ( .A(n11114), .B(n11115), .Z(n11116) );
  XNOR U11460 ( .A(n11117), .B(n11116), .Z(n11013) );
  XOR U11461 ( .A(n11015), .B(n11014), .Z(n11069) );
  XNOR U11462 ( .A(n11068), .B(n11069), .Z(n11126) );
  XNOR U11463 ( .A(n11127), .B(n11126), .Z(n11129) );
  XNOR U11464 ( .A(n11128), .B(n11129), .Z(n11138) );
  XNOR U11465 ( .A(n11139), .B(n11138), .Z(n11140) );
  XOR U11466 ( .A(n11141), .B(n11140), .Z(n11135) );
  NAND U11467 ( .A(n10980), .B(n10979), .Z(n10984) );
  NANDN U11468 ( .A(n10982), .B(n10981), .Z(n10983) );
  AND U11469 ( .A(n10984), .B(n10983), .Z(n11132) );
  XNOR U11470 ( .A(n11133), .B(n11132), .Z(n11134) );
  XNOR U11471 ( .A(n11135), .B(n11134), .Z(n11009) );
  NANDN U11472 ( .A(n10986), .B(n10985), .Z(n10990) );
  NAND U11473 ( .A(n10988), .B(n10987), .Z(n10989) );
  NAND U11474 ( .A(n10990), .B(n10989), .Z(n11006) );
  NANDN U11475 ( .A(n10992), .B(n10991), .Z(n10996) );
  NANDN U11476 ( .A(n10994), .B(n10993), .Z(n10995) );
  NAND U11477 ( .A(n10996), .B(n10995), .Z(n11007) );
  XNOR U11478 ( .A(n11006), .B(n11007), .Z(n11008) );
  XNOR U11479 ( .A(n11009), .B(n11008), .Z(n11002) );
  XOR U11480 ( .A(n11003), .B(n11002), .Z(n11004) );
  XNOR U11481 ( .A(n11005), .B(n11004), .Z(n11144) );
  XNOR U11482 ( .A(n11144), .B(sreg[183]), .Z(n11146) );
  NAND U11483 ( .A(n10997), .B(sreg[182]), .Z(n11001) );
  OR U11484 ( .A(n10999), .B(n10998), .Z(n11000) );
  AND U11485 ( .A(n11001), .B(n11000), .Z(n11145) );
  XOR U11486 ( .A(n11146), .B(n11145), .Z(c[183]) );
  NANDN U11487 ( .A(n11007), .B(n11006), .Z(n11011) );
  NANDN U11488 ( .A(n11009), .B(n11008), .Z(n11010) );
  NAND U11489 ( .A(n11011), .B(n11010), .Z(n11150) );
  OR U11490 ( .A(n11013), .B(n11012), .Z(n11017) );
  NANDN U11491 ( .A(n11015), .B(n11014), .Z(n11016) );
  NAND U11492 ( .A(n11017), .B(n11016), .Z(n11280) );
  OR U11493 ( .A(n11019), .B(n11018), .Z(n11023) );
  NAND U11494 ( .A(n11021), .B(n11020), .Z(n11022) );
  NAND U11495 ( .A(n11023), .B(n11022), .Z(n11219) );
  OR U11496 ( .A(n11025), .B(n11024), .Z(n11029) );
  NANDN U11497 ( .A(n11027), .B(n11026), .Z(n11028) );
  NAND U11498 ( .A(n11029), .B(n11028), .Z(n11218) );
  OR U11499 ( .A(n11031), .B(n11030), .Z(n11035) );
  NANDN U11500 ( .A(n11033), .B(n11032), .Z(n11034) );
  NAND U11501 ( .A(n11035), .B(n11034), .Z(n11217) );
  XOR U11502 ( .A(n11219), .B(n11220), .Z(n11278) );
  OR U11503 ( .A(n11037), .B(n11036), .Z(n11041) );
  NANDN U11504 ( .A(n11039), .B(n11038), .Z(n11040) );
  NAND U11505 ( .A(n11041), .B(n11040), .Z(n11231) );
  NANDN U11506 ( .A(n11042), .B(n18832), .Z(n11044) );
  XNOR U11507 ( .A(b[19]), .B(a[70]), .Z(n11177) );
  NANDN U11508 ( .A(n11177), .B(n18834), .Z(n11043) );
  NAND U11509 ( .A(n11044), .B(n11043), .Z(n11244) );
  XNOR U11510 ( .A(b[27]), .B(a[62]), .Z(n11180) );
  NANDN U11511 ( .A(n11180), .B(n19336), .Z(n11047) );
  NANDN U11512 ( .A(n11045), .B(n19337), .Z(n11046) );
  NAND U11513 ( .A(n11047), .B(n11046), .Z(n11241) );
  XNOR U11514 ( .A(b[5]), .B(a[84]), .Z(n11183) );
  NANDN U11515 ( .A(n11183), .B(n17310), .Z(n11050) );
  NAND U11516 ( .A(n11048), .B(n17311), .Z(n11049) );
  AND U11517 ( .A(n11050), .B(n11049), .Z(n11242) );
  XNOR U11518 ( .A(n11241), .B(n11242), .Z(n11243) );
  XNOR U11519 ( .A(n11244), .B(n11243), .Z(n11230) );
  XOR U11520 ( .A(b[17]), .B(a[72]), .Z(n11186) );
  NAND U11521 ( .A(n11186), .B(n18673), .Z(n11053) );
  NAND U11522 ( .A(n11051), .B(n18674), .Z(n11052) );
  NAND U11523 ( .A(n11053), .B(n11052), .Z(n11204) );
  XNOR U11524 ( .A(b[31]), .B(a[58]), .Z(n11189) );
  NANDN U11525 ( .A(n11189), .B(n19472), .Z(n11056) );
  NANDN U11526 ( .A(n11054), .B(n19473), .Z(n11055) );
  NAND U11527 ( .A(n11056), .B(n11055), .Z(n11201) );
  OR U11528 ( .A(n11057), .B(n16988), .Z(n11059) );
  XOR U11529 ( .A(b[3]), .B(n15429), .Z(n11192) );
  NANDN U11530 ( .A(n11192), .B(n16990), .Z(n11058) );
  AND U11531 ( .A(n11059), .B(n11058), .Z(n11202) );
  XNOR U11532 ( .A(n11201), .B(n11202), .Z(n11203) );
  XOR U11533 ( .A(n11204), .B(n11203), .Z(n11229) );
  XOR U11534 ( .A(n11230), .B(n11229), .Z(n11232) );
  XOR U11535 ( .A(n11231), .B(n11232), .Z(n11277) );
  XOR U11536 ( .A(n11278), .B(n11277), .Z(n11279) );
  XNOR U11537 ( .A(n11280), .B(n11279), .Z(n11168) );
  OR U11538 ( .A(n11061), .B(n11060), .Z(n11065) );
  NANDN U11539 ( .A(n11063), .B(n11062), .Z(n11064) );
  NAND U11540 ( .A(n11065), .B(n11064), .Z(n11166) );
  NANDN U11541 ( .A(n11067), .B(n11066), .Z(n11071) );
  NANDN U11542 ( .A(n11069), .B(n11068), .Z(n11070) );
  NAND U11543 ( .A(n11071), .B(n11070), .Z(n11286) );
  OR U11544 ( .A(n11073), .B(n11072), .Z(n11077) );
  NAND U11545 ( .A(n11075), .B(n11074), .Z(n11076) );
  NAND U11546 ( .A(n11077), .B(n11076), .Z(n11283) );
  XOR U11547 ( .A(b[9]), .B(n14551), .Z(n11247) );
  NANDN U11548 ( .A(n11247), .B(n17814), .Z(n11080) );
  NAND U11549 ( .A(n17815), .B(n11078), .Z(n11079) );
  NAND U11550 ( .A(n11080), .B(n11079), .Z(n11209) );
  XNOR U11551 ( .A(b[15]), .B(a[74]), .Z(n11250) );
  OR U11552 ( .A(n11250), .B(n18512), .Z(n11083) );
  NAND U11553 ( .A(n11081), .B(n18513), .Z(n11082) );
  NAND U11554 ( .A(n11083), .B(n11082), .Z(n11207) );
  XNOR U11555 ( .A(b[21]), .B(a[68]), .Z(n11253) );
  NANDN U11556 ( .A(n11253), .B(n19015), .Z(n11086) );
  NAND U11557 ( .A(n19013), .B(n11084), .Z(n11085) );
  NAND U11558 ( .A(n11086), .B(n11085), .Z(n11208) );
  XNOR U11559 ( .A(n11207), .B(n11208), .Z(n11210) );
  XOR U11560 ( .A(n11209), .B(n11210), .Z(n11198) );
  XNOR U11561 ( .A(b[11]), .B(a[78]), .Z(n11256) );
  OR U11562 ( .A(n11256), .B(n18194), .Z(n11089) );
  NANDN U11563 ( .A(n11087), .B(n18104), .Z(n11088) );
  NAND U11564 ( .A(n11089), .B(n11088), .Z(n11196) );
  XOR U11565 ( .A(n580), .B(a[76]), .Z(n11259) );
  NANDN U11566 ( .A(n11259), .B(n18336), .Z(n11092) );
  NANDN U11567 ( .A(n11090), .B(n18337), .Z(n11091) );
  AND U11568 ( .A(n11092), .B(n11091), .Z(n11195) );
  XNOR U11569 ( .A(n11196), .B(n11195), .Z(n11197) );
  XNOR U11570 ( .A(n11198), .B(n11197), .Z(n11214) );
  NANDN U11571 ( .A(n577), .B(a[88]), .Z(n11093) );
  XOR U11572 ( .A(n17151), .B(n11093), .Z(n11095) );
  NANDN U11573 ( .A(b[0]), .B(a[87]), .Z(n11094) );
  AND U11574 ( .A(n11095), .B(n11094), .Z(n11173) );
  NAND U11575 ( .A(n11096), .B(n19406), .Z(n11098) );
  XNOR U11576 ( .A(n584), .B(a[60]), .Z(n11265) );
  NANDN U11577 ( .A(n576), .B(n11265), .Z(n11097) );
  NAND U11578 ( .A(n11098), .B(n11097), .Z(n11171) );
  NANDN U11579 ( .A(n585), .B(a[56]), .Z(n11172) );
  XNOR U11580 ( .A(n11171), .B(n11172), .Z(n11174) );
  XNOR U11581 ( .A(n11173), .B(n11174), .Z(n11212) );
  XOR U11582 ( .A(b[23]), .B(a[66]), .Z(n11268) );
  NANDN U11583 ( .A(n19127), .B(n11268), .Z(n11101) );
  NANDN U11584 ( .A(n11099), .B(n19128), .Z(n11100) );
  NAND U11585 ( .A(n11101), .B(n11100), .Z(n11238) );
  NAND U11586 ( .A(n11102), .B(n17553), .Z(n11104) );
  XOR U11587 ( .A(b[7]), .B(a[82]), .Z(n11271) );
  NAND U11588 ( .A(n11271), .B(n17555), .Z(n11103) );
  NAND U11589 ( .A(n11104), .B(n11103), .Z(n11235) );
  XOR U11590 ( .A(b[25]), .B(a[64]), .Z(n11274) );
  NAND U11591 ( .A(n11274), .B(n19240), .Z(n11107) );
  NAND U11592 ( .A(n11105), .B(n19242), .Z(n11106) );
  AND U11593 ( .A(n11107), .B(n11106), .Z(n11236) );
  XNOR U11594 ( .A(n11235), .B(n11236), .Z(n11237) );
  XOR U11595 ( .A(n11238), .B(n11237), .Z(n11211) );
  XOR U11596 ( .A(n11214), .B(n11213), .Z(n11226) );
  NANDN U11597 ( .A(n11109), .B(n11108), .Z(n11113) );
  NAND U11598 ( .A(n11111), .B(n11110), .Z(n11112) );
  NAND U11599 ( .A(n11113), .B(n11112), .Z(n11224) );
  NANDN U11600 ( .A(n11115), .B(n11114), .Z(n11119) );
  NAND U11601 ( .A(n11117), .B(n11116), .Z(n11118) );
  AND U11602 ( .A(n11119), .B(n11118), .Z(n11223) );
  XNOR U11603 ( .A(n11224), .B(n11223), .Z(n11225) );
  XNOR U11604 ( .A(n11226), .B(n11225), .Z(n11284) );
  XNOR U11605 ( .A(n11283), .B(n11284), .Z(n11285) );
  XOR U11606 ( .A(n11286), .B(n11285), .Z(n11165) );
  XNOR U11607 ( .A(n11166), .B(n11165), .Z(n11167) );
  XOR U11608 ( .A(n11168), .B(n11167), .Z(n11162) );
  NANDN U11609 ( .A(n11121), .B(n11120), .Z(n11125) );
  NAND U11610 ( .A(n11123), .B(n11122), .Z(n11124) );
  NAND U11611 ( .A(n11125), .B(n11124), .Z(n11160) );
  NAND U11612 ( .A(n11127), .B(n11126), .Z(n11131) );
  NANDN U11613 ( .A(n11129), .B(n11128), .Z(n11130) );
  AND U11614 ( .A(n11131), .B(n11130), .Z(n11159) );
  XNOR U11615 ( .A(n11160), .B(n11159), .Z(n11161) );
  XNOR U11616 ( .A(n11162), .B(n11161), .Z(n11156) );
  NANDN U11617 ( .A(n11133), .B(n11132), .Z(n11137) );
  NAND U11618 ( .A(n11135), .B(n11134), .Z(n11136) );
  NAND U11619 ( .A(n11137), .B(n11136), .Z(n11153) );
  NANDN U11620 ( .A(n11139), .B(n11138), .Z(n11143) );
  NANDN U11621 ( .A(n11141), .B(n11140), .Z(n11142) );
  NAND U11622 ( .A(n11143), .B(n11142), .Z(n11154) );
  XNOR U11623 ( .A(n11153), .B(n11154), .Z(n11155) );
  XNOR U11624 ( .A(n11156), .B(n11155), .Z(n11149) );
  XOR U11625 ( .A(n11150), .B(n11149), .Z(n11151) );
  XNOR U11626 ( .A(n11152), .B(n11151), .Z(n11289) );
  XNOR U11627 ( .A(n11289), .B(sreg[184]), .Z(n11291) );
  NAND U11628 ( .A(n11144), .B(sreg[183]), .Z(n11148) );
  OR U11629 ( .A(n11146), .B(n11145), .Z(n11147) );
  AND U11630 ( .A(n11148), .B(n11147), .Z(n11290) );
  XOR U11631 ( .A(n11291), .B(n11290), .Z(c[184]) );
  NANDN U11632 ( .A(n11154), .B(n11153), .Z(n11158) );
  NANDN U11633 ( .A(n11156), .B(n11155), .Z(n11157) );
  NAND U11634 ( .A(n11158), .B(n11157), .Z(n11295) );
  NANDN U11635 ( .A(n11160), .B(n11159), .Z(n11164) );
  NAND U11636 ( .A(n11162), .B(n11161), .Z(n11163) );
  NAND U11637 ( .A(n11164), .B(n11163), .Z(n11300) );
  NANDN U11638 ( .A(n11166), .B(n11165), .Z(n11170) );
  NANDN U11639 ( .A(n11168), .B(n11167), .Z(n11169) );
  NAND U11640 ( .A(n11170), .B(n11169), .Z(n11301) );
  XNOR U11641 ( .A(n11300), .B(n11301), .Z(n11302) );
  NANDN U11642 ( .A(n11172), .B(n11171), .Z(n11176) );
  NAND U11643 ( .A(n11174), .B(n11173), .Z(n11175) );
  NAND U11644 ( .A(n11176), .B(n11175), .Z(n11375) );
  NANDN U11645 ( .A(n11177), .B(n18832), .Z(n11179) );
  XNOR U11646 ( .A(b[19]), .B(a[71]), .Z(n11320) );
  NANDN U11647 ( .A(n11320), .B(n18834), .Z(n11178) );
  NAND U11648 ( .A(n11179), .B(n11178), .Z(n11385) );
  XNOR U11649 ( .A(b[27]), .B(a[63]), .Z(n11323) );
  NANDN U11650 ( .A(n11323), .B(n19336), .Z(n11182) );
  NANDN U11651 ( .A(n11180), .B(n19337), .Z(n11181) );
  NAND U11652 ( .A(n11182), .B(n11181), .Z(n11382) );
  XOR U11653 ( .A(b[5]), .B(a[85]), .Z(n11326) );
  NAND U11654 ( .A(n11326), .B(n17310), .Z(n11185) );
  NANDN U11655 ( .A(n11183), .B(n17311), .Z(n11184) );
  AND U11656 ( .A(n11185), .B(n11184), .Z(n11383) );
  XNOR U11657 ( .A(n11382), .B(n11383), .Z(n11384) );
  XNOR U11658 ( .A(n11385), .B(n11384), .Z(n11373) );
  XOR U11659 ( .A(b[17]), .B(a[73]), .Z(n11329) );
  NAND U11660 ( .A(n11329), .B(n18673), .Z(n11188) );
  NAND U11661 ( .A(n11186), .B(n18674), .Z(n11187) );
  NAND U11662 ( .A(n11188), .B(n11187), .Z(n11347) );
  XNOR U11663 ( .A(b[31]), .B(a[59]), .Z(n11332) );
  NANDN U11664 ( .A(n11332), .B(n19472), .Z(n11191) );
  NANDN U11665 ( .A(n11189), .B(n19473), .Z(n11190) );
  NAND U11666 ( .A(n11191), .B(n11190), .Z(n11344) );
  OR U11667 ( .A(n11192), .B(n16988), .Z(n11194) );
  XNOR U11668 ( .A(b[3]), .B(a[87]), .Z(n11335) );
  NANDN U11669 ( .A(n11335), .B(n16990), .Z(n11193) );
  AND U11670 ( .A(n11194), .B(n11193), .Z(n11345) );
  XNOR U11671 ( .A(n11344), .B(n11345), .Z(n11346) );
  XOR U11672 ( .A(n11347), .B(n11346), .Z(n11372) );
  XNOR U11673 ( .A(n11373), .B(n11372), .Z(n11374) );
  XNOR U11674 ( .A(n11375), .B(n11374), .Z(n11311) );
  NANDN U11675 ( .A(n11196), .B(n11195), .Z(n11200) );
  NAND U11676 ( .A(n11198), .B(n11197), .Z(n11199) );
  NAND U11677 ( .A(n11200), .B(n11199), .Z(n11364) );
  NANDN U11678 ( .A(n11202), .B(n11201), .Z(n11206) );
  NAND U11679 ( .A(n11204), .B(n11203), .Z(n11205) );
  NAND U11680 ( .A(n11206), .B(n11205), .Z(n11363) );
  XNOR U11681 ( .A(n11363), .B(n11362), .Z(n11365) );
  XOR U11682 ( .A(n11364), .B(n11365), .Z(n11310) );
  XOR U11683 ( .A(n11311), .B(n11310), .Z(n11312) );
  NANDN U11684 ( .A(n11212), .B(n11211), .Z(n11216) );
  NAND U11685 ( .A(n11214), .B(n11213), .Z(n11215) );
  NAND U11686 ( .A(n11216), .B(n11215), .Z(n11313) );
  XNOR U11687 ( .A(n11312), .B(n11313), .Z(n11426) );
  OR U11688 ( .A(n11218), .B(n11217), .Z(n11222) );
  NANDN U11689 ( .A(n11220), .B(n11219), .Z(n11221) );
  NAND U11690 ( .A(n11222), .B(n11221), .Z(n11425) );
  NANDN U11691 ( .A(n11224), .B(n11223), .Z(n11228) );
  NANDN U11692 ( .A(n11226), .B(n11225), .Z(n11227) );
  NAND U11693 ( .A(n11228), .B(n11227), .Z(n11308) );
  NANDN U11694 ( .A(n11230), .B(n11229), .Z(n11234) );
  OR U11695 ( .A(n11232), .B(n11231), .Z(n11233) );
  NAND U11696 ( .A(n11234), .B(n11233), .Z(n11307) );
  NANDN U11697 ( .A(n11236), .B(n11235), .Z(n11240) );
  NAND U11698 ( .A(n11238), .B(n11237), .Z(n11239) );
  NAND U11699 ( .A(n11240), .B(n11239), .Z(n11366) );
  NANDN U11700 ( .A(n11242), .B(n11241), .Z(n11246) );
  NAND U11701 ( .A(n11244), .B(n11243), .Z(n11245) );
  AND U11702 ( .A(n11246), .B(n11245), .Z(n11367) );
  XNOR U11703 ( .A(n11366), .B(n11367), .Z(n11368) );
  XNOR U11704 ( .A(n579), .B(a[81]), .Z(n11394) );
  NAND U11705 ( .A(n17814), .B(n11394), .Z(n11249) );
  NANDN U11706 ( .A(n11247), .B(n17815), .Z(n11248) );
  NAND U11707 ( .A(n11249), .B(n11248), .Z(n11352) );
  NANDN U11708 ( .A(n11250), .B(n18513), .Z(n11252) );
  XOR U11709 ( .A(b[15]), .B(a[75]), .Z(n11391) );
  NANDN U11710 ( .A(n18512), .B(n11391), .Z(n11251) );
  AND U11711 ( .A(n11252), .B(n11251), .Z(n11350) );
  NANDN U11712 ( .A(n11253), .B(n19013), .Z(n11255) );
  XNOR U11713 ( .A(n582), .B(a[69]), .Z(n11388) );
  NAND U11714 ( .A(n11388), .B(n19015), .Z(n11254) );
  AND U11715 ( .A(n11255), .B(n11254), .Z(n11351) );
  XOR U11716 ( .A(n11352), .B(n11353), .Z(n11341) );
  XNOR U11717 ( .A(b[11]), .B(a[79]), .Z(n11397) );
  OR U11718 ( .A(n11397), .B(n18194), .Z(n11258) );
  NANDN U11719 ( .A(n11256), .B(n18104), .Z(n11257) );
  NAND U11720 ( .A(n11258), .B(n11257), .Z(n11339) );
  XOR U11721 ( .A(n580), .B(a[77]), .Z(n11400) );
  NANDN U11722 ( .A(n11400), .B(n18336), .Z(n11261) );
  NANDN U11723 ( .A(n11259), .B(n18337), .Z(n11260) );
  AND U11724 ( .A(n11261), .B(n11260), .Z(n11338) );
  XNOR U11725 ( .A(n11339), .B(n11338), .Z(n11340) );
  XOR U11726 ( .A(n11341), .B(n11340), .Z(n11358) );
  NANDN U11727 ( .A(n577), .B(a[89]), .Z(n11262) );
  XOR U11728 ( .A(n17151), .B(n11262), .Z(n11264) );
  NANDN U11729 ( .A(b[0]), .B(a[88]), .Z(n11263) );
  AND U11730 ( .A(n11264), .B(n11263), .Z(n11316) );
  NAND U11731 ( .A(n19406), .B(n11265), .Z(n11267) );
  XNOR U11732 ( .A(n584), .B(a[61]), .Z(n11406) );
  NANDN U11733 ( .A(n576), .B(n11406), .Z(n11266) );
  NAND U11734 ( .A(n11267), .B(n11266), .Z(n11314) );
  NANDN U11735 ( .A(n585), .B(a[57]), .Z(n11315) );
  XNOR U11736 ( .A(n11314), .B(n11315), .Z(n11317) );
  XOR U11737 ( .A(n11316), .B(n11317), .Z(n11356) );
  XOR U11738 ( .A(b[23]), .B(a[67]), .Z(n11409) );
  NANDN U11739 ( .A(n19127), .B(n11409), .Z(n11270) );
  NAND U11740 ( .A(n11268), .B(n19128), .Z(n11269) );
  NAND U11741 ( .A(n11270), .B(n11269), .Z(n11379) );
  NAND U11742 ( .A(n11271), .B(n17553), .Z(n11273) );
  XOR U11743 ( .A(b[7]), .B(a[83]), .Z(n11412) );
  NAND U11744 ( .A(n11412), .B(n17555), .Z(n11272) );
  NAND U11745 ( .A(n11273), .B(n11272), .Z(n11376) );
  XNOR U11746 ( .A(b[25]), .B(a[65]), .Z(n11415) );
  NANDN U11747 ( .A(n11415), .B(n19240), .Z(n11276) );
  NAND U11748 ( .A(n11274), .B(n19242), .Z(n11275) );
  AND U11749 ( .A(n11276), .B(n11275), .Z(n11377) );
  XNOR U11750 ( .A(n11376), .B(n11377), .Z(n11378) );
  XNOR U11751 ( .A(n11379), .B(n11378), .Z(n11357) );
  XOR U11752 ( .A(n11356), .B(n11357), .Z(n11359) );
  XNOR U11753 ( .A(n11358), .B(n11359), .Z(n11369) );
  XNOR U11754 ( .A(n11368), .B(n11369), .Z(n11306) );
  XNOR U11755 ( .A(n11307), .B(n11306), .Z(n11309) );
  XOR U11756 ( .A(n11308), .B(n11309), .Z(n11424) );
  XOR U11757 ( .A(n11425), .B(n11424), .Z(n11427) );
  NAND U11758 ( .A(n11278), .B(n11277), .Z(n11282) );
  NAND U11759 ( .A(n11280), .B(n11279), .Z(n11281) );
  NAND U11760 ( .A(n11282), .B(n11281), .Z(n11419) );
  NANDN U11761 ( .A(n11284), .B(n11283), .Z(n11288) );
  NAND U11762 ( .A(n11286), .B(n11285), .Z(n11287) );
  AND U11763 ( .A(n11288), .B(n11287), .Z(n11418) );
  XNOR U11764 ( .A(n11419), .B(n11418), .Z(n11420) );
  XOR U11765 ( .A(n11421), .B(n11420), .Z(n11303) );
  XOR U11766 ( .A(n11302), .B(n11303), .Z(n11294) );
  XOR U11767 ( .A(n11295), .B(n11294), .Z(n11296) );
  XNOR U11768 ( .A(n11297), .B(n11296), .Z(n11430) );
  XNOR U11769 ( .A(n11430), .B(sreg[185]), .Z(n11432) );
  NAND U11770 ( .A(n11289), .B(sreg[184]), .Z(n11293) );
  OR U11771 ( .A(n11291), .B(n11290), .Z(n11292) );
  AND U11772 ( .A(n11293), .B(n11292), .Z(n11431) );
  XOR U11773 ( .A(n11432), .B(n11431), .Z(c[185]) );
  NAND U11774 ( .A(n11295), .B(n11294), .Z(n11299) );
  NAND U11775 ( .A(n11297), .B(n11296), .Z(n11298) );
  NAND U11776 ( .A(n11299), .B(n11298), .Z(n11438) );
  NANDN U11777 ( .A(n11301), .B(n11300), .Z(n11305) );
  NAND U11778 ( .A(n11303), .B(n11302), .Z(n11304) );
  NAND U11779 ( .A(n11305), .B(n11304), .Z(n11435) );
  XNOR U11780 ( .A(n11563), .B(n11564), .Z(n11565) );
  NANDN U11781 ( .A(n11315), .B(n11314), .Z(n11319) );
  NAND U11782 ( .A(n11317), .B(n11316), .Z(n11318) );
  NAND U11783 ( .A(n11319), .B(n11318), .Z(n11508) );
  NANDN U11784 ( .A(n11320), .B(n18832), .Z(n11322) );
  XNOR U11785 ( .A(b[19]), .B(a[72]), .Z(n11453) );
  NANDN U11786 ( .A(n11453), .B(n18834), .Z(n11321) );
  NAND U11787 ( .A(n11322), .B(n11321), .Z(n11518) );
  XNOR U11788 ( .A(b[27]), .B(a[64]), .Z(n11456) );
  NANDN U11789 ( .A(n11456), .B(n19336), .Z(n11325) );
  NANDN U11790 ( .A(n11323), .B(n19337), .Z(n11324) );
  NAND U11791 ( .A(n11325), .B(n11324), .Z(n11515) );
  XNOR U11792 ( .A(b[5]), .B(a[86]), .Z(n11459) );
  NANDN U11793 ( .A(n11459), .B(n17310), .Z(n11328) );
  NAND U11794 ( .A(n11326), .B(n17311), .Z(n11327) );
  AND U11795 ( .A(n11328), .B(n11327), .Z(n11516) );
  XNOR U11796 ( .A(n11515), .B(n11516), .Z(n11517) );
  XNOR U11797 ( .A(n11518), .B(n11517), .Z(n11506) );
  XOR U11798 ( .A(b[17]), .B(a[74]), .Z(n11462) );
  NAND U11799 ( .A(n11462), .B(n18673), .Z(n11331) );
  NAND U11800 ( .A(n11329), .B(n18674), .Z(n11330) );
  NAND U11801 ( .A(n11331), .B(n11330), .Z(n11480) );
  XNOR U11802 ( .A(b[31]), .B(a[60]), .Z(n11465) );
  NANDN U11803 ( .A(n11465), .B(n19472), .Z(n11334) );
  NANDN U11804 ( .A(n11332), .B(n19473), .Z(n11333) );
  NAND U11805 ( .A(n11334), .B(n11333), .Z(n11477) );
  OR U11806 ( .A(n11335), .B(n16988), .Z(n11337) );
  XNOR U11807 ( .A(b[3]), .B(a[88]), .Z(n11468) );
  NANDN U11808 ( .A(n11468), .B(n16990), .Z(n11336) );
  AND U11809 ( .A(n11337), .B(n11336), .Z(n11478) );
  XNOR U11810 ( .A(n11477), .B(n11478), .Z(n11479) );
  XOR U11811 ( .A(n11480), .B(n11479), .Z(n11505) );
  XNOR U11812 ( .A(n11506), .B(n11505), .Z(n11507) );
  XNOR U11813 ( .A(n11508), .B(n11507), .Z(n11551) );
  NANDN U11814 ( .A(n11339), .B(n11338), .Z(n11343) );
  NAND U11815 ( .A(n11341), .B(n11340), .Z(n11342) );
  NAND U11816 ( .A(n11343), .B(n11342), .Z(n11496) );
  NANDN U11817 ( .A(n11345), .B(n11344), .Z(n11349) );
  NAND U11818 ( .A(n11347), .B(n11346), .Z(n11348) );
  NAND U11819 ( .A(n11349), .B(n11348), .Z(n11494) );
  OR U11820 ( .A(n11351), .B(n11350), .Z(n11355) );
  NANDN U11821 ( .A(n11353), .B(n11352), .Z(n11354) );
  NAND U11822 ( .A(n11355), .B(n11354), .Z(n11493) );
  XNOR U11823 ( .A(n11496), .B(n11495), .Z(n11552) );
  XNOR U11824 ( .A(n11551), .B(n11552), .Z(n11553) );
  NANDN U11825 ( .A(n11357), .B(n11356), .Z(n11361) );
  OR U11826 ( .A(n11359), .B(n11358), .Z(n11360) );
  AND U11827 ( .A(n11361), .B(n11360), .Z(n11554) );
  XOR U11828 ( .A(n11553), .B(n11554), .Z(n11571) );
  NANDN U11829 ( .A(n11367), .B(n11366), .Z(n11371) );
  NANDN U11830 ( .A(n11369), .B(n11368), .Z(n11370) );
  NAND U11831 ( .A(n11371), .B(n11370), .Z(n11560) );
  NANDN U11832 ( .A(n11377), .B(n11376), .Z(n11381) );
  NAND U11833 ( .A(n11379), .B(n11378), .Z(n11380) );
  NAND U11834 ( .A(n11381), .B(n11380), .Z(n11499) );
  NANDN U11835 ( .A(n11383), .B(n11382), .Z(n11387) );
  NAND U11836 ( .A(n11385), .B(n11384), .Z(n11386) );
  AND U11837 ( .A(n11387), .B(n11386), .Z(n11500) );
  XNOR U11838 ( .A(n11499), .B(n11500), .Z(n11501) );
  XNOR U11839 ( .A(b[21]), .B(a[70]), .Z(n11527) );
  NANDN U11840 ( .A(n11527), .B(n19015), .Z(n11390) );
  NAND U11841 ( .A(n19013), .B(n11388), .Z(n11389) );
  NAND U11842 ( .A(n11390), .B(n11389), .Z(n11489) );
  NAND U11843 ( .A(n11391), .B(n18513), .Z(n11393) );
  XOR U11844 ( .A(b[15]), .B(a[76]), .Z(n11524) );
  NANDN U11845 ( .A(n18512), .B(n11524), .Z(n11392) );
  AND U11846 ( .A(n11393), .B(n11392), .Z(n11490) );
  XNOR U11847 ( .A(n11489), .B(n11490), .Z(n11492) );
  XNOR U11848 ( .A(b[9]), .B(a[82]), .Z(n11521) );
  NANDN U11849 ( .A(n11521), .B(n17814), .Z(n11396) );
  NAND U11850 ( .A(n17815), .B(n11394), .Z(n11395) );
  NAND U11851 ( .A(n11396), .B(n11395), .Z(n11491) );
  XNOR U11852 ( .A(n11492), .B(n11491), .Z(n11485) );
  XOR U11853 ( .A(b[11]), .B(n14551), .Z(n11530) );
  OR U11854 ( .A(n11530), .B(n18194), .Z(n11399) );
  NANDN U11855 ( .A(n11397), .B(n18104), .Z(n11398) );
  NAND U11856 ( .A(n11399), .B(n11398), .Z(n11484) );
  XOR U11857 ( .A(n580), .B(a[78]), .Z(n11533) );
  NANDN U11858 ( .A(n11533), .B(n18336), .Z(n11402) );
  NANDN U11859 ( .A(n11400), .B(n18337), .Z(n11401) );
  NAND U11860 ( .A(n11402), .B(n11401), .Z(n11483) );
  XNOR U11861 ( .A(n11484), .B(n11483), .Z(n11486) );
  XNOR U11862 ( .A(n11485), .B(n11486), .Z(n11474) );
  NANDN U11863 ( .A(n577), .B(a[90]), .Z(n11403) );
  XOR U11864 ( .A(n17151), .B(n11403), .Z(n11405) );
  NANDN U11865 ( .A(b[0]), .B(a[89]), .Z(n11404) );
  AND U11866 ( .A(n11405), .B(n11404), .Z(n11449) );
  NAND U11867 ( .A(n19406), .B(n11406), .Z(n11408) );
  XNOR U11868 ( .A(n584), .B(a[62]), .Z(n11539) );
  NANDN U11869 ( .A(n576), .B(n11539), .Z(n11407) );
  NAND U11870 ( .A(n11408), .B(n11407), .Z(n11447) );
  NANDN U11871 ( .A(n585), .B(a[58]), .Z(n11448) );
  XNOR U11872 ( .A(n11447), .B(n11448), .Z(n11450) );
  XNOR U11873 ( .A(n11449), .B(n11450), .Z(n11472) );
  XOR U11874 ( .A(b[23]), .B(a[68]), .Z(n11542) );
  NANDN U11875 ( .A(n19127), .B(n11542), .Z(n11411) );
  NAND U11876 ( .A(n11409), .B(n19128), .Z(n11410) );
  NAND U11877 ( .A(n11411), .B(n11410), .Z(n11512) );
  NAND U11878 ( .A(n11412), .B(n17553), .Z(n11414) );
  XNOR U11879 ( .A(b[7]), .B(a[84]), .Z(n11545) );
  NANDN U11880 ( .A(n11545), .B(n17555), .Z(n11413) );
  NAND U11881 ( .A(n11414), .B(n11413), .Z(n11509) );
  XOR U11882 ( .A(b[25]), .B(a[66]), .Z(n11548) );
  NAND U11883 ( .A(n11548), .B(n19240), .Z(n11417) );
  NANDN U11884 ( .A(n11415), .B(n19242), .Z(n11416) );
  AND U11885 ( .A(n11417), .B(n11416), .Z(n11510) );
  XNOR U11886 ( .A(n11509), .B(n11510), .Z(n11511) );
  XOR U11887 ( .A(n11512), .B(n11511), .Z(n11471) );
  XOR U11888 ( .A(n11474), .B(n11473), .Z(n11502) );
  XNOR U11889 ( .A(n11501), .B(n11502), .Z(n11557) );
  XOR U11890 ( .A(n11558), .B(n11557), .Z(n11559) );
  XNOR U11891 ( .A(n11560), .B(n11559), .Z(n11569) );
  XNOR U11892 ( .A(n11570), .B(n11569), .Z(n11572) );
  XNOR U11893 ( .A(n11571), .B(n11572), .Z(n11566) );
  XOR U11894 ( .A(n11565), .B(n11566), .Z(n11444) );
  NANDN U11895 ( .A(n11419), .B(n11418), .Z(n11423) );
  NAND U11896 ( .A(n11421), .B(n11420), .Z(n11422) );
  NAND U11897 ( .A(n11423), .B(n11422), .Z(n11441) );
  NANDN U11898 ( .A(n11425), .B(n11424), .Z(n11429) );
  OR U11899 ( .A(n11427), .B(n11426), .Z(n11428) );
  NAND U11900 ( .A(n11429), .B(n11428), .Z(n11442) );
  XNOR U11901 ( .A(n11441), .B(n11442), .Z(n11443) );
  XNOR U11902 ( .A(n11444), .B(n11443), .Z(n11436) );
  XNOR U11903 ( .A(n11435), .B(n11436), .Z(n11437) );
  XNOR U11904 ( .A(n11438), .B(n11437), .Z(n11575) );
  XNOR U11905 ( .A(n11575), .B(sreg[186]), .Z(n11577) );
  NAND U11906 ( .A(n11430), .B(sreg[185]), .Z(n11434) );
  OR U11907 ( .A(n11432), .B(n11431), .Z(n11433) );
  AND U11908 ( .A(n11434), .B(n11433), .Z(n11576) );
  XOR U11909 ( .A(n11577), .B(n11576), .Z(c[186]) );
  NANDN U11910 ( .A(n11436), .B(n11435), .Z(n11440) );
  NAND U11911 ( .A(n11438), .B(n11437), .Z(n11439) );
  NAND U11912 ( .A(n11440), .B(n11439), .Z(n11583) );
  NANDN U11913 ( .A(n11442), .B(n11441), .Z(n11446) );
  NAND U11914 ( .A(n11444), .B(n11443), .Z(n11445) );
  NAND U11915 ( .A(n11446), .B(n11445), .Z(n11581) );
  NANDN U11916 ( .A(n11448), .B(n11447), .Z(n11452) );
  NAND U11917 ( .A(n11450), .B(n11449), .Z(n11451) );
  NAND U11918 ( .A(n11452), .B(n11451), .Z(n11653) );
  NANDN U11919 ( .A(n11453), .B(n18832), .Z(n11455) );
  XNOR U11920 ( .A(b[19]), .B(a[73]), .Z(n11598) );
  NANDN U11921 ( .A(n11598), .B(n18834), .Z(n11454) );
  NAND U11922 ( .A(n11455), .B(n11454), .Z(n11663) );
  XOR U11923 ( .A(b[27]), .B(n12055), .Z(n11601) );
  NANDN U11924 ( .A(n11601), .B(n19336), .Z(n11458) );
  NANDN U11925 ( .A(n11456), .B(n19337), .Z(n11457) );
  NAND U11926 ( .A(n11458), .B(n11457), .Z(n11660) );
  XOR U11927 ( .A(b[5]), .B(a[87]), .Z(n11604) );
  NAND U11928 ( .A(n11604), .B(n17310), .Z(n11461) );
  NANDN U11929 ( .A(n11459), .B(n17311), .Z(n11460) );
  AND U11930 ( .A(n11461), .B(n11460), .Z(n11661) );
  XNOR U11931 ( .A(n11660), .B(n11661), .Z(n11662) );
  XNOR U11932 ( .A(n11663), .B(n11662), .Z(n11651) );
  XOR U11933 ( .A(b[17]), .B(a[75]), .Z(n11607) );
  NAND U11934 ( .A(n11607), .B(n18673), .Z(n11464) );
  NAND U11935 ( .A(n11462), .B(n18674), .Z(n11463) );
  NAND U11936 ( .A(n11464), .B(n11463), .Z(n11625) );
  XNOR U11937 ( .A(b[31]), .B(a[61]), .Z(n11610) );
  NANDN U11938 ( .A(n11610), .B(n19472), .Z(n11467) );
  NANDN U11939 ( .A(n11465), .B(n19473), .Z(n11466) );
  NAND U11940 ( .A(n11467), .B(n11466), .Z(n11622) );
  OR U11941 ( .A(n11468), .B(n16988), .Z(n11470) );
  XNOR U11942 ( .A(b[3]), .B(a[89]), .Z(n11613) );
  NANDN U11943 ( .A(n11613), .B(n16990), .Z(n11469) );
  AND U11944 ( .A(n11470), .B(n11469), .Z(n11623) );
  XNOR U11945 ( .A(n11622), .B(n11623), .Z(n11624) );
  XOR U11946 ( .A(n11625), .B(n11624), .Z(n11650) );
  XNOR U11947 ( .A(n11651), .B(n11650), .Z(n11652) );
  XNOR U11948 ( .A(n11653), .B(n11652), .Z(n11702) );
  NANDN U11949 ( .A(n11472), .B(n11471), .Z(n11476) );
  NANDN U11950 ( .A(n11474), .B(n11473), .Z(n11475) );
  NAND U11951 ( .A(n11476), .B(n11475), .Z(n11703) );
  XNOR U11952 ( .A(n11702), .B(n11703), .Z(n11704) );
  NANDN U11953 ( .A(n11478), .B(n11477), .Z(n11482) );
  NAND U11954 ( .A(n11480), .B(n11479), .Z(n11481) );
  NAND U11955 ( .A(n11482), .B(n11481), .Z(n11643) );
  OR U11956 ( .A(n11484), .B(n11483), .Z(n11488) );
  NANDN U11957 ( .A(n11486), .B(n11485), .Z(n11487) );
  NAND U11958 ( .A(n11488), .B(n11487), .Z(n11641) );
  XNOR U11959 ( .A(n11641), .B(n11640), .Z(n11642) );
  XOR U11960 ( .A(n11643), .B(n11642), .Z(n11705) );
  XOR U11961 ( .A(n11704), .B(n11705), .Z(n11715) );
  OR U11962 ( .A(n11494), .B(n11493), .Z(n11498) );
  NAND U11963 ( .A(n11496), .B(n11495), .Z(n11497) );
  NAND U11964 ( .A(n11498), .B(n11497), .Z(n11713) );
  NANDN U11965 ( .A(n11500), .B(n11499), .Z(n11504) );
  NANDN U11966 ( .A(n11502), .B(n11501), .Z(n11503) );
  NAND U11967 ( .A(n11504), .B(n11503), .Z(n11698) );
  NANDN U11968 ( .A(n11510), .B(n11509), .Z(n11514) );
  NAND U11969 ( .A(n11512), .B(n11511), .Z(n11513) );
  NAND U11970 ( .A(n11514), .B(n11513), .Z(n11644) );
  NANDN U11971 ( .A(n11516), .B(n11515), .Z(n11520) );
  NAND U11972 ( .A(n11518), .B(n11517), .Z(n11519) );
  AND U11973 ( .A(n11520), .B(n11519), .Z(n11645) );
  XNOR U11974 ( .A(n11644), .B(n11645), .Z(n11646) );
  XNOR U11975 ( .A(b[9]), .B(a[83]), .Z(n11666) );
  NANDN U11976 ( .A(n11666), .B(n17814), .Z(n11523) );
  NANDN U11977 ( .A(n11521), .B(n17815), .Z(n11522) );
  NAND U11978 ( .A(n11523), .B(n11522), .Z(n11630) );
  NAND U11979 ( .A(n11524), .B(n18513), .Z(n11526) );
  XOR U11980 ( .A(b[15]), .B(a[77]), .Z(n11669) );
  NANDN U11981 ( .A(n18512), .B(n11669), .Z(n11525) );
  AND U11982 ( .A(n11526), .B(n11525), .Z(n11628) );
  NANDN U11983 ( .A(n11527), .B(n19013), .Z(n11529) );
  XNOR U11984 ( .A(b[21]), .B(a[71]), .Z(n11672) );
  NANDN U11985 ( .A(n11672), .B(n19015), .Z(n11528) );
  AND U11986 ( .A(n11529), .B(n11528), .Z(n11629) );
  XOR U11987 ( .A(n11630), .B(n11631), .Z(n11619) );
  XNOR U11988 ( .A(b[11]), .B(a[81]), .Z(n11675) );
  OR U11989 ( .A(n11675), .B(n18194), .Z(n11532) );
  NANDN U11990 ( .A(n11530), .B(n18104), .Z(n11531) );
  NAND U11991 ( .A(n11532), .B(n11531), .Z(n11617) );
  XOR U11992 ( .A(n580), .B(a[79]), .Z(n11678) );
  NANDN U11993 ( .A(n11678), .B(n18336), .Z(n11535) );
  NANDN U11994 ( .A(n11533), .B(n18337), .Z(n11534) );
  AND U11995 ( .A(n11535), .B(n11534), .Z(n11616) );
  XNOR U11996 ( .A(n11617), .B(n11616), .Z(n11618) );
  XOR U11997 ( .A(n11619), .B(n11618), .Z(n11636) );
  NANDN U11998 ( .A(n577), .B(a[91]), .Z(n11536) );
  XOR U11999 ( .A(n17151), .B(n11536), .Z(n11538) );
  NANDN U12000 ( .A(b[0]), .B(a[90]), .Z(n11537) );
  AND U12001 ( .A(n11538), .B(n11537), .Z(n11594) );
  NAND U12002 ( .A(n19406), .B(n11539), .Z(n11541) );
  XNOR U12003 ( .A(n584), .B(a[63]), .Z(n11684) );
  NANDN U12004 ( .A(n576), .B(n11684), .Z(n11540) );
  NAND U12005 ( .A(n11541), .B(n11540), .Z(n11592) );
  NANDN U12006 ( .A(n585), .B(a[59]), .Z(n11593) );
  XNOR U12007 ( .A(n11592), .B(n11593), .Z(n11595) );
  XOR U12008 ( .A(n11594), .B(n11595), .Z(n11634) );
  XOR U12009 ( .A(b[23]), .B(a[69]), .Z(n11687) );
  NANDN U12010 ( .A(n19127), .B(n11687), .Z(n11544) );
  NAND U12011 ( .A(n11542), .B(n19128), .Z(n11543) );
  NAND U12012 ( .A(n11544), .B(n11543), .Z(n11657) );
  NANDN U12013 ( .A(n11545), .B(n17553), .Z(n11547) );
  XOR U12014 ( .A(b[7]), .B(a[85]), .Z(n11690) );
  NAND U12015 ( .A(n11690), .B(n17555), .Z(n11546) );
  NAND U12016 ( .A(n11547), .B(n11546), .Z(n11654) );
  XOR U12017 ( .A(b[25]), .B(a[67]), .Z(n11693) );
  NAND U12018 ( .A(n11693), .B(n19240), .Z(n11550) );
  NAND U12019 ( .A(n11548), .B(n19242), .Z(n11549) );
  AND U12020 ( .A(n11550), .B(n11549), .Z(n11655) );
  XNOR U12021 ( .A(n11654), .B(n11655), .Z(n11656) );
  XNOR U12022 ( .A(n11657), .B(n11656), .Z(n11635) );
  XOR U12023 ( .A(n11634), .B(n11635), .Z(n11637) );
  XNOR U12024 ( .A(n11636), .B(n11637), .Z(n11647) );
  XNOR U12025 ( .A(n11646), .B(n11647), .Z(n11696) );
  XNOR U12026 ( .A(n11697), .B(n11696), .Z(n11699) );
  XNOR U12027 ( .A(n11698), .B(n11699), .Z(n11712) );
  XOR U12028 ( .A(n11713), .B(n11712), .Z(n11714) );
  XNOR U12029 ( .A(n11715), .B(n11714), .Z(n11709) );
  NANDN U12030 ( .A(n11552), .B(n11551), .Z(n11556) );
  NAND U12031 ( .A(n11554), .B(n11553), .Z(n11555) );
  NAND U12032 ( .A(n11556), .B(n11555), .Z(n11706) );
  NAND U12033 ( .A(n11558), .B(n11557), .Z(n11562) );
  NAND U12034 ( .A(n11560), .B(n11559), .Z(n11561) );
  NAND U12035 ( .A(n11562), .B(n11561), .Z(n11707) );
  XNOR U12036 ( .A(n11706), .B(n11707), .Z(n11708) );
  XOR U12037 ( .A(n11709), .B(n11708), .Z(n11588) );
  NANDN U12038 ( .A(n11564), .B(n11563), .Z(n11568) );
  NANDN U12039 ( .A(n11566), .B(n11565), .Z(n11567) );
  NAND U12040 ( .A(n11568), .B(n11567), .Z(n11587) );
  OR U12041 ( .A(n11570), .B(n11569), .Z(n11574) );
  OR U12042 ( .A(n11572), .B(n11571), .Z(n11573) );
  AND U12043 ( .A(n11574), .B(n11573), .Z(n11586) );
  XNOR U12044 ( .A(n11587), .B(n11586), .Z(n11589) );
  XOR U12045 ( .A(n11588), .B(n11589), .Z(n11580) );
  XOR U12046 ( .A(n11581), .B(n11580), .Z(n11582) );
  XNOR U12047 ( .A(n11583), .B(n11582), .Z(n11718) );
  XNOR U12048 ( .A(n11718), .B(sreg[187]), .Z(n11720) );
  NAND U12049 ( .A(n11575), .B(sreg[186]), .Z(n11579) );
  OR U12050 ( .A(n11577), .B(n11576), .Z(n11578) );
  AND U12051 ( .A(n11579), .B(n11578), .Z(n11719) );
  XOR U12052 ( .A(n11720), .B(n11719), .Z(c[187]) );
  NAND U12053 ( .A(n11581), .B(n11580), .Z(n11585) );
  NAND U12054 ( .A(n11583), .B(n11582), .Z(n11584) );
  NAND U12055 ( .A(n11585), .B(n11584), .Z(n11726) );
  NANDN U12056 ( .A(n11587), .B(n11586), .Z(n11591) );
  NAND U12057 ( .A(n11589), .B(n11588), .Z(n11590) );
  NAND U12058 ( .A(n11591), .B(n11590), .Z(n11724) );
  NANDN U12059 ( .A(n11593), .B(n11592), .Z(n11597) );
  NAND U12060 ( .A(n11595), .B(n11594), .Z(n11596) );
  NAND U12061 ( .A(n11597), .B(n11596), .Z(n11806) );
  NANDN U12062 ( .A(n11598), .B(n18832), .Z(n11600) );
  XNOR U12063 ( .A(b[19]), .B(a[74]), .Z(n11773) );
  NANDN U12064 ( .A(n11773), .B(n18834), .Z(n11599) );
  NAND U12065 ( .A(n11600), .B(n11599), .Z(n11818) );
  XNOR U12066 ( .A(b[27]), .B(a[66]), .Z(n11776) );
  NANDN U12067 ( .A(n11776), .B(n19336), .Z(n11603) );
  NANDN U12068 ( .A(n11601), .B(n19337), .Z(n11602) );
  NAND U12069 ( .A(n11603), .B(n11602), .Z(n11815) );
  XOR U12070 ( .A(b[5]), .B(a[88]), .Z(n11779) );
  NAND U12071 ( .A(n11779), .B(n17310), .Z(n11606) );
  NAND U12072 ( .A(n11604), .B(n17311), .Z(n11605) );
  AND U12073 ( .A(n11606), .B(n11605), .Z(n11816) );
  XNOR U12074 ( .A(n11815), .B(n11816), .Z(n11817) );
  XNOR U12075 ( .A(n11818), .B(n11817), .Z(n11803) );
  XOR U12076 ( .A(b[17]), .B(a[76]), .Z(n11782) );
  NAND U12077 ( .A(n11782), .B(n18673), .Z(n11609) );
  NAND U12078 ( .A(n11607), .B(n18674), .Z(n11608) );
  NAND U12079 ( .A(n11609), .B(n11608), .Z(n11757) );
  XNOR U12080 ( .A(b[31]), .B(a[62]), .Z(n11785) );
  NANDN U12081 ( .A(n11785), .B(n19472), .Z(n11612) );
  NANDN U12082 ( .A(n11610), .B(n19473), .Z(n11611) );
  AND U12083 ( .A(n11612), .B(n11611), .Z(n11755) );
  OR U12084 ( .A(n11613), .B(n16988), .Z(n11615) );
  XNOR U12085 ( .A(b[3]), .B(a[90]), .Z(n11788) );
  NANDN U12086 ( .A(n11788), .B(n16990), .Z(n11614) );
  AND U12087 ( .A(n11615), .B(n11614), .Z(n11756) );
  XOR U12088 ( .A(n11757), .B(n11758), .Z(n11804) );
  XOR U12089 ( .A(n11803), .B(n11804), .Z(n11805) );
  XNOR U12090 ( .A(n11806), .B(n11805), .Z(n11851) );
  NANDN U12091 ( .A(n11617), .B(n11616), .Z(n11621) );
  NAND U12092 ( .A(n11619), .B(n11618), .Z(n11620) );
  NAND U12093 ( .A(n11621), .B(n11620), .Z(n11794) );
  NANDN U12094 ( .A(n11623), .B(n11622), .Z(n11627) );
  NAND U12095 ( .A(n11625), .B(n11624), .Z(n11626) );
  NAND U12096 ( .A(n11627), .B(n11626), .Z(n11792) );
  OR U12097 ( .A(n11629), .B(n11628), .Z(n11633) );
  NANDN U12098 ( .A(n11631), .B(n11630), .Z(n11632) );
  NAND U12099 ( .A(n11633), .B(n11632), .Z(n11791) );
  XNOR U12100 ( .A(n11794), .B(n11793), .Z(n11852) );
  XNOR U12101 ( .A(n11851), .B(n11852), .Z(n11853) );
  NANDN U12102 ( .A(n11635), .B(n11634), .Z(n11639) );
  OR U12103 ( .A(n11637), .B(n11636), .Z(n11638) );
  AND U12104 ( .A(n11639), .B(n11638), .Z(n11854) );
  XNOR U12105 ( .A(n11853), .B(n11854), .Z(n11736) );
  NANDN U12106 ( .A(n11645), .B(n11644), .Z(n11649) );
  NANDN U12107 ( .A(n11647), .B(n11646), .Z(n11648) );
  NAND U12108 ( .A(n11649), .B(n11648), .Z(n11860) );
  NANDN U12109 ( .A(n11655), .B(n11654), .Z(n11659) );
  NAND U12110 ( .A(n11657), .B(n11656), .Z(n11658) );
  NAND U12111 ( .A(n11659), .B(n11658), .Z(n11797) );
  NANDN U12112 ( .A(n11661), .B(n11660), .Z(n11665) );
  NAND U12113 ( .A(n11663), .B(n11662), .Z(n11664) );
  AND U12114 ( .A(n11665), .B(n11664), .Z(n11798) );
  XNOR U12115 ( .A(n11797), .B(n11798), .Z(n11799) );
  XOR U12116 ( .A(n579), .B(n15134), .Z(n11821) );
  NAND U12117 ( .A(n17814), .B(n11821), .Z(n11668) );
  NANDN U12118 ( .A(n11666), .B(n17815), .Z(n11667) );
  NAND U12119 ( .A(n11668), .B(n11667), .Z(n11763) );
  NAND U12120 ( .A(n11669), .B(n18513), .Z(n11671) );
  XOR U12121 ( .A(b[15]), .B(a[78]), .Z(n11824) );
  NANDN U12122 ( .A(n18512), .B(n11824), .Z(n11670) );
  AND U12123 ( .A(n11671), .B(n11670), .Z(n11761) );
  NANDN U12124 ( .A(n11672), .B(n19013), .Z(n11674) );
  XNOR U12125 ( .A(n582), .B(a[72]), .Z(n11827) );
  NAND U12126 ( .A(n11827), .B(n19015), .Z(n11673) );
  AND U12127 ( .A(n11674), .B(n11673), .Z(n11762) );
  XOR U12128 ( .A(n11763), .B(n11764), .Z(n11752) );
  XNOR U12129 ( .A(b[11]), .B(a[82]), .Z(n11830) );
  OR U12130 ( .A(n11830), .B(n18194), .Z(n11677) );
  NANDN U12131 ( .A(n11675), .B(n18104), .Z(n11676) );
  NAND U12132 ( .A(n11677), .B(n11676), .Z(n11750) );
  XOR U12133 ( .A(n580), .B(a[80]), .Z(n11833) );
  NANDN U12134 ( .A(n11833), .B(n18336), .Z(n11680) );
  NANDN U12135 ( .A(n11678), .B(n18337), .Z(n11679) );
  NAND U12136 ( .A(n11680), .B(n11679), .Z(n11749) );
  XOR U12137 ( .A(n11752), .B(n11751), .Z(n11746) );
  NANDN U12138 ( .A(n577), .B(a[92]), .Z(n11681) );
  XOR U12139 ( .A(n17151), .B(n11681), .Z(n11683) );
  NANDN U12140 ( .A(b[0]), .B(a[91]), .Z(n11682) );
  AND U12141 ( .A(n11683), .B(n11682), .Z(n11769) );
  NAND U12142 ( .A(n19406), .B(n11684), .Z(n11686) );
  XNOR U12143 ( .A(n584), .B(a[64]), .Z(n11839) );
  NANDN U12144 ( .A(n576), .B(n11839), .Z(n11685) );
  NAND U12145 ( .A(n11686), .B(n11685), .Z(n11767) );
  NANDN U12146 ( .A(n585), .B(a[60]), .Z(n11768) );
  XNOR U12147 ( .A(n11767), .B(n11768), .Z(n11770) );
  XNOR U12148 ( .A(n11769), .B(n11770), .Z(n11744) );
  XOR U12149 ( .A(b[23]), .B(a[70]), .Z(n11842) );
  NANDN U12150 ( .A(n19127), .B(n11842), .Z(n11689) );
  NAND U12151 ( .A(n11687), .B(n19128), .Z(n11688) );
  NAND U12152 ( .A(n11689), .B(n11688), .Z(n11812) );
  NAND U12153 ( .A(n11690), .B(n17553), .Z(n11692) );
  XNOR U12154 ( .A(b[7]), .B(a[86]), .Z(n11845) );
  NANDN U12155 ( .A(n11845), .B(n17555), .Z(n11691) );
  NAND U12156 ( .A(n11692), .B(n11691), .Z(n11809) );
  XOR U12157 ( .A(b[25]), .B(a[68]), .Z(n11848) );
  NAND U12158 ( .A(n11848), .B(n19240), .Z(n11695) );
  NAND U12159 ( .A(n11693), .B(n19242), .Z(n11694) );
  AND U12160 ( .A(n11695), .B(n11694), .Z(n11810) );
  XNOR U12161 ( .A(n11809), .B(n11810), .Z(n11811) );
  XOR U12162 ( .A(n11812), .B(n11811), .Z(n11743) );
  XOR U12163 ( .A(n11746), .B(n11745), .Z(n11800) );
  XNOR U12164 ( .A(n11799), .B(n11800), .Z(n11857) );
  XOR U12165 ( .A(n11858), .B(n11857), .Z(n11859) );
  XOR U12166 ( .A(n11860), .B(n11859), .Z(n11734) );
  XNOR U12167 ( .A(n11733), .B(n11734), .Z(n11735) );
  XNOR U12168 ( .A(n11736), .B(n11735), .Z(n11740) );
  NAND U12169 ( .A(n11697), .B(n11696), .Z(n11701) );
  NANDN U12170 ( .A(n11699), .B(n11698), .Z(n11700) );
  NAND U12171 ( .A(n11701), .B(n11700), .Z(n11737) );
  XNOR U12172 ( .A(n11737), .B(n11738), .Z(n11739) );
  XNOR U12173 ( .A(n11740), .B(n11739), .Z(n11730) );
  NANDN U12174 ( .A(n11707), .B(n11706), .Z(n11711) );
  NAND U12175 ( .A(n11709), .B(n11708), .Z(n11710) );
  NAND U12176 ( .A(n11711), .B(n11710), .Z(n11727) );
  NANDN U12177 ( .A(n11713), .B(n11712), .Z(n11717) );
  OR U12178 ( .A(n11715), .B(n11714), .Z(n11716) );
  NAND U12179 ( .A(n11717), .B(n11716), .Z(n11728) );
  XNOR U12180 ( .A(n11727), .B(n11728), .Z(n11729) );
  XNOR U12181 ( .A(n11730), .B(n11729), .Z(n11723) );
  XOR U12182 ( .A(n11724), .B(n11723), .Z(n11725) );
  XNOR U12183 ( .A(n11726), .B(n11725), .Z(n11863) );
  XNOR U12184 ( .A(n11863), .B(sreg[188]), .Z(n11865) );
  NAND U12185 ( .A(n11718), .B(sreg[187]), .Z(n11722) );
  OR U12186 ( .A(n11720), .B(n11719), .Z(n11721) );
  AND U12187 ( .A(n11722), .B(n11721), .Z(n11864) );
  XOR U12188 ( .A(n11865), .B(n11864), .Z(c[188]) );
  NANDN U12189 ( .A(n11728), .B(n11727), .Z(n11732) );
  NANDN U12190 ( .A(n11730), .B(n11729), .Z(n11731) );
  NAND U12191 ( .A(n11732), .B(n11731), .Z(n11869) );
  NANDN U12192 ( .A(n11738), .B(n11737), .Z(n11742) );
  NANDN U12193 ( .A(n11740), .B(n11739), .Z(n11741) );
  NAND U12194 ( .A(n11742), .B(n11741), .Z(n11875) );
  XNOR U12195 ( .A(n11874), .B(n11875), .Z(n11876) );
  NANDN U12196 ( .A(n11744), .B(n11743), .Z(n11748) );
  NANDN U12197 ( .A(n11746), .B(n11745), .Z(n11747) );
  NAND U12198 ( .A(n11748), .B(n11747), .Z(n11989) );
  OR U12199 ( .A(n11750), .B(n11749), .Z(n11754) );
  NAND U12200 ( .A(n11752), .B(n11751), .Z(n11753) );
  NAND U12201 ( .A(n11754), .B(n11753), .Z(n11928) );
  OR U12202 ( .A(n11756), .B(n11755), .Z(n11760) );
  NANDN U12203 ( .A(n11758), .B(n11757), .Z(n11759) );
  NAND U12204 ( .A(n11760), .B(n11759), .Z(n11927) );
  OR U12205 ( .A(n11762), .B(n11761), .Z(n11766) );
  NANDN U12206 ( .A(n11764), .B(n11763), .Z(n11765) );
  NAND U12207 ( .A(n11766), .B(n11765), .Z(n11926) );
  XOR U12208 ( .A(n11928), .B(n11929), .Z(n11986) );
  NANDN U12209 ( .A(n11768), .B(n11767), .Z(n11772) );
  NAND U12210 ( .A(n11770), .B(n11769), .Z(n11771) );
  NAND U12211 ( .A(n11772), .B(n11771), .Z(n11941) );
  NANDN U12212 ( .A(n11773), .B(n18832), .Z(n11775) );
  XNOR U12213 ( .A(b[19]), .B(a[75]), .Z(n11886) );
  NANDN U12214 ( .A(n11886), .B(n18834), .Z(n11774) );
  NAND U12215 ( .A(n11775), .B(n11774), .Z(n11953) );
  XNOR U12216 ( .A(b[27]), .B(a[67]), .Z(n11889) );
  NANDN U12217 ( .A(n11889), .B(n19336), .Z(n11778) );
  NANDN U12218 ( .A(n11776), .B(n19337), .Z(n11777) );
  NAND U12219 ( .A(n11778), .B(n11777), .Z(n11950) );
  XOR U12220 ( .A(b[5]), .B(a[89]), .Z(n11892) );
  NAND U12221 ( .A(n11892), .B(n17310), .Z(n11781) );
  NAND U12222 ( .A(n11779), .B(n17311), .Z(n11780) );
  AND U12223 ( .A(n11781), .B(n11780), .Z(n11951) );
  XNOR U12224 ( .A(n11950), .B(n11951), .Z(n11952) );
  XNOR U12225 ( .A(n11953), .B(n11952), .Z(n11939) );
  XOR U12226 ( .A(b[17]), .B(a[77]), .Z(n11895) );
  NAND U12227 ( .A(n11895), .B(n18673), .Z(n11784) );
  NAND U12228 ( .A(n11782), .B(n18674), .Z(n11783) );
  NAND U12229 ( .A(n11784), .B(n11783), .Z(n11913) );
  XNOR U12230 ( .A(b[31]), .B(a[63]), .Z(n11898) );
  NANDN U12231 ( .A(n11898), .B(n19472), .Z(n11787) );
  NANDN U12232 ( .A(n11785), .B(n19473), .Z(n11786) );
  NAND U12233 ( .A(n11787), .B(n11786), .Z(n11910) );
  OR U12234 ( .A(n11788), .B(n16988), .Z(n11790) );
  XNOR U12235 ( .A(b[3]), .B(a[91]), .Z(n11901) );
  NANDN U12236 ( .A(n11901), .B(n16990), .Z(n11789) );
  AND U12237 ( .A(n11790), .B(n11789), .Z(n11911) );
  XNOR U12238 ( .A(n11910), .B(n11911), .Z(n11912) );
  XOR U12239 ( .A(n11913), .B(n11912), .Z(n11938) );
  XNOR U12240 ( .A(n11939), .B(n11938), .Z(n11940) );
  XNOR U12241 ( .A(n11941), .B(n11940), .Z(n11987) );
  XNOR U12242 ( .A(n11986), .B(n11987), .Z(n11988) );
  XNOR U12243 ( .A(n11989), .B(n11988), .Z(n12007) );
  OR U12244 ( .A(n11792), .B(n11791), .Z(n11796) );
  NAND U12245 ( .A(n11794), .B(n11793), .Z(n11795) );
  NAND U12246 ( .A(n11796), .B(n11795), .Z(n12005) );
  NANDN U12247 ( .A(n11798), .B(n11797), .Z(n11802) );
  NANDN U12248 ( .A(n11800), .B(n11799), .Z(n11801) );
  NAND U12249 ( .A(n11802), .B(n11801), .Z(n11994) );
  OR U12250 ( .A(n11804), .B(n11803), .Z(n11808) );
  NAND U12251 ( .A(n11806), .B(n11805), .Z(n11807) );
  NAND U12252 ( .A(n11808), .B(n11807), .Z(n11993) );
  NANDN U12253 ( .A(n11810), .B(n11809), .Z(n11814) );
  NAND U12254 ( .A(n11812), .B(n11811), .Z(n11813) );
  NAND U12255 ( .A(n11814), .B(n11813), .Z(n11932) );
  NANDN U12256 ( .A(n11816), .B(n11815), .Z(n11820) );
  NAND U12257 ( .A(n11818), .B(n11817), .Z(n11819) );
  AND U12258 ( .A(n11820), .B(n11819), .Z(n11933) );
  XNOR U12259 ( .A(n11932), .B(n11933), .Z(n11934) );
  XNOR U12260 ( .A(b[9]), .B(a[85]), .Z(n11956) );
  NANDN U12261 ( .A(n11956), .B(n17814), .Z(n11823) );
  NAND U12262 ( .A(n17815), .B(n11821), .Z(n11822) );
  NAND U12263 ( .A(n11823), .B(n11822), .Z(n11918) );
  XNOR U12264 ( .A(b[15]), .B(a[79]), .Z(n11959) );
  OR U12265 ( .A(n11959), .B(n18512), .Z(n11826) );
  NAND U12266 ( .A(n11824), .B(n18513), .Z(n11825) );
  NAND U12267 ( .A(n11826), .B(n11825), .Z(n11916) );
  XNOR U12268 ( .A(b[21]), .B(a[73]), .Z(n11962) );
  NANDN U12269 ( .A(n11962), .B(n19015), .Z(n11829) );
  NAND U12270 ( .A(n19013), .B(n11827), .Z(n11828) );
  NAND U12271 ( .A(n11829), .B(n11828), .Z(n11917) );
  XNOR U12272 ( .A(n11916), .B(n11917), .Z(n11919) );
  XOR U12273 ( .A(n11918), .B(n11919), .Z(n11907) );
  XNOR U12274 ( .A(b[11]), .B(a[83]), .Z(n11965) );
  OR U12275 ( .A(n11965), .B(n18194), .Z(n11832) );
  NANDN U12276 ( .A(n11830), .B(n18104), .Z(n11831) );
  NAND U12277 ( .A(n11832), .B(n11831), .Z(n11905) );
  XOR U12278 ( .A(n580), .B(a[81]), .Z(n11968) );
  NANDN U12279 ( .A(n11968), .B(n18336), .Z(n11835) );
  NANDN U12280 ( .A(n11833), .B(n18337), .Z(n11834) );
  AND U12281 ( .A(n11835), .B(n11834), .Z(n11904) );
  XNOR U12282 ( .A(n11905), .B(n11904), .Z(n11906) );
  XNOR U12283 ( .A(n11907), .B(n11906), .Z(n11923) );
  NANDN U12284 ( .A(n577), .B(a[93]), .Z(n11836) );
  XOR U12285 ( .A(n17151), .B(n11836), .Z(n11838) );
  NANDN U12286 ( .A(b[0]), .B(a[92]), .Z(n11837) );
  AND U12287 ( .A(n11838), .B(n11837), .Z(n11882) );
  NAND U12288 ( .A(n19406), .B(n11839), .Z(n11841) );
  XOR U12289 ( .A(n584), .B(n12055), .Z(n11974) );
  NANDN U12290 ( .A(n576), .B(n11974), .Z(n11840) );
  NAND U12291 ( .A(n11841), .B(n11840), .Z(n11880) );
  NANDN U12292 ( .A(n585), .B(a[61]), .Z(n11881) );
  XNOR U12293 ( .A(n11880), .B(n11881), .Z(n11883) );
  XNOR U12294 ( .A(n11882), .B(n11883), .Z(n11921) );
  XOR U12295 ( .A(b[23]), .B(a[71]), .Z(n11977) );
  NANDN U12296 ( .A(n19127), .B(n11977), .Z(n11844) );
  NAND U12297 ( .A(n11842), .B(n19128), .Z(n11843) );
  NAND U12298 ( .A(n11844), .B(n11843), .Z(n11947) );
  NANDN U12299 ( .A(n11845), .B(n17553), .Z(n11847) );
  XOR U12300 ( .A(b[7]), .B(a[87]), .Z(n11980) );
  NAND U12301 ( .A(n11980), .B(n17555), .Z(n11846) );
  NAND U12302 ( .A(n11847), .B(n11846), .Z(n11944) );
  XOR U12303 ( .A(b[25]), .B(a[69]), .Z(n11983) );
  NAND U12304 ( .A(n11983), .B(n19240), .Z(n11850) );
  NAND U12305 ( .A(n11848), .B(n19242), .Z(n11849) );
  AND U12306 ( .A(n11850), .B(n11849), .Z(n11945) );
  XNOR U12307 ( .A(n11944), .B(n11945), .Z(n11946) );
  XOR U12308 ( .A(n11947), .B(n11946), .Z(n11920) );
  XOR U12309 ( .A(n11923), .B(n11922), .Z(n11935) );
  XOR U12310 ( .A(n11934), .B(n11935), .Z(n11992) );
  XNOR U12311 ( .A(n11993), .B(n11992), .Z(n11995) );
  XNOR U12312 ( .A(n11994), .B(n11995), .Z(n12004) );
  XNOR U12313 ( .A(n12005), .B(n12004), .Z(n12006) );
  XOR U12314 ( .A(n12007), .B(n12006), .Z(n12001) );
  NANDN U12315 ( .A(n11852), .B(n11851), .Z(n11856) );
  NAND U12316 ( .A(n11854), .B(n11853), .Z(n11855) );
  NAND U12317 ( .A(n11856), .B(n11855), .Z(n11998) );
  NAND U12318 ( .A(n11858), .B(n11857), .Z(n11862) );
  NAND U12319 ( .A(n11860), .B(n11859), .Z(n11861) );
  NAND U12320 ( .A(n11862), .B(n11861), .Z(n11999) );
  XNOR U12321 ( .A(n11998), .B(n11999), .Z(n12000) );
  XOR U12322 ( .A(n12001), .B(n12000), .Z(n11877) );
  XOR U12323 ( .A(n11876), .B(n11877), .Z(n11868) );
  XOR U12324 ( .A(n11869), .B(n11868), .Z(n11870) );
  XNOR U12325 ( .A(n11871), .B(n11870), .Z(n12010) );
  XNOR U12326 ( .A(n12010), .B(sreg[189]), .Z(n12012) );
  NAND U12327 ( .A(n11863), .B(sreg[188]), .Z(n11867) );
  OR U12328 ( .A(n11865), .B(n11864), .Z(n11866) );
  AND U12329 ( .A(n11867), .B(n11866), .Z(n12011) );
  XOR U12330 ( .A(n12012), .B(n12011), .Z(c[189]) );
  NAND U12331 ( .A(n11869), .B(n11868), .Z(n11873) );
  NAND U12332 ( .A(n11871), .B(n11870), .Z(n11872) );
  NAND U12333 ( .A(n11873), .B(n11872), .Z(n12018) );
  NANDN U12334 ( .A(n11875), .B(n11874), .Z(n11879) );
  NAND U12335 ( .A(n11877), .B(n11876), .Z(n11878) );
  NAND U12336 ( .A(n11879), .B(n11878), .Z(n12016) );
  NANDN U12337 ( .A(n11881), .B(n11880), .Z(n11885) );
  NAND U12338 ( .A(n11883), .B(n11882), .Z(n11884) );
  NAND U12339 ( .A(n11885), .B(n11884), .Z(n12099) );
  NANDN U12340 ( .A(n11886), .B(n18832), .Z(n11888) );
  XNOR U12341 ( .A(b[19]), .B(a[76]), .Z(n12043) );
  NANDN U12342 ( .A(n12043), .B(n18834), .Z(n11887) );
  NAND U12343 ( .A(n11888), .B(n11887), .Z(n12109) );
  XNOR U12344 ( .A(b[27]), .B(a[68]), .Z(n12046) );
  NANDN U12345 ( .A(n12046), .B(n19336), .Z(n11891) );
  NANDN U12346 ( .A(n11889), .B(n19337), .Z(n11890) );
  NAND U12347 ( .A(n11891), .B(n11890), .Z(n12106) );
  XOR U12348 ( .A(b[5]), .B(a[90]), .Z(n12049) );
  NAND U12349 ( .A(n12049), .B(n17310), .Z(n11894) );
  NAND U12350 ( .A(n11892), .B(n17311), .Z(n11893) );
  AND U12351 ( .A(n11894), .B(n11893), .Z(n12107) );
  XNOR U12352 ( .A(n12106), .B(n12107), .Z(n12108) );
  XNOR U12353 ( .A(n12109), .B(n12108), .Z(n12097) );
  XOR U12354 ( .A(b[17]), .B(a[78]), .Z(n12052) );
  NAND U12355 ( .A(n12052), .B(n18673), .Z(n11897) );
  NAND U12356 ( .A(n11895), .B(n18674), .Z(n11896) );
  NAND U12357 ( .A(n11897), .B(n11896), .Z(n12071) );
  XNOR U12358 ( .A(b[31]), .B(a[64]), .Z(n12056) );
  NANDN U12359 ( .A(n12056), .B(n19472), .Z(n11900) );
  NANDN U12360 ( .A(n11898), .B(n19473), .Z(n11899) );
  NAND U12361 ( .A(n11900), .B(n11899), .Z(n12068) );
  OR U12362 ( .A(n11901), .B(n16988), .Z(n11903) );
  XNOR U12363 ( .A(b[3]), .B(a[92]), .Z(n12059) );
  NANDN U12364 ( .A(n12059), .B(n16990), .Z(n11902) );
  AND U12365 ( .A(n11903), .B(n11902), .Z(n12069) );
  XNOR U12366 ( .A(n12068), .B(n12069), .Z(n12070) );
  XOR U12367 ( .A(n12071), .B(n12070), .Z(n12096) );
  XNOR U12368 ( .A(n12097), .B(n12096), .Z(n12098) );
  XNOR U12369 ( .A(n12099), .B(n12098), .Z(n12034) );
  NANDN U12370 ( .A(n11905), .B(n11904), .Z(n11909) );
  NAND U12371 ( .A(n11907), .B(n11906), .Z(n11908) );
  NAND U12372 ( .A(n11909), .B(n11908), .Z(n12088) );
  NANDN U12373 ( .A(n11911), .B(n11910), .Z(n11915) );
  NAND U12374 ( .A(n11913), .B(n11912), .Z(n11914) );
  NAND U12375 ( .A(n11915), .B(n11914), .Z(n12087) );
  XNOR U12376 ( .A(n12087), .B(n12086), .Z(n12089) );
  XOR U12377 ( .A(n12088), .B(n12089), .Z(n12033) );
  XOR U12378 ( .A(n12034), .B(n12033), .Z(n12035) );
  NANDN U12379 ( .A(n11921), .B(n11920), .Z(n11925) );
  NAND U12380 ( .A(n11923), .B(n11922), .Z(n11924) );
  NAND U12381 ( .A(n11925), .B(n11924), .Z(n12036) );
  XNOR U12382 ( .A(n12035), .B(n12036), .Z(n12150) );
  OR U12383 ( .A(n11927), .B(n11926), .Z(n11931) );
  NANDN U12384 ( .A(n11929), .B(n11928), .Z(n11930) );
  NAND U12385 ( .A(n11931), .B(n11930), .Z(n12149) );
  NANDN U12386 ( .A(n11933), .B(n11932), .Z(n11937) );
  NAND U12387 ( .A(n11935), .B(n11934), .Z(n11936) );
  NAND U12388 ( .A(n11937), .B(n11936), .Z(n12029) );
  NANDN U12389 ( .A(n11939), .B(n11938), .Z(n11943) );
  NAND U12390 ( .A(n11941), .B(n11940), .Z(n11942) );
  NAND U12391 ( .A(n11943), .B(n11942), .Z(n12028) );
  NANDN U12392 ( .A(n11945), .B(n11944), .Z(n11949) );
  NAND U12393 ( .A(n11947), .B(n11946), .Z(n11948) );
  NAND U12394 ( .A(n11949), .B(n11948), .Z(n12090) );
  NANDN U12395 ( .A(n11951), .B(n11950), .Z(n11955) );
  NAND U12396 ( .A(n11953), .B(n11952), .Z(n11954) );
  AND U12397 ( .A(n11955), .B(n11954), .Z(n12091) );
  XNOR U12398 ( .A(n12090), .B(n12091), .Z(n12092) );
  XOR U12399 ( .A(b[9]), .B(n15429), .Z(n12112) );
  NANDN U12400 ( .A(n12112), .B(n17814), .Z(n11958) );
  NANDN U12401 ( .A(n11956), .B(n17815), .Z(n11957) );
  NAND U12402 ( .A(n11958), .B(n11957), .Z(n12082) );
  NANDN U12403 ( .A(n11959), .B(n18513), .Z(n11961) );
  XNOR U12404 ( .A(b[15]), .B(a[80]), .Z(n12115) );
  OR U12405 ( .A(n12115), .B(n18512), .Z(n11960) );
  AND U12406 ( .A(n11961), .B(n11960), .Z(n12080) );
  NANDN U12407 ( .A(n11962), .B(n19013), .Z(n11964) );
  XNOR U12408 ( .A(b[21]), .B(a[74]), .Z(n12118) );
  NANDN U12409 ( .A(n12118), .B(n19015), .Z(n11963) );
  AND U12410 ( .A(n11964), .B(n11963), .Z(n12081) );
  XOR U12411 ( .A(n12082), .B(n12083), .Z(n12077) );
  XOR U12412 ( .A(b[11]), .B(n15134), .Z(n12121) );
  OR U12413 ( .A(n12121), .B(n18194), .Z(n11967) );
  NANDN U12414 ( .A(n11965), .B(n18104), .Z(n11966) );
  NAND U12415 ( .A(n11967), .B(n11966), .Z(n12075) );
  XOR U12416 ( .A(n580), .B(a[82]), .Z(n12124) );
  NANDN U12417 ( .A(n12124), .B(n18336), .Z(n11970) );
  NANDN U12418 ( .A(n11968), .B(n18337), .Z(n11969) );
  AND U12419 ( .A(n11970), .B(n11969), .Z(n12074) );
  XNOR U12420 ( .A(n12075), .B(n12074), .Z(n12076) );
  XOR U12421 ( .A(n12077), .B(n12076), .Z(n12064) );
  NANDN U12422 ( .A(n577), .B(a[94]), .Z(n11971) );
  XOR U12423 ( .A(n17151), .B(n11971), .Z(n11973) );
  NANDN U12424 ( .A(b[0]), .B(a[93]), .Z(n11972) );
  AND U12425 ( .A(n11973), .B(n11972), .Z(n12039) );
  NAND U12426 ( .A(n19406), .B(n11974), .Z(n11976) );
  XNOR U12427 ( .A(n584), .B(a[66]), .Z(n12130) );
  NANDN U12428 ( .A(n576), .B(n12130), .Z(n11975) );
  NAND U12429 ( .A(n11976), .B(n11975), .Z(n12037) );
  NANDN U12430 ( .A(n585), .B(a[62]), .Z(n12038) );
  XNOR U12431 ( .A(n12037), .B(n12038), .Z(n12040) );
  XOR U12432 ( .A(n12039), .B(n12040), .Z(n12062) );
  XOR U12433 ( .A(b[23]), .B(a[72]), .Z(n12133) );
  NANDN U12434 ( .A(n19127), .B(n12133), .Z(n11979) );
  NAND U12435 ( .A(n11977), .B(n19128), .Z(n11978) );
  NAND U12436 ( .A(n11979), .B(n11978), .Z(n12103) );
  NAND U12437 ( .A(n11980), .B(n17553), .Z(n11982) );
  XOR U12438 ( .A(b[7]), .B(a[88]), .Z(n12136) );
  NAND U12439 ( .A(n12136), .B(n17555), .Z(n11981) );
  NAND U12440 ( .A(n11982), .B(n11981), .Z(n12100) );
  XOR U12441 ( .A(b[25]), .B(a[70]), .Z(n12139) );
  NAND U12442 ( .A(n12139), .B(n19240), .Z(n11985) );
  NAND U12443 ( .A(n11983), .B(n19242), .Z(n11984) );
  AND U12444 ( .A(n11985), .B(n11984), .Z(n12101) );
  XNOR U12445 ( .A(n12100), .B(n12101), .Z(n12102) );
  XNOR U12446 ( .A(n12103), .B(n12102), .Z(n12063) );
  XOR U12447 ( .A(n12062), .B(n12063), .Z(n12065) );
  XNOR U12448 ( .A(n12064), .B(n12065), .Z(n12093) );
  XNOR U12449 ( .A(n12092), .B(n12093), .Z(n12027) );
  XNOR U12450 ( .A(n12028), .B(n12027), .Z(n12030) );
  XNOR U12451 ( .A(n12029), .B(n12030), .Z(n12148) );
  XOR U12452 ( .A(n12149), .B(n12148), .Z(n12151) );
  NANDN U12453 ( .A(n11987), .B(n11986), .Z(n11991) );
  NAND U12454 ( .A(n11989), .B(n11988), .Z(n11990) );
  NAND U12455 ( .A(n11991), .B(n11990), .Z(n12143) );
  NAND U12456 ( .A(n11993), .B(n11992), .Z(n11997) );
  NANDN U12457 ( .A(n11995), .B(n11994), .Z(n11996) );
  AND U12458 ( .A(n11997), .B(n11996), .Z(n12142) );
  XNOR U12459 ( .A(n12143), .B(n12142), .Z(n12144) );
  XOR U12460 ( .A(n12145), .B(n12144), .Z(n12023) );
  NANDN U12461 ( .A(n11999), .B(n11998), .Z(n12003) );
  NAND U12462 ( .A(n12001), .B(n12000), .Z(n12002) );
  NAND U12463 ( .A(n12003), .B(n12002), .Z(n12021) );
  NANDN U12464 ( .A(n12005), .B(n12004), .Z(n12009) );
  NANDN U12465 ( .A(n12007), .B(n12006), .Z(n12008) );
  NAND U12466 ( .A(n12009), .B(n12008), .Z(n12022) );
  XNOR U12467 ( .A(n12021), .B(n12022), .Z(n12024) );
  XOR U12468 ( .A(n12023), .B(n12024), .Z(n12015) );
  XOR U12469 ( .A(n12016), .B(n12015), .Z(n12017) );
  XNOR U12470 ( .A(n12018), .B(n12017), .Z(n12154) );
  XNOR U12471 ( .A(n12154), .B(sreg[190]), .Z(n12156) );
  NAND U12472 ( .A(n12010), .B(sreg[189]), .Z(n12014) );
  OR U12473 ( .A(n12012), .B(n12011), .Z(n12013) );
  AND U12474 ( .A(n12014), .B(n12013), .Z(n12155) );
  XOR U12475 ( .A(n12156), .B(n12155), .Z(c[190]) );
  NAND U12476 ( .A(n12016), .B(n12015), .Z(n12020) );
  NAND U12477 ( .A(n12018), .B(n12017), .Z(n12019) );
  NAND U12478 ( .A(n12020), .B(n12019), .Z(n12162) );
  NANDN U12479 ( .A(n12022), .B(n12021), .Z(n12026) );
  NAND U12480 ( .A(n12024), .B(n12023), .Z(n12025) );
  NAND U12481 ( .A(n12026), .B(n12025), .Z(n12159) );
  NAND U12482 ( .A(n12028), .B(n12027), .Z(n12032) );
  NANDN U12483 ( .A(n12030), .B(n12029), .Z(n12031) );
  NAND U12484 ( .A(n12032), .B(n12031), .Z(n12291) );
  XNOR U12485 ( .A(n12291), .B(n12292), .Z(n12293) );
  NANDN U12486 ( .A(n12038), .B(n12037), .Z(n12042) );
  NAND U12487 ( .A(n12040), .B(n12039), .Z(n12041) );
  NAND U12488 ( .A(n12042), .B(n12041), .Z(n12246) );
  NANDN U12489 ( .A(n12043), .B(n18832), .Z(n12045) );
  XNOR U12490 ( .A(b[19]), .B(a[77]), .Z(n12213) );
  NANDN U12491 ( .A(n12213), .B(n18834), .Z(n12044) );
  NAND U12492 ( .A(n12045), .B(n12044), .Z(n12258) );
  XNOR U12493 ( .A(b[27]), .B(a[69]), .Z(n12216) );
  NANDN U12494 ( .A(n12216), .B(n19336), .Z(n12048) );
  NANDN U12495 ( .A(n12046), .B(n19337), .Z(n12047) );
  NAND U12496 ( .A(n12048), .B(n12047), .Z(n12255) );
  XOR U12497 ( .A(b[5]), .B(a[91]), .Z(n12219) );
  NAND U12498 ( .A(n12219), .B(n17310), .Z(n12051) );
  NAND U12499 ( .A(n12049), .B(n17311), .Z(n12050) );
  AND U12500 ( .A(n12051), .B(n12050), .Z(n12256) );
  XNOR U12501 ( .A(n12255), .B(n12256), .Z(n12257) );
  XNOR U12502 ( .A(n12258), .B(n12257), .Z(n12243) );
  XOR U12503 ( .A(b[17]), .B(a[79]), .Z(n12222) );
  NAND U12504 ( .A(n12222), .B(n18673), .Z(n12054) );
  NAND U12505 ( .A(n12052), .B(n18674), .Z(n12053) );
  NAND U12506 ( .A(n12054), .B(n12053), .Z(n12197) );
  XOR U12507 ( .A(b[31]), .B(n12055), .Z(n12225) );
  NANDN U12508 ( .A(n12225), .B(n19472), .Z(n12058) );
  NANDN U12509 ( .A(n12056), .B(n19473), .Z(n12057) );
  AND U12510 ( .A(n12058), .B(n12057), .Z(n12195) );
  OR U12511 ( .A(n12059), .B(n16988), .Z(n12061) );
  XNOR U12512 ( .A(b[3]), .B(a[93]), .Z(n12228) );
  NANDN U12513 ( .A(n12228), .B(n16990), .Z(n12060) );
  AND U12514 ( .A(n12061), .B(n12060), .Z(n12196) );
  XOR U12515 ( .A(n12197), .B(n12198), .Z(n12244) );
  XOR U12516 ( .A(n12243), .B(n12244), .Z(n12245) );
  XNOR U12517 ( .A(n12246), .B(n12245), .Z(n12171) );
  NANDN U12518 ( .A(n12063), .B(n12062), .Z(n12067) );
  OR U12519 ( .A(n12065), .B(n12064), .Z(n12066) );
  NAND U12520 ( .A(n12067), .B(n12066), .Z(n12172) );
  XNOR U12521 ( .A(n12171), .B(n12172), .Z(n12173) );
  NANDN U12522 ( .A(n12069), .B(n12068), .Z(n12073) );
  NAND U12523 ( .A(n12071), .B(n12070), .Z(n12072) );
  NAND U12524 ( .A(n12073), .B(n12072), .Z(n12234) );
  NANDN U12525 ( .A(n12075), .B(n12074), .Z(n12079) );
  NAND U12526 ( .A(n12077), .B(n12076), .Z(n12078) );
  NAND U12527 ( .A(n12079), .B(n12078), .Z(n12231) );
  OR U12528 ( .A(n12081), .B(n12080), .Z(n12085) );
  NANDN U12529 ( .A(n12083), .B(n12082), .Z(n12084) );
  NAND U12530 ( .A(n12085), .B(n12084), .Z(n12232) );
  XNOR U12531 ( .A(n12231), .B(n12232), .Z(n12233) );
  XOR U12532 ( .A(n12234), .B(n12233), .Z(n12174) );
  XNOR U12533 ( .A(n12173), .B(n12174), .Z(n12299) );
  NANDN U12534 ( .A(n12091), .B(n12090), .Z(n12095) );
  NANDN U12535 ( .A(n12093), .B(n12092), .Z(n12094) );
  NAND U12536 ( .A(n12095), .B(n12094), .Z(n12180) );
  NANDN U12537 ( .A(n12101), .B(n12100), .Z(n12105) );
  NAND U12538 ( .A(n12103), .B(n12102), .Z(n12104) );
  NAND U12539 ( .A(n12105), .B(n12104), .Z(n12237) );
  NANDN U12540 ( .A(n12107), .B(n12106), .Z(n12111) );
  NAND U12541 ( .A(n12109), .B(n12108), .Z(n12110) );
  AND U12542 ( .A(n12111), .B(n12110), .Z(n12238) );
  XNOR U12543 ( .A(n12237), .B(n12238), .Z(n12239) );
  XNOR U12544 ( .A(n579), .B(a[87]), .Z(n12267) );
  NAND U12545 ( .A(n17814), .B(n12267), .Z(n12114) );
  NANDN U12546 ( .A(n12112), .B(n17815), .Z(n12113) );
  NAND U12547 ( .A(n12114), .B(n12113), .Z(n12203) );
  NANDN U12548 ( .A(n12115), .B(n18513), .Z(n12117) );
  XOR U12549 ( .A(b[15]), .B(a[81]), .Z(n12264) );
  NANDN U12550 ( .A(n18512), .B(n12264), .Z(n12116) );
  AND U12551 ( .A(n12117), .B(n12116), .Z(n12201) );
  NANDN U12552 ( .A(n12118), .B(n19013), .Z(n12120) );
  XNOR U12553 ( .A(n582), .B(a[75]), .Z(n12261) );
  NAND U12554 ( .A(n12261), .B(n19015), .Z(n12119) );
  AND U12555 ( .A(n12120), .B(n12119), .Z(n12202) );
  XOR U12556 ( .A(n12203), .B(n12204), .Z(n12192) );
  XNOR U12557 ( .A(b[11]), .B(a[85]), .Z(n12270) );
  OR U12558 ( .A(n12270), .B(n18194), .Z(n12123) );
  NANDN U12559 ( .A(n12121), .B(n18104), .Z(n12122) );
  NAND U12560 ( .A(n12123), .B(n12122), .Z(n12190) );
  XOR U12561 ( .A(n580), .B(a[83]), .Z(n12273) );
  NANDN U12562 ( .A(n12273), .B(n18336), .Z(n12126) );
  NANDN U12563 ( .A(n12124), .B(n18337), .Z(n12125) );
  NAND U12564 ( .A(n12126), .B(n12125), .Z(n12189) );
  XOR U12565 ( .A(n12192), .B(n12191), .Z(n12186) );
  NANDN U12566 ( .A(n577), .B(a[95]), .Z(n12127) );
  XOR U12567 ( .A(n17151), .B(n12127), .Z(n12129) );
  IV U12568 ( .A(a[94]), .Z(n16590) );
  NANDN U12569 ( .A(n16590), .B(n577), .Z(n12128) );
  AND U12570 ( .A(n12129), .B(n12128), .Z(n12209) );
  NAND U12571 ( .A(n19406), .B(n12130), .Z(n12132) );
  XNOR U12572 ( .A(n584), .B(a[67]), .Z(n12279) );
  NANDN U12573 ( .A(n576), .B(n12279), .Z(n12131) );
  NAND U12574 ( .A(n12132), .B(n12131), .Z(n12207) );
  NANDN U12575 ( .A(n585), .B(a[63]), .Z(n12208) );
  XNOR U12576 ( .A(n12207), .B(n12208), .Z(n12210) );
  XNOR U12577 ( .A(n12209), .B(n12210), .Z(n12184) );
  XOR U12578 ( .A(b[23]), .B(a[73]), .Z(n12282) );
  NANDN U12579 ( .A(n19127), .B(n12282), .Z(n12135) );
  NAND U12580 ( .A(n12133), .B(n19128), .Z(n12134) );
  NAND U12581 ( .A(n12135), .B(n12134), .Z(n12252) );
  NAND U12582 ( .A(n12136), .B(n17553), .Z(n12138) );
  XOR U12583 ( .A(b[7]), .B(a[89]), .Z(n12285) );
  NAND U12584 ( .A(n12285), .B(n17555), .Z(n12137) );
  NAND U12585 ( .A(n12138), .B(n12137), .Z(n12249) );
  XOR U12586 ( .A(b[25]), .B(a[71]), .Z(n12288) );
  NAND U12587 ( .A(n12288), .B(n19240), .Z(n12141) );
  NAND U12588 ( .A(n12139), .B(n19242), .Z(n12140) );
  AND U12589 ( .A(n12141), .B(n12140), .Z(n12250) );
  XNOR U12590 ( .A(n12249), .B(n12250), .Z(n12251) );
  XOR U12591 ( .A(n12252), .B(n12251), .Z(n12183) );
  XOR U12592 ( .A(n12186), .B(n12185), .Z(n12240) );
  XNOR U12593 ( .A(n12239), .B(n12240), .Z(n12177) );
  XOR U12594 ( .A(n12178), .B(n12177), .Z(n12179) );
  XNOR U12595 ( .A(n12180), .B(n12179), .Z(n12297) );
  XNOR U12596 ( .A(n12298), .B(n12297), .Z(n12300) );
  XNOR U12597 ( .A(n12299), .B(n12300), .Z(n12294) );
  XOR U12598 ( .A(n12293), .B(n12294), .Z(n12168) );
  NANDN U12599 ( .A(n12143), .B(n12142), .Z(n12147) );
  NAND U12600 ( .A(n12145), .B(n12144), .Z(n12146) );
  NAND U12601 ( .A(n12147), .B(n12146), .Z(n12165) );
  NANDN U12602 ( .A(n12149), .B(n12148), .Z(n12153) );
  OR U12603 ( .A(n12151), .B(n12150), .Z(n12152) );
  NAND U12604 ( .A(n12153), .B(n12152), .Z(n12166) );
  XNOR U12605 ( .A(n12165), .B(n12166), .Z(n12167) );
  XNOR U12606 ( .A(n12168), .B(n12167), .Z(n12160) );
  XNOR U12607 ( .A(n12159), .B(n12160), .Z(n12161) );
  XNOR U12608 ( .A(n12162), .B(n12161), .Z(n12303) );
  XNOR U12609 ( .A(n12303), .B(sreg[191]), .Z(n12305) );
  NAND U12610 ( .A(n12154), .B(sreg[190]), .Z(n12158) );
  OR U12611 ( .A(n12156), .B(n12155), .Z(n12157) );
  AND U12612 ( .A(n12158), .B(n12157), .Z(n12304) );
  XOR U12613 ( .A(n12305), .B(n12304), .Z(c[191]) );
  NANDN U12614 ( .A(n12160), .B(n12159), .Z(n12164) );
  NAND U12615 ( .A(n12162), .B(n12161), .Z(n12163) );
  NAND U12616 ( .A(n12164), .B(n12163), .Z(n12311) );
  NANDN U12617 ( .A(n12166), .B(n12165), .Z(n12170) );
  NAND U12618 ( .A(n12168), .B(n12167), .Z(n12169) );
  NAND U12619 ( .A(n12170), .B(n12169), .Z(n12309) );
  NANDN U12620 ( .A(n12172), .B(n12171), .Z(n12176) );
  NANDN U12621 ( .A(n12174), .B(n12173), .Z(n12175) );
  NAND U12622 ( .A(n12176), .B(n12175), .Z(n12442) );
  NAND U12623 ( .A(n12178), .B(n12177), .Z(n12182) );
  NAND U12624 ( .A(n12180), .B(n12179), .Z(n12181) );
  NAND U12625 ( .A(n12182), .B(n12181), .Z(n12443) );
  XNOR U12626 ( .A(n12442), .B(n12443), .Z(n12444) );
  NANDN U12627 ( .A(n12184), .B(n12183), .Z(n12188) );
  NANDN U12628 ( .A(n12186), .B(n12185), .Z(n12187) );
  NAND U12629 ( .A(n12188), .B(n12187), .Z(n12429) );
  OR U12630 ( .A(n12190), .B(n12189), .Z(n12194) );
  NAND U12631 ( .A(n12192), .B(n12191), .Z(n12193) );
  NAND U12632 ( .A(n12194), .B(n12193), .Z(n12368) );
  OR U12633 ( .A(n12196), .B(n12195), .Z(n12200) );
  NANDN U12634 ( .A(n12198), .B(n12197), .Z(n12199) );
  NAND U12635 ( .A(n12200), .B(n12199), .Z(n12367) );
  OR U12636 ( .A(n12202), .B(n12201), .Z(n12206) );
  NANDN U12637 ( .A(n12204), .B(n12203), .Z(n12205) );
  NAND U12638 ( .A(n12206), .B(n12205), .Z(n12366) );
  XOR U12639 ( .A(n12368), .B(n12369), .Z(n12426) );
  NANDN U12640 ( .A(n12208), .B(n12207), .Z(n12212) );
  NAND U12641 ( .A(n12210), .B(n12209), .Z(n12211) );
  NAND U12642 ( .A(n12212), .B(n12211), .Z(n12381) );
  NANDN U12643 ( .A(n12213), .B(n18832), .Z(n12215) );
  XNOR U12644 ( .A(b[19]), .B(a[78]), .Z(n12326) );
  NANDN U12645 ( .A(n12326), .B(n18834), .Z(n12214) );
  NAND U12646 ( .A(n12215), .B(n12214), .Z(n12393) );
  XNOR U12647 ( .A(b[27]), .B(a[70]), .Z(n12329) );
  NANDN U12648 ( .A(n12329), .B(n19336), .Z(n12218) );
  NANDN U12649 ( .A(n12216), .B(n19337), .Z(n12217) );
  NAND U12650 ( .A(n12218), .B(n12217), .Z(n12390) );
  XOR U12651 ( .A(b[5]), .B(a[92]), .Z(n12332) );
  NAND U12652 ( .A(n12332), .B(n17310), .Z(n12221) );
  NAND U12653 ( .A(n12219), .B(n17311), .Z(n12220) );
  AND U12654 ( .A(n12221), .B(n12220), .Z(n12391) );
  XNOR U12655 ( .A(n12390), .B(n12391), .Z(n12392) );
  XNOR U12656 ( .A(n12393), .B(n12392), .Z(n12379) );
  XNOR U12657 ( .A(b[17]), .B(a[80]), .Z(n12335) );
  NANDN U12658 ( .A(n12335), .B(n18673), .Z(n12224) );
  NAND U12659 ( .A(n12222), .B(n18674), .Z(n12223) );
  NAND U12660 ( .A(n12224), .B(n12223), .Z(n12353) );
  XNOR U12661 ( .A(b[31]), .B(a[66]), .Z(n12338) );
  NANDN U12662 ( .A(n12338), .B(n19472), .Z(n12227) );
  NANDN U12663 ( .A(n12225), .B(n19473), .Z(n12226) );
  NAND U12664 ( .A(n12227), .B(n12226), .Z(n12350) );
  OR U12665 ( .A(n12228), .B(n16988), .Z(n12230) );
  XOR U12666 ( .A(b[3]), .B(n16590), .Z(n12341) );
  NANDN U12667 ( .A(n12341), .B(n16990), .Z(n12229) );
  AND U12668 ( .A(n12230), .B(n12229), .Z(n12351) );
  XNOR U12669 ( .A(n12350), .B(n12351), .Z(n12352) );
  XOR U12670 ( .A(n12353), .B(n12352), .Z(n12378) );
  XNOR U12671 ( .A(n12379), .B(n12378), .Z(n12380) );
  XNOR U12672 ( .A(n12381), .B(n12380), .Z(n12427) );
  XNOR U12673 ( .A(n12426), .B(n12427), .Z(n12428) );
  XNOR U12674 ( .A(n12429), .B(n12428), .Z(n12439) );
  NANDN U12675 ( .A(n12232), .B(n12231), .Z(n12236) );
  NANDN U12676 ( .A(n12234), .B(n12233), .Z(n12235) );
  NAND U12677 ( .A(n12236), .B(n12235), .Z(n12436) );
  NANDN U12678 ( .A(n12238), .B(n12237), .Z(n12242) );
  NANDN U12679 ( .A(n12240), .B(n12239), .Z(n12241) );
  NAND U12680 ( .A(n12242), .B(n12241), .Z(n12433) );
  OR U12681 ( .A(n12244), .B(n12243), .Z(n12248) );
  NAND U12682 ( .A(n12246), .B(n12245), .Z(n12247) );
  NAND U12683 ( .A(n12248), .B(n12247), .Z(n12431) );
  NANDN U12684 ( .A(n12250), .B(n12249), .Z(n12254) );
  NAND U12685 ( .A(n12252), .B(n12251), .Z(n12253) );
  NAND U12686 ( .A(n12254), .B(n12253), .Z(n12372) );
  NANDN U12687 ( .A(n12256), .B(n12255), .Z(n12260) );
  NAND U12688 ( .A(n12258), .B(n12257), .Z(n12259) );
  AND U12689 ( .A(n12260), .B(n12259), .Z(n12373) );
  XNOR U12690 ( .A(n12372), .B(n12373), .Z(n12374) );
  XNOR U12691 ( .A(b[21]), .B(a[76]), .Z(n12402) );
  NANDN U12692 ( .A(n12402), .B(n19015), .Z(n12263) );
  NAND U12693 ( .A(n19013), .B(n12261), .Z(n12262) );
  NAND U12694 ( .A(n12263), .B(n12262), .Z(n12362) );
  NAND U12695 ( .A(n12264), .B(n18513), .Z(n12266) );
  XOR U12696 ( .A(b[15]), .B(a[82]), .Z(n12399) );
  NANDN U12697 ( .A(n18512), .B(n12399), .Z(n12265) );
  AND U12698 ( .A(n12266), .B(n12265), .Z(n12363) );
  XNOR U12699 ( .A(n12362), .B(n12363), .Z(n12365) );
  XNOR U12700 ( .A(b[9]), .B(a[88]), .Z(n12396) );
  NANDN U12701 ( .A(n12396), .B(n17814), .Z(n12269) );
  NAND U12702 ( .A(n17815), .B(n12267), .Z(n12268) );
  NAND U12703 ( .A(n12269), .B(n12268), .Z(n12364) );
  XNOR U12704 ( .A(n12365), .B(n12364), .Z(n12358) );
  XOR U12705 ( .A(b[11]), .B(n15429), .Z(n12405) );
  OR U12706 ( .A(n12405), .B(n18194), .Z(n12272) );
  NANDN U12707 ( .A(n12270), .B(n18104), .Z(n12271) );
  NAND U12708 ( .A(n12272), .B(n12271), .Z(n12357) );
  XOR U12709 ( .A(n580), .B(a[84]), .Z(n12408) );
  NANDN U12710 ( .A(n12408), .B(n18336), .Z(n12275) );
  NANDN U12711 ( .A(n12273), .B(n18337), .Z(n12274) );
  NAND U12712 ( .A(n12275), .B(n12274), .Z(n12356) );
  XNOR U12713 ( .A(n12357), .B(n12356), .Z(n12359) );
  XNOR U12714 ( .A(n12358), .B(n12359), .Z(n12347) );
  NANDN U12715 ( .A(n577), .B(a[96]), .Z(n12276) );
  XOR U12716 ( .A(n17151), .B(n12276), .Z(n12278) );
  NANDN U12717 ( .A(b[0]), .B(a[95]), .Z(n12277) );
  AND U12718 ( .A(n12278), .B(n12277), .Z(n12322) );
  NAND U12719 ( .A(n19406), .B(n12279), .Z(n12281) );
  XNOR U12720 ( .A(n584), .B(a[68]), .Z(n12411) );
  NANDN U12721 ( .A(n576), .B(n12411), .Z(n12280) );
  NAND U12722 ( .A(n12281), .B(n12280), .Z(n12320) );
  NANDN U12723 ( .A(n585), .B(a[64]), .Z(n12321) );
  XNOR U12724 ( .A(n12320), .B(n12321), .Z(n12323) );
  XNOR U12725 ( .A(n12322), .B(n12323), .Z(n12345) );
  XOR U12726 ( .A(b[23]), .B(a[74]), .Z(n12417) );
  NANDN U12727 ( .A(n19127), .B(n12417), .Z(n12284) );
  NAND U12728 ( .A(n12282), .B(n19128), .Z(n12283) );
  NAND U12729 ( .A(n12284), .B(n12283), .Z(n12387) );
  NAND U12730 ( .A(n12285), .B(n17553), .Z(n12287) );
  XOR U12731 ( .A(b[7]), .B(a[90]), .Z(n12420) );
  NAND U12732 ( .A(n12420), .B(n17555), .Z(n12286) );
  NAND U12733 ( .A(n12287), .B(n12286), .Z(n12384) );
  XOR U12734 ( .A(b[25]), .B(a[72]), .Z(n12423) );
  NAND U12735 ( .A(n12423), .B(n19240), .Z(n12290) );
  NAND U12736 ( .A(n12288), .B(n19242), .Z(n12289) );
  AND U12737 ( .A(n12290), .B(n12289), .Z(n12385) );
  XNOR U12738 ( .A(n12384), .B(n12385), .Z(n12386) );
  XOR U12739 ( .A(n12387), .B(n12386), .Z(n12344) );
  XOR U12740 ( .A(n12347), .B(n12346), .Z(n12375) );
  XNOR U12741 ( .A(n12374), .B(n12375), .Z(n12430) );
  XOR U12742 ( .A(n12431), .B(n12430), .Z(n12432) );
  XOR U12743 ( .A(n12433), .B(n12432), .Z(n12437) );
  XNOR U12744 ( .A(n12436), .B(n12437), .Z(n12438) );
  XOR U12745 ( .A(n12439), .B(n12438), .Z(n12445) );
  XOR U12746 ( .A(n12444), .B(n12445), .Z(n12316) );
  NANDN U12747 ( .A(n12292), .B(n12291), .Z(n12296) );
  NANDN U12748 ( .A(n12294), .B(n12293), .Z(n12295) );
  NAND U12749 ( .A(n12296), .B(n12295), .Z(n12315) );
  OR U12750 ( .A(n12298), .B(n12297), .Z(n12302) );
  OR U12751 ( .A(n12300), .B(n12299), .Z(n12301) );
  AND U12752 ( .A(n12302), .B(n12301), .Z(n12314) );
  XNOR U12753 ( .A(n12315), .B(n12314), .Z(n12317) );
  XOR U12754 ( .A(n12316), .B(n12317), .Z(n12308) );
  XOR U12755 ( .A(n12309), .B(n12308), .Z(n12310) );
  XNOR U12756 ( .A(n12311), .B(n12310), .Z(n12448) );
  XNOR U12757 ( .A(n12448), .B(sreg[192]), .Z(n12450) );
  NAND U12758 ( .A(n12303), .B(sreg[191]), .Z(n12307) );
  OR U12759 ( .A(n12305), .B(n12304), .Z(n12306) );
  AND U12760 ( .A(n12307), .B(n12306), .Z(n12449) );
  XOR U12761 ( .A(n12450), .B(n12449), .Z(c[192]) );
  NAND U12762 ( .A(n12309), .B(n12308), .Z(n12313) );
  NAND U12763 ( .A(n12311), .B(n12310), .Z(n12312) );
  NAND U12764 ( .A(n12313), .B(n12312), .Z(n12456) );
  NANDN U12765 ( .A(n12315), .B(n12314), .Z(n12319) );
  NAND U12766 ( .A(n12317), .B(n12316), .Z(n12318) );
  NAND U12767 ( .A(n12319), .B(n12318), .Z(n12454) );
  NANDN U12768 ( .A(n12321), .B(n12320), .Z(n12325) );
  NAND U12769 ( .A(n12323), .B(n12322), .Z(n12324) );
  NAND U12770 ( .A(n12325), .B(n12324), .Z(n12478) );
  NANDN U12771 ( .A(n12326), .B(n18832), .Z(n12328) );
  XNOR U12772 ( .A(b[19]), .B(a[79]), .Z(n12527) );
  NANDN U12773 ( .A(n12527), .B(n18834), .Z(n12327) );
  NAND U12774 ( .A(n12328), .B(n12327), .Z(n12488) );
  XNOR U12775 ( .A(b[27]), .B(a[71]), .Z(n12530) );
  NANDN U12776 ( .A(n12530), .B(n19336), .Z(n12331) );
  NANDN U12777 ( .A(n12329), .B(n19337), .Z(n12330) );
  NAND U12778 ( .A(n12331), .B(n12330), .Z(n12485) );
  XOR U12779 ( .A(b[5]), .B(a[93]), .Z(n12533) );
  NAND U12780 ( .A(n12533), .B(n17310), .Z(n12334) );
  NAND U12781 ( .A(n12332), .B(n17311), .Z(n12333) );
  AND U12782 ( .A(n12334), .B(n12333), .Z(n12486) );
  XNOR U12783 ( .A(n12485), .B(n12486), .Z(n12487) );
  XNOR U12784 ( .A(n12488), .B(n12487), .Z(n12476) );
  XOR U12785 ( .A(b[17]), .B(a[81]), .Z(n12536) );
  NAND U12786 ( .A(n12536), .B(n18673), .Z(n12337) );
  NANDN U12787 ( .A(n12335), .B(n18674), .Z(n12336) );
  NAND U12788 ( .A(n12337), .B(n12336), .Z(n12554) );
  XNOR U12789 ( .A(b[31]), .B(a[67]), .Z(n12539) );
  NANDN U12790 ( .A(n12539), .B(n19472), .Z(n12340) );
  NANDN U12791 ( .A(n12338), .B(n19473), .Z(n12339) );
  NAND U12792 ( .A(n12340), .B(n12339), .Z(n12551) );
  OR U12793 ( .A(n12341), .B(n16988), .Z(n12343) );
  XNOR U12794 ( .A(b[3]), .B(a[95]), .Z(n12542) );
  NANDN U12795 ( .A(n12542), .B(n16990), .Z(n12342) );
  AND U12796 ( .A(n12343), .B(n12342), .Z(n12552) );
  XNOR U12797 ( .A(n12551), .B(n12552), .Z(n12553) );
  XOR U12798 ( .A(n12554), .B(n12553), .Z(n12475) );
  XNOR U12799 ( .A(n12476), .B(n12475), .Z(n12477) );
  XNOR U12800 ( .A(n12478), .B(n12477), .Z(n12575) );
  NANDN U12801 ( .A(n12345), .B(n12344), .Z(n12349) );
  NANDN U12802 ( .A(n12347), .B(n12346), .Z(n12348) );
  NAND U12803 ( .A(n12349), .B(n12348), .Z(n12576) );
  XNOR U12804 ( .A(n12575), .B(n12576), .Z(n12577) );
  NANDN U12805 ( .A(n12351), .B(n12350), .Z(n12355) );
  NAND U12806 ( .A(n12353), .B(n12352), .Z(n12354) );
  NAND U12807 ( .A(n12355), .B(n12354), .Z(n12468) );
  OR U12808 ( .A(n12357), .B(n12356), .Z(n12361) );
  NANDN U12809 ( .A(n12359), .B(n12358), .Z(n12360) );
  NAND U12810 ( .A(n12361), .B(n12360), .Z(n12466) );
  XNOR U12811 ( .A(n12466), .B(n12465), .Z(n12467) );
  XOR U12812 ( .A(n12468), .B(n12467), .Z(n12578) );
  XOR U12813 ( .A(n12577), .B(n12578), .Z(n12588) );
  OR U12814 ( .A(n12367), .B(n12366), .Z(n12371) );
  NANDN U12815 ( .A(n12369), .B(n12368), .Z(n12370) );
  NAND U12816 ( .A(n12371), .B(n12370), .Z(n12586) );
  NANDN U12817 ( .A(n12373), .B(n12372), .Z(n12377) );
  NANDN U12818 ( .A(n12375), .B(n12374), .Z(n12376) );
  NAND U12819 ( .A(n12377), .B(n12376), .Z(n12571) );
  NANDN U12820 ( .A(n12379), .B(n12378), .Z(n12383) );
  NAND U12821 ( .A(n12381), .B(n12380), .Z(n12382) );
  NAND U12822 ( .A(n12383), .B(n12382), .Z(n12570) );
  NANDN U12823 ( .A(n12385), .B(n12384), .Z(n12389) );
  NAND U12824 ( .A(n12387), .B(n12386), .Z(n12388) );
  NAND U12825 ( .A(n12389), .B(n12388), .Z(n12469) );
  NANDN U12826 ( .A(n12391), .B(n12390), .Z(n12395) );
  NAND U12827 ( .A(n12393), .B(n12392), .Z(n12394) );
  AND U12828 ( .A(n12395), .B(n12394), .Z(n12470) );
  XNOR U12829 ( .A(n12469), .B(n12470), .Z(n12471) );
  XNOR U12830 ( .A(b[9]), .B(a[89]), .Z(n12491) );
  NANDN U12831 ( .A(n12491), .B(n17814), .Z(n12398) );
  NANDN U12832 ( .A(n12396), .B(n17815), .Z(n12397) );
  NAND U12833 ( .A(n12398), .B(n12397), .Z(n12565) );
  NAND U12834 ( .A(n12399), .B(n18513), .Z(n12401) );
  XOR U12835 ( .A(b[15]), .B(a[83]), .Z(n12494) );
  NANDN U12836 ( .A(n18512), .B(n12494), .Z(n12400) );
  AND U12837 ( .A(n12401), .B(n12400), .Z(n12563) );
  NANDN U12838 ( .A(n12402), .B(n19013), .Z(n12404) );
  XNOR U12839 ( .A(b[21]), .B(a[77]), .Z(n12497) );
  NANDN U12840 ( .A(n12497), .B(n19015), .Z(n12403) );
  AND U12841 ( .A(n12404), .B(n12403), .Z(n12564) );
  XOR U12842 ( .A(n12565), .B(n12566), .Z(n12560) );
  XNOR U12843 ( .A(b[11]), .B(a[87]), .Z(n12500) );
  OR U12844 ( .A(n12500), .B(n18194), .Z(n12407) );
  NANDN U12845 ( .A(n12405), .B(n18104), .Z(n12406) );
  NAND U12846 ( .A(n12407), .B(n12406), .Z(n12558) );
  XOR U12847 ( .A(n580), .B(a[85]), .Z(n12503) );
  NANDN U12848 ( .A(n12503), .B(n18336), .Z(n12410) );
  NANDN U12849 ( .A(n12408), .B(n18337), .Z(n12409) );
  AND U12850 ( .A(n12410), .B(n12409), .Z(n12557) );
  XNOR U12851 ( .A(n12558), .B(n12557), .Z(n12559) );
  XOR U12852 ( .A(n12560), .B(n12559), .Z(n12547) );
  NAND U12853 ( .A(n19406), .B(n12411), .Z(n12413) );
  XNOR U12854 ( .A(n584), .B(a[69]), .Z(n12509) );
  NANDN U12855 ( .A(n576), .B(n12509), .Z(n12412) );
  NAND U12856 ( .A(n12413), .B(n12412), .Z(n12521) );
  NANDN U12857 ( .A(n585), .B(a[65]), .Z(n12522) );
  XNOR U12858 ( .A(n12521), .B(n12522), .Z(n12524) );
  NANDN U12859 ( .A(n577), .B(a[97]), .Z(n12414) );
  XOR U12860 ( .A(n17151), .B(n12414), .Z(n12416) );
  NANDN U12861 ( .A(b[0]), .B(a[96]), .Z(n12415) );
  AND U12862 ( .A(n12416), .B(n12415), .Z(n12523) );
  XOR U12863 ( .A(n12524), .B(n12523), .Z(n12545) );
  XOR U12864 ( .A(b[23]), .B(a[75]), .Z(n12512) );
  NANDN U12865 ( .A(n19127), .B(n12512), .Z(n12419) );
  NAND U12866 ( .A(n12417), .B(n19128), .Z(n12418) );
  NAND U12867 ( .A(n12419), .B(n12418), .Z(n12482) );
  NAND U12868 ( .A(n12420), .B(n17553), .Z(n12422) );
  XOR U12869 ( .A(b[7]), .B(a[91]), .Z(n12515) );
  NAND U12870 ( .A(n12515), .B(n17555), .Z(n12421) );
  NAND U12871 ( .A(n12422), .B(n12421), .Z(n12479) );
  XOR U12872 ( .A(b[25]), .B(a[73]), .Z(n12518) );
  NAND U12873 ( .A(n12518), .B(n19240), .Z(n12425) );
  NAND U12874 ( .A(n12423), .B(n19242), .Z(n12424) );
  AND U12875 ( .A(n12425), .B(n12424), .Z(n12480) );
  XNOR U12876 ( .A(n12479), .B(n12480), .Z(n12481) );
  XNOR U12877 ( .A(n12482), .B(n12481), .Z(n12546) );
  XOR U12878 ( .A(n12545), .B(n12546), .Z(n12548) );
  XNOR U12879 ( .A(n12547), .B(n12548), .Z(n12472) );
  XNOR U12880 ( .A(n12471), .B(n12472), .Z(n12569) );
  XNOR U12881 ( .A(n12570), .B(n12569), .Z(n12572) );
  XNOR U12882 ( .A(n12571), .B(n12572), .Z(n12585) );
  XOR U12883 ( .A(n12586), .B(n12585), .Z(n12587) );
  XNOR U12884 ( .A(n12588), .B(n12587), .Z(n12582) );
  NAND U12885 ( .A(n12431), .B(n12430), .Z(n12435) );
  NAND U12886 ( .A(n12433), .B(n12432), .Z(n12434) );
  AND U12887 ( .A(n12435), .B(n12434), .Z(n12579) );
  XNOR U12888 ( .A(n12580), .B(n12579), .Z(n12581) );
  XOR U12889 ( .A(n12582), .B(n12581), .Z(n12461) );
  NANDN U12890 ( .A(n12437), .B(n12436), .Z(n12441) );
  NAND U12891 ( .A(n12439), .B(n12438), .Z(n12440) );
  NAND U12892 ( .A(n12441), .B(n12440), .Z(n12459) );
  NANDN U12893 ( .A(n12443), .B(n12442), .Z(n12447) );
  NAND U12894 ( .A(n12445), .B(n12444), .Z(n12446) );
  AND U12895 ( .A(n12447), .B(n12446), .Z(n12460) );
  XNOR U12896 ( .A(n12459), .B(n12460), .Z(n12462) );
  XOR U12897 ( .A(n12461), .B(n12462), .Z(n12453) );
  XOR U12898 ( .A(n12454), .B(n12453), .Z(n12455) );
  XNOR U12899 ( .A(n12456), .B(n12455), .Z(n12591) );
  XNOR U12900 ( .A(n12591), .B(sreg[193]), .Z(n12593) );
  NAND U12901 ( .A(n12448), .B(sreg[192]), .Z(n12452) );
  OR U12902 ( .A(n12450), .B(n12449), .Z(n12451) );
  AND U12903 ( .A(n12452), .B(n12451), .Z(n12592) );
  XOR U12904 ( .A(n12593), .B(n12592), .Z(c[193]) );
  NAND U12905 ( .A(n12454), .B(n12453), .Z(n12458) );
  NAND U12906 ( .A(n12456), .B(n12455), .Z(n12457) );
  NAND U12907 ( .A(n12458), .B(n12457), .Z(n12599) );
  NANDN U12908 ( .A(n12460), .B(n12459), .Z(n12464) );
  NAND U12909 ( .A(n12462), .B(n12461), .Z(n12463) );
  NAND U12910 ( .A(n12464), .B(n12463), .Z(n12597) );
  NANDN U12911 ( .A(n12470), .B(n12469), .Z(n12474) );
  NANDN U12912 ( .A(n12472), .B(n12471), .Z(n12473) );
  NAND U12913 ( .A(n12474), .B(n12473), .Z(n12613) );
  NANDN U12914 ( .A(n12480), .B(n12479), .Z(n12484) );
  NAND U12915 ( .A(n12482), .B(n12481), .Z(n12483) );
  NAND U12916 ( .A(n12484), .B(n12483), .Z(n12670) );
  NANDN U12917 ( .A(n12486), .B(n12485), .Z(n12490) );
  NAND U12918 ( .A(n12488), .B(n12487), .Z(n12489) );
  AND U12919 ( .A(n12490), .B(n12489), .Z(n12671) );
  XNOR U12920 ( .A(n12670), .B(n12671), .Z(n12672) );
  XNOR U12921 ( .A(n579), .B(a[90]), .Z(n12694) );
  NAND U12922 ( .A(n17814), .B(n12694), .Z(n12493) );
  NANDN U12923 ( .A(n12491), .B(n17815), .Z(n12492) );
  NAND U12924 ( .A(n12493), .B(n12492), .Z(n12636) );
  NAND U12925 ( .A(n12494), .B(n18513), .Z(n12496) );
  XNOR U12926 ( .A(b[15]), .B(a[84]), .Z(n12697) );
  OR U12927 ( .A(n12697), .B(n18512), .Z(n12495) );
  AND U12928 ( .A(n12496), .B(n12495), .Z(n12634) );
  NANDN U12929 ( .A(n12497), .B(n19013), .Z(n12499) );
  XNOR U12930 ( .A(n582), .B(a[78]), .Z(n12700) );
  NAND U12931 ( .A(n12700), .B(n19015), .Z(n12498) );
  AND U12932 ( .A(n12499), .B(n12498), .Z(n12635) );
  XOR U12933 ( .A(n12636), .B(n12637), .Z(n12625) );
  XNOR U12934 ( .A(b[11]), .B(a[88]), .Z(n12703) );
  OR U12935 ( .A(n12703), .B(n18194), .Z(n12502) );
  NANDN U12936 ( .A(n12500), .B(n18104), .Z(n12501) );
  NAND U12937 ( .A(n12502), .B(n12501), .Z(n12623) );
  XOR U12938 ( .A(n580), .B(a[86]), .Z(n12706) );
  NANDN U12939 ( .A(n12706), .B(n18336), .Z(n12505) );
  NANDN U12940 ( .A(n12503), .B(n18337), .Z(n12504) );
  NAND U12941 ( .A(n12505), .B(n12504), .Z(n12622) );
  XOR U12942 ( .A(n12625), .B(n12624), .Z(n12619) );
  NANDN U12943 ( .A(n577), .B(a[98]), .Z(n12506) );
  XOR U12944 ( .A(n17151), .B(n12506), .Z(n12508) );
  IV U12945 ( .A(a[97]), .Z(n17038) );
  NANDN U12946 ( .A(n17038), .B(n577), .Z(n12507) );
  AND U12947 ( .A(n12508), .B(n12507), .Z(n12642) );
  NAND U12948 ( .A(n19406), .B(n12509), .Z(n12511) );
  XNOR U12949 ( .A(n584), .B(a[70]), .Z(n12709) );
  NANDN U12950 ( .A(n576), .B(n12709), .Z(n12510) );
  NAND U12951 ( .A(n12511), .B(n12510), .Z(n12640) );
  NANDN U12952 ( .A(n585), .B(a[66]), .Z(n12641) );
  XNOR U12953 ( .A(n12640), .B(n12641), .Z(n12643) );
  XNOR U12954 ( .A(n12642), .B(n12643), .Z(n12617) );
  XOR U12955 ( .A(b[23]), .B(a[76]), .Z(n12715) );
  NANDN U12956 ( .A(n19127), .B(n12715), .Z(n12514) );
  NAND U12957 ( .A(n12512), .B(n19128), .Z(n12513) );
  NAND U12958 ( .A(n12514), .B(n12513), .Z(n12685) );
  NAND U12959 ( .A(n12515), .B(n17553), .Z(n12517) );
  XOR U12960 ( .A(b[7]), .B(a[92]), .Z(n12718) );
  NAND U12961 ( .A(n12718), .B(n17555), .Z(n12516) );
  NAND U12962 ( .A(n12517), .B(n12516), .Z(n12682) );
  XOR U12963 ( .A(b[25]), .B(a[74]), .Z(n12721) );
  NAND U12964 ( .A(n12721), .B(n19240), .Z(n12520) );
  NAND U12965 ( .A(n12518), .B(n19242), .Z(n12519) );
  AND U12966 ( .A(n12520), .B(n12519), .Z(n12683) );
  XNOR U12967 ( .A(n12682), .B(n12683), .Z(n12684) );
  XOR U12968 ( .A(n12685), .B(n12684), .Z(n12616) );
  XOR U12969 ( .A(n12619), .B(n12618), .Z(n12673) );
  XNOR U12970 ( .A(n12672), .B(n12673), .Z(n12610) );
  XOR U12971 ( .A(n12611), .B(n12610), .Z(n12612) );
  XOR U12972 ( .A(n12613), .B(n12612), .Z(n12725) );
  XNOR U12973 ( .A(n12724), .B(n12725), .Z(n12727) );
  NANDN U12974 ( .A(n12522), .B(n12521), .Z(n12526) );
  NAND U12975 ( .A(n12524), .B(n12523), .Z(n12525) );
  NAND U12976 ( .A(n12526), .B(n12525), .Z(n12679) );
  NANDN U12977 ( .A(n12527), .B(n18832), .Z(n12529) );
  XOR U12978 ( .A(b[19]), .B(n14551), .Z(n12646) );
  NANDN U12979 ( .A(n12646), .B(n18834), .Z(n12528) );
  NAND U12980 ( .A(n12529), .B(n12528), .Z(n12691) );
  XNOR U12981 ( .A(b[27]), .B(a[72]), .Z(n12649) );
  NANDN U12982 ( .A(n12649), .B(n19336), .Z(n12532) );
  NANDN U12983 ( .A(n12530), .B(n19337), .Z(n12531) );
  NAND U12984 ( .A(n12532), .B(n12531), .Z(n12688) );
  XNOR U12985 ( .A(b[5]), .B(a[94]), .Z(n12652) );
  NANDN U12986 ( .A(n12652), .B(n17310), .Z(n12535) );
  NAND U12987 ( .A(n12533), .B(n17311), .Z(n12534) );
  AND U12988 ( .A(n12535), .B(n12534), .Z(n12689) );
  XNOR U12989 ( .A(n12688), .B(n12689), .Z(n12690) );
  XNOR U12990 ( .A(n12691), .B(n12690), .Z(n12676) );
  XOR U12991 ( .A(b[17]), .B(a[82]), .Z(n12655) );
  NAND U12992 ( .A(n12655), .B(n18673), .Z(n12538) );
  NAND U12993 ( .A(n12536), .B(n18674), .Z(n12537) );
  NAND U12994 ( .A(n12538), .B(n12537), .Z(n12630) );
  XNOR U12995 ( .A(b[31]), .B(a[68]), .Z(n12658) );
  NANDN U12996 ( .A(n12658), .B(n19472), .Z(n12541) );
  NANDN U12997 ( .A(n12539), .B(n19473), .Z(n12540) );
  AND U12998 ( .A(n12541), .B(n12540), .Z(n12628) );
  OR U12999 ( .A(n12542), .B(n16988), .Z(n12544) );
  XNOR U13000 ( .A(b[3]), .B(a[96]), .Z(n12661) );
  NANDN U13001 ( .A(n12661), .B(n16990), .Z(n12543) );
  AND U13002 ( .A(n12544), .B(n12543), .Z(n12629) );
  XOR U13003 ( .A(n12630), .B(n12631), .Z(n12677) );
  XOR U13004 ( .A(n12676), .B(n12677), .Z(n12678) );
  XNOR U13005 ( .A(n12679), .B(n12678), .Z(n12606) );
  NANDN U13006 ( .A(n12546), .B(n12545), .Z(n12550) );
  OR U13007 ( .A(n12548), .B(n12547), .Z(n12549) );
  NAND U13008 ( .A(n12550), .B(n12549), .Z(n12607) );
  XNOR U13009 ( .A(n12606), .B(n12607), .Z(n12608) );
  NANDN U13010 ( .A(n12552), .B(n12551), .Z(n12556) );
  NAND U13011 ( .A(n12554), .B(n12553), .Z(n12555) );
  NAND U13012 ( .A(n12556), .B(n12555), .Z(n12667) );
  NANDN U13013 ( .A(n12558), .B(n12557), .Z(n12562) );
  NAND U13014 ( .A(n12560), .B(n12559), .Z(n12561) );
  NAND U13015 ( .A(n12562), .B(n12561), .Z(n12664) );
  OR U13016 ( .A(n12564), .B(n12563), .Z(n12568) );
  NANDN U13017 ( .A(n12566), .B(n12565), .Z(n12567) );
  NAND U13018 ( .A(n12568), .B(n12567), .Z(n12665) );
  XNOR U13019 ( .A(n12664), .B(n12665), .Z(n12666) );
  XOR U13020 ( .A(n12667), .B(n12666), .Z(n12609) );
  XNOR U13021 ( .A(n12608), .B(n12609), .Z(n12726) );
  XOR U13022 ( .A(n12727), .B(n12726), .Z(n12731) );
  NAND U13023 ( .A(n12570), .B(n12569), .Z(n12574) );
  NANDN U13024 ( .A(n12572), .B(n12571), .Z(n12573) );
  NAND U13025 ( .A(n12574), .B(n12573), .Z(n12728) );
  XNOR U13026 ( .A(n12728), .B(n12729), .Z(n12730) );
  XNOR U13027 ( .A(n12731), .B(n12730), .Z(n12603) );
  NANDN U13028 ( .A(n12580), .B(n12579), .Z(n12584) );
  NAND U13029 ( .A(n12582), .B(n12581), .Z(n12583) );
  NAND U13030 ( .A(n12584), .B(n12583), .Z(n12600) );
  NANDN U13031 ( .A(n12586), .B(n12585), .Z(n12590) );
  OR U13032 ( .A(n12588), .B(n12587), .Z(n12589) );
  NAND U13033 ( .A(n12590), .B(n12589), .Z(n12601) );
  XNOR U13034 ( .A(n12600), .B(n12601), .Z(n12602) );
  XNOR U13035 ( .A(n12603), .B(n12602), .Z(n12596) );
  XOR U13036 ( .A(n12597), .B(n12596), .Z(n12598) );
  XNOR U13037 ( .A(n12599), .B(n12598), .Z(n12734) );
  XNOR U13038 ( .A(n12734), .B(sreg[194]), .Z(n12736) );
  NAND U13039 ( .A(n12591), .B(sreg[193]), .Z(n12595) );
  OR U13040 ( .A(n12593), .B(n12592), .Z(n12594) );
  AND U13041 ( .A(n12595), .B(n12594), .Z(n12735) );
  XOR U13042 ( .A(n12736), .B(n12735), .Z(c[194]) );
  NANDN U13043 ( .A(n12601), .B(n12600), .Z(n12605) );
  NANDN U13044 ( .A(n12603), .B(n12602), .Z(n12604) );
  NAND U13045 ( .A(n12605), .B(n12604), .Z(n12740) );
  NAND U13046 ( .A(n12611), .B(n12610), .Z(n12615) );
  NAND U13047 ( .A(n12613), .B(n12612), .Z(n12614) );
  NAND U13048 ( .A(n12615), .B(n12614), .Z(n12874) );
  XNOR U13049 ( .A(n12873), .B(n12874), .Z(n12875) );
  NANDN U13050 ( .A(n12617), .B(n12616), .Z(n12621) );
  NANDN U13051 ( .A(n12619), .B(n12618), .Z(n12620) );
  NAND U13052 ( .A(n12621), .B(n12620), .Z(n12860) );
  OR U13053 ( .A(n12623), .B(n12622), .Z(n12627) );
  NAND U13054 ( .A(n12625), .B(n12624), .Z(n12626) );
  NAND U13055 ( .A(n12627), .B(n12626), .Z(n12799) );
  OR U13056 ( .A(n12629), .B(n12628), .Z(n12633) );
  NANDN U13057 ( .A(n12631), .B(n12630), .Z(n12632) );
  NAND U13058 ( .A(n12633), .B(n12632), .Z(n12798) );
  OR U13059 ( .A(n12635), .B(n12634), .Z(n12639) );
  NANDN U13060 ( .A(n12637), .B(n12636), .Z(n12638) );
  NAND U13061 ( .A(n12639), .B(n12638), .Z(n12797) );
  XOR U13062 ( .A(n12799), .B(n12800), .Z(n12857) );
  NANDN U13063 ( .A(n12641), .B(n12640), .Z(n12645) );
  NAND U13064 ( .A(n12643), .B(n12642), .Z(n12644) );
  NAND U13065 ( .A(n12645), .B(n12644), .Z(n12812) );
  NANDN U13066 ( .A(n12646), .B(n18832), .Z(n12648) );
  XNOR U13067 ( .A(b[19]), .B(a[81]), .Z(n12757) );
  NANDN U13068 ( .A(n12757), .B(n18834), .Z(n12647) );
  NAND U13069 ( .A(n12648), .B(n12647), .Z(n12824) );
  XNOR U13070 ( .A(b[27]), .B(a[73]), .Z(n12760) );
  NANDN U13071 ( .A(n12760), .B(n19336), .Z(n12651) );
  NANDN U13072 ( .A(n12649), .B(n19337), .Z(n12650) );
  NAND U13073 ( .A(n12651), .B(n12650), .Z(n12821) );
  XOR U13074 ( .A(b[5]), .B(a[95]), .Z(n12763) );
  NAND U13075 ( .A(n12763), .B(n17310), .Z(n12654) );
  NANDN U13076 ( .A(n12652), .B(n17311), .Z(n12653) );
  AND U13077 ( .A(n12654), .B(n12653), .Z(n12822) );
  XNOR U13078 ( .A(n12821), .B(n12822), .Z(n12823) );
  XNOR U13079 ( .A(n12824), .B(n12823), .Z(n12810) );
  XOR U13080 ( .A(b[17]), .B(a[83]), .Z(n12766) );
  NAND U13081 ( .A(n12766), .B(n18673), .Z(n12657) );
  NAND U13082 ( .A(n12655), .B(n18674), .Z(n12656) );
  NAND U13083 ( .A(n12657), .B(n12656), .Z(n12784) );
  XNOR U13084 ( .A(b[31]), .B(a[69]), .Z(n12769) );
  NANDN U13085 ( .A(n12769), .B(n19472), .Z(n12660) );
  NANDN U13086 ( .A(n12658), .B(n19473), .Z(n12659) );
  NAND U13087 ( .A(n12660), .B(n12659), .Z(n12781) );
  OR U13088 ( .A(n12661), .B(n16988), .Z(n12663) );
  XOR U13089 ( .A(b[3]), .B(n17038), .Z(n12772) );
  NANDN U13090 ( .A(n12772), .B(n16990), .Z(n12662) );
  AND U13091 ( .A(n12663), .B(n12662), .Z(n12782) );
  XNOR U13092 ( .A(n12781), .B(n12782), .Z(n12783) );
  XOR U13093 ( .A(n12784), .B(n12783), .Z(n12809) );
  XNOR U13094 ( .A(n12810), .B(n12809), .Z(n12811) );
  XNOR U13095 ( .A(n12812), .B(n12811), .Z(n12858) );
  XNOR U13096 ( .A(n12857), .B(n12858), .Z(n12859) );
  XNOR U13097 ( .A(n12860), .B(n12859), .Z(n12870) );
  NANDN U13098 ( .A(n12665), .B(n12664), .Z(n12669) );
  NANDN U13099 ( .A(n12667), .B(n12666), .Z(n12668) );
  NAND U13100 ( .A(n12669), .B(n12668), .Z(n12867) );
  NANDN U13101 ( .A(n12671), .B(n12670), .Z(n12675) );
  NANDN U13102 ( .A(n12673), .B(n12672), .Z(n12674) );
  NAND U13103 ( .A(n12675), .B(n12674), .Z(n12864) );
  OR U13104 ( .A(n12677), .B(n12676), .Z(n12681) );
  NAND U13105 ( .A(n12679), .B(n12678), .Z(n12680) );
  NAND U13106 ( .A(n12681), .B(n12680), .Z(n12862) );
  NANDN U13107 ( .A(n12683), .B(n12682), .Z(n12687) );
  NAND U13108 ( .A(n12685), .B(n12684), .Z(n12686) );
  NAND U13109 ( .A(n12687), .B(n12686), .Z(n12803) );
  NANDN U13110 ( .A(n12689), .B(n12688), .Z(n12693) );
  NAND U13111 ( .A(n12691), .B(n12690), .Z(n12692) );
  AND U13112 ( .A(n12693), .B(n12692), .Z(n12804) );
  XNOR U13113 ( .A(n12803), .B(n12804), .Z(n12805) );
  XOR U13114 ( .A(n579), .B(a[91]), .Z(n12833) );
  NANDN U13115 ( .A(n12833), .B(n17814), .Z(n12696) );
  NAND U13116 ( .A(n17815), .B(n12694), .Z(n12695) );
  NAND U13117 ( .A(n12696), .B(n12695), .Z(n12789) );
  XNOR U13118 ( .A(b[15]), .B(a[85]), .Z(n12830) );
  OR U13119 ( .A(n12830), .B(n18512), .Z(n12699) );
  NANDN U13120 ( .A(n12697), .B(n18513), .Z(n12698) );
  NAND U13121 ( .A(n12699), .B(n12698), .Z(n12787) );
  XOR U13122 ( .A(n582), .B(a[79]), .Z(n12827) );
  NANDN U13123 ( .A(n12827), .B(n19015), .Z(n12702) );
  NAND U13124 ( .A(n19013), .B(n12700), .Z(n12701) );
  NAND U13125 ( .A(n12702), .B(n12701), .Z(n12788) );
  XNOR U13126 ( .A(n12787), .B(n12788), .Z(n12790) );
  XOR U13127 ( .A(n12789), .B(n12790), .Z(n12778) );
  XNOR U13128 ( .A(b[11]), .B(a[89]), .Z(n12836) );
  OR U13129 ( .A(n12836), .B(n18194), .Z(n12705) );
  NANDN U13130 ( .A(n12703), .B(n18104), .Z(n12704) );
  NAND U13131 ( .A(n12705), .B(n12704), .Z(n12776) );
  XOR U13132 ( .A(n580), .B(a[87]), .Z(n12839) );
  NANDN U13133 ( .A(n12839), .B(n18336), .Z(n12708) );
  NANDN U13134 ( .A(n12706), .B(n18337), .Z(n12707) );
  AND U13135 ( .A(n12708), .B(n12707), .Z(n12775) );
  XNOR U13136 ( .A(n12776), .B(n12775), .Z(n12777) );
  XNOR U13137 ( .A(n12778), .B(n12777), .Z(n12794) );
  NAND U13138 ( .A(n19406), .B(n12709), .Z(n12711) );
  XNOR U13139 ( .A(n584), .B(a[71]), .Z(n12845) );
  NANDN U13140 ( .A(n576), .B(n12845), .Z(n12710) );
  NAND U13141 ( .A(n12711), .B(n12710), .Z(n12751) );
  NANDN U13142 ( .A(n585), .B(a[67]), .Z(n12752) );
  XNOR U13143 ( .A(n12751), .B(n12752), .Z(n12754) );
  NANDN U13144 ( .A(n577), .B(a[99]), .Z(n12712) );
  XOR U13145 ( .A(n17151), .B(n12712), .Z(n12714) );
  NANDN U13146 ( .A(b[0]), .B(a[98]), .Z(n12713) );
  AND U13147 ( .A(n12714), .B(n12713), .Z(n12753) );
  XNOR U13148 ( .A(n12754), .B(n12753), .Z(n12792) );
  XOR U13149 ( .A(b[23]), .B(a[77]), .Z(n12848) );
  NANDN U13150 ( .A(n19127), .B(n12848), .Z(n12717) );
  NAND U13151 ( .A(n12715), .B(n19128), .Z(n12716) );
  NAND U13152 ( .A(n12717), .B(n12716), .Z(n12818) );
  NAND U13153 ( .A(n12718), .B(n17553), .Z(n12720) );
  XOR U13154 ( .A(b[7]), .B(a[93]), .Z(n12851) );
  NAND U13155 ( .A(n12851), .B(n17555), .Z(n12719) );
  NAND U13156 ( .A(n12720), .B(n12719), .Z(n12815) );
  XOR U13157 ( .A(b[25]), .B(a[75]), .Z(n12854) );
  NAND U13158 ( .A(n12854), .B(n19240), .Z(n12723) );
  NAND U13159 ( .A(n12721), .B(n19242), .Z(n12722) );
  AND U13160 ( .A(n12723), .B(n12722), .Z(n12816) );
  XNOR U13161 ( .A(n12815), .B(n12816), .Z(n12817) );
  XOR U13162 ( .A(n12818), .B(n12817), .Z(n12791) );
  XOR U13163 ( .A(n12794), .B(n12793), .Z(n12806) );
  XOR U13164 ( .A(n12805), .B(n12806), .Z(n12861) );
  XOR U13165 ( .A(n12862), .B(n12861), .Z(n12863) );
  XOR U13166 ( .A(n12864), .B(n12863), .Z(n12868) );
  XNOR U13167 ( .A(n12867), .B(n12868), .Z(n12869) );
  XOR U13168 ( .A(n12870), .B(n12869), .Z(n12876) );
  XOR U13169 ( .A(n12875), .B(n12876), .Z(n12747) );
  NANDN U13170 ( .A(n12729), .B(n12728), .Z(n12733) );
  NANDN U13171 ( .A(n12731), .B(n12730), .Z(n12732) );
  NAND U13172 ( .A(n12733), .B(n12732), .Z(n12746) );
  XNOR U13173 ( .A(n12745), .B(n12746), .Z(n12748) );
  XOR U13174 ( .A(n12747), .B(n12748), .Z(n12739) );
  XOR U13175 ( .A(n12740), .B(n12739), .Z(n12741) );
  XNOR U13176 ( .A(n12742), .B(n12741), .Z(n12879) );
  XNOR U13177 ( .A(n12879), .B(sreg[195]), .Z(n12881) );
  NAND U13178 ( .A(n12734), .B(sreg[194]), .Z(n12738) );
  OR U13179 ( .A(n12736), .B(n12735), .Z(n12737) );
  AND U13180 ( .A(n12738), .B(n12737), .Z(n12880) );
  XOR U13181 ( .A(n12881), .B(n12880), .Z(c[195]) );
  NAND U13182 ( .A(n12740), .B(n12739), .Z(n12744) );
  NAND U13183 ( .A(n12742), .B(n12741), .Z(n12743) );
  NAND U13184 ( .A(n12744), .B(n12743), .Z(n12887) );
  NANDN U13185 ( .A(n12746), .B(n12745), .Z(n12750) );
  NAND U13186 ( .A(n12748), .B(n12747), .Z(n12749) );
  NAND U13187 ( .A(n12750), .B(n12749), .Z(n12885) );
  NANDN U13188 ( .A(n12752), .B(n12751), .Z(n12756) );
  NAND U13189 ( .A(n12754), .B(n12753), .Z(n12755) );
  NAND U13190 ( .A(n12756), .B(n12755), .Z(n12965) );
  NANDN U13191 ( .A(n12757), .B(n18832), .Z(n12759) );
  XNOR U13192 ( .A(b[19]), .B(a[82]), .Z(n12912) );
  NANDN U13193 ( .A(n12912), .B(n18834), .Z(n12758) );
  NAND U13194 ( .A(n12759), .B(n12758), .Z(n12975) );
  XNOR U13195 ( .A(b[27]), .B(a[74]), .Z(n12915) );
  NANDN U13196 ( .A(n12915), .B(n19336), .Z(n12762) );
  NANDN U13197 ( .A(n12760), .B(n19337), .Z(n12761) );
  NAND U13198 ( .A(n12762), .B(n12761), .Z(n12972) );
  XOR U13199 ( .A(b[5]), .B(a[96]), .Z(n12918) );
  NAND U13200 ( .A(n12918), .B(n17310), .Z(n12765) );
  NAND U13201 ( .A(n12763), .B(n17311), .Z(n12764) );
  AND U13202 ( .A(n12765), .B(n12764), .Z(n12973) );
  XNOR U13203 ( .A(n12972), .B(n12973), .Z(n12974) );
  XNOR U13204 ( .A(n12975), .B(n12974), .Z(n12963) );
  XNOR U13205 ( .A(b[17]), .B(a[84]), .Z(n12921) );
  NANDN U13206 ( .A(n12921), .B(n18673), .Z(n12768) );
  NAND U13207 ( .A(n12766), .B(n18674), .Z(n12767) );
  NAND U13208 ( .A(n12768), .B(n12767), .Z(n12939) );
  XNOR U13209 ( .A(b[31]), .B(a[70]), .Z(n12924) );
  NANDN U13210 ( .A(n12924), .B(n19472), .Z(n12771) );
  NANDN U13211 ( .A(n12769), .B(n19473), .Z(n12770) );
  NAND U13212 ( .A(n12771), .B(n12770), .Z(n12936) );
  OR U13213 ( .A(n12772), .B(n16988), .Z(n12774) );
  XNOR U13214 ( .A(b[3]), .B(a[98]), .Z(n12927) );
  NANDN U13215 ( .A(n12927), .B(n16990), .Z(n12773) );
  AND U13216 ( .A(n12774), .B(n12773), .Z(n12937) );
  XNOR U13217 ( .A(n12936), .B(n12937), .Z(n12938) );
  XOR U13218 ( .A(n12939), .B(n12938), .Z(n12962) );
  XNOR U13219 ( .A(n12963), .B(n12962), .Z(n12964) );
  XNOR U13220 ( .A(n12965), .B(n12964), .Z(n12903) );
  NANDN U13221 ( .A(n12776), .B(n12775), .Z(n12780) );
  NAND U13222 ( .A(n12778), .B(n12777), .Z(n12779) );
  NAND U13223 ( .A(n12780), .B(n12779), .Z(n12954) );
  NANDN U13224 ( .A(n12782), .B(n12781), .Z(n12786) );
  NAND U13225 ( .A(n12784), .B(n12783), .Z(n12785) );
  NAND U13226 ( .A(n12786), .B(n12785), .Z(n12953) );
  XNOR U13227 ( .A(n12953), .B(n12952), .Z(n12955) );
  XOR U13228 ( .A(n12954), .B(n12955), .Z(n12902) );
  XOR U13229 ( .A(n12903), .B(n12902), .Z(n12904) );
  NANDN U13230 ( .A(n12792), .B(n12791), .Z(n12796) );
  NAND U13231 ( .A(n12794), .B(n12793), .Z(n12795) );
  NAND U13232 ( .A(n12796), .B(n12795), .Z(n12905) );
  XNOR U13233 ( .A(n12904), .B(n12905), .Z(n13016) );
  OR U13234 ( .A(n12798), .B(n12797), .Z(n12802) );
  NANDN U13235 ( .A(n12800), .B(n12799), .Z(n12801) );
  NAND U13236 ( .A(n12802), .B(n12801), .Z(n13015) );
  NANDN U13237 ( .A(n12804), .B(n12803), .Z(n12808) );
  NAND U13238 ( .A(n12806), .B(n12805), .Z(n12807) );
  NAND U13239 ( .A(n12808), .B(n12807), .Z(n12898) );
  NANDN U13240 ( .A(n12810), .B(n12809), .Z(n12814) );
  NAND U13241 ( .A(n12812), .B(n12811), .Z(n12813) );
  NAND U13242 ( .A(n12814), .B(n12813), .Z(n12897) );
  NANDN U13243 ( .A(n12816), .B(n12815), .Z(n12820) );
  NAND U13244 ( .A(n12818), .B(n12817), .Z(n12819) );
  NAND U13245 ( .A(n12820), .B(n12819), .Z(n12956) );
  NANDN U13246 ( .A(n12822), .B(n12821), .Z(n12826) );
  NAND U13247 ( .A(n12824), .B(n12823), .Z(n12825) );
  AND U13248 ( .A(n12826), .B(n12825), .Z(n12957) );
  XNOR U13249 ( .A(n12956), .B(n12957), .Z(n12958) );
  XOR U13250 ( .A(n582), .B(a[80]), .Z(n12984) );
  NANDN U13251 ( .A(n12984), .B(n19015), .Z(n12829) );
  NANDN U13252 ( .A(n12827), .B(n19013), .Z(n12828) );
  NAND U13253 ( .A(n12829), .B(n12828), .Z(n12948) );
  NANDN U13254 ( .A(n12830), .B(n18513), .Z(n12832) );
  XNOR U13255 ( .A(b[15]), .B(a[86]), .Z(n12981) );
  OR U13256 ( .A(n12981), .B(n18512), .Z(n12831) );
  AND U13257 ( .A(n12832), .B(n12831), .Z(n12949) );
  XNOR U13258 ( .A(n12948), .B(n12949), .Z(n12951) );
  XOR U13259 ( .A(n579), .B(a[92]), .Z(n12978) );
  NANDN U13260 ( .A(n12978), .B(n17814), .Z(n12835) );
  NANDN U13261 ( .A(n12833), .B(n17815), .Z(n12834) );
  NAND U13262 ( .A(n12835), .B(n12834), .Z(n12950) );
  XNOR U13263 ( .A(n12951), .B(n12950), .Z(n12944) );
  XNOR U13264 ( .A(b[11]), .B(a[90]), .Z(n12987) );
  OR U13265 ( .A(n12987), .B(n18194), .Z(n12838) );
  NANDN U13266 ( .A(n12836), .B(n18104), .Z(n12837) );
  NAND U13267 ( .A(n12838), .B(n12837), .Z(n12943) );
  XOR U13268 ( .A(n580), .B(a[88]), .Z(n12990) );
  NANDN U13269 ( .A(n12990), .B(n18336), .Z(n12841) );
  NANDN U13270 ( .A(n12839), .B(n18337), .Z(n12840) );
  NAND U13271 ( .A(n12841), .B(n12840), .Z(n12942) );
  XNOR U13272 ( .A(n12943), .B(n12942), .Z(n12945) );
  XNOR U13273 ( .A(n12944), .B(n12945), .Z(n12933) );
  NANDN U13274 ( .A(n577), .B(a[100]), .Z(n12842) );
  XOR U13275 ( .A(n17151), .B(n12842), .Z(n12844) );
  NANDN U13276 ( .A(b[0]), .B(a[99]), .Z(n12843) );
  AND U13277 ( .A(n12844), .B(n12843), .Z(n12908) );
  NAND U13278 ( .A(n19406), .B(n12845), .Z(n12847) );
  XNOR U13279 ( .A(n584), .B(a[72]), .Z(n12996) );
  NANDN U13280 ( .A(n576), .B(n12996), .Z(n12846) );
  NAND U13281 ( .A(n12847), .B(n12846), .Z(n12906) );
  NANDN U13282 ( .A(n585), .B(a[68]), .Z(n12907) );
  XNOR U13283 ( .A(n12906), .B(n12907), .Z(n12909) );
  XNOR U13284 ( .A(n12908), .B(n12909), .Z(n12931) );
  XOR U13285 ( .A(b[23]), .B(a[78]), .Z(n12999) );
  NANDN U13286 ( .A(n19127), .B(n12999), .Z(n12850) );
  NAND U13287 ( .A(n12848), .B(n19128), .Z(n12849) );
  NAND U13288 ( .A(n12850), .B(n12849), .Z(n12969) );
  NAND U13289 ( .A(n12851), .B(n17553), .Z(n12853) );
  XNOR U13290 ( .A(b[7]), .B(a[94]), .Z(n13002) );
  NANDN U13291 ( .A(n13002), .B(n17555), .Z(n12852) );
  NAND U13292 ( .A(n12853), .B(n12852), .Z(n12966) );
  XOR U13293 ( .A(b[25]), .B(a[76]), .Z(n13005) );
  NAND U13294 ( .A(n13005), .B(n19240), .Z(n12856) );
  NAND U13295 ( .A(n12854), .B(n19242), .Z(n12855) );
  AND U13296 ( .A(n12856), .B(n12855), .Z(n12967) );
  XNOR U13297 ( .A(n12966), .B(n12967), .Z(n12968) );
  XOR U13298 ( .A(n12969), .B(n12968), .Z(n12930) );
  XOR U13299 ( .A(n12933), .B(n12932), .Z(n12959) );
  XNOR U13300 ( .A(n12958), .B(n12959), .Z(n12896) );
  XNOR U13301 ( .A(n12897), .B(n12896), .Z(n12899) );
  XNOR U13302 ( .A(n12898), .B(n12899), .Z(n13014) );
  XOR U13303 ( .A(n13015), .B(n13014), .Z(n13017) );
  NAND U13304 ( .A(n12862), .B(n12861), .Z(n12866) );
  NAND U13305 ( .A(n12864), .B(n12863), .Z(n12865) );
  AND U13306 ( .A(n12866), .B(n12865), .Z(n13008) );
  XNOR U13307 ( .A(n13009), .B(n13008), .Z(n13010) );
  XOR U13308 ( .A(n13011), .B(n13010), .Z(n12892) );
  NANDN U13309 ( .A(n12868), .B(n12867), .Z(n12872) );
  NAND U13310 ( .A(n12870), .B(n12869), .Z(n12871) );
  NAND U13311 ( .A(n12872), .B(n12871), .Z(n12890) );
  NANDN U13312 ( .A(n12874), .B(n12873), .Z(n12878) );
  NAND U13313 ( .A(n12876), .B(n12875), .Z(n12877) );
  AND U13314 ( .A(n12878), .B(n12877), .Z(n12891) );
  XNOR U13315 ( .A(n12890), .B(n12891), .Z(n12893) );
  XOR U13316 ( .A(n12892), .B(n12893), .Z(n12884) );
  XOR U13317 ( .A(n12885), .B(n12884), .Z(n12886) );
  XNOR U13318 ( .A(n12887), .B(n12886), .Z(n13020) );
  XNOR U13319 ( .A(n13020), .B(sreg[196]), .Z(n13022) );
  NAND U13320 ( .A(n12879), .B(sreg[195]), .Z(n12883) );
  OR U13321 ( .A(n12881), .B(n12880), .Z(n12882) );
  AND U13322 ( .A(n12883), .B(n12882), .Z(n13021) );
  XOR U13323 ( .A(n13022), .B(n13021), .Z(c[196]) );
  NAND U13324 ( .A(n12885), .B(n12884), .Z(n12889) );
  NAND U13325 ( .A(n12887), .B(n12886), .Z(n12888) );
  NAND U13326 ( .A(n12889), .B(n12888), .Z(n13028) );
  NANDN U13327 ( .A(n12891), .B(n12890), .Z(n12895) );
  NAND U13328 ( .A(n12893), .B(n12892), .Z(n12894) );
  NAND U13329 ( .A(n12895), .B(n12894), .Z(n13025) );
  NAND U13330 ( .A(n12897), .B(n12896), .Z(n12901) );
  NANDN U13331 ( .A(n12899), .B(n12898), .Z(n12900) );
  NAND U13332 ( .A(n12901), .B(n12900), .Z(n13151) );
  XNOR U13333 ( .A(n13151), .B(n13152), .Z(n13153) );
  NANDN U13334 ( .A(n12907), .B(n12906), .Z(n12911) );
  NAND U13335 ( .A(n12909), .B(n12908), .Z(n12910) );
  NAND U13336 ( .A(n12911), .B(n12910), .Z(n13096) );
  NANDN U13337 ( .A(n12912), .B(n18832), .Z(n12914) );
  XNOR U13338 ( .A(b[19]), .B(a[83]), .Z(n13043) );
  NANDN U13339 ( .A(n13043), .B(n18834), .Z(n12913) );
  NAND U13340 ( .A(n12914), .B(n12913), .Z(n13106) );
  XNOR U13341 ( .A(b[27]), .B(a[75]), .Z(n13046) );
  NANDN U13342 ( .A(n13046), .B(n19336), .Z(n12917) );
  NANDN U13343 ( .A(n12915), .B(n19337), .Z(n12916) );
  NAND U13344 ( .A(n12917), .B(n12916), .Z(n13103) );
  XNOR U13345 ( .A(b[5]), .B(a[97]), .Z(n13049) );
  NANDN U13346 ( .A(n13049), .B(n17310), .Z(n12920) );
  NAND U13347 ( .A(n12918), .B(n17311), .Z(n12919) );
  AND U13348 ( .A(n12920), .B(n12919), .Z(n13104) );
  XNOR U13349 ( .A(n13103), .B(n13104), .Z(n13105) );
  XNOR U13350 ( .A(n13106), .B(n13105), .Z(n13094) );
  XOR U13351 ( .A(b[17]), .B(a[85]), .Z(n13052) );
  NAND U13352 ( .A(n13052), .B(n18673), .Z(n12923) );
  NANDN U13353 ( .A(n12921), .B(n18674), .Z(n12922) );
  NAND U13354 ( .A(n12923), .B(n12922), .Z(n13070) );
  XNOR U13355 ( .A(b[31]), .B(a[71]), .Z(n13055) );
  NANDN U13356 ( .A(n13055), .B(n19472), .Z(n12926) );
  NANDN U13357 ( .A(n12924), .B(n19473), .Z(n12925) );
  NAND U13358 ( .A(n12926), .B(n12925), .Z(n13067) );
  OR U13359 ( .A(n12927), .B(n16988), .Z(n12929) );
  XNOR U13360 ( .A(b[3]), .B(a[99]), .Z(n13058) );
  NANDN U13361 ( .A(n13058), .B(n16990), .Z(n12928) );
  AND U13362 ( .A(n12929), .B(n12928), .Z(n13068) );
  XNOR U13363 ( .A(n13067), .B(n13068), .Z(n13069) );
  XOR U13364 ( .A(n13070), .B(n13069), .Z(n13093) );
  XNOR U13365 ( .A(n13094), .B(n13093), .Z(n13095) );
  XNOR U13366 ( .A(n13096), .B(n13095), .Z(n13145) );
  NANDN U13367 ( .A(n12931), .B(n12930), .Z(n12935) );
  NANDN U13368 ( .A(n12933), .B(n12932), .Z(n12934) );
  NAND U13369 ( .A(n12935), .B(n12934), .Z(n13146) );
  XNOR U13370 ( .A(n13145), .B(n13146), .Z(n13147) );
  NANDN U13371 ( .A(n12937), .B(n12936), .Z(n12941) );
  NAND U13372 ( .A(n12939), .B(n12938), .Z(n12940) );
  NAND U13373 ( .A(n12941), .B(n12940), .Z(n13086) );
  OR U13374 ( .A(n12943), .B(n12942), .Z(n12947) );
  NANDN U13375 ( .A(n12945), .B(n12944), .Z(n12946) );
  NAND U13376 ( .A(n12947), .B(n12946), .Z(n13084) );
  XNOR U13377 ( .A(n13084), .B(n13083), .Z(n13085) );
  XOR U13378 ( .A(n13086), .B(n13085), .Z(n13148) );
  XOR U13379 ( .A(n13147), .B(n13148), .Z(n13159) );
  NANDN U13380 ( .A(n12957), .B(n12956), .Z(n12961) );
  NANDN U13381 ( .A(n12959), .B(n12958), .Z(n12960) );
  NAND U13382 ( .A(n12961), .B(n12960), .Z(n13142) );
  NANDN U13383 ( .A(n12967), .B(n12966), .Z(n12971) );
  NAND U13384 ( .A(n12969), .B(n12968), .Z(n12970) );
  NAND U13385 ( .A(n12971), .B(n12970), .Z(n13087) );
  NANDN U13386 ( .A(n12973), .B(n12972), .Z(n12977) );
  NAND U13387 ( .A(n12975), .B(n12974), .Z(n12976) );
  AND U13388 ( .A(n12977), .B(n12976), .Z(n13088) );
  XNOR U13389 ( .A(n13087), .B(n13088), .Z(n13089) );
  XNOR U13390 ( .A(b[9]), .B(a[93]), .Z(n13109) );
  NANDN U13391 ( .A(n13109), .B(n17814), .Z(n12980) );
  NANDN U13392 ( .A(n12978), .B(n17815), .Z(n12979) );
  NAND U13393 ( .A(n12980), .B(n12979), .Z(n13075) );
  XNOR U13394 ( .A(b[15]), .B(a[87]), .Z(n13112) );
  OR U13395 ( .A(n13112), .B(n18512), .Z(n12983) );
  NANDN U13396 ( .A(n12981), .B(n18513), .Z(n12982) );
  NAND U13397 ( .A(n12983), .B(n12982), .Z(n13073) );
  XNOR U13398 ( .A(b[21]), .B(a[81]), .Z(n13115) );
  NANDN U13399 ( .A(n13115), .B(n19015), .Z(n12986) );
  NANDN U13400 ( .A(n12984), .B(n19013), .Z(n12985) );
  NAND U13401 ( .A(n12986), .B(n12985), .Z(n13074) );
  XNOR U13402 ( .A(n13073), .B(n13074), .Z(n13076) );
  XOR U13403 ( .A(n13075), .B(n13076), .Z(n13064) );
  XNOR U13404 ( .A(b[11]), .B(a[91]), .Z(n13118) );
  OR U13405 ( .A(n13118), .B(n18194), .Z(n12989) );
  NANDN U13406 ( .A(n12987), .B(n18104), .Z(n12988) );
  NAND U13407 ( .A(n12989), .B(n12988), .Z(n13062) );
  XOR U13408 ( .A(n580), .B(a[89]), .Z(n13121) );
  NANDN U13409 ( .A(n13121), .B(n18336), .Z(n12992) );
  NANDN U13410 ( .A(n12990), .B(n18337), .Z(n12991) );
  AND U13411 ( .A(n12992), .B(n12991), .Z(n13061) );
  XNOR U13412 ( .A(n13062), .B(n13061), .Z(n13063) );
  XNOR U13413 ( .A(n13064), .B(n13063), .Z(n13080) );
  NANDN U13414 ( .A(n577), .B(a[101]), .Z(n12993) );
  XOR U13415 ( .A(n17151), .B(n12993), .Z(n12995) );
  IV U13416 ( .A(a[100]), .Z(n17447) );
  NANDN U13417 ( .A(n17447), .B(n577), .Z(n12994) );
  AND U13418 ( .A(n12995), .B(n12994), .Z(n13039) );
  NAND U13419 ( .A(n19406), .B(n12996), .Z(n12998) );
  XNOR U13420 ( .A(n584), .B(a[73]), .Z(n13127) );
  NANDN U13421 ( .A(n576), .B(n13127), .Z(n12997) );
  NAND U13422 ( .A(n12998), .B(n12997), .Z(n13037) );
  NANDN U13423 ( .A(n585), .B(a[69]), .Z(n13038) );
  XNOR U13424 ( .A(n13037), .B(n13038), .Z(n13040) );
  XNOR U13425 ( .A(n13039), .B(n13040), .Z(n13078) );
  XOR U13426 ( .A(b[23]), .B(a[79]), .Z(n13130) );
  NANDN U13427 ( .A(n19127), .B(n13130), .Z(n13001) );
  NAND U13428 ( .A(n12999), .B(n19128), .Z(n13000) );
  NAND U13429 ( .A(n13001), .B(n13000), .Z(n13100) );
  NANDN U13430 ( .A(n13002), .B(n17553), .Z(n13004) );
  XOR U13431 ( .A(b[7]), .B(a[95]), .Z(n13133) );
  NAND U13432 ( .A(n13133), .B(n17555), .Z(n13003) );
  NAND U13433 ( .A(n13004), .B(n13003), .Z(n13097) );
  XOR U13434 ( .A(b[25]), .B(a[77]), .Z(n13136) );
  NAND U13435 ( .A(n13136), .B(n19240), .Z(n13007) );
  NAND U13436 ( .A(n13005), .B(n19242), .Z(n13006) );
  AND U13437 ( .A(n13007), .B(n13006), .Z(n13098) );
  XNOR U13438 ( .A(n13097), .B(n13098), .Z(n13099) );
  XOR U13439 ( .A(n13100), .B(n13099), .Z(n13077) );
  XOR U13440 ( .A(n13080), .B(n13079), .Z(n13090) );
  XOR U13441 ( .A(n13089), .B(n13090), .Z(n13139) );
  XOR U13442 ( .A(n13140), .B(n13139), .Z(n13141) );
  XNOR U13443 ( .A(n13142), .B(n13141), .Z(n13157) );
  XNOR U13444 ( .A(n13158), .B(n13157), .Z(n13160) );
  XNOR U13445 ( .A(n13159), .B(n13160), .Z(n13154) );
  XOR U13446 ( .A(n13153), .B(n13154), .Z(n13034) );
  NANDN U13447 ( .A(n13009), .B(n13008), .Z(n13013) );
  NAND U13448 ( .A(n13011), .B(n13010), .Z(n13012) );
  NAND U13449 ( .A(n13013), .B(n13012), .Z(n13031) );
  NANDN U13450 ( .A(n13015), .B(n13014), .Z(n13019) );
  OR U13451 ( .A(n13017), .B(n13016), .Z(n13018) );
  NAND U13452 ( .A(n13019), .B(n13018), .Z(n13032) );
  XNOR U13453 ( .A(n13031), .B(n13032), .Z(n13033) );
  XNOR U13454 ( .A(n13034), .B(n13033), .Z(n13026) );
  XNOR U13455 ( .A(n13025), .B(n13026), .Z(n13027) );
  XNOR U13456 ( .A(n13028), .B(n13027), .Z(n13163) );
  XNOR U13457 ( .A(n13163), .B(sreg[197]), .Z(n13165) );
  NAND U13458 ( .A(n13020), .B(sreg[196]), .Z(n13024) );
  OR U13459 ( .A(n13022), .B(n13021), .Z(n13023) );
  AND U13460 ( .A(n13024), .B(n13023), .Z(n13164) );
  XOR U13461 ( .A(n13165), .B(n13164), .Z(c[197]) );
  NANDN U13462 ( .A(n13026), .B(n13025), .Z(n13030) );
  NAND U13463 ( .A(n13028), .B(n13027), .Z(n13029) );
  NAND U13464 ( .A(n13030), .B(n13029), .Z(n13171) );
  NANDN U13465 ( .A(n13032), .B(n13031), .Z(n13036) );
  NAND U13466 ( .A(n13034), .B(n13033), .Z(n13035) );
  NAND U13467 ( .A(n13036), .B(n13035), .Z(n13169) );
  NANDN U13468 ( .A(n13038), .B(n13037), .Z(n13042) );
  NAND U13469 ( .A(n13040), .B(n13039), .Z(n13041) );
  NAND U13470 ( .A(n13042), .B(n13041), .Z(n13249) );
  NANDN U13471 ( .A(n13043), .B(n18832), .Z(n13045) );
  XOR U13472 ( .A(b[19]), .B(n15134), .Z(n13194) );
  NANDN U13473 ( .A(n13194), .B(n18834), .Z(n13044) );
  NAND U13474 ( .A(n13045), .B(n13044), .Z(n13259) );
  XNOR U13475 ( .A(b[27]), .B(a[76]), .Z(n13197) );
  NANDN U13476 ( .A(n13197), .B(n19336), .Z(n13048) );
  NANDN U13477 ( .A(n13046), .B(n19337), .Z(n13047) );
  NAND U13478 ( .A(n13048), .B(n13047), .Z(n13256) );
  XOR U13479 ( .A(b[5]), .B(a[98]), .Z(n13200) );
  NAND U13480 ( .A(n13200), .B(n17310), .Z(n13051) );
  NANDN U13481 ( .A(n13049), .B(n17311), .Z(n13050) );
  AND U13482 ( .A(n13051), .B(n13050), .Z(n13257) );
  XNOR U13483 ( .A(n13256), .B(n13257), .Z(n13258) );
  XNOR U13484 ( .A(n13259), .B(n13258), .Z(n13247) );
  XNOR U13485 ( .A(b[17]), .B(a[86]), .Z(n13203) );
  NANDN U13486 ( .A(n13203), .B(n18673), .Z(n13054) );
  NAND U13487 ( .A(n13052), .B(n18674), .Z(n13053) );
  NAND U13488 ( .A(n13054), .B(n13053), .Z(n13221) );
  XNOR U13489 ( .A(b[31]), .B(a[72]), .Z(n13206) );
  NANDN U13490 ( .A(n13206), .B(n19472), .Z(n13057) );
  NANDN U13491 ( .A(n13055), .B(n19473), .Z(n13056) );
  NAND U13492 ( .A(n13057), .B(n13056), .Z(n13218) );
  OR U13493 ( .A(n13058), .B(n16988), .Z(n13060) );
  XOR U13494 ( .A(b[3]), .B(n17447), .Z(n13209) );
  NANDN U13495 ( .A(n13209), .B(n16990), .Z(n13059) );
  AND U13496 ( .A(n13060), .B(n13059), .Z(n13219) );
  XNOR U13497 ( .A(n13218), .B(n13219), .Z(n13220) );
  XOR U13498 ( .A(n13221), .B(n13220), .Z(n13246) );
  XNOR U13499 ( .A(n13247), .B(n13246), .Z(n13248) );
  XNOR U13500 ( .A(n13249), .B(n13248), .Z(n13185) );
  NANDN U13501 ( .A(n13062), .B(n13061), .Z(n13066) );
  NAND U13502 ( .A(n13064), .B(n13063), .Z(n13065) );
  NAND U13503 ( .A(n13066), .B(n13065), .Z(n13238) );
  NANDN U13504 ( .A(n13068), .B(n13067), .Z(n13072) );
  NAND U13505 ( .A(n13070), .B(n13069), .Z(n13071) );
  NAND U13506 ( .A(n13072), .B(n13071), .Z(n13237) );
  XNOR U13507 ( .A(n13237), .B(n13236), .Z(n13239) );
  XOR U13508 ( .A(n13238), .B(n13239), .Z(n13184) );
  XOR U13509 ( .A(n13185), .B(n13184), .Z(n13186) );
  NANDN U13510 ( .A(n13078), .B(n13077), .Z(n13082) );
  NAND U13511 ( .A(n13080), .B(n13079), .Z(n13081) );
  AND U13512 ( .A(n13082), .B(n13081), .Z(n13187) );
  XNOR U13513 ( .A(n13186), .B(n13187), .Z(n13295) );
  NANDN U13514 ( .A(n13088), .B(n13087), .Z(n13092) );
  NAND U13515 ( .A(n13090), .B(n13089), .Z(n13091) );
  NAND U13516 ( .A(n13092), .B(n13091), .Z(n13181) );
  NANDN U13517 ( .A(n13098), .B(n13097), .Z(n13102) );
  NAND U13518 ( .A(n13100), .B(n13099), .Z(n13101) );
  NAND U13519 ( .A(n13102), .B(n13101), .Z(n13240) );
  NANDN U13520 ( .A(n13104), .B(n13103), .Z(n13108) );
  NAND U13521 ( .A(n13106), .B(n13105), .Z(n13107) );
  AND U13522 ( .A(n13108), .B(n13107), .Z(n13241) );
  XNOR U13523 ( .A(n13240), .B(n13241), .Z(n13242) );
  XOR U13524 ( .A(n579), .B(n16590), .Z(n13262) );
  NAND U13525 ( .A(n17814), .B(n13262), .Z(n13111) );
  NANDN U13526 ( .A(n13109), .B(n17815), .Z(n13110) );
  NAND U13527 ( .A(n13111), .B(n13110), .Z(n13226) );
  NANDN U13528 ( .A(n13112), .B(n18513), .Z(n13114) );
  XOR U13529 ( .A(b[15]), .B(a[88]), .Z(n13265) );
  NANDN U13530 ( .A(n18512), .B(n13265), .Z(n13113) );
  AND U13531 ( .A(n13114), .B(n13113), .Z(n13224) );
  NANDN U13532 ( .A(n13115), .B(n19013), .Z(n13117) );
  XNOR U13533 ( .A(n582), .B(a[82]), .Z(n13268) );
  NAND U13534 ( .A(n13268), .B(n19015), .Z(n13116) );
  AND U13535 ( .A(n13117), .B(n13116), .Z(n13225) );
  XOR U13536 ( .A(n13226), .B(n13227), .Z(n13215) );
  XNOR U13537 ( .A(b[11]), .B(a[92]), .Z(n13271) );
  OR U13538 ( .A(n13271), .B(n18194), .Z(n13120) );
  NANDN U13539 ( .A(n13118), .B(n18104), .Z(n13119) );
  NAND U13540 ( .A(n13120), .B(n13119), .Z(n13213) );
  XOR U13541 ( .A(n580), .B(a[90]), .Z(n13274) );
  NANDN U13542 ( .A(n13274), .B(n18336), .Z(n13123) );
  NANDN U13543 ( .A(n13121), .B(n18337), .Z(n13122) );
  AND U13544 ( .A(n13123), .B(n13122), .Z(n13212) );
  XNOR U13545 ( .A(n13213), .B(n13212), .Z(n13214) );
  XOR U13546 ( .A(n13215), .B(n13214), .Z(n13232) );
  NANDN U13547 ( .A(n577), .B(a[102]), .Z(n13124) );
  XOR U13548 ( .A(n17151), .B(n13124), .Z(n13126) );
  NANDN U13549 ( .A(b[0]), .B(a[101]), .Z(n13125) );
  AND U13550 ( .A(n13126), .B(n13125), .Z(n13190) );
  NAND U13551 ( .A(n19406), .B(n13127), .Z(n13129) );
  XNOR U13552 ( .A(n584), .B(a[74]), .Z(n13280) );
  NANDN U13553 ( .A(n576), .B(n13280), .Z(n13128) );
  NAND U13554 ( .A(n13129), .B(n13128), .Z(n13188) );
  NANDN U13555 ( .A(n585), .B(a[70]), .Z(n13189) );
  XNOR U13556 ( .A(n13188), .B(n13189), .Z(n13191) );
  XOR U13557 ( .A(n13190), .B(n13191), .Z(n13230) );
  XNOR U13558 ( .A(b[23]), .B(a[80]), .Z(n13283) );
  OR U13559 ( .A(n13283), .B(n19127), .Z(n13132) );
  NAND U13560 ( .A(n13130), .B(n19128), .Z(n13131) );
  NAND U13561 ( .A(n13132), .B(n13131), .Z(n13253) );
  NAND U13562 ( .A(n13133), .B(n17553), .Z(n13135) );
  XOR U13563 ( .A(b[7]), .B(a[96]), .Z(n13286) );
  NAND U13564 ( .A(n13286), .B(n17555), .Z(n13134) );
  NAND U13565 ( .A(n13135), .B(n13134), .Z(n13250) );
  XOR U13566 ( .A(b[25]), .B(a[78]), .Z(n13289) );
  NAND U13567 ( .A(n13289), .B(n19240), .Z(n13138) );
  NAND U13568 ( .A(n13136), .B(n19242), .Z(n13137) );
  AND U13569 ( .A(n13138), .B(n13137), .Z(n13251) );
  XNOR U13570 ( .A(n13250), .B(n13251), .Z(n13252) );
  XNOR U13571 ( .A(n13253), .B(n13252), .Z(n13231) );
  XOR U13572 ( .A(n13230), .B(n13231), .Z(n13233) );
  XNOR U13573 ( .A(n13232), .B(n13233), .Z(n13243) );
  XOR U13574 ( .A(n13242), .B(n13243), .Z(n13179) );
  XNOR U13575 ( .A(n13178), .B(n13179), .Z(n13180) );
  XOR U13576 ( .A(n13181), .B(n13180), .Z(n13293) );
  XNOR U13577 ( .A(n13292), .B(n13293), .Z(n13294) );
  XNOR U13578 ( .A(n13295), .B(n13294), .Z(n13299) );
  NAND U13579 ( .A(n13140), .B(n13139), .Z(n13144) );
  NAND U13580 ( .A(n13142), .B(n13141), .Z(n13143) );
  NAND U13581 ( .A(n13144), .B(n13143), .Z(n13296) );
  NANDN U13582 ( .A(n13146), .B(n13145), .Z(n13150) );
  NAND U13583 ( .A(n13148), .B(n13147), .Z(n13149) );
  NAND U13584 ( .A(n13150), .B(n13149), .Z(n13297) );
  XNOR U13585 ( .A(n13296), .B(n13297), .Z(n13298) );
  XNOR U13586 ( .A(n13299), .B(n13298), .Z(n13175) );
  NANDN U13587 ( .A(n13152), .B(n13151), .Z(n13156) );
  NANDN U13588 ( .A(n13154), .B(n13153), .Z(n13155) );
  NAND U13589 ( .A(n13156), .B(n13155), .Z(n13173) );
  OR U13590 ( .A(n13158), .B(n13157), .Z(n13162) );
  OR U13591 ( .A(n13160), .B(n13159), .Z(n13161) );
  AND U13592 ( .A(n13162), .B(n13161), .Z(n13172) );
  XNOR U13593 ( .A(n13173), .B(n13172), .Z(n13174) );
  XNOR U13594 ( .A(n13175), .B(n13174), .Z(n13168) );
  XOR U13595 ( .A(n13169), .B(n13168), .Z(n13170) );
  XNOR U13596 ( .A(n13171), .B(n13170), .Z(n13302) );
  XNOR U13597 ( .A(n13302), .B(sreg[198]), .Z(n13304) );
  NAND U13598 ( .A(n13163), .B(sreg[197]), .Z(n13167) );
  OR U13599 ( .A(n13165), .B(n13164), .Z(n13166) );
  AND U13600 ( .A(n13167), .B(n13166), .Z(n13303) );
  XOR U13601 ( .A(n13304), .B(n13303), .Z(c[198]) );
  NANDN U13602 ( .A(n13173), .B(n13172), .Z(n13177) );
  NANDN U13603 ( .A(n13175), .B(n13174), .Z(n13176) );
  NAND U13604 ( .A(n13177), .B(n13176), .Z(n13307) );
  NANDN U13605 ( .A(n13179), .B(n13178), .Z(n13183) );
  NAND U13606 ( .A(n13181), .B(n13180), .Z(n13182) );
  NAND U13607 ( .A(n13183), .B(n13182), .Z(n13319) );
  XNOR U13608 ( .A(n13319), .B(n13320), .Z(n13321) );
  NANDN U13609 ( .A(n13189), .B(n13188), .Z(n13193) );
  NAND U13610 ( .A(n13191), .B(n13190), .Z(n13192) );
  NAND U13611 ( .A(n13193), .B(n13192), .Z(n13392) );
  NANDN U13612 ( .A(n13194), .B(n18832), .Z(n13196) );
  XNOR U13613 ( .A(b[19]), .B(a[85]), .Z(n13337) );
  NANDN U13614 ( .A(n13337), .B(n18834), .Z(n13195) );
  NAND U13615 ( .A(n13196), .B(n13195), .Z(n13402) );
  XNOR U13616 ( .A(b[27]), .B(a[77]), .Z(n13340) );
  NANDN U13617 ( .A(n13340), .B(n19336), .Z(n13199) );
  NANDN U13618 ( .A(n13197), .B(n19337), .Z(n13198) );
  NAND U13619 ( .A(n13199), .B(n13198), .Z(n13399) );
  XOR U13620 ( .A(b[5]), .B(a[99]), .Z(n13343) );
  NAND U13621 ( .A(n13343), .B(n17310), .Z(n13202) );
  NAND U13622 ( .A(n13200), .B(n17311), .Z(n13201) );
  AND U13623 ( .A(n13202), .B(n13201), .Z(n13400) );
  XNOR U13624 ( .A(n13399), .B(n13400), .Z(n13401) );
  XNOR U13625 ( .A(n13402), .B(n13401), .Z(n13390) );
  XOR U13626 ( .A(b[17]), .B(a[87]), .Z(n13346) );
  NAND U13627 ( .A(n13346), .B(n18673), .Z(n13205) );
  NANDN U13628 ( .A(n13203), .B(n18674), .Z(n13204) );
  NAND U13629 ( .A(n13205), .B(n13204), .Z(n13364) );
  XNOR U13630 ( .A(b[31]), .B(a[73]), .Z(n13349) );
  NANDN U13631 ( .A(n13349), .B(n19472), .Z(n13208) );
  NANDN U13632 ( .A(n13206), .B(n19473), .Z(n13207) );
  NAND U13633 ( .A(n13208), .B(n13207), .Z(n13361) );
  OR U13634 ( .A(n13209), .B(n16988), .Z(n13211) );
  XNOR U13635 ( .A(b[3]), .B(a[101]), .Z(n13352) );
  NANDN U13636 ( .A(n13352), .B(n16990), .Z(n13210) );
  AND U13637 ( .A(n13211), .B(n13210), .Z(n13362) );
  XNOR U13638 ( .A(n13361), .B(n13362), .Z(n13363) );
  XOR U13639 ( .A(n13364), .B(n13363), .Z(n13389) );
  XNOR U13640 ( .A(n13390), .B(n13389), .Z(n13391) );
  XNOR U13641 ( .A(n13392), .B(n13391), .Z(n13435) );
  NANDN U13642 ( .A(n13213), .B(n13212), .Z(n13217) );
  NAND U13643 ( .A(n13215), .B(n13214), .Z(n13216) );
  NAND U13644 ( .A(n13217), .B(n13216), .Z(n13380) );
  NANDN U13645 ( .A(n13219), .B(n13218), .Z(n13223) );
  NAND U13646 ( .A(n13221), .B(n13220), .Z(n13222) );
  NAND U13647 ( .A(n13223), .B(n13222), .Z(n13378) );
  OR U13648 ( .A(n13225), .B(n13224), .Z(n13229) );
  NANDN U13649 ( .A(n13227), .B(n13226), .Z(n13228) );
  NAND U13650 ( .A(n13229), .B(n13228), .Z(n13377) );
  XNOR U13651 ( .A(n13380), .B(n13379), .Z(n13436) );
  XNOR U13652 ( .A(n13435), .B(n13436), .Z(n13437) );
  NANDN U13653 ( .A(n13231), .B(n13230), .Z(n13235) );
  OR U13654 ( .A(n13233), .B(n13232), .Z(n13234) );
  AND U13655 ( .A(n13235), .B(n13234), .Z(n13438) );
  XOR U13656 ( .A(n13437), .B(n13438), .Z(n13327) );
  NANDN U13657 ( .A(n13241), .B(n13240), .Z(n13245) );
  NANDN U13658 ( .A(n13243), .B(n13242), .Z(n13244) );
  NAND U13659 ( .A(n13245), .B(n13244), .Z(n13444) );
  NANDN U13660 ( .A(n13251), .B(n13250), .Z(n13255) );
  NAND U13661 ( .A(n13253), .B(n13252), .Z(n13254) );
  NAND U13662 ( .A(n13255), .B(n13254), .Z(n13383) );
  NANDN U13663 ( .A(n13257), .B(n13256), .Z(n13261) );
  NAND U13664 ( .A(n13259), .B(n13258), .Z(n13260) );
  AND U13665 ( .A(n13261), .B(n13260), .Z(n13384) );
  XNOR U13666 ( .A(n13383), .B(n13384), .Z(n13385) );
  XNOR U13667 ( .A(b[9]), .B(a[95]), .Z(n13405) );
  NANDN U13668 ( .A(n13405), .B(n17814), .Z(n13264) );
  NAND U13669 ( .A(n17815), .B(n13262), .Z(n13263) );
  NAND U13670 ( .A(n13264), .B(n13263), .Z(n13369) );
  XNOR U13671 ( .A(b[15]), .B(a[89]), .Z(n13408) );
  OR U13672 ( .A(n13408), .B(n18512), .Z(n13267) );
  NAND U13673 ( .A(n13265), .B(n18513), .Z(n13266) );
  NAND U13674 ( .A(n13267), .B(n13266), .Z(n13367) );
  XNOR U13675 ( .A(b[21]), .B(a[83]), .Z(n13411) );
  NANDN U13676 ( .A(n13411), .B(n19015), .Z(n13270) );
  NAND U13677 ( .A(n19013), .B(n13268), .Z(n13269) );
  NAND U13678 ( .A(n13270), .B(n13269), .Z(n13368) );
  XNOR U13679 ( .A(n13367), .B(n13368), .Z(n13370) );
  XOR U13680 ( .A(n13369), .B(n13370), .Z(n13358) );
  XNOR U13681 ( .A(b[11]), .B(a[93]), .Z(n13414) );
  OR U13682 ( .A(n13414), .B(n18194), .Z(n13273) );
  NANDN U13683 ( .A(n13271), .B(n18104), .Z(n13272) );
  NAND U13684 ( .A(n13273), .B(n13272), .Z(n13356) );
  XOR U13685 ( .A(n580), .B(a[91]), .Z(n13417) );
  NANDN U13686 ( .A(n13417), .B(n18336), .Z(n13276) );
  NANDN U13687 ( .A(n13274), .B(n18337), .Z(n13275) );
  AND U13688 ( .A(n13276), .B(n13275), .Z(n13355) );
  XNOR U13689 ( .A(n13356), .B(n13355), .Z(n13357) );
  XNOR U13690 ( .A(n13358), .B(n13357), .Z(n13374) );
  NANDN U13691 ( .A(n577), .B(a[103]), .Z(n13277) );
  XOR U13692 ( .A(n17151), .B(n13277), .Z(n13279) );
  IV U13693 ( .A(a[102]), .Z(n17208) );
  NANDN U13694 ( .A(n17208), .B(n577), .Z(n13278) );
  AND U13695 ( .A(n13279), .B(n13278), .Z(n13333) );
  NAND U13696 ( .A(n19406), .B(n13280), .Z(n13282) );
  XNOR U13697 ( .A(n584), .B(a[75]), .Z(n13423) );
  NANDN U13698 ( .A(n576), .B(n13423), .Z(n13281) );
  NAND U13699 ( .A(n13282), .B(n13281), .Z(n13331) );
  NANDN U13700 ( .A(n585), .B(a[71]), .Z(n13332) );
  XNOR U13701 ( .A(n13331), .B(n13332), .Z(n13334) );
  XNOR U13702 ( .A(n13333), .B(n13334), .Z(n13372) );
  XOR U13703 ( .A(b[23]), .B(a[81]), .Z(n13426) );
  NANDN U13704 ( .A(n19127), .B(n13426), .Z(n13285) );
  NANDN U13705 ( .A(n13283), .B(n19128), .Z(n13284) );
  NAND U13706 ( .A(n13285), .B(n13284), .Z(n13396) );
  NAND U13707 ( .A(n13286), .B(n17553), .Z(n13288) );
  XNOR U13708 ( .A(b[7]), .B(a[97]), .Z(n13429) );
  NANDN U13709 ( .A(n13429), .B(n17555), .Z(n13287) );
  NAND U13710 ( .A(n13288), .B(n13287), .Z(n13393) );
  XOR U13711 ( .A(b[25]), .B(a[79]), .Z(n13432) );
  NAND U13712 ( .A(n13432), .B(n19240), .Z(n13291) );
  NAND U13713 ( .A(n13289), .B(n19242), .Z(n13290) );
  AND U13714 ( .A(n13291), .B(n13290), .Z(n13394) );
  XNOR U13715 ( .A(n13393), .B(n13394), .Z(n13395) );
  XOR U13716 ( .A(n13396), .B(n13395), .Z(n13371) );
  XOR U13717 ( .A(n13374), .B(n13373), .Z(n13386) );
  XOR U13718 ( .A(n13385), .B(n13386), .Z(n13441) );
  XOR U13719 ( .A(n13442), .B(n13441), .Z(n13443) );
  XNOR U13720 ( .A(n13444), .B(n13443), .Z(n13325) );
  XNOR U13721 ( .A(n13326), .B(n13325), .Z(n13328) );
  XNOR U13722 ( .A(n13327), .B(n13328), .Z(n13322) );
  XOR U13723 ( .A(n13321), .B(n13322), .Z(n13316) );
  NANDN U13724 ( .A(n13297), .B(n13296), .Z(n13301) );
  NANDN U13725 ( .A(n13299), .B(n13298), .Z(n13300) );
  NAND U13726 ( .A(n13301), .B(n13300), .Z(n13314) );
  XNOR U13727 ( .A(n13313), .B(n13314), .Z(n13315) );
  XNOR U13728 ( .A(n13316), .B(n13315), .Z(n13308) );
  XNOR U13729 ( .A(n13307), .B(n13308), .Z(n13309) );
  XNOR U13730 ( .A(n13310), .B(n13309), .Z(n13447) );
  XNOR U13731 ( .A(n13447), .B(sreg[199]), .Z(n13449) );
  NAND U13732 ( .A(n13302), .B(sreg[198]), .Z(n13306) );
  OR U13733 ( .A(n13304), .B(n13303), .Z(n13305) );
  AND U13734 ( .A(n13306), .B(n13305), .Z(n13448) );
  XOR U13735 ( .A(n13449), .B(n13448), .Z(c[199]) );
  NANDN U13736 ( .A(n13308), .B(n13307), .Z(n13312) );
  NAND U13737 ( .A(n13310), .B(n13309), .Z(n13311) );
  NAND U13738 ( .A(n13312), .B(n13311), .Z(n13455) );
  NANDN U13739 ( .A(n13314), .B(n13313), .Z(n13318) );
  NAND U13740 ( .A(n13316), .B(n13315), .Z(n13317) );
  NAND U13741 ( .A(n13318), .B(n13317), .Z(n13453) );
  NANDN U13742 ( .A(n13320), .B(n13319), .Z(n13324) );
  NANDN U13743 ( .A(n13322), .B(n13321), .Z(n13323) );
  NAND U13744 ( .A(n13324), .B(n13323), .Z(n13459) );
  OR U13745 ( .A(n13326), .B(n13325), .Z(n13330) );
  OR U13746 ( .A(n13328), .B(n13327), .Z(n13329) );
  AND U13747 ( .A(n13330), .B(n13329), .Z(n13458) );
  XNOR U13748 ( .A(n13459), .B(n13458), .Z(n13460) );
  NANDN U13749 ( .A(n13332), .B(n13331), .Z(n13336) );
  NAND U13750 ( .A(n13334), .B(n13333), .Z(n13335) );
  NAND U13751 ( .A(n13336), .B(n13335), .Z(n13535) );
  NANDN U13752 ( .A(n13337), .B(n18832), .Z(n13339) );
  XOR U13753 ( .A(b[19]), .B(n15429), .Z(n13480) );
  NANDN U13754 ( .A(n13480), .B(n18834), .Z(n13338) );
  NAND U13755 ( .A(n13339), .B(n13338), .Z(n13545) );
  XNOR U13756 ( .A(b[27]), .B(a[78]), .Z(n13483) );
  NANDN U13757 ( .A(n13483), .B(n19336), .Z(n13342) );
  NANDN U13758 ( .A(n13340), .B(n19337), .Z(n13341) );
  NAND U13759 ( .A(n13342), .B(n13341), .Z(n13542) );
  XNOR U13760 ( .A(b[5]), .B(a[100]), .Z(n13486) );
  NANDN U13761 ( .A(n13486), .B(n17310), .Z(n13345) );
  NAND U13762 ( .A(n13343), .B(n17311), .Z(n13344) );
  AND U13763 ( .A(n13345), .B(n13344), .Z(n13543) );
  XNOR U13764 ( .A(n13542), .B(n13543), .Z(n13544) );
  XNOR U13765 ( .A(n13545), .B(n13544), .Z(n13533) );
  XOR U13766 ( .A(b[17]), .B(a[88]), .Z(n13489) );
  NAND U13767 ( .A(n13489), .B(n18673), .Z(n13348) );
  NAND U13768 ( .A(n13346), .B(n18674), .Z(n13347) );
  NAND U13769 ( .A(n13348), .B(n13347), .Z(n13507) );
  XNOR U13770 ( .A(b[31]), .B(a[74]), .Z(n13492) );
  NANDN U13771 ( .A(n13492), .B(n19472), .Z(n13351) );
  NANDN U13772 ( .A(n13349), .B(n19473), .Z(n13350) );
  NAND U13773 ( .A(n13351), .B(n13350), .Z(n13504) );
  OR U13774 ( .A(n13352), .B(n16988), .Z(n13354) );
  XOR U13775 ( .A(a[102]), .B(n578), .Z(n13495) );
  NANDN U13776 ( .A(n13495), .B(n16990), .Z(n13353) );
  AND U13777 ( .A(n13354), .B(n13353), .Z(n13505) );
  XNOR U13778 ( .A(n13504), .B(n13505), .Z(n13506) );
  XOR U13779 ( .A(n13507), .B(n13506), .Z(n13532) );
  XNOR U13780 ( .A(n13533), .B(n13532), .Z(n13534) );
  XNOR U13781 ( .A(n13535), .B(n13534), .Z(n13471) );
  NANDN U13782 ( .A(n13356), .B(n13355), .Z(n13360) );
  NAND U13783 ( .A(n13358), .B(n13357), .Z(n13359) );
  NAND U13784 ( .A(n13360), .B(n13359), .Z(n13524) );
  NANDN U13785 ( .A(n13362), .B(n13361), .Z(n13366) );
  NAND U13786 ( .A(n13364), .B(n13363), .Z(n13365) );
  NAND U13787 ( .A(n13366), .B(n13365), .Z(n13523) );
  XNOR U13788 ( .A(n13523), .B(n13522), .Z(n13525) );
  XOR U13789 ( .A(n13524), .B(n13525), .Z(n13470) );
  XOR U13790 ( .A(n13471), .B(n13470), .Z(n13472) );
  NANDN U13791 ( .A(n13372), .B(n13371), .Z(n13376) );
  NAND U13792 ( .A(n13374), .B(n13373), .Z(n13375) );
  NAND U13793 ( .A(n13376), .B(n13375), .Z(n13473) );
  XNOR U13794 ( .A(n13472), .B(n13473), .Z(n13586) );
  OR U13795 ( .A(n13378), .B(n13377), .Z(n13382) );
  NAND U13796 ( .A(n13380), .B(n13379), .Z(n13381) );
  NAND U13797 ( .A(n13382), .B(n13381), .Z(n13585) );
  NANDN U13798 ( .A(n13384), .B(n13383), .Z(n13388) );
  NAND U13799 ( .A(n13386), .B(n13385), .Z(n13387) );
  NAND U13800 ( .A(n13388), .B(n13387), .Z(n13466) );
  NANDN U13801 ( .A(n13394), .B(n13393), .Z(n13398) );
  NAND U13802 ( .A(n13396), .B(n13395), .Z(n13397) );
  NAND U13803 ( .A(n13398), .B(n13397), .Z(n13526) );
  NANDN U13804 ( .A(n13400), .B(n13399), .Z(n13404) );
  NAND U13805 ( .A(n13402), .B(n13401), .Z(n13403) );
  AND U13806 ( .A(n13404), .B(n13403), .Z(n13527) );
  XNOR U13807 ( .A(n13526), .B(n13527), .Z(n13528) );
  XNOR U13808 ( .A(b[9]), .B(a[96]), .Z(n13548) );
  NANDN U13809 ( .A(n13548), .B(n17814), .Z(n13407) );
  NANDN U13810 ( .A(n13405), .B(n17815), .Z(n13406) );
  NAND U13811 ( .A(n13407), .B(n13406), .Z(n13512) );
  NANDN U13812 ( .A(n13408), .B(n18513), .Z(n13410) );
  XOR U13813 ( .A(b[15]), .B(a[90]), .Z(n13551) );
  NANDN U13814 ( .A(n18512), .B(n13551), .Z(n13409) );
  AND U13815 ( .A(n13410), .B(n13409), .Z(n13510) );
  NANDN U13816 ( .A(n13411), .B(n19013), .Z(n13413) );
  XOR U13817 ( .A(b[21]), .B(n15134), .Z(n13554) );
  NANDN U13818 ( .A(n13554), .B(n19015), .Z(n13412) );
  AND U13819 ( .A(n13413), .B(n13412), .Z(n13511) );
  XOR U13820 ( .A(n13512), .B(n13513), .Z(n13501) );
  XOR U13821 ( .A(b[11]), .B(n16590), .Z(n13557) );
  OR U13822 ( .A(n13557), .B(n18194), .Z(n13416) );
  NANDN U13823 ( .A(n13414), .B(n18104), .Z(n13415) );
  NAND U13824 ( .A(n13416), .B(n13415), .Z(n13499) );
  XOR U13825 ( .A(n580), .B(a[92]), .Z(n13560) );
  NANDN U13826 ( .A(n13560), .B(n18336), .Z(n13419) );
  NANDN U13827 ( .A(n13417), .B(n18337), .Z(n13418) );
  AND U13828 ( .A(n13419), .B(n13418), .Z(n13498) );
  XNOR U13829 ( .A(n13499), .B(n13498), .Z(n13500) );
  XOR U13830 ( .A(n13501), .B(n13500), .Z(n13518) );
  NANDN U13831 ( .A(n577), .B(a[104]), .Z(n13420) );
  XOR U13832 ( .A(n17151), .B(n13420), .Z(n13422) );
  NANDN U13833 ( .A(b[0]), .B(a[103]), .Z(n13421) );
  AND U13834 ( .A(n13422), .B(n13421), .Z(n13476) );
  NAND U13835 ( .A(n19406), .B(n13423), .Z(n13425) );
  XNOR U13836 ( .A(n584), .B(a[76]), .Z(n13563) );
  NANDN U13837 ( .A(n576), .B(n13563), .Z(n13424) );
  NAND U13838 ( .A(n13425), .B(n13424), .Z(n13474) );
  NANDN U13839 ( .A(n585), .B(a[72]), .Z(n13475) );
  XNOR U13840 ( .A(n13474), .B(n13475), .Z(n13477) );
  XOR U13841 ( .A(n13476), .B(n13477), .Z(n13516) );
  XOR U13842 ( .A(b[23]), .B(a[82]), .Z(n13569) );
  NANDN U13843 ( .A(n19127), .B(n13569), .Z(n13428) );
  NAND U13844 ( .A(n13426), .B(n19128), .Z(n13427) );
  NAND U13845 ( .A(n13428), .B(n13427), .Z(n13539) );
  NANDN U13846 ( .A(n13429), .B(n17553), .Z(n13431) );
  XOR U13847 ( .A(b[7]), .B(a[98]), .Z(n13572) );
  NAND U13848 ( .A(n13572), .B(n17555), .Z(n13430) );
  NAND U13849 ( .A(n13431), .B(n13430), .Z(n13536) );
  XNOR U13850 ( .A(b[25]), .B(a[80]), .Z(n13575) );
  NANDN U13851 ( .A(n13575), .B(n19240), .Z(n13434) );
  NAND U13852 ( .A(n13432), .B(n19242), .Z(n13433) );
  AND U13853 ( .A(n13434), .B(n13433), .Z(n13537) );
  XNOR U13854 ( .A(n13536), .B(n13537), .Z(n13538) );
  XNOR U13855 ( .A(n13539), .B(n13538), .Z(n13517) );
  XOR U13856 ( .A(n13516), .B(n13517), .Z(n13519) );
  XNOR U13857 ( .A(n13518), .B(n13519), .Z(n13529) );
  XNOR U13858 ( .A(n13528), .B(n13529), .Z(n13464) );
  XNOR U13859 ( .A(n13465), .B(n13464), .Z(n13467) );
  XNOR U13860 ( .A(n13466), .B(n13467), .Z(n13584) );
  XOR U13861 ( .A(n13585), .B(n13584), .Z(n13587) );
  NANDN U13862 ( .A(n13436), .B(n13435), .Z(n13440) );
  NAND U13863 ( .A(n13438), .B(n13437), .Z(n13439) );
  NAND U13864 ( .A(n13440), .B(n13439), .Z(n13578) );
  NAND U13865 ( .A(n13442), .B(n13441), .Z(n13446) );
  NAND U13866 ( .A(n13444), .B(n13443), .Z(n13445) );
  NAND U13867 ( .A(n13446), .B(n13445), .Z(n13579) );
  XNOR U13868 ( .A(n13578), .B(n13579), .Z(n13580) );
  XOR U13869 ( .A(n13581), .B(n13580), .Z(n13461) );
  XOR U13870 ( .A(n13460), .B(n13461), .Z(n13452) );
  XOR U13871 ( .A(n13453), .B(n13452), .Z(n13454) );
  XNOR U13872 ( .A(n13455), .B(n13454), .Z(n13590) );
  XNOR U13873 ( .A(n13590), .B(sreg[200]), .Z(n13592) );
  NAND U13874 ( .A(n13447), .B(sreg[199]), .Z(n13451) );
  OR U13875 ( .A(n13449), .B(n13448), .Z(n13450) );
  AND U13876 ( .A(n13451), .B(n13450), .Z(n13591) );
  XOR U13877 ( .A(n13592), .B(n13591), .Z(c[200]) );
  NAND U13878 ( .A(n13453), .B(n13452), .Z(n13457) );
  NAND U13879 ( .A(n13455), .B(n13454), .Z(n13456) );
  NAND U13880 ( .A(n13457), .B(n13456), .Z(n13598) );
  NANDN U13881 ( .A(n13459), .B(n13458), .Z(n13463) );
  NAND U13882 ( .A(n13461), .B(n13460), .Z(n13462) );
  NAND U13883 ( .A(n13463), .B(n13462), .Z(n13595) );
  NAND U13884 ( .A(n13465), .B(n13464), .Z(n13469) );
  NANDN U13885 ( .A(n13467), .B(n13466), .Z(n13468) );
  NAND U13886 ( .A(n13469), .B(n13468), .Z(n13725) );
  XNOR U13887 ( .A(n13725), .B(n13726), .Z(n13727) );
  NANDN U13888 ( .A(n13475), .B(n13474), .Z(n13479) );
  NAND U13889 ( .A(n13477), .B(n13476), .Z(n13478) );
  NAND U13890 ( .A(n13479), .B(n13478), .Z(n13670) );
  NANDN U13891 ( .A(n13480), .B(n18832), .Z(n13482) );
  XNOR U13892 ( .A(b[19]), .B(a[87]), .Z(n13613) );
  NANDN U13893 ( .A(n13613), .B(n18834), .Z(n13481) );
  NAND U13894 ( .A(n13482), .B(n13481), .Z(n13680) );
  XNOR U13895 ( .A(b[27]), .B(a[79]), .Z(n13616) );
  NANDN U13896 ( .A(n13616), .B(n19336), .Z(n13485) );
  NANDN U13897 ( .A(n13483), .B(n19337), .Z(n13484) );
  NAND U13898 ( .A(n13485), .B(n13484), .Z(n13677) );
  XOR U13899 ( .A(b[5]), .B(a[101]), .Z(n13619) );
  NAND U13900 ( .A(n13619), .B(n17310), .Z(n13488) );
  NANDN U13901 ( .A(n13486), .B(n17311), .Z(n13487) );
  AND U13902 ( .A(n13488), .B(n13487), .Z(n13678) );
  XNOR U13903 ( .A(n13677), .B(n13678), .Z(n13679) );
  XNOR U13904 ( .A(n13680), .B(n13679), .Z(n13668) );
  XOR U13905 ( .A(b[17]), .B(a[89]), .Z(n13622) );
  NAND U13906 ( .A(n13622), .B(n18673), .Z(n13491) );
  NAND U13907 ( .A(n13489), .B(n18674), .Z(n13490) );
  NAND U13908 ( .A(n13491), .B(n13490), .Z(n13640) );
  XNOR U13909 ( .A(b[31]), .B(a[75]), .Z(n13625) );
  NANDN U13910 ( .A(n13625), .B(n19472), .Z(n13494) );
  NANDN U13911 ( .A(n13492), .B(n19473), .Z(n13493) );
  NAND U13912 ( .A(n13494), .B(n13493), .Z(n13637) );
  OR U13913 ( .A(n13495), .B(n16988), .Z(n13497) );
  XNOR U13914 ( .A(a[103]), .B(b[3]), .Z(n13628) );
  NANDN U13915 ( .A(n13628), .B(n16990), .Z(n13496) );
  AND U13916 ( .A(n13497), .B(n13496), .Z(n13638) );
  XNOR U13917 ( .A(n13637), .B(n13638), .Z(n13639) );
  XOR U13918 ( .A(n13640), .B(n13639), .Z(n13667) );
  XNOR U13919 ( .A(n13668), .B(n13667), .Z(n13669) );
  XNOR U13920 ( .A(n13670), .B(n13669), .Z(n13713) );
  NANDN U13921 ( .A(n13499), .B(n13498), .Z(n13503) );
  NAND U13922 ( .A(n13501), .B(n13500), .Z(n13502) );
  NAND U13923 ( .A(n13503), .B(n13502), .Z(n13658) );
  NANDN U13924 ( .A(n13505), .B(n13504), .Z(n13509) );
  NAND U13925 ( .A(n13507), .B(n13506), .Z(n13508) );
  NAND U13926 ( .A(n13509), .B(n13508), .Z(n13656) );
  OR U13927 ( .A(n13511), .B(n13510), .Z(n13515) );
  NANDN U13928 ( .A(n13513), .B(n13512), .Z(n13514) );
  NAND U13929 ( .A(n13515), .B(n13514), .Z(n13655) );
  XNOR U13930 ( .A(n13658), .B(n13657), .Z(n13714) );
  XNOR U13931 ( .A(n13713), .B(n13714), .Z(n13715) );
  NANDN U13932 ( .A(n13517), .B(n13516), .Z(n13521) );
  OR U13933 ( .A(n13519), .B(n13518), .Z(n13520) );
  AND U13934 ( .A(n13521), .B(n13520), .Z(n13716) );
  XOR U13935 ( .A(n13715), .B(n13716), .Z(n13733) );
  NANDN U13936 ( .A(n13527), .B(n13526), .Z(n13531) );
  NANDN U13937 ( .A(n13529), .B(n13528), .Z(n13530) );
  NAND U13938 ( .A(n13531), .B(n13530), .Z(n13722) );
  NANDN U13939 ( .A(n13537), .B(n13536), .Z(n13541) );
  NAND U13940 ( .A(n13539), .B(n13538), .Z(n13540) );
  NAND U13941 ( .A(n13541), .B(n13540), .Z(n13661) );
  NANDN U13942 ( .A(n13543), .B(n13542), .Z(n13547) );
  NAND U13943 ( .A(n13545), .B(n13544), .Z(n13546) );
  AND U13944 ( .A(n13547), .B(n13546), .Z(n13662) );
  XNOR U13945 ( .A(n13661), .B(n13662), .Z(n13663) );
  XOR U13946 ( .A(n579), .B(n17038), .Z(n13689) );
  NAND U13947 ( .A(n17814), .B(n13689), .Z(n13550) );
  NANDN U13948 ( .A(n13548), .B(n17815), .Z(n13549) );
  NAND U13949 ( .A(n13550), .B(n13549), .Z(n13645) );
  NAND U13950 ( .A(n13551), .B(n18513), .Z(n13553) );
  XOR U13951 ( .A(b[15]), .B(a[91]), .Z(n13686) );
  NANDN U13952 ( .A(n18512), .B(n13686), .Z(n13552) );
  AND U13953 ( .A(n13553), .B(n13552), .Z(n13643) );
  NANDN U13954 ( .A(n13554), .B(n19013), .Z(n13556) );
  XNOR U13955 ( .A(n582), .B(a[85]), .Z(n13683) );
  NAND U13956 ( .A(n13683), .B(n19015), .Z(n13555) );
  AND U13957 ( .A(n13556), .B(n13555), .Z(n13644) );
  XOR U13958 ( .A(n13645), .B(n13646), .Z(n13634) );
  XNOR U13959 ( .A(b[11]), .B(a[95]), .Z(n13692) );
  OR U13960 ( .A(n13692), .B(n18194), .Z(n13559) );
  NANDN U13961 ( .A(n13557), .B(n18104), .Z(n13558) );
  NAND U13962 ( .A(n13559), .B(n13558), .Z(n13632) );
  XOR U13963 ( .A(n580), .B(a[93]), .Z(n13695) );
  NANDN U13964 ( .A(n13695), .B(n18336), .Z(n13562) );
  NANDN U13965 ( .A(n13560), .B(n18337), .Z(n13561) );
  AND U13966 ( .A(n13562), .B(n13561), .Z(n13631) );
  XNOR U13967 ( .A(n13632), .B(n13631), .Z(n13633) );
  XOR U13968 ( .A(n13634), .B(n13633), .Z(n13651) );
  NAND U13969 ( .A(n19406), .B(n13563), .Z(n13565) );
  XNOR U13970 ( .A(n584), .B(a[77]), .Z(n13701) );
  NANDN U13971 ( .A(n576), .B(n13701), .Z(n13564) );
  NAND U13972 ( .A(n13565), .B(n13564), .Z(n13607) );
  NANDN U13973 ( .A(n585), .B(a[73]), .Z(n13608) );
  XNOR U13974 ( .A(n13607), .B(n13608), .Z(n13610) );
  NANDN U13975 ( .A(n577), .B(a[105]), .Z(n13566) );
  XOR U13976 ( .A(n17151), .B(n13566), .Z(n13568) );
  IV U13977 ( .A(a[104]), .Z(n17716) );
  NANDN U13978 ( .A(n17716), .B(n577), .Z(n13567) );
  AND U13979 ( .A(n13568), .B(n13567), .Z(n13609) );
  XOR U13980 ( .A(n13610), .B(n13609), .Z(n13649) );
  XOR U13981 ( .A(b[23]), .B(a[83]), .Z(n13704) );
  NANDN U13982 ( .A(n19127), .B(n13704), .Z(n13571) );
  NAND U13983 ( .A(n13569), .B(n19128), .Z(n13570) );
  NAND U13984 ( .A(n13571), .B(n13570), .Z(n13674) );
  NAND U13985 ( .A(n13572), .B(n17553), .Z(n13574) );
  XOR U13986 ( .A(b[7]), .B(a[99]), .Z(n13707) );
  NAND U13987 ( .A(n13707), .B(n17555), .Z(n13573) );
  NAND U13988 ( .A(n13574), .B(n13573), .Z(n13671) );
  XOR U13989 ( .A(b[25]), .B(a[81]), .Z(n13710) );
  NAND U13990 ( .A(n13710), .B(n19240), .Z(n13577) );
  NANDN U13991 ( .A(n13575), .B(n19242), .Z(n13576) );
  AND U13992 ( .A(n13577), .B(n13576), .Z(n13672) );
  XNOR U13993 ( .A(n13671), .B(n13672), .Z(n13673) );
  XNOR U13994 ( .A(n13674), .B(n13673), .Z(n13650) );
  XOR U13995 ( .A(n13649), .B(n13650), .Z(n13652) );
  XNOR U13996 ( .A(n13651), .B(n13652), .Z(n13664) );
  XOR U13997 ( .A(n13663), .B(n13664), .Z(n13720) );
  XNOR U13998 ( .A(n13719), .B(n13720), .Z(n13721) );
  XNOR U13999 ( .A(n13722), .B(n13721), .Z(n13731) );
  XNOR U14000 ( .A(n13732), .B(n13731), .Z(n13734) );
  XNOR U14001 ( .A(n13733), .B(n13734), .Z(n13728) );
  XOR U14002 ( .A(n13727), .B(n13728), .Z(n13604) );
  NANDN U14003 ( .A(n13579), .B(n13578), .Z(n13583) );
  NAND U14004 ( .A(n13581), .B(n13580), .Z(n13582) );
  NAND U14005 ( .A(n13583), .B(n13582), .Z(n13601) );
  NANDN U14006 ( .A(n13585), .B(n13584), .Z(n13589) );
  OR U14007 ( .A(n13587), .B(n13586), .Z(n13588) );
  NAND U14008 ( .A(n13589), .B(n13588), .Z(n13602) );
  XNOR U14009 ( .A(n13601), .B(n13602), .Z(n13603) );
  XNOR U14010 ( .A(n13604), .B(n13603), .Z(n13596) );
  XNOR U14011 ( .A(n13595), .B(n13596), .Z(n13597) );
  XNOR U14012 ( .A(n13598), .B(n13597), .Z(n13737) );
  XNOR U14013 ( .A(n13737), .B(sreg[201]), .Z(n13739) );
  NAND U14014 ( .A(n13590), .B(sreg[200]), .Z(n13594) );
  OR U14015 ( .A(n13592), .B(n13591), .Z(n13593) );
  AND U14016 ( .A(n13594), .B(n13593), .Z(n13738) );
  XOR U14017 ( .A(n13739), .B(n13738), .Z(c[201]) );
  NANDN U14018 ( .A(n13596), .B(n13595), .Z(n13600) );
  NAND U14019 ( .A(n13598), .B(n13597), .Z(n13599) );
  NAND U14020 ( .A(n13600), .B(n13599), .Z(n13745) );
  NANDN U14021 ( .A(n13602), .B(n13601), .Z(n13606) );
  NAND U14022 ( .A(n13604), .B(n13603), .Z(n13605) );
  NAND U14023 ( .A(n13606), .B(n13605), .Z(n13743) );
  NANDN U14024 ( .A(n13608), .B(n13607), .Z(n13612) );
  NAND U14025 ( .A(n13610), .B(n13609), .Z(n13611) );
  NAND U14026 ( .A(n13612), .B(n13611), .Z(n13815) );
  NANDN U14027 ( .A(n13613), .B(n18832), .Z(n13615) );
  XNOR U14028 ( .A(b[19]), .B(a[88]), .Z(n13760) );
  NANDN U14029 ( .A(n13760), .B(n18834), .Z(n13614) );
  NAND U14030 ( .A(n13615), .B(n13614), .Z(n13825) );
  XOR U14031 ( .A(b[27]), .B(n14551), .Z(n13763) );
  NANDN U14032 ( .A(n13763), .B(n19336), .Z(n13618) );
  NANDN U14033 ( .A(n13616), .B(n19337), .Z(n13617) );
  NAND U14034 ( .A(n13618), .B(n13617), .Z(n13822) );
  XNOR U14035 ( .A(b[5]), .B(a[102]), .Z(n13766) );
  NANDN U14036 ( .A(n13766), .B(n17310), .Z(n13621) );
  NAND U14037 ( .A(n13619), .B(n17311), .Z(n13620) );
  AND U14038 ( .A(n13621), .B(n13620), .Z(n13823) );
  XNOR U14039 ( .A(n13822), .B(n13823), .Z(n13824) );
  XNOR U14040 ( .A(n13825), .B(n13824), .Z(n13813) );
  XOR U14041 ( .A(b[17]), .B(a[90]), .Z(n13769) );
  NAND U14042 ( .A(n13769), .B(n18673), .Z(n13624) );
  NAND U14043 ( .A(n13622), .B(n18674), .Z(n13623) );
  NAND U14044 ( .A(n13624), .B(n13623), .Z(n13787) );
  XNOR U14045 ( .A(b[31]), .B(a[76]), .Z(n13772) );
  NANDN U14046 ( .A(n13772), .B(n19472), .Z(n13627) );
  NANDN U14047 ( .A(n13625), .B(n19473), .Z(n13626) );
  NAND U14048 ( .A(n13627), .B(n13626), .Z(n13784) );
  OR U14049 ( .A(n13628), .B(n16988), .Z(n13630) );
  XOR U14050 ( .A(a[104]), .B(n578), .Z(n13775) );
  NANDN U14051 ( .A(n13775), .B(n16990), .Z(n13629) );
  AND U14052 ( .A(n13630), .B(n13629), .Z(n13785) );
  XNOR U14053 ( .A(n13784), .B(n13785), .Z(n13786) );
  XOR U14054 ( .A(n13787), .B(n13786), .Z(n13812) );
  XNOR U14055 ( .A(n13813), .B(n13812), .Z(n13814) );
  XNOR U14056 ( .A(n13815), .B(n13814), .Z(n13858) );
  NANDN U14057 ( .A(n13632), .B(n13631), .Z(n13636) );
  NAND U14058 ( .A(n13634), .B(n13633), .Z(n13635) );
  NAND U14059 ( .A(n13636), .B(n13635), .Z(n13803) );
  NANDN U14060 ( .A(n13638), .B(n13637), .Z(n13642) );
  NAND U14061 ( .A(n13640), .B(n13639), .Z(n13641) );
  NAND U14062 ( .A(n13642), .B(n13641), .Z(n13801) );
  OR U14063 ( .A(n13644), .B(n13643), .Z(n13648) );
  NANDN U14064 ( .A(n13646), .B(n13645), .Z(n13647) );
  NAND U14065 ( .A(n13648), .B(n13647), .Z(n13800) );
  XNOR U14066 ( .A(n13803), .B(n13802), .Z(n13859) );
  XOR U14067 ( .A(n13858), .B(n13859), .Z(n13861) );
  NANDN U14068 ( .A(n13650), .B(n13649), .Z(n13654) );
  OR U14069 ( .A(n13652), .B(n13651), .Z(n13653) );
  NAND U14070 ( .A(n13654), .B(n13653), .Z(n13860) );
  XOR U14071 ( .A(n13861), .B(n13860), .Z(n13878) );
  OR U14072 ( .A(n13656), .B(n13655), .Z(n13660) );
  NAND U14073 ( .A(n13658), .B(n13657), .Z(n13659) );
  NAND U14074 ( .A(n13660), .B(n13659), .Z(n13877) );
  NANDN U14075 ( .A(n13662), .B(n13661), .Z(n13666) );
  NANDN U14076 ( .A(n13664), .B(n13663), .Z(n13665) );
  NAND U14077 ( .A(n13666), .B(n13665), .Z(n13866) );
  NANDN U14078 ( .A(n13672), .B(n13671), .Z(n13676) );
  NAND U14079 ( .A(n13674), .B(n13673), .Z(n13675) );
  NAND U14080 ( .A(n13676), .B(n13675), .Z(n13806) );
  NANDN U14081 ( .A(n13678), .B(n13677), .Z(n13682) );
  NAND U14082 ( .A(n13680), .B(n13679), .Z(n13681) );
  AND U14083 ( .A(n13682), .B(n13681), .Z(n13807) );
  XNOR U14084 ( .A(n13806), .B(n13807), .Z(n13808) );
  XOR U14085 ( .A(n582), .B(a[86]), .Z(n13834) );
  NANDN U14086 ( .A(n13834), .B(n19015), .Z(n13685) );
  NAND U14087 ( .A(n19013), .B(n13683), .Z(n13684) );
  NAND U14088 ( .A(n13685), .B(n13684), .Z(n13796) );
  NAND U14089 ( .A(n13686), .B(n18513), .Z(n13688) );
  XOR U14090 ( .A(b[15]), .B(a[92]), .Z(n13831) );
  NANDN U14091 ( .A(n18512), .B(n13831), .Z(n13687) );
  AND U14092 ( .A(n13688), .B(n13687), .Z(n13797) );
  XNOR U14093 ( .A(n13796), .B(n13797), .Z(n13799) );
  XOR U14094 ( .A(n579), .B(a[98]), .Z(n13828) );
  NANDN U14095 ( .A(n13828), .B(n17814), .Z(n13691) );
  NAND U14096 ( .A(n17815), .B(n13689), .Z(n13690) );
  NAND U14097 ( .A(n13691), .B(n13690), .Z(n13798) );
  XNOR U14098 ( .A(n13799), .B(n13798), .Z(n13792) );
  XNOR U14099 ( .A(b[11]), .B(a[96]), .Z(n13837) );
  OR U14100 ( .A(n13837), .B(n18194), .Z(n13694) );
  NANDN U14101 ( .A(n13692), .B(n18104), .Z(n13693) );
  NAND U14102 ( .A(n13694), .B(n13693), .Z(n13791) );
  XOR U14103 ( .A(n580), .B(a[94]), .Z(n13840) );
  NANDN U14104 ( .A(n13840), .B(n18336), .Z(n13697) );
  NANDN U14105 ( .A(n13695), .B(n18337), .Z(n13696) );
  NAND U14106 ( .A(n13697), .B(n13696), .Z(n13790) );
  XNOR U14107 ( .A(n13791), .B(n13790), .Z(n13793) );
  XNOR U14108 ( .A(n13792), .B(n13793), .Z(n13781) );
  NANDN U14109 ( .A(n577), .B(a[106]), .Z(n13698) );
  XOR U14110 ( .A(n17151), .B(n13698), .Z(n13700) );
  NANDN U14111 ( .A(b[0]), .B(a[105]), .Z(n13699) );
  AND U14112 ( .A(n13700), .B(n13699), .Z(n13756) );
  NAND U14113 ( .A(n19406), .B(n13701), .Z(n13703) );
  XNOR U14114 ( .A(n584), .B(a[78]), .Z(n13846) );
  NANDN U14115 ( .A(n576), .B(n13846), .Z(n13702) );
  NAND U14116 ( .A(n13703), .B(n13702), .Z(n13754) );
  NANDN U14117 ( .A(n585), .B(a[74]), .Z(n13755) );
  XNOR U14118 ( .A(n13754), .B(n13755), .Z(n13757) );
  XNOR U14119 ( .A(n13756), .B(n13757), .Z(n13779) );
  XNOR U14120 ( .A(b[23]), .B(a[84]), .Z(n13849) );
  OR U14121 ( .A(n13849), .B(n19127), .Z(n13706) );
  NAND U14122 ( .A(n13704), .B(n19128), .Z(n13705) );
  NAND U14123 ( .A(n13706), .B(n13705), .Z(n13819) );
  NAND U14124 ( .A(n13707), .B(n17553), .Z(n13709) );
  XNOR U14125 ( .A(b[7]), .B(a[100]), .Z(n13852) );
  NANDN U14126 ( .A(n13852), .B(n17555), .Z(n13708) );
  NAND U14127 ( .A(n13709), .B(n13708), .Z(n13816) );
  XOR U14128 ( .A(b[25]), .B(a[82]), .Z(n13855) );
  NAND U14129 ( .A(n13855), .B(n19240), .Z(n13712) );
  NAND U14130 ( .A(n13710), .B(n19242), .Z(n13711) );
  AND U14131 ( .A(n13712), .B(n13711), .Z(n13817) );
  XNOR U14132 ( .A(n13816), .B(n13817), .Z(n13818) );
  XOR U14133 ( .A(n13819), .B(n13818), .Z(n13778) );
  XOR U14134 ( .A(n13781), .B(n13780), .Z(n13809) );
  XNOR U14135 ( .A(n13808), .B(n13809), .Z(n13864) );
  XNOR U14136 ( .A(n13865), .B(n13864), .Z(n13867) );
  XNOR U14137 ( .A(n13866), .B(n13867), .Z(n13876) );
  XOR U14138 ( .A(n13877), .B(n13876), .Z(n13879) );
  NANDN U14139 ( .A(n13714), .B(n13713), .Z(n13718) );
  NAND U14140 ( .A(n13716), .B(n13715), .Z(n13717) );
  NAND U14141 ( .A(n13718), .B(n13717), .Z(n13870) );
  NANDN U14142 ( .A(n13720), .B(n13719), .Z(n13724) );
  NAND U14143 ( .A(n13722), .B(n13721), .Z(n13723) );
  NAND U14144 ( .A(n13724), .B(n13723), .Z(n13871) );
  XNOR U14145 ( .A(n13870), .B(n13871), .Z(n13872) );
  XOR U14146 ( .A(n13873), .B(n13872), .Z(n13750) );
  NANDN U14147 ( .A(n13726), .B(n13725), .Z(n13730) );
  NANDN U14148 ( .A(n13728), .B(n13727), .Z(n13729) );
  NAND U14149 ( .A(n13730), .B(n13729), .Z(n13749) );
  OR U14150 ( .A(n13732), .B(n13731), .Z(n13736) );
  OR U14151 ( .A(n13734), .B(n13733), .Z(n13735) );
  AND U14152 ( .A(n13736), .B(n13735), .Z(n13748) );
  XNOR U14153 ( .A(n13749), .B(n13748), .Z(n13751) );
  XOR U14154 ( .A(n13750), .B(n13751), .Z(n13742) );
  XOR U14155 ( .A(n13743), .B(n13742), .Z(n13744) );
  XNOR U14156 ( .A(n13745), .B(n13744), .Z(n13882) );
  XNOR U14157 ( .A(n13882), .B(sreg[202]), .Z(n13884) );
  NAND U14158 ( .A(n13737), .B(sreg[201]), .Z(n13741) );
  OR U14159 ( .A(n13739), .B(n13738), .Z(n13740) );
  AND U14160 ( .A(n13741), .B(n13740), .Z(n13883) );
  XOR U14161 ( .A(n13884), .B(n13883), .Z(c[202]) );
  NAND U14162 ( .A(n13743), .B(n13742), .Z(n13747) );
  NAND U14163 ( .A(n13745), .B(n13744), .Z(n13746) );
  NAND U14164 ( .A(n13747), .B(n13746), .Z(n13890) );
  NANDN U14165 ( .A(n13749), .B(n13748), .Z(n13753) );
  NAND U14166 ( .A(n13751), .B(n13750), .Z(n13752) );
  NAND U14167 ( .A(n13753), .B(n13752), .Z(n13888) );
  NANDN U14168 ( .A(n13755), .B(n13754), .Z(n13759) );
  NAND U14169 ( .A(n13757), .B(n13756), .Z(n13758) );
  NAND U14170 ( .A(n13759), .B(n13758), .Z(n13958) );
  NANDN U14171 ( .A(n13760), .B(n18832), .Z(n13762) );
  XNOR U14172 ( .A(b[19]), .B(a[89]), .Z(n13905) );
  NANDN U14173 ( .A(n13905), .B(n18834), .Z(n13761) );
  NAND U14174 ( .A(n13762), .B(n13761), .Z(n13968) );
  XNOR U14175 ( .A(b[27]), .B(a[81]), .Z(n13908) );
  NANDN U14176 ( .A(n13908), .B(n19336), .Z(n13765) );
  NANDN U14177 ( .A(n13763), .B(n19337), .Z(n13764) );
  NAND U14178 ( .A(n13765), .B(n13764), .Z(n13965) );
  XOR U14179 ( .A(b[5]), .B(a[103]), .Z(n13911) );
  NAND U14180 ( .A(n13911), .B(n17310), .Z(n13768) );
  NANDN U14181 ( .A(n13766), .B(n17311), .Z(n13767) );
  AND U14182 ( .A(n13768), .B(n13767), .Z(n13966) );
  XNOR U14183 ( .A(n13965), .B(n13966), .Z(n13967) );
  XNOR U14184 ( .A(n13968), .B(n13967), .Z(n13956) );
  XOR U14185 ( .A(b[17]), .B(a[91]), .Z(n13914) );
  NAND U14186 ( .A(n13914), .B(n18673), .Z(n13771) );
  NAND U14187 ( .A(n13769), .B(n18674), .Z(n13770) );
  NAND U14188 ( .A(n13771), .B(n13770), .Z(n13932) );
  XNOR U14189 ( .A(b[31]), .B(a[77]), .Z(n13917) );
  NANDN U14190 ( .A(n13917), .B(n19472), .Z(n13774) );
  NANDN U14191 ( .A(n13772), .B(n19473), .Z(n13773) );
  NAND U14192 ( .A(n13774), .B(n13773), .Z(n13929) );
  OR U14193 ( .A(n13775), .B(n16988), .Z(n13777) );
  XNOR U14194 ( .A(a[105]), .B(b[3]), .Z(n13920) );
  NANDN U14195 ( .A(n13920), .B(n16990), .Z(n13776) );
  AND U14196 ( .A(n13777), .B(n13776), .Z(n13930) );
  XNOR U14197 ( .A(n13929), .B(n13930), .Z(n13931) );
  XOR U14198 ( .A(n13932), .B(n13931), .Z(n13955) );
  XNOR U14199 ( .A(n13956), .B(n13955), .Z(n13957) );
  XNOR U14200 ( .A(n13958), .B(n13957), .Z(n14007) );
  NANDN U14201 ( .A(n13779), .B(n13778), .Z(n13783) );
  NANDN U14202 ( .A(n13781), .B(n13780), .Z(n13782) );
  NAND U14203 ( .A(n13783), .B(n13782), .Z(n14008) );
  XNOR U14204 ( .A(n14007), .B(n14008), .Z(n14009) );
  NANDN U14205 ( .A(n13785), .B(n13784), .Z(n13789) );
  NAND U14206 ( .A(n13787), .B(n13786), .Z(n13788) );
  NAND U14207 ( .A(n13789), .B(n13788), .Z(n13948) );
  OR U14208 ( .A(n13791), .B(n13790), .Z(n13795) );
  NANDN U14209 ( .A(n13793), .B(n13792), .Z(n13794) );
  NAND U14210 ( .A(n13795), .B(n13794), .Z(n13946) );
  XNOR U14211 ( .A(n13946), .B(n13945), .Z(n13947) );
  XOR U14212 ( .A(n13948), .B(n13947), .Z(n14010) );
  XOR U14213 ( .A(n14009), .B(n14010), .Z(n14020) );
  OR U14214 ( .A(n13801), .B(n13800), .Z(n13805) );
  NAND U14215 ( .A(n13803), .B(n13802), .Z(n13804) );
  NAND U14216 ( .A(n13805), .B(n13804), .Z(n14018) );
  NANDN U14217 ( .A(n13807), .B(n13806), .Z(n13811) );
  NANDN U14218 ( .A(n13809), .B(n13808), .Z(n13810) );
  NAND U14219 ( .A(n13811), .B(n13810), .Z(n14003) );
  NANDN U14220 ( .A(n13817), .B(n13816), .Z(n13821) );
  NAND U14221 ( .A(n13819), .B(n13818), .Z(n13820) );
  NAND U14222 ( .A(n13821), .B(n13820), .Z(n13949) );
  NANDN U14223 ( .A(n13823), .B(n13822), .Z(n13827) );
  NAND U14224 ( .A(n13825), .B(n13824), .Z(n13826) );
  AND U14225 ( .A(n13827), .B(n13826), .Z(n13950) );
  XNOR U14226 ( .A(n13949), .B(n13950), .Z(n13951) );
  XOR U14227 ( .A(n579), .B(a[99]), .Z(n13971) );
  NANDN U14228 ( .A(n13971), .B(n17814), .Z(n13830) );
  NANDN U14229 ( .A(n13828), .B(n17815), .Z(n13829) );
  NAND U14230 ( .A(n13830), .B(n13829), .Z(n13937) );
  XNOR U14231 ( .A(b[15]), .B(a[93]), .Z(n13974) );
  OR U14232 ( .A(n13974), .B(n18512), .Z(n13833) );
  NAND U14233 ( .A(n13831), .B(n18513), .Z(n13832) );
  NAND U14234 ( .A(n13833), .B(n13832), .Z(n13935) );
  XOR U14235 ( .A(n582), .B(a[87]), .Z(n13977) );
  NANDN U14236 ( .A(n13977), .B(n19015), .Z(n13836) );
  NANDN U14237 ( .A(n13834), .B(n19013), .Z(n13835) );
  NAND U14238 ( .A(n13836), .B(n13835), .Z(n13936) );
  XNOR U14239 ( .A(n13935), .B(n13936), .Z(n13938) );
  XOR U14240 ( .A(n13937), .B(n13938), .Z(n13926) );
  XOR U14241 ( .A(b[11]), .B(n17038), .Z(n13980) );
  OR U14242 ( .A(n13980), .B(n18194), .Z(n13839) );
  NANDN U14243 ( .A(n13837), .B(n18104), .Z(n13838) );
  NAND U14244 ( .A(n13839), .B(n13838), .Z(n13924) );
  XOR U14245 ( .A(n580), .B(a[95]), .Z(n13983) );
  NANDN U14246 ( .A(n13983), .B(n18336), .Z(n13842) );
  NANDN U14247 ( .A(n13840), .B(n18337), .Z(n13841) );
  AND U14248 ( .A(n13842), .B(n13841), .Z(n13923) );
  XNOR U14249 ( .A(n13924), .B(n13923), .Z(n13925) );
  XNOR U14250 ( .A(n13926), .B(n13925), .Z(n13942) );
  NANDN U14251 ( .A(n577), .B(a[107]), .Z(n13843) );
  XOR U14252 ( .A(n17151), .B(n13843), .Z(n13845) );
  IV U14253 ( .A(a[106]), .Z(n17690) );
  NANDN U14254 ( .A(n17690), .B(n577), .Z(n13844) );
  AND U14255 ( .A(n13845), .B(n13844), .Z(n13901) );
  NAND U14256 ( .A(n19406), .B(n13846), .Z(n13848) );
  XNOR U14257 ( .A(n584), .B(a[79]), .Z(n13986) );
  NANDN U14258 ( .A(n576), .B(n13986), .Z(n13847) );
  NAND U14259 ( .A(n13848), .B(n13847), .Z(n13899) );
  NANDN U14260 ( .A(n585), .B(a[75]), .Z(n13900) );
  XNOR U14261 ( .A(n13899), .B(n13900), .Z(n13902) );
  XNOR U14262 ( .A(n13901), .B(n13902), .Z(n13940) );
  XOR U14263 ( .A(b[23]), .B(a[85]), .Z(n13992) );
  NANDN U14264 ( .A(n19127), .B(n13992), .Z(n13851) );
  NANDN U14265 ( .A(n13849), .B(n19128), .Z(n13850) );
  NAND U14266 ( .A(n13851), .B(n13850), .Z(n13962) );
  NANDN U14267 ( .A(n13852), .B(n17553), .Z(n13854) );
  XOR U14268 ( .A(b[7]), .B(a[101]), .Z(n13995) );
  NAND U14269 ( .A(n13995), .B(n17555), .Z(n13853) );
  NAND U14270 ( .A(n13854), .B(n13853), .Z(n13959) );
  XOR U14271 ( .A(b[25]), .B(a[83]), .Z(n13998) );
  NAND U14272 ( .A(n13998), .B(n19240), .Z(n13857) );
  NAND U14273 ( .A(n13855), .B(n19242), .Z(n13856) );
  AND U14274 ( .A(n13857), .B(n13856), .Z(n13960) );
  XNOR U14275 ( .A(n13959), .B(n13960), .Z(n13961) );
  XOR U14276 ( .A(n13962), .B(n13961), .Z(n13939) );
  XOR U14277 ( .A(n13942), .B(n13941), .Z(n13952) );
  XOR U14278 ( .A(n13951), .B(n13952), .Z(n14001) );
  XNOR U14279 ( .A(n14002), .B(n14001), .Z(n14004) );
  XNOR U14280 ( .A(n14003), .B(n14004), .Z(n14017) );
  XOR U14281 ( .A(n14018), .B(n14017), .Z(n14019) );
  XNOR U14282 ( .A(n14020), .B(n14019), .Z(n14014) );
  NANDN U14283 ( .A(n13859), .B(n13858), .Z(n13863) );
  OR U14284 ( .A(n13861), .B(n13860), .Z(n13862) );
  NAND U14285 ( .A(n13863), .B(n13862), .Z(n14011) );
  NAND U14286 ( .A(n13865), .B(n13864), .Z(n13869) );
  NANDN U14287 ( .A(n13867), .B(n13866), .Z(n13868) );
  NAND U14288 ( .A(n13869), .B(n13868), .Z(n14012) );
  XNOR U14289 ( .A(n14011), .B(n14012), .Z(n14013) );
  XOR U14290 ( .A(n14014), .B(n14013), .Z(n13895) );
  NANDN U14291 ( .A(n13871), .B(n13870), .Z(n13875) );
  NAND U14292 ( .A(n13873), .B(n13872), .Z(n13874) );
  NAND U14293 ( .A(n13875), .B(n13874), .Z(n13893) );
  NANDN U14294 ( .A(n13877), .B(n13876), .Z(n13881) );
  OR U14295 ( .A(n13879), .B(n13878), .Z(n13880) );
  NAND U14296 ( .A(n13881), .B(n13880), .Z(n13894) );
  XNOR U14297 ( .A(n13893), .B(n13894), .Z(n13896) );
  XOR U14298 ( .A(n13895), .B(n13896), .Z(n13887) );
  XOR U14299 ( .A(n13888), .B(n13887), .Z(n13889) );
  XNOR U14300 ( .A(n13890), .B(n13889), .Z(n14023) );
  XNOR U14301 ( .A(n14023), .B(sreg[203]), .Z(n14025) );
  NAND U14302 ( .A(n13882), .B(sreg[202]), .Z(n13886) );
  OR U14303 ( .A(n13884), .B(n13883), .Z(n13885) );
  AND U14304 ( .A(n13886), .B(n13885), .Z(n14024) );
  XOR U14305 ( .A(n14025), .B(n14024), .Z(c[203]) );
  NAND U14306 ( .A(n13888), .B(n13887), .Z(n13892) );
  NAND U14307 ( .A(n13890), .B(n13889), .Z(n13891) );
  NAND U14308 ( .A(n13892), .B(n13891), .Z(n14031) );
  NANDN U14309 ( .A(n13894), .B(n13893), .Z(n13898) );
  NAND U14310 ( .A(n13896), .B(n13895), .Z(n13897) );
  NAND U14311 ( .A(n13898), .B(n13897), .Z(n14029) );
  NANDN U14312 ( .A(n13900), .B(n13899), .Z(n13904) );
  NAND U14313 ( .A(n13902), .B(n13901), .Z(n13903) );
  NAND U14314 ( .A(n13904), .B(n13903), .Z(n14107) );
  NANDN U14315 ( .A(n13905), .B(n18832), .Z(n13907) );
  XNOR U14316 ( .A(b[19]), .B(a[90]), .Z(n14054) );
  NANDN U14317 ( .A(n14054), .B(n18834), .Z(n13906) );
  NAND U14318 ( .A(n13907), .B(n13906), .Z(n14117) );
  XNOR U14319 ( .A(b[27]), .B(a[82]), .Z(n14057) );
  NANDN U14320 ( .A(n14057), .B(n19336), .Z(n13910) );
  NANDN U14321 ( .A(n13908), .B(n19337), .Z(n13909) );
  NAND U14322 ( .A(n13910), .B(n13909), .Z(n14114) );
  XNOR U14323 ( .A(a[104]), .B(b[5]), .Z(n14060) );
  NANDN U14324 ( .A(n14060), .B(n17310), .Z(n13913) );
  NAND U14325 ( .A(n13911), .B(n17311), .Z(n13912) );
  AND U14326 ( .A(n13913), .B(n13912), .Z(n14115) );
  XNOR U14327 ( .A(n14114), .B(n14115), .Z(n14116) );
  XNOR U14328 ( .A(n14117), .B(n14116), .Z(n14105) );
  XOR U14329 ( .A(b[17]), .B(a[92]), .Z(n14063) );
  NAND U14330 ( .A(n14063), .B(n18673), .Z(n13916) );
  NAND U14331 ( .A(n13914), .B(n18674), .Z(n13915) );
  NAND U14332 ( .A(n13916), .B(n13915), .Z(n14081) );
  XNOR U14333 ( .A(b[31]), .B(a[78]), .Z(n14066) );
  NANDN U14334 ( .A(n14066), .B(n19472), .Z(n13919) );
  NANDN U14335 ( .A(n13917), .B(n19473), .Z(n13918) );
  NAND U14336 ( .A(n13919), .B(n13918), .Z(n14078) );
  OR U14337 ( .A(n13920), .B(n16988), .Z(n13922) );
  XOR U14338 ( .A(a[106]), .B(n578), .Z(n14069) );
  NANDN U14339 ( .A(n14069), .B(n16990), .Z(n13921) );
  AND U14340 ( .A(n13922), .B(n13921), .Z(n14079) );
  XNOR U14341 ( .A(n14078), .B(n14079), .Z(n14080) );
  XOR U14342 ( .A(n14081), .B(n14080), .Z(n14104) );
  XNOR U14343 ( .A(n14105), .B(n14104), .Z(n14106) );
  XNOR U14344 ( .A(n14107), .B(n14106), .Z(n14045) );
  NANDN U14345 ( .A(n13924), .B(n13923), .Z(n13928) );
  NAND U14346 ( .A(n13926), .B(n13925), .Z(n13927) );
  NAND U14347 ( .A(n13928), .B(n13927), .Z(n14096) );
  NANDN U14348 ( .A(n13930), .B(n13929), .Z(n13934) );
  NAND U14349 ( .A(n13932), .B(n13931), .Z(n13933) );
  NAND U14350 ( .A(n13934), .B(n13933), .Z(n14095) );
  XNOR U14351 ( .A(n14095), .B(n14094), .Z(n14097) );
  XOR U14352 ( .A(n14096), .B(n14097), .Z(n14044) );
  XOR U14353 ( .A(n14045), .B(n14044), .Z(n14046) );
  NANDN U14354 ( .A(n13940), .B(n13939), .Z(n13944) );
  NAND U14355 ( .A(n13942), .B(n13941), .Z(n13943) );
  AND U14356 ( .A(n13944), .B(n13943), .Z(n14047) );
  XNOR U14357 ( .A(n14046), .B(n14047), .Z(n14153) );
  NANDN U14358 ( .A(n13950), .B(n13949), .Z(n13954) );
  NAND U14359 ( .A(n13952), .B(n13951), .Z(n13953) );
  NAND U14360 ( .A(n13954), .B(n13953), .Z(n14041) );
  NANDN U14361 ( .A(n13960), .B(n13959), .Z(n13964) );
  NAND U14362 ( .A(n13962), .B(n13961), .Z(n13963) );
  NAND U14363 ( .A(n13964), .B(n13963), .Z(n14098) );
  NANDN U14364 ( .A(n13966), .B(n13965), .Z(n13970) );
  NAND U14365 ( .A(n13968), .B(n13967), .Z(n13969) );
  AND U14366 ( .A(n13970), .B(n13969), .Z(n14099) );
  XNOR U14367 ( .A(n14098), .B(n14099), .Z(n14100) );
  XOR U14368 ( .A(n579), .B(a[100]), .Z(n14126) );
  NANDN U14369 ( .A(n14126), .B(n17814), .Z(n13973) );
  NANDN U14370 ( .A(n13971), .B(n17815), .Z(n13972) );
  NAND U14371 ( .A(n13973), .B(n13972), .Z(n14086) );
  XNOR U14372 ( .A(b[15]), .B(a[94]), .Z(n14123) );
  OR U14373 ( .A(n14123), .B(n18512), .Z(n13976) );
  NANDN U14374 ( .A(n13974), .B(n18513), .Z(n13975) );
  NAND U14375 ( .A(n13976), .B(n13975), .Z(n14084) );
  XOR U14376 ( .A(n582), .B(a[88]), .Z(n14120) );
  NANDN U14377 ( .A(n14120), .B(n19015), .Z(n13979) );
  NANDN U14378 ( .A(n13977), .B(n19013), .Z(n13978) );
  NAND U14379 ( .A(n13979), .B(n13978), .Z(n14085) );
  XNOR U14380 ( .A(n14084), .B(n14085), .Z(n14087) );
  XOR U14381 ( .A(n14086), .B(n14087), .Z(n14075) );
  XNOR U14382 ( .A(b[11]), .B(a[98]), .Z(n14129) );
  OR U14383 ( .A(n14129), .B(n18194), .Z(n13982) );
  NANDN U14384 ( .A(n13980), .B(n18104), .Z(n13981) );
  NAND U14385 ( .A(n13982), .B(n13981), .Z(n14073) );
  XOR U14386 ( .A(n580), .B(a[96]), .Z(n14132) );
  NANDN U14387 ( .A(n14132), .B(n18336), .Z(n13985) );
  NANDN U14388 ( .A(n13983), .B(n18337), .Z(n13984) );
  AND U14389 ( .A(n13985), .B(n13984), .Z(n14072) );
  XNOR U14390 ( .A(n14073), .B(n14072), .Z(n14074) );
  XNOR U14391 ( .A(n14075), .B(n14074), .Z(n14091) );
  NAND U14392 ( .A(n19406), .B(n13986), .Z(n13988) );
  XOR U14393 ( .A(n584), .B(n14551), .Z(n14138) );
  NANDN U14394 ( .A(n576), .B(n14138), .Z(n13987) );
  NAND U14395 ( .A(n13988), .B(n13987), .Z(n14048) );
  NANDN U14396 ( .A(n585), .B(a[76]), .Z(n14049) );
  XNOR U14397 ( .A(n14048), .B(n14049), .Z(n14051) );
  NANDN U14398 ( .A(n577), .B(a[108]), .Z(n13989) );
  XOR U14399 ( .A(n17151), .B(n13989), .Z(n13991) );
  NANDN U14400 ( .A(b[0]), .B(a[107]), .Z(n13990) );
  AND U14401 ( .A(n13991), .B(n13990), .Z(n14050) );
  XNOR U14402 ( .A(n14051), .B(n14050), .Z(n14089) );
  XNOR U14403 ( .A(b[23]), .B(a[86]), .Z(n14141) );
  OR U14404 ( .A(n14141), .B(n19127), .Z(n13994) );
  NAND U14405 ( .A(n13992), .B(n19128), .Z(n13993) );
  NAND U14406 ( .A(n13994), .B(n13993), .Z(n14111) );
  NAND U14407 ( .A(n13995), .B(n17553), .Z(n13997) );
  XNOR U14408 ( .A(b[7]), .B(a[102]), .Z(n14144) );
  NANDN U14409 ( .A(n14144), .B(n17555), .Z(n13996) );
  NAND U14410 ( .A(n13997), .B(n13996), .Z(n14108) );
  XNOR U14411 ( .A(b[25]), .B(a[84]), .Z(n14147) );
  NANDN U14412 ( .A(n14147), .B(n19240), .Z(n14000) );
  NAND U14413 ( .A(n13998), .B(n19242), .Z(n13999) );
  AND U14414 ( .A(n14000), .B(n13999), .Z(n14109) );
  XNOR U14415 ( .A(n14108), .B(n14109), .Z(n14110) );
  XOR U14416 ( .A(n14111), .B(n14110), .Z(n14088) );
  XOR U14417 ( .A(n14091), .B(n14090), .Z(n14101) );
  XOR U14418 ( .A(n14100), .B(n14101), .Z(n14038) );
  XOR U14419 ( .A(n14039), .B(n14038), .Z(n14040) );
  XOR U14420 ( .A(n14041), .B(n14040), .Z(n14151) );
  XNOR U14421 ( .A(n14150), .B(n14151), .Z(n14152) );
  XNOR U14422 ( .A(n14153), .B(n14152), .Z(n14157) );
  NAND U14423 ( .A(n14002), .B(n14001), .Z(n14006) );
  NANDN U14424 ( .A(n14004), .B(n14003), .Z(n14005) );
  NAND U14425 ( .A(n14006), .B(n14005), .Z(n14154) );
  XNOR U14426 ( .A(n14154), .B(n14155), .Z(n14156) );
  XNOR U14427 ( .A(n14157), .B(n14156), .Z(n14035) );
  NANDN U14428 ( .A(n14012), .B(n14011), .Z(n14016) );
  NAND U14429 ( .A(n14014), .B(n14013), .Z(n14015) );
  NAND U14430 ( .A(n14016), .B(n14015), .Z(n14032) );
  NANDN U14431 ( .A(n14018), .B(n14017), .Z(n14022) );
  OR U14432 ( .A(n14020), .B(n14019), .Z(n14021) );
  NAND U14433 ( .A(n14022), .B(n14021), .Z(n14033) );
  XNOR U14434 ( .A(n14032), .B(n14033), .Z(n14034) );
  XNOR U14435 ( .A(n14035), .B(n14034), .Z(n14028) );
  XOR U14436 ( .A(n14029), .B(n14028), .Z(n14030) );
  XNOR U14437 ( .A(n14031), .B(n14030), .Z(n14160) );
  XNOR U14438 ( .A(n14160), .B(sreg[204]), .Z(n14162) );
  NAND U14439 ( .A(n14023), .B(sreg[203]), .Z(n14027) );
  OR U14440 ( .A(n14025), .B(n14024), .Z(n14026) );
  AND U14441 ( .A(n14027), .B(n14026), .Z(n14161) );
  XOR U14442 ( .A(n14162), .B(n14161), .Z(c[204]) );
  NANDN U14443 ( .A(n14033), .B(n14032), .Z(n14037) );
  NANDN U14444 ( .A(n14035), .B(n14034), .Z(n14036) );
  NAND U14445 ( .A(n14037), .B(n14036), .Z(n14165) );
  NAND U14446 ( .A(n14039), .B(n14038), .Z(n14043) );
  NAND U14447 ( .A(n14041), .B(n14040), .Z(n14042) );
  NAND U14448 ( .A(n14043), .B(n14042), .Z(n14289) );
  XNOR U14449 ( .A(n14289), .B(n14290), .Z(n14291) );
  NANDN U14450 ( .A(n14049), .B(n14048), .Z(n14053) );
  NAND U14451 ( .A(n14051), .B(n14050), .Z(n14052) );
  NAND U14452 ( .A(n14053), .B(n14052), .Z(n14246) );
  NANDN U14453 ( .A(n14054), .B(n18832), .Z(n14056) );
  XNOR U14454 ( .A(b[19]), .B(a[91]), .Z(n14193) );
  NANDN U14455 ( .A(n14193), .B(n18834), .Z(n14055) );
  NAND U14456 ( .A(n14056), .B(n14055), .Z(n14256) );
  XNOR U14457 ( .A(b[27]), .B(a[83]), .Z(n14196) );
  NANDN U14458 ( .A(n14196), .B(n19336), .Z(n14059) );
  NANDN U14459 ( .A(n14057), .B(n19337), .Z(n14058) );
  NAND U14460 ( .A(n14059), .B(n14058), .Z(n14253) );
  XOR U14461 ( .A(a[105]), .B(b[5]), .Z(n14199) );
  NAND U14462 ( .A(n14199), .B(n17310), .Z(n14062) );
  NANDN U14463 ( .A(n14060), .B(n17311), .Z(n14061) );
  AND U14464 ( .A(n14062), .B(n14061), .Z(n14254) );
  XNOR U14465 ( .A(n14253), .B(n14254), .Z(n14255) );
  XNOR U14466 ( .A(n14256), .B(n14255), .Z(n14244) );
  XOR U14467 ( .A(b[17]), .B(a[93]), .Z(n14202) );
  NAND U14468 ( .A(n14202), .B(n18673), .Z(n14065) );
  NAND U14469 ( .A(n14063), .B(n18674), .Z(n14064) );
  NAND U14470 ( .A(n14065), .B(n14064), .Z(n14220) );
  XNOR U14471 ( .A(b[31]), .B(a[79]), .Z(n14205) );
  NANDN U14472 ( .A(n14205), .B(n19472), .Z(n14068) );
  NANDN U14473 ( .A(n14066), .B(n19473), .Z(n14067) );
  NAND U14474 ( .A(n14068), .B(n14067), .Z(n14217) );
  OR U14475 ( .A(n14069), .B(n16988), .Z(n14071) );
  XNOR U14476 ( .A(a[107]), .B(b[3]), .Z(n14208) );
  NANDN U14477 ( .A(n14208), .B(n16990), .Z(n14070) );
  AND U14478 ( .A(n14071), .B(n14070), .Z(n14218) );
  XNOR U14479 ( .A(n14217), .B(n14218), .Z(n14219) );
  XOR U14480 ( .A(n14220), .B(n14219), .Z(n14243) );
  XNOR U14481 ( .A(n14244), .B(n14243), .Z(n14245) );
  XNOR U14482 ( .A(n14246), .B(n14245), .Z(n14184) );
  NANDN U14483 ( .A(n14073), .B(n14072), .Z(n14077) );
  NAND U14484 ( .A(n14075), .B(n14074), .Z(n14076) );
  NAND U14485 ( .A(n14077), .B(n14076), .Z(n14235) );
  NANDN U14486 ( .A(n14079), .B(n14078), .Z(n14083) );
  NAND U14487 ( .A(n14081), .B(n14080), .Z(n14082) );
  NAND U14488 ( .A(n14083), .B(n14082), .Z(n14234) );
  XNOR U14489 ( .A(n14234), .B(n14233), .Z(n14236) );
  XOR U14490 ( .A(n14235), .B(n14236), .Z(n14183) );
  XOR U14491 ( .A(n14184), .B(n14183), .Z(n14185) );
  NANDN U14492 ( .A(n14089), .B(n14088), .Z(n14093) );
  NAND U14493 ( .A(n14091), .B(n14090), .Z(n14092) );
  AND U14494 ( .A(n14093), .B(n14092), .Z(n14186) );
  XOR U14495 ( .A(n14185), .B(n14186), .Z(n14297) );
  NANDN U14496 ( .A(n14099), .B(n14098), .Z(n14103) );
  NAND U14497 ( .A(n14101), .B(n14100), .Z(n14102) );
  NAND U14498 ( .A(n14103), .B(n14102), .Z(n14180) );
  NANDN U14499 ( .A(n14109), .B(n14108), .Z(n14113) );
  NAND U14500 ( .A(n14111), .B(n14110), .Z(n14112) );
  NAND U14501 ( .A(n14113), .B(n14112), .Z(n14237) );
  NANDN U14502 ( .A(n14115), .B(n14114), .Z(n14119) );
  NAND U14503 ( .A(n14117), .B(n14116), .Z(n14118) );
  AND U14504 ( .A(n14119), .B(n14118), .Z(n14238) );
  XNOR U14505 ( .A(n14237), .B(n14238), .Z(n14239) );
  XOR U14506 ( .A(n582), .B(a[89]), .Z(n14259) );
  NANDN U14507 ( .A(n14259), .B(n19015), .Z(n14122) );
  NANDN U14508 ( .A(n14120), .B(n19013), .Z(n14121) );
  NAND U14509 ( .A(n14122), .B(n14121), .Z(n14229) );
  NANDN U14510 ( .A(n14123), .B(n18513), .Z(n14125) );
  XOR U14511 ( .A(b[15]), .B(a[95]), .Z(n14262) );
  NANDN U14512 ( .A(n18512), .B(n14262), .Z(n14124) );
  AND U14513 ( .A(n14125), .B(n14124), .Z(n14230) );
  XNOR U14514 ( .A(n14229), .B(n14230), .Z(n14232) );
  XOR U14515 ( .A(n579), .B(a[101]), .Z(n14265) );
  NANDN U14516 ( .A(n14265), .B(n17814), .Z(n14128) );
  NANDN U14517 ( .A(n14126), .B(n17815), .Z(n14127) );
  NAND U14518 ( .A(n14128), .B(n14127), .Z(n14231) );
  XNOR U14519 ( .A(n14232), .B(n14231), .Z(n14225) );
  XNOR U14520 ( .A(b[11]), .B(a[99]), .Z(n14268) );
  OR U14521 ( .A(n14268), .B(n18194), .Z(n14131) );
  NANDN U14522 ( .A(n14129), .B(n18104), .Z(n14130) );
  NAND U14523 ( .A(n14131), .B(n14130), .Z(n14224) );
  XOR U14524 ( .A(n580), .B(a[97]), .Z(n14271) );
  NANDN U14525 ( .A(n14271), .B(n18336), .Z(n14134) );
  NANDN U14526 ( .A(n14132), .B(n18337), .Z(n14133) );
  NAND U14527 ( .A(n14134), .B(n14133), .Z(n14223) );
  XNOR U14528 ( .A(n14224), .B(n14223), .Z(n14226) );
  XNOR U14529 ( .A(n14225), .B(n14226), .Z(n14214) );
  NANDN U14530 ( .A(n577), .B(a[109]), .Z(n14135) );
  XOR U14531 ( .A(n17151), .B(n14135), .Z(n14137) );
  IV U14532 ( .A(a[108]), .Z(n18198) );
  NANDN U14533 ( .A(n18198), .B(n577), .Z(n14136) );
  AND U14534 ( .A(n14137), .B(n14136), .Z(n14189) );
  NAND U14535 ( .A(n19406), .B(n14138), .Z(n14140) );
  XNOR U14536 ( .A(n584), .B(a[81]), .Z(n14277) );
  NANDN U14537 ( .A(n576), .B(n14277), .Z(n14139) );
  NAND U14538 ( .A(n14140), .B(n14139), .Z(n14187) );
  NANDN U14539 ( .A(n585), .B(a[77]), .Z(n14188) );
  XNOR U14540 ( .A(n14187), .B(n14188), .Z(n14190) );
  XNOR U14541 ( .A(n14189), .B(n14190), .Z(n14212) );
  XOR U14542 ( .A(b[23]), .B(a[87]), .Z(n14280) );
  NANDN U14543 ( .A(n19127), .B(n14280), .Z(n14143) );
  NANDN U14544 ( .A(n14141), .B(n19128), .Z(n14142) );
  NAND U14545 ( .A(n14143), .B(n14142), .Z(n14250) );
  NANDN U14546 ( .A(n14144), .B(n17553), .Z(n14146) );
  XOR U14547 ( .A(b[7]), .B(a[103]), .Z(n14283) );
  NAND U14548 ( .A(n14283), .B(n17555), .Z(n14145) );
  NAND U14549 ( .A(n14146), .B(n14145), .Z(n14247) );
  XOR U14550 ( .A(b[25]), .B(a[85]), .Z(n14286) );
  NAND U14551 ( .A(n14286), .B(n19240), .Z(n14149) );
  NANDN U14552 ( .A(n14147), .B(n19242), .Z(n14148) );
  AND U14553 ( .A(n14149), .B(n14148), .Z(n14248) );
  XNOR U14554 ( .A(n14247), .B(n14248), .Z(n14249) );
  XOR U14555 ( .A(n14250), .B(n14249), .Z(n14211) );
  XOR U14556 ( .A(n14214), .B(n14213), .Z(n14240) );
  XNOR U14557 ( .A(n14239), .B(n14240), .Z(n14177) );
  XOR U14558 ( .A(n14178), .B(n14177), .Z(n14179) );
  XNOR U14559 ( .A(n14180), .B(n14179), .Z(n14295) );
  XNOR U14560 ( .A(n14296), .B(n14295), .Z(n14298) );
  XNOR U14561 ( .A(n14297), .B(n14298), .Z(n14292) );
  XOR U14562 ( .A(n14291), .B(n14292), .Z(n14174) );
  NANDN U14563 ( .A(n14155), .B(n14154), .Z(n14159) );
  NANDN U14564 ( .A(n14157), .B(n14156), .Z(n14158) );
  NAND U14565 ( .A(n14159), .B(n14158), .Z(n14172) );
  XNOR U14566 ( .A(n14171), .B(n14172), .Z(n14173) );
  XNOR U14567 ( .A(n14174), .B(n14173), .Z(n14166) );
  XNOR U14568 ( .A(n14165), .B(n14166), .Z(n14167) );
  XNOR U14569 ( .A(n14168), .B(n14167), .Z(n14301) );
  XNOR U14570 ( .A(n14301), .B(sreg[205]), .Z(n14303) );
  NAND U14571 ( .A(n14160), .B(sreg[204]), .Z(n14164) );
  OR U14572 ( .A(n14162), .B(n14161), .Z(n14163) );
  AND U14573 ( .A(n14164), .B(n14163), .Z(n14302) );
  XOR U14574 ( .A(n14303), .B(n14302), .Z(c[205]) );
  NANDN U14575 ( .A(n14166), .B(n14165), .Z(n14170) );
  NAND U14576 ( .A(n14168), .B(n14167), .Z(n14169) );
  NAND U14577 ( .A(n14170), .B(n14169), .Z(n14309) );
  NANDN U14578 ( .A(n14172), .B(n14171), .Z(n14176) );
  NAND U14579 ( .A(n14174), .B(n14173), .Z(n14175) );
  NAND U14580 ( .A(n14176), .B(n14175), .Z(n14306) );
  NAND U14581 ( .A(n14178), .B(n14177), .Z(n14182) );
  NAND U14582 ( .A(n14180), .B(n14179), .Z(n14181) );
  NAND U14583 ( .A(n14182), .B(n14181), .Z(n14432) );
  XNOR U14584 ( .A(n14432), .B(n14433), .Z(n14434) );
  NANDN U14585 ( .A(n14188), .B(n14187), .Z(n14192) );
  NAND U14586 ( .A(n14190), .B(n14189), .Z(n14191) );
  NAND U14587 ( .A(n14192), .B(n14191), .Z(n14331) );
  NANDN U14588 ( .A(n14193), .B(n18832), .Z(n14195) );
  XNOR U14589 ( .A(b[19]), .B(a[92]), .Z(n14380) );
  NANDN U14590 ( .A(n14380), .B(n18834), .Z(n14194) );
  NAND U14591 ( .A(n14195), .B(n14194), .Z(n14341) );
  XOR U14592 ( .A(b[27]), .B(n15134), .Z(n14383) );
  NANDN U14593 ( .A(n14383), .B(n19336), .Z(n14198) );
  NANDN U14594 ( .A(n14196), .B(n19337), .Z(n14197) );
  NAND U14595 ( .A(n14198), .B(n14197), .Z(n14338) );
  XNOR U14596 ( .A(a[106]), .B(b[5]), .Z(n14386) );
  NANDN U14597 ( .A(n14386), .B(n17310), .Z(n14201) );
  NAND U14598 ( .A(n14199), .B(n17311), .Z(n14200) );
  AND U14599 ( .A(n14201), .B(n14200), .Z(n14339) );
  XNOR U14600 ( .A(n14338), .B(n14339), .Z(n14340) );
  XNOR U14601 ( .A(n14341), .B(n14340), .Z(n14329) );
  XNOR U14602 ( .A(b[17]), .B(a[94]), .Z(n14389) );
  NANDN U14603 ( .A(n14389), .B(n18673), .Z(n14204) );
  NAND U14604 ( .A(n14202), .B(n18674), .Z(n14203) );
  NAND U14605 ( .A(n14204), .B(n14203), .Z(n14407) );
  XOR U14606 ( .A(b[31]), .B(n14551), .Z(n14392) );
  NANDN U14607 ( .A(n14392), .B(n19472), .Z(n14207) );
  NANDN U14608 ( .A(n14205), .B(n19473), .Z(n14206) );
  NAND U14609 ( .A(n14207), .B(n14206), .Z(n14404) );
  OR U14610 ( .A(n14208), .B(n16988), .Z(n14210) );
  XOR U14611 ( .A(a[108]), .B(n578), .Z(n14395) );
  NANDN U14612 ( .A(n14395), .B(n16990), .Z(n14209) );
  AND U14613 ( .A(n14210), .B(n14209), .Z(n14405) );
  XNOR U14614 ( .A(n14404), .B(n14405), .Z(n14406) );
  XOR U14615 ( .A(n14407), .B(n14406), .Z(n14328) );
  XNOR U14616 ( .A(n14329), .B(n14328), .Z(n14330) );
  XNOR U14617 ( .A(n14331), .B(n14330), .Z(n14426) );
  NANDN U14618 ( .A(n14212), .B(n14211), .Z(n14216) );
  NANDN U14619 ( .A(n14214), .B(n14213), .Z(n14215) );
  NAND U14620 ( .A(n14216), .B(n14215), .Z(n14427) );
  XNOR U14621 ( .A(n14426), .B(n14427), .Z(n14428) );
  NANDN U14622 ( .A(n14218), .B(n14217), .Z(n14222) );
  NAND U14623 ( .A(n14220), .B(n14219), .Z(n14221) );
  NAND U14624 ( .A(n14222), .B(n14221), .Z(n14321) );
  OR U14625 ( .A(n14224), .B(n14223), .Z(n14228) );
  NANDN U14626 ( .A(n14226), .B(n14225), .Z(n14227) );
  NAND U14627 ( .A(n14228), .B(n14227), .Z(n14319) );
  XNOR U14628 ( .A(n14319), .B(n14318), .Z(n14320) );
  XOR U14629 ( .A(n14321), .B(n14320), .Z(n14429) );
  XOR U14630 ( .A(n14428), .B(n14429), .Z(n14440) );
  NANDN U14631 ( .A(n14238), .B(n14237), .Z(n14242) );
  NANDN U14632 ( .A(n14240), .B(n14239), .Z(n14241) );
  NAND U14633 ( .A(n14242), .B(n14241), .Z(n14423) );
  NANDN U14634 ( .A(n14248), .B(n14247), .Z(n14252) );
  NAND U14635 ( .A(n14250), .B(n14249), .Z(n14251) );
  NAND U14636 ( .A(n14252), .B(n14251), .Z(n14322) );
  NANDN U14637 ( .A(n14254), .B(n14253), .Z(n14258) );
  NAND U14638 ( .A(n14256), .B(n14255), .Z(n14257) );
  AND U14639 ( .A(n14258), .B(n14257), .Z(n14323) );
  XNOR U14640 ( .A(n14322), .B(n14323), .Z(n14324) );
  XNOR U14641 ( .A(b[21]), .B(a[90]), .Z(n14350) );
  NANDN U14642 ( .A(n14350), .B(n19015), .Z(n14261) );
  NANDN U14643 ( .A(n14259), .B(n19013), .Z(n14260) );
  NAND U14644 ( .A(n14261), .B(n14260), .Z(n14416) );
  NAND U14645 ( .A(n14262), .B(n18513), .Z(n14264) );
  XOR U14646 ( .A(b[15]), .B(a[96]), .Z(n14347) );
  NANDN U14647 ( .A(n18512), .B(n14347), .Z(n14263) );
  AND U14648 ( .A(n14264), .B(n14263), .Z(n14417) );
  XNOR U14649 ( .A(n14416), .B(n14417), .Z(n14419) );
  XOR U14650 ( .A(b[9]), .B(n17208), .Z(n14344) );
  NANDN U14651 ( .A(n14344), .B(n17814), .Z(n14267) );
  NANDN U14652 ( .A(n14265), .B(n17815), .Z(n14266) );
  NAND U14653 ( .A(n14267), .B(n14266), .Z(n14418) );
  XNOR U14654 ( .A(n14419), .B(n14418), .Z(n14412) );
  XOR U14655 ( .A(b[11]), .B(n17447), .Z(n14353) );
  OR U14656 ( .A(n14353), .B(n18194), .Z(n14270) );
  NANDN U14657 ( .A(n14268), .B(n18104), .Z(n14269) );
  NAND U14658 ( .A(n14270), .B(n14269), .Z(n14411) );
  XOR U14659 ( .A(n580), .B(a[98]), .Z(n14356) );
  NANDN U14660 ( .A(n14356), .B(n18336), .Z(n14273) );
  NANDN U14661 ( .A(n14271), .B(n18337), .Z(n14272) );
  NAND U14662 ( .A(n14273), .B(n14272), .Z(n14410) );
  XNOR U14663 ( .A(n14411), .B(n14410), .Z(n14413) );
  XNOR U14664 ( .A(n14412), .B(n14413), .Z(n14401) );
  NANDN U14665 ( .A(n577), .B(a[110]), .Z(n14274) );
  XOR U14666 ( .A(n17151), .B(n14274), .Z(n14276) );
  NANDN U14667 ( .A(b[0]), .B(a[109]), .Z(n14275) );
  AND U14668 ( .A(n14276), .B(n14275), .Z(n14376) );
  NAND U14669 ( .A(n19406), .B(n14277), .Z(n14279) );
  XNOR U14670 ( .A(n584), .B(a[82]), .Z(n14359) );
  NANDN U14671 ( .A(n576), .B(n14359), .Z(n14278) );
  NAND U14672 ( .A(n14279), .B(n14278), .Z(n14374) );
  NANDN U14673 ( .A(n585), .B(a[78]), .Z(n14375) );
  XNOR U14674 ( .A(n14374), .B(n14375), .Z(n14377) );
  XNOR U14675 ( .A(n14376), .B(n14377), .Z(n14399) );
  XOR U14676 ( .A(b[23]), .B(a[88]), .Z(n14365) );
  NANDN U14677 ( .A(n19127), .B(n14365), .Z(n14282) );
  NAND U14678 ( .A(n14280), .B(n19128), .Z(n14281) );
  NAND U14679 ( .A(n14282), .B(n14281), .Z(n14335) );
  NAND U14680 ( .A(n14283), .B(n17553), .Z(n14285) );
  XNOR U14681 ( .A(a[104]), .B(b[7]), .Z(n14368) );
  NANDN U14682 ( .A(n14368), .B(n17555), .Z(n14284) );
  NAND U14683 ( .A(n14285), .B(n14284), .Z(n14332) );
  XNOR U14684 ( .A(b[25]), .B(a[86]), .Z(n14371) );
  NANDN U14685 ( .A(n14371), .B(n19240), .Z(n14288) );
  NAND U14686 ( .A(n14286), .B(n19242), .Z(n14287) );
  AND U14687 ( .A(n14288), .B(n14287), .Z(n14333) );
  XNOR U14688 ( .A(n14332), .B(n14333), .Z(n14334) );
  XOR U14689 ( .A(n14335), .B(n14334), .Z(n14398) );
  XOR U14690 ( .A(n14401), .B(n14400), .Z(n14325) );
  XNOR U14691 ( .A(n14324), .B(n14325), .Z(n14420) );
  XOR U14692 ( .A(n14421), .B(n14420), .Z(n14422) );
  XNOR U14693 ( .A(n14423), .B(n14422), .Z(n14438) );
  XNOR U14694 ( .A(n14439), .B(n14438), .Z(n14441) );
  XNOR U14695 ( .A(n14440), .B(n14441), .Z(n14435) );
  XOR U14696 ( .A(n14434), .B(n14435), .Z(n14315) );
  NANDN U14697 ( .A(n14290), .B(n14289), .Z(n14294) );
  NANDN U14698 ( .A(n14292), .B(n14291), .Z(n14293) );
  NAND U14699 ( .A(n14294), .B(n14293), .Z(n14313) );
  OR U14700 ( .A(n14296), .B(n14295), .Z(n14300) );
  OR U14701 ( .A(n14298), .B(n14297), .Z(n14299) );
  AND U14702 ( .A(n14300), .B(n14299), .Z(n14312) );
  XNOR U14703 ( .A(n14313), .B(n14312), .Z(n14314) );
  XNOR U14704 ( .A(n14315), .B(n14314), .Z(n14307) );
  XNOR U14705 ( .A(n14306), .B(n14307), .Z(n14308) );
  XNOR U14706 ( .A(n14309), .B(n14308), .Z(n14444) );
  XNOR U14707 ( .A(n14444), .B(sreg[206]), .Z(n14446) );
  NAND U14708 ( .A(n14301), .B(sreg[205]), .Z(n14305) );
  OR U14709 ( .A(n14303), .B(n14302), .Z(n14304) );
  AND U14710 ( .A(n14305), .B(n14304), .Z(n14445) );
  XOR U14711 ( .A(n14446), .B(n14445), .Z(c[206]) );
  NANDN U14712 ( .A(n14307), .B(n14306), .Z(n14311) );
  NAND U14713 ( .A(n14309), .B(n14308), .Z(n14310) );
  NAND U14714 ( .A(n14311), .B(n14310), .Z(n14452) );
  NANDN U14715 ( .A(n14313), .B(n14312), .Z(n14317) );
  NAND U14716 ( .A(n14315), .B(n14314), .Z(n14316) );
  NAND U14717 ( .A(n14317), .B(n14316), .Z(n14450) );
  NANDN U14718 ( .A(n14323), .B(n14322), .Z(n14327) );
  NANDN U14719 ( .A(n14325), .B(n14324), .Z(n14326) );
  NAND U14720 ( .A(n14327), .B(n14326), .Z(n14567) );
  NANDN U14721 ( .A(n14333), .B(n14332), .Z(n14337) );
  NAND U14722 ( .A(n14335), .B(n14334), .Z(n14336) );
  NAND U14723 ( .A(n14337), .B(n14336), .Z(n14511) );
  NANDN U14724 ( .A(n14339), .B(n14338), .Z(n14343) );
  NAND U14725 ( .A(n14341), .B(n14340), .Z(n14342) );
  AND U14726 ( .A(n14343), .B(n14342), .Z(n14512) );
  XNOR U14727 ( .A(n14511), .B(n14512), .Z(n14513) );
  XNOR U14728 ( .A(n579), .B(a[103]), .Z(n14533) );
  NAND U14729 ( .A(n17814), .B(n14533), .Z(n14346) );
  NANDN U14730 ( .A(n14344), .B(n17815), .Z(n14345) );
  NAND U14731 ( .A(n14346), .B(n14345), .Z(n14497) );
  NAND U14732 ( .A(n14347), .B(n18513), .Z(n14349) );
  XNOR U14733 ( .A(b[15]), .B(a[97]), .Z(n14536) );
  OR U14734 ( .A(n14536), .B(n18512), .Z(n14348) );
  AND U14735 ( .A(n14349), .B(n14348), .Z(n14495) );
  NANDN U14736 ( .A(n14350), .B(n19013), .Z(n14352) );
  XNOR U14737 ( .A(n582), .B(a[91]), .Z(n14539) );
  NAND U14738 ( .A(n14539), .B(n19015), .Z(n14351) );
  AND U14739 ( .A(n14352), .B(n14351), .Z(n14496) );
  XOR U14740 ( .A(n14497), .B(n14498), .Z(n14486) );
  XNOR U14741 ( .A(b[11]), .B(a[101]), .Z(n14542) );
  OR U14742 ( .A(n14542), .B(n18194), .Z(n14355) );
  NANDN U14743 ( .A(n14353), .B(n18104), .Z(n14354) );
  NAND U14744 ( .A(n14355), .B(n14354), .Z(n14484) );
  XOR U14745 ( .A(n580), .B(a[99]), .Z(n14545) );
  NANDN U14746 ( .A(n14545), .B(n18336), .Z(n14358) );
  NANDN U14747 ( .A(n14356), .B(n18337), .Z(n14357) );
  AND U14748 ( .A(n14358), .B(n14357), .Z(n14483) );
  XNOR U14749 ( .A(n14484), .B(n14483), .Z(n14485) );
  XOR U14750 ( .A(n14486), .B(n14485), .Z(n14503) );
  NAND U14751 ( .A(n19406), .B(n14359), .Z(n14361) );
  XNOR U14752 ( .A(b[29]), .B(a[83]), .Z(n14552) );
  OR U14753 ( .A(n14552), .B(n576), .Z(n14360) );
  NAND U14754 ( .A(n14361), .B(n14360), .Z(n14459) );
  NANDN U14755 ( .A(n585), .B(a[79]), .Z(n14460) );
  XNOR U14756 ( .A(n14459), .B(n14460), .Z(n14462) );
  NANDN U14757 ( .A(n577), .B(a[111]), .Z(n14362) );
  XOR U14758 ( .A(n17151), .B(n14362), .Z(n14364) );
  IV U14759 ( .A(a[110]), .Z(n18415) );
  NANDN U14760 ( .A(n18415), .B(n577), .Z(n14363) );
  AND U14761 ( .A(n14364), .B(n14363), .Z(n14461) );
  XOR U14762 ( .A(n14462), .B(n14461), .Z(n14501) );
  XOR U14763 ( .A(b[23]), .B(a[89]), .Z(n14555) );
  NANDN U14764 ( .A(n19127), .B(n14555), .Z(n14367) );
  NAND U14765 ( .A(n14365), .B(n19128), .Z(n14366) );
  NAND U14766 ( .A(n14367), .B(n14366), .Z(n14524) );
  NANDN U14767 ( .A(n14368), .B(n17553), .Z(n14370) );
  XOR U14768 ( .A(b[7]), .B(a[105]), .Z(n14558) );
  NAND U14769 ( .A(n14558), .B(n17555), .Z(n14369) );
  NAND U14770 ( .A(n14370), .B(n14369), .Z(n14521) );
  XOR U14771 ( .A(b[25]), .B(a[87]), .Z(n14561) );
  NAND U14772 ( .A(n14561), .B(n19240), .Z(n14373) );
  NANDN U14773 ( .A(n14371), .B(n19242), .Z(n14372) );
  AND U14774 ( .A(n14373), .B(n14372), .Z(n14522) );
  XNOR U14775 ( .A(n14521), .B(n14522), .Z(n14523) );
  XNOR U14776 ( .A(n14524), .B(n14523), .Z(n14502) );
  XOR U14777 ( .A(n14501), .B(n14502), .Z(n14504) );
  XNOR U14778 ( .A(n14503), .B(n14504), .Z(n14514) );
  XOR U14779 ( .A(n14513), .B(n14514), .Z(n14565) );
  XNOR U14780 ( .A(n14564), .B(n14565), .Z(n14566) );
  XOR U14781 ( .A(n14567), .B(n14566), .Z(n14575) );
  XNOR U14782 ( .A(n14574), .B(n14575), .Z(n14577) );
  NANDN U14783 ( .A(n14375), .B(n14374), .Z(n14379) );
  NAND U14784 ( .A(n14377), .B(n14376), .Z(n14378) );
  NAND U14785 ( .A(n14379), .B(n14378), .Z(n14520) );
  NANDN U14786 ( .A(n14380), .B(n18832), .Z(n14382) );
  XNOR U14787 ( .A(b[19]), .B(a[93]), .Z(n14465) );
  NANDN U14788 ( .A(n14465), .B(n18834), .Z(n14381) );
  NAND U14789 ( .A(n14382), .B(n14381), .Z(n14530) );
  XNOR U14790 ( .A(b[27]), .B(a[85]), .Z(n14468) );
  NANDN U14791 ( .A(n14468), .B(n19336), .Z(n14385) );
  NANDN U14792 ( .A(n14383), .B(n19337), .Z(n14384) );
  NAND U14793 ( .A(n14385), .B(n14384), .Z(n14527) );
  XOR U14794 ( .A(a[107]), .B(b[5]), .Z(n14471) );
  NAND U14795 ( .A(n14471), .B(n17310), .Z(n14388) );
  NANDN U14796 ( .A(n14386), .B(n17311), .Z(n14387) );
  AND U14797 ( .A(n14388), .B(n14387), .Z(n14528) );
  XNOR U14798 ( .A(n14527), .B(n14528), .Z(n14529) );
  XNOR U14799 ( .A(n14530), .B(n14529), .Z(n14518) );
  XOR U14800 ( .A(b[17]), .B(a[95]), .Z(n14474) );
  NAND U14801 ( .A(n14474), .B(n18673), .Z(n14391) );
  NANDN U14802 ( .A(n14389), .B(n18674), .Z(n14390) );
  NAND U14803 ( .A(n14391), .B(n14390), .Z(n14492) );
  XNOR U14804 ( .A(b[31]), .B(a[81]), .Z(n14477) );
  NANDN U14805 ( .A(n14477), .B(n19472), .Z(n14394) );
  NANDN U14806 ( .A(n14392), .B(n19473), .Z(n14393) );
  NAND U14807 ( .A(n14394), .B(n14393), .Z(n14489) );
  OR U14808 ( .A(n14395), .B(n16988), .Z(n14397) );
  XNOR U14809 ( .A(a[109]), .B(b[3]), .Z(n14480) );
  NANDN U14810 ( .A(n14480), .B(n16990), .Z(n14396) );
  AND U14811 ( .A(n14397), .B(n14396), .Z(n14490) );
  XNOR U14812 ( .A(n14489), .B(n14490), .Z(n14491) );
  XOR U14813 ( .A(n14492), .B(n14491), .Z(n14517) );
  XNOR U14814 ( .A(n14518), .B(n14517), .Z(n14519) );
  XNOR U14815 ( .A(n14520), .B(n14519), .Z(n14570) );
  NANDN U14816 ( .A(n14399), .B(n14398), .Z(n14403) );
  NANDN U14817 ( .A(n14401), .B(n14400), .Z(n14402) );
  NAND U14818 ( .A(n14403), .B(n14402), .Z(n14571) );
  XNOR U14819 ( .A(n14570), .B(n14571), .Z(n14572) );
  NANDN U14820 ( .A(n14405), .B(n14404), .Z(n14409) );
  NAND U14821 ( .A(n14407), .B(n14406), .Z(n14408) );
  NAND U14822 ( .A(n14409), .B(n14408), .Z(n14510) );
  OR U14823 ( .A(n14411), .B(n14410), .Z(n14415) );
  NANDN U14824 ( .A(n14413), .B(n14412), .Z(n14414) );
  NAND U14825 ( .A(n14415), .B(n14414), .Z(n14508) );
  XNOR U14826 ( .A(n14508), .B(n14507), .Z(n14509) );
  XOR U14827 ( .A(n14510), .B(n14509), .Z(n14573) );
  XOR U14828 ( .A(n14572), .B(n14573), .Z(n14576) );
  XOR U14829 ( .A(n14577), .B(n14576), .Z(n14581) );
  NAND U14830 ( .A(n14421), .B(n14420), .Z(n14425) );
  NAND U14831 ( .A(n14423), .B(n14422), .Z(n14424) );
  NAND U14832 ( .A(n14425), .B(n14424), .Z(n14578) );
  NANDN U14833 ( .A(n14427), .B(n14426), .Z(n14431) );
  NAND U14834 ( .A(n14429), .B(n14428), .Z(n14430) );
  NAND U14835 ( .A(n14431), .B(n14430), .Z(n14579) );
  XNOR U14836 ( .A(n14578), .B(n14579), .Z(n14580) );
  XNOR U14837 ( .A(n14581), .B(n14580), .Z(n14456) );
  NANDN U14838 ( .A(n14433), .B(n14432), .Z(n14437) );
  NANDN U14839 ( .A(n14435), .B(n14434), .Z(n14436) );
  NAND U14840 ( .A(n14437), .B(n14436), .Z(n14454) );
  OR U14841 ( .A(n14439), .B(n14438), .Z(n14443) );
  OR U14842 ( .A(n14441), .B(n14440), .Z(n14442) );
  AND U14843 ( .A(n14443), .B(n14442), .Z(n14453) );
  XNOR U14844 ( .A(n14454), .B(n14453), .Z(n14455) );
  XNOR U14845 ( .A(n14456), .B(n14455), .Z(n14449) );
  XOR U14846 ( .A(n14450), .B(n14449), .Z(n14451) );
  XNOR U14847 ( .A(n14452), .B(n14451), .Z(n14584) );
  XNOR U14848 ( .A(n14584), .B(sreg[207]), .Z(n14586) );
  NAND U14849 ( .A(n14444), .B(sreg[206]), .Z(n14448) );
  OR U14850 ( .A(n14446), .B(n14445), .Z(n14447) );
  AND U14851 ( .A(n14448), .B(n14447), .Z(n14585) );
  XOR U14852 ( .A(n14586), .B(n14585), .Z(c[207]) );
  NANDN U14853 ( .A(n14454), .B(n14453), .Z(n14458) );
  NANDN U14854 ( .A(n14456), .B(n14455), .Z(n14457) );
  NAND U14855 ( .A(n14458), .B(n14457), .Z(n14590) );
  NANDN U14856 ( .A(n14460), .B(n14459), .Z(n14464) );
  NAND U14857 ( .A(n14462), .B(n14461), .Z(n14463) );
  NAND U14858 ( .A(n14464), .B(n14463), .Z(n14670) );
  NANDN U14859 ( .A(n14465), .B(n18832), .Z(n14467) );
  XOR U14860 ( .A(b[19]), .B(n16590), .Z(n14615) );
  NANDN U14861 ( .A(n14615), .B(n18834), .Z(n14466) );
  NAND U14862 ( .A(n14467), .B(n14466), .Z(n14680) );
  XOR U14863 ( .A(b[27]), .B(n15429), .Z(n14618) );
  NANDN U14864 ( .A(n14618), .B(n19336), .Z(n14470) );
  NANDN U14865 ( .A(n14468), .B(n19337), .Z(n14469) );
  NAND U14866 ( .A(n14470), .B(n14469), .Z(n14677) );
  XNOR U14867 ( .A(a[108]), .B(b[5]), .Z(n14621) );
  NANDN U14868 ( .A(n14621), .B(n17310), .Z(n14473) );
  NAND U14869 ( .A(n14471), .B(n17311), .Z(n14472) );
  AND U14870 ( .A(n14473), .B(n14472), .Z(n14678) );
  XNOR U14871 ( .A(n14677), .B(n14678), .Z(n14679) );
  XNOR U14872 ( .A(n14680), .B(n14679), .Z(n14668) );
  XOR U14873 ( .A(b[17]), .B(a[96]), .Z(n14624) );
  NAND U14874 ( .A(n14624), .B(n18673), .Z(n14476) );
  NAND U14875 ( .A(n14474), .B(n18674), .Z(n14475) );
  NAND U14876 ( .A(n14476), .B(n14475), .Z(n14642) );
  XNOR U14877 ( .A(b[31]), .B(a[82]), .Z(n14627) );
  NANDN U14878 ( .A(n14627), .B(n19472), .Z(n14479) );
  NANDN U14879 ( .A(n14477), .B(n19473), .Z(n14478) );
  NAND U14880 ( .A(n14479), .B(n14478), .Z(n14639) );
  OR U14881 ( .A(n14480), .B(n16988), .Z(n14482) );
  XOR U14882 ( .A(a[110]), .B(n578), .Z(n14630) );
  NANDN U14883 ( .A(n14630), .B(n16990), .Z(n14481) );
  AND U14884 ( .A(n14482), .B(n14481), .Z(n14640) );
  XNOR U14885 ( .A(n14639), .B(n14640), .Z(n14641) );
  XOR U14886 ( .A(n14642), .B(n14641), .Z(n14667) );
  XNOR U14887 ( .A(n14668), .B(n14667), .Z(n14669) );
  XNOR U14888 ( .A(n14670), .B(n14669), .Z(n14713) );
  NANDN U14889 ( .A(n14484), .B(n14483), .Z(n14488) );
  NAND U14890 ( .A(n14486), .B(n14485), .Z(n14487) );
  NAND U14891 ( .A(n14488), .B(n14487), .Z(n14658) );
  NANDN U14892 ( .A(n14490), .B(n14489), .Z(n14494) );
  NAND U14893 ( .A(n14492), .B(n14491), .Z(n14493) );
  NAND U14894 ( .A(n14494), .B(n14493), .Z(n14656) );
  OR U14895 ( .A(n14496), .B(n14495), .Z(n14500) );
  NANDN U14896 ( .A(n14498), .B(n14497), .Z(n14499) );
  NAND U14897 ( .A(n14500), .B(n14499), .Z(n14655) );
  XNOR U14898 ( .A(n14658), .B(n14657), .Z(n14714) );
  XNOR U14899 ( .A(n14713), .B(n14714), .Z(n14715) );
  NANDN U14900 ( .A(n14502), .B(n14501), .Z(n14506) );
  OR U14901 ( .A(n14504), .B(n14503), .Z(n14505) );
  AND U14902 ( .A(n14506), .B(n14505), .Z(n14716) );
  XNOR U14903 ( .A(n14715), .B(n14716), .Z(n14602) );
  NANDN U14904 ( .A(n14512), .B(n14511), .Z(n14516) );
  NANDN U14905 ( .A(n14514), .B(n14513), .Z(n14515) );
  NAND U14906 ( .A(n14516), .B(n14515), .Z(n14722) );
  NANDN U14907 ( .A(n14522), .B(n14521), .Z(n14526) );
  NAND U14908 ( .A(n14524), .B(n14523), .Z(n14525) );
  NAND U14909 ( .A(n14526), .B(n14525), .Z(n14661) );
  NANDN U14910 ( .A(n14528), .B(n14527), .Z(n14532) );
  NAND U14911 ( .A(n14530), .B(n14529), .Z(n14531) );
  AND U14912 ( .A(n14532), .B(n14531), .Z(n14662) );
  XNOR U14913 ( .A(n14661), .B(n14662), .Z(n14663) );
  XOR U14914 ( .A(b[9]), .B(n17716), .Z(n14683) );
  NANDN U14915 ( .A(n14683), .B(n17814), .Z(n14535) );
  NAND U14916 ( .A(n17815), .B(n14533), .Z(n14534) );
  NAND U14917 ( .A(n14535), .B(n14534), .Z(n14647) );
  XNOR U14918 ( .A(b[15]), .B(a[98]), .Z(n14686) );
  OR U14919 ( .A(n14686), .B(n18512), .Z(n14538) );
  NANDN U14920 ( .A(n14536), .B(n18513), .Z(n14537) );
  NAND U14921 ( .A(n14538), .B(n14537), .Z(n14645) );
  XNOR U14922 ( .A(b[21]), .B(a[92]), .Z(n14689) );
  NANDN U14923 ( .A(n14689), .B(n19015), .Z(n14541) );
  NAND U14924 ( .A(n19013), .B(n14539), .Z(n14540) );
  NAND U14925 ( .A(n14541), .B(n14540), .Z(n14646) );
  XNOR U14926 ( .A(n14645), .B(n14646), .Z(n14648) );
  XOR U14927 ( .A(n14647), .B(n14648), .Z(n14636) );
  XOR U14928 ( .A(b[11]), .B(n17208), .Z(n14692) );
  OR U14929 ( .A(n14692), .B(n18194), .Z(n14544) );
  NANDN U14930 ( .A(n14542), .B(n18104), .Z(n14543) );
  NAND U14931 ( .A(n14544), .B(n14543), .Z(n14634) );
  XOR U14932 ( .A(n580), .B(a[100]), .Z(n14695) );
  NANDN U14933 ( .A(n14695), .B(n18336), .Z(n14547) );
  NANDN U14934 ( .A(n14545), .B(n18337), .Z(n14546) );
  AND U14935 ( .A(n14547), .B(n14546), .Z(n14633) );
  XNOR U14936 ( .A(n14634), .B(n14633), .Z(n14635) );
  XNOR U14937 ( .A(n14636), .B(n14635), .Z(n14651) );
  NANDN U14938 ( .A(n577), .B(a[112]), .Z(n14548) );
  XOR U14939 ( .A(n17151), .B(n14548), .Z(n14550) );
  NANDN U14940 ( .A(b[0]), .B(a[111]), .Z(n14549) );
  AND U14941 ( .A(n14550), .B(n14549), .Z(n14612) );
  ANDN U14942 ( .B(b[31]), .A(n14551), .Z(n14609) );
  NANDN U14943 ( .A(n14552), .B(n19406), .Z(n14554) );
  XNOR U14944 ( .A(n584), .B(a[84]), .Z(n14698) );
  NANDN U14945 ( .A(n576), .B(n14698), .Z(n14553) );
  NAND U14946 ( .A(n14554), .B(n14553), .Z(n14610) );
  XOR U14947 ( .A(n14609), .B(n14610), .Z(n14611) );
  XNOR U14948 ( .A(n14612), .B(n14611), .Z(n14649) );
  XOR U14949 ( .A(b[23]), .B(a[90]), .Z(n14704) );
  NANDN U14950 ( .A(n19127), .B(n14704), .Z(n14557) );
  NAND U14951 ( .A(n14555), .B(n19128), .Z(n14556) );
  NAND U14952 ( .A(n14557), .B(n14556), .Z(n14674) );
  NAND U14953 ( .A(n14558), .B(n17553), .Z(n14560) );
  XNOR U14954 ( .A(a[106]), .B(b[7]), .Z(n14707) );
  NANDN U14955 ( .A(n14707), .B(n17555), .Z(n14559) );
  NAND U14956 ( .A(n14560), .B(n14559), .Z(n14671) );
  XOR U14957 ( .A(b[25]), .B(a[88]), .Z(n14710) );
  NAND U14958 ( .A(n14710), .B(n19240), .Z(n14563) );
  NAND U14959 ( .A(n14561), .B(n19242), .Z(n14562) );
  AND U14960 ( .A(n14563), .B(n14562), .Z(n14672) );
  XNOR U14961 ( .A(n14671), .B(n14672), .Z(n14673) );
  XNOR U14962 ( .A(n14674), .B(n14673), .Z(n14650) );
  XOR U14963 ( .A(n14663), .B(n14664), .Z(n14719) );
  XOR U14964 ( .A(n14720), .B(n14719), .Z(n14721) );
  XOR U14965 ( .A(n14722), .B(n14721), .Z(n14600) );
  XNOR U14966 ( .A(n14599), .B(n14600), .Z(n14601) );
  XNOR U14967 ( .A(n14602), .B(n14601), .Z(n14606) );
  NANDN U14968 ( .A(n14565), .B(n14564), .Z(n14569) );
  NAND U14969 ( .A(n14567), .B(n14566), .Z(n14568) );
  NAND U14970 ( .A(n14569), .B(n14568), .Z(n14603) );
  XNOR U14971 ( .A(n14603), .B(n14604), .Z(n14605) );
  XNOR U14972 ( .A(n14606), .B(n14605), .Z(n14596) );
  NANDN U14973 ( .A(n14579), .B(n14578), .Z(n14583) );
  NANDN U14974 ( .A(n14581), .B(n14580), .Z(n14582) );
  NAND U14975 ( .A(n14583), .B(n14582), .Z(n14594) );
  XNOR U14976 ( .A(n14593), .B(n14594), .Z(n14595) );
  XNOR U14977 ( .A(n14596), .B(n14595), .Z(n14589) );
  XOR U14978 ( .A(n14590), .B(n14589), .Z(n14591) );
  XNOR U14979 ( .A(n14592), .B(n14591), .Z(n14725) );
  XNOR U14980 ( .A(n14725), .B(sreg[208]), .Z(n14727) );
  NAND U14981 ( .A(n14584), .B(sreg[207]), .Z(n14588) );
  OR U14982 ( .A(n14586), .B(n14585), .Z(n14587) );
  AND U14983 ( .A(n14588), .B(n14587), .Z(n14726) );
  XOR U14984 ( .A(n14727), .B(n14726), .Z(c[208]) );
  NANDN U14985 ( .A(n14594), .B(n14593), .Z(n14598) );
  NANDN U14986 ( .A(n14596), .B(n14595), .Z(n14597) );
  NAND U14987 ( .A(n14598), .B(n14597), .Z(n14731) );
  NANDN U14988 ( .A(n14604), .B(n14603), .Z(n14608) );
  NANDN U14989 ( .A(n14606), .B(n14605), .Z(n14607) );
  NAND U14990 ( .A(n14608), .B(n14607), .Z(n14737) );
  XNOR U14991 ( .A(n14736), .B(n14737), .Z(n14738) );
  OR U14992 ( .A(n14610), .B(n14609), .Z(n14614) );
  NANDN U14993 ( .A(n14612), .B(n14611), .Z(n14613) );
  NAND U14994 ( .A(n14614), .B(n14613), .Z(n14814) );
  NANDN U14995 ( .A(n14615), .B(n18832), .Z(n14617) );
  XNOR U14996 ( .A(b[19]), .B(a[95]), .Z(n14760) );
  NANDN U14997 ( .A(n14760), .B(n18834), .Z(n14616) );
  NAND U14998 ( .A(n14617), .B(n14616), .Z(n14827) );
  XNOR U14999 ( .A(b[27]), .B(a[87]), .Z(n14763) );
  NANDN U15000 ( .A(n14763), .B(n19336), .Z(n14620) );
  NANDN U15001 ( .A(n14618), .B(n19337), .Z(n14619) );
  NAND U15002 ( .A(n14620), .B(n14619), .Z(n14824) );
  XOR U15003 ( .A(a[109]), .B(b[5]), .Z(n14766) );
  NAND U15004 ( .A(n14766), .B(n17310), .Z(n14623) );
  NANDN U15005 ( .A(n14621), .B(n17311), .Z(n14622) );
  AND U15006 ( .A(n14623), .B(n14622), .Z(n14825) );
  XNOR U15007 ( .A(n14824), .B(n14825), .Z(n14826) );
  XNOR U15008 ( .A(n14827), .B(n14826), .Z(n14813) );
  XNOR U15009 ( .A(b[17]), .B(a[97]), .Z(n14769) );
  NANDN U15010 ( .A(n14769), .B(n18673), .Z(n14626) );
  NAND U15011 ( .A(n14624), .B(n18674), .Z(n14625) );
  NAND U15012 ( .A(n14626), .B(n14625), .Z(n14787) );
  XNOR U15013 ( .A(b[31]), .B(a[83]), .Z(n14772) );
  NANDN U15014 ( .A(n14772), .B(n19472), .Z(n14629) );
  NANDN U15015 ( .A(n14627), .B(n19473), .Z(n14628) );
  NAND U15016 ( .A(n14629), .B(n14628), .Z(n14784) );
  OR U15017 ( .A(n14630), .B(n16988), .Z(n14632) );
  XNOR U15018 ( .A(a[111]), .B(b[3]), .Z(n14775) );
  NANDN U15019 ( .A(n14775), .B(n16990), .Z(n14631) );
  AND U15020 ( .A(n14632), .B(n14631), .Z(n14785) );
  XNOR U15021 ( .A(n14784), .B(n14785), .Z(n14786) );
  XOR U15022 ( .A(n14787), .B(n14786), .Z(n14812) );
  XOR U15023 ( .A(n14813), .B(n14812), .Z(n14815) );
  XNOR U15024 ( .A(n14814), .B(n14815), .Z(n14749) );
  NANDN U15025 ( .A(n14634), .B(n14633), .Z(n14638) );
  NAND U15026 ( .A(n14636), .B(n14635), .Z(n14637) );
  AND U15027 ( .A(n14638), .B(n14637), .Z(n14805) );
  NANDN U15028 ( .A(n14640), .B(n14639), .Z(n14644) );
  NAND U15029 ( .A(n14642), .B(n14641), .Z(n14643) );
  NAND U15030 ( .A(n14644), .B(n14643), .Z(n14803) );
  XNOR U15031 ( .A(n14803), .B(n14802), .Z(n14804) );
  XNOR U15032 ( .A(n14805), .B(n14804), .Z(n14748) );
  XNOR U15033 ( .A(n14749), .B(n14748), .Z(n14751) );
  OR U15034 ( .A(n14650), .B(n14649), .Z(n14654) );
  NANDN U15035 ( .A(n14652), .B(n14651), .Z(n14653) );
  NAND U15036 ( .A(n14654), .B(n14653), .Z(n14750) );
  XOR U15037 ( .A(n14751), .B(n14750), .Z(n14868) );
  OR U15038 ( .A(n14656), .B(n14655), .Z(n14660) );
  NAND U15039 ( .A(n14658), .B(n14657), .Z(n14659) );
  NAND U15040 ( .A(n14660), .B(n14659), .Z(n14867) );
  NANDN U15041 ( .A(n14662), .B(n14661), .Z(n14666) );
  NAND U15042 ( .A(n14664), .B(n14663), .Z(n14665) );
  NAND U15043 ( .A(n14666), .B(n14665), .Z(n14744) );
  NANDN U15044 ( .A(n14672), .B(n14671), .Z(n14676) );
  NAND U15045 ( .A(n14674), .B(n14673), .Z(n14675) );
  NAND U15046 ( .A(n14676), .B(n14675), .Z(n14806) );
  NANDN U15047 ( .A(n14678), .B(n14677), .Z(n14682) );
  NAND U15048 ( .A(n14680), .B(n14679), .Z(n14681) );
  AND U15049 ( .A(n14682), .B(n14681), .Z(n14807) );
  XNOR U15050 ( .A(n14806), .B(n14807), .Z(n14808) );
  XNOR U15051 ( .A(b[9]), .B(a[105]), .Z(n14830) );
  NANDN U15052 ( .A(n14830), .B(n17814), .Z(n14685) );
  NANDN U15053 ( .A(n14683), .B(n17815), .Z(n14684) );
  NAND U15054 ( .A(n14685), .B(n14684), .Z(n14798) );
  NANDN U15055 ( .A(n14686), .B(n18513), .Z(n14688) );
  XOR U15056 ( .A(b[15]), .B(a[99]), .Z(n14833) );
  NANDN U15057 ( .A(n18512), .B(n14833), .Z(n14687) );
  AND U15058 ( .A(n14688), .B(n14687), .Z(n14796) );
  NANDN U15059 ( .A(n14689), .B(n19013), .Z(n14691) );
  XNOR U15060 ( .A(b[21]), .B(a[93]), .Z(n14836) );
  NANDN U15061 ( .A(n14836), .B(n19015), .Z(n14690) );
  AND U15062 ( .A(n14691), .B(n14690), .Z(n14797) );
  XOR U15063 ( .A(n14798), .B(n14799), .Z(n14793) );
  XNOR U15064 ( .A(b[11]), .B(a[103]), .Z(n14839) );
  OR U15065 ( .A(n14839), .B(n18194), .Z(n14694) );
  NANDN U15066 ( .A(n14692), .B(n18104), .Z(n14693) );
  NAND U15067 ( .A(n14694), .B(n14693), .Z(n14791) );
  XOR U15068 ( .A(n580), .B(a[101]), .Z(n14842) );
  NANDN U15069 ( .A(n14842), .B(n18336), .Z(n14697) );
  NANDN U15070 ( .A(n14695), .B(n18337), .Z(n14696) );
  AND U15071 ( .A(n14697), .B(n14696), .Z(n14790) );
  XNOR U15072 ( .A(n14791), .B(n14790), .Z(n14792) );
  XOR U15073 ( .A(n14793), .B(n14792), .Z(n14780) );
  NAND U15074 ( .A(n14698), .B(n19406), .Z(n14700) );
  XNOR U15075 ( .A(n584), .B(a[85]), .Z(n14848) );
  NANDN U15076 ( .A(n576), .B(n14848), .Z(n14699) );
  NAND U15077 ( .A(n14700), .B(n14699), .Z(n14754) );
  NANDN U15078 ( .A(n585), .B(a[81]), .Z(n14755) );
  XNOR U15079 ( .A(n14754), .B(n14755), .Z(n14757) );
  NANDN U15080 ( .A(n577), .B(a[113]), .Z(n14701) );
  XOR U15081 ( .A(n17151), .B(n14701), .Z(n14703) );
  IV U15082 ( .A(a[112]), .Z(n18582) );
  NANDN U15083 ( .A(n18582), .B(n577), .Z(n14702) );
  AND U15084 ( .A(n14703), .B(n14702), .Z(n14756) );
  XOR U15085 ( .A(n14757), .B(n14756), .Z(n14778) );
  XOR U15086 ( .A(b[23]), .B(a[91]), .Z(n14851) );
  NANDN U15087 ( .A(n19127), .B(n14851), .Z(n14706) );
  NAND U15088 ( .A(n14704), .B(n19128), .Z(n14705) );
  NAND U15089 ( .A(n14706), .B(n14705), .Z(n14821) );
  NANDN U15090 ( .A(n14707), .B(n17553), .Z(n14709) );
  XOR U15091 ( .A(a[107]), .B(b[7]), .Z(n14854) );
  NAND U15092 ( .A(n14854), .B(n17555), .Z(n14708) );
  NAND U15093 ( .A(n14709), .B(n14708), .Z(n14818) );
  XOR U15094 ( .A(b[25]), .B(a[89]), .Z(n14857) );
  NAND U15095 ( .A(n14857), .B(n19240), .Z(n14712) );
  NAND U15096 ( .A(n14710), .B(n19242), .Z(n14711) );
  AND U15097 ( .A(n14712), .B(n14711), .Z(n14819) );
  XNOR U15098 ( .A(n14818), .B(n14819), .Z(n14820) );
  XNOR U15099 ( .A(n14821), .B(n14820), .Z(n14779) );
  XOR U15100 ( .A(n14778), .B(n14779), .Z(n14781) );
  XNOR U15101 ( .A(n14780), .B(n14781), .Z(n14809) );
  XNOR U15102 ( .A(n14808), .B(n14809), .Z(n14742) );
  XNOR U15103 ( .A(n14743), .B(n14742), .Z(n14745) );
  XNOR U15104 ( .A(n14744), .B(n14745), .Z(n14866) );
  XOR U15105 ( .A(n14867), .B(n14866), .Z(n14869) );
  NANDN U15106 ( .A(n14714), .B(n14713), .Z(n14718) );
  NAND U15107 ( .A(n14716), .B(n14715), .Z(n14717) );
  NAND U15108 ( .A(n14718), .B(n14717), .Z(n14860) );
  NAND U15109 ( .A(n14720), .B(n14719), .Z(n14724) );
  NAND U15110 ( .A(n14722), .B(n14721), .Z(n14723) );
  NAND U15111 ( .A(n14724), .B(n14723), .Z(n14861) );
  XNOR U15112 ( .A(n14860), .B(n14861), .Z(n14862) );
  XOR U15113 ( .A(n14863), .B(n14862), .Z(n14739) );
  XOR U15114 ( .A(n14738), .B(n14739), .Z(n14730) );
  XOR U15115 ( .A(n14731), .B(n14730), .Z(n14732) );
  XNOR U15116 ( .A(n14733), .B(n14732), .Z(n14872) );
  XNOR U15117 ( .A(n14872), .B(sreg[209]), .Z(n14874) );
  NAND U15118 ( .A(n14725), .B(sreg[208]), .Z(n14729) );
  OR U15119 ( .A(n14727), .B(n14726), .Z(n14728) );
  AND U15120 ( .A(n14729), .B(n14728), .Z(n14873) );
  XOR U15121 ( .A(n14874), .B(n14873), .Z(c[209]) );
  NAND U15122 ( .A(n14731), .B(n14730), .Z(n14735) );
  NAND U15123 ( .A(n14733), .B(n14732), .Z(n14734) );
  NAND U15124 ( .A(n14735), .B(n14734), .Z(n14880) );
  NANDN U15125 ( .A(n14737), .B(n14736), .Z(n14741) );
  NAND U15126 ( .A(n14739), .B(n14738), .Z(n14740) );
  NAND U15127 ( .A(n14741), .B(n14740), .Z(n14877) );
  NAND U15128 ( .A(n14743), .B(n14742), .Z(n14747) );
  NANDN U15129 ( .A(n14745), .B(n14744), .Z(n14746) );
  NAND U15130 ( .A(n14747), .B(n14746), .Z(n15009) );
  NAND U15131 ( .A(n14749), .B(n14748), .Z(n14753) );
  OR U15132 ( .A(n14751), .B(n14750), .Z(n14752) );
  NAND U15133 ( .A(n14753), .B(n14752), .Z(n15010) );
  XNOR U15134 ( .A(n15009), .B(n15010), .Z(n15011) );
  NANDN U15135 ( .A(n14755), .B(n14754), .Z(n14759) );
  NAND U15136 ( .A(n14757), .B(n14756), .Z(n14758) );
  NAND U15137 ( .A(n14759), .B(n14758), .Z(n14964) );
  NANDN U15138 ( .A(n14760), .B(n18832), .Z(n14762) );
  XNOR U15139 ( .A(b[19]), .B(a[96]), .Z(n14931) );
  NANDN U15140 ( .A(n14931), .B(n18834), .Z(n14761) );
  NAND U15141 ( .A(n14762), .B(n14761), .Z(n14976) );
  XNOR U15142 ( .A(b[27]), .B(a[88]), .Z(n14934) );
  NANDN U15143 ( .A(n14934), .B(n19336), .Z(n14765) );
  NANDN U15144 ( .A(n14763), .B(n19337), .Z(n14764) );
  NAND U15145 ( .A(n14765), .B(n14764), .Z(n14973) );
  XNOR U15146 ( .A(a[110]), .B(b[5]), .Z(n14937) );
  NANDN U15147 ( .A(n14937), .B(n17310), .Z(n14768) );
  NAND U15148 ( .A(n14766), .B(n17311), .Z(n14767) );
  AND U15149 ( .A(n14768), .B(n14767), .Z(n14974) );
  XNOR U15150 ( .A(n14973), .B(n14974), .Z(n14975) );
  XNOR U15151 ( .A(n14976), .B(n14975), .Z(n14961) );
  XOR U15152 ( .A(b[17]), .B(a[98]), .Z(n14940) );
  NAND U15153 ( .A(n14940), .B(n18673), .Z(n14771) );
  NANDN U15154 ( .A(n14769), .B(n18674), .Z(n14770) );
  NAND U15155 ( .A(n14771), .B(n14770), .Z(n14915) );
  XOR U15156 ( .A(b[31]), .B(n15134), .Z(n14943) );
  NANDN U15157 ( .A(n14943), .B(n19472), .Z(n14774) );
  NANDN U15158 ( .A(n14772), .B(n19473), .Z(n14773) );
  AND U15159 ( .A(n14774), .B(n14773), .Z(n14913) );
  OR U15160 ( .A(n14775), .B(n16988), .Z(n14777) );
  XOR U15161 ( .A(a[112]), .B(n578), .Z(n14946) );
  NANDN U15162 ( .A(n14946), .B(n16990), .Z(n14776) );
  AND U15163 ( .A(n14777), .B(n14776), .Z(n14914) );
  XOR U15164 ( .A(n14915), .B(n14916), .Z(n14962) );
  XOR U15165 ( .A(n14961), .B(n14962), .Z(n14963) );
  XNOR U15166 ( .A(n14964), .B(n14963), .Z(n14889) );
  NANDN U15167 ( .A(n14779), .B(n14778), .Z(n14783) );
  OR U15168 ( .A(n14781), .B(n14780), .Z(n14782) );
  NAND U15169 ( .A(n14783), .B(n14782), .Z(n14890) );
  XNOR U15170 ( .A(n14889), .B(n14890), .Z(n14891) );
  NANDN U15171 ( .A(n14785), .B(n14784), .Z(n14789) );
  NAND U15172 ( .A(n14787), .B(n14786), .Z(n14788) );
  NAND U15173 ( .A(n14789), .B(n14788), .Z(n14952) );
  NANDN U15174 ( .A(n14791), .B(n14790), .Z(n14795) );
  NAND U15175 ( .A(n14793), .B(n14792), .Z(n14794) );
  NAND U15176 ( .A(n14795), .B(n14794), .Z(n14949) );
  OR U15177 ( .A(n14797), .B(n14796), .Z(n14801) );
  NANDN U15178 ( .A(n14799), .B(n14798), .Z(n14800) );
  NAND U15179 ( .A(n14801), .B(n14800), .Z(n14950) );
  XNOR U15180 ( .A(n14949), .B(n14950), .Z(n14951) );
  XOR U15181 ( .A(n14952), .B(n14951), .Z(n14892) );
  XNOR U15182 ( .A(n14891), .B(n14892), .Z(n15017) );
  NANDN U15183 ( .A(n14807), .B(n14806), .Z(n14811) );
  NANDN U15184 ( .A(n14809), .B(n14808), .Z(n14810) );
  NAND U15185 ( .A(n14811), .B(n14810), .Z(n14898) );
  NANDN U15186 ( .A(n14813), .B(n14812), .Z(n14817) );
  OR U15187 ( .A(n14815), .B(n14814), .Z(n14816) );
  NAND U15188 ( .A(n14817), .B(n14816), .Z(n14896) );
  NANDN U15189 ( .A(n14819), .B(n14818), .Z(n14823) );
  NAND U15190 ( .A(n14821), .B(n14820), .Z(n14822) );
  NAND U15191 ( .A(n14823), .B(n14822), .Z(n14955) );
  NANDN U15192 ( .A(n14825), .B(n14824), .Z(n14829) );
  NAND U15193 ( .A(n14827), .B(n14826), .Z(n14828) );
  AND U15194 ( .A(n14829), .B(n14828), .Z(n14956) );
  XNOR U15195 ( .A(n14955), .B(n14956), .Z(n14957) );
  XOR U15196 ( .A(b[9]), .B(n17690), .Z(n14979) );
  NANDN U15197 ( .A(n14979), .B(n17814), .Z(n14832) );
  NANDN U15198 ( .A(n14830), .B(n17815), .Z(n14831) );
  NAND U15199 ( .A(n14832), .B(n14831), .Z(n14921) );
  NAND U15200 ( .A(n14833), .B(n18513), .Z(n14835) );
  XNOR U15201 ( .A(b[15]), .B(a[100]), .Z(n14982) );
  OR U15202 ( .A(n14982), .B(n18512), .Z(n14834) );
  AND U15203 ( .A(n14835), .B(n14834), .Z(n14919) );
  NANDN U15204 ( .A(n14836), .B(n19013), .Z(n14838) );
  XOR U15205 ( .A(b[21]), .B(n16590), .Z(n14985) );
  NANDN U15206 ( .A(n14985), .B(n19015), .Z(n14837) );
  AND U15207 ( .A(n14838), .B(n14837), .Z(n14920) );
  XOR U15208 ( .A(n14921), .B(n14922), .Z(n14910) );
  XOR U15209 ( .A(b[11]), .B(n17716), .Z(n14988) );
  OR U15210 ( .A(n14988), .B(n18194), .Z(n14841) );
  NANDN U15211 ( .A(n14839), .B(n18104), .Z(n14840) );
  NAND U15212 ( .A(n14841), .B(n14840), .Z(n14908) );
  XOR U15213 ( .A(n580), .B(a[102]), .Z(n14991) );
  NANDN U15214 ( .A(n14991), .B(n18336), .Z(n14844) );
  NANDN U15215 ( .A(n14842), .B(n18337), .Z(n14843) );
  NAND U15216 ( .A(n14844), .B(n14843), .Z(n14907) );
  XOR U15217 ( .A(n14910), .B(n14909), .Z(n14904) );
  NANDN U15218 ( .A(n577), .B(a[114]), .Z(n14845) );
  XOR U15219 ( .A(n17151), .B(n14845), .Z(n14847) );
  NANDN U15220 ( .A(b[0]), .B(a[113]), .Z(n14846) );
  AND U15221 ( .A(n14847), .B(n14846), .Z(n14927) );
  NAND U15222 ( .A(n19406), .B(n14848), .Z(n14850) );
  XOR U15223 ( .A(n584), .B(n15429), .Z(n14994) );
  NANDN U15224 ( .A(n576), .B(n14994), .Z(n14849) );
  NAND U15225 ( .A(n14850), .B(n14849), .Z(n14925) );
  NANDN U15226 ( .A(n585), .B(a[82]), .Z(n14926) );
  XNOR U15227 ( .A(n14925), .B(n14926), .Z(n14928) );
  XNOR U15228 ( .A(n14927), .B(n14928), .Z(n14902) );
  XOR U15229 ( .A(b[23]), .B(a[92]), .Z(n15000) );
  NANDN U15230 ( .A(n19127), .B(n15000), .Z(n14853) );
  NAND U15231 ( .A(n14851), .B(n19128), .Z(n14852) );
  NAND U15232 ( .A(n14853), .B(n14852), .Z(n14970) );
  NAND U15233 ( .A(n14854), .B(n17553), .Z(n14856) );
  XNOR U15234 ( .A(a[108]), .B(b[7]), .Z(n15003) );
  NANDN U15235 ( .A(n15003), .B(n17555), .Z(n14855) );
  NAND U15236 ( .A(n14856), .B(n14855), .Z(n14967) );
  XOR U15237 ( .A(b[25]), .B(a[90]), .Z(n15006) );
  NAND U15238 ( .A(n15006), .B(n19240), .Z(n14859) );
  NAND U15239 ( .A(n14857), .B(n19242), .Z(n14858) );
  AND U15240 ( .A(n14859), .B(n14858), .Z(n14968) );
  XNOR U15241 ( .A(n14967), .B(n14968), .Z(n14969) );
  XOR U15242 ( .A(n14970), .B(n14969), .Z(n14901) );
  XOR U15243 ( .A(n14904), .B(n14903), .Z(n14958) );
  XNOR U15244 ( .A(n14957), .B(n14958), .Z(n14895) );
  XOR U15245 ( .A(n14896), .B(n14895), .Z(n14897) );
  XNOR U15246 ( .A(n14898), .B(n14897), .Z(n15015) );
  XNOR U15247 ( .A(n15016), .B(n15015), .Z(n15018) );
  XNOR U15248 ( .A(n15017), .B(n15018), .Z(n15012) );
  XOR U15249 ( .A(n15011), .B(n15012), .Z(n14886) );
  NANDN U15250 ( .A(n14861), .B(n14860), .Z(n14865) );
  NAND U15251 ( .A(n14863), .B(n14862), .Z(n14864) );
  NAND U15252 ( .A(n14865), .B(n14864), .Z(n14883) );
  NANDN U15253 ( .A(n14867), .B(n14866), .Z(n14871) );
  OR U15254 ( .A(n14869), .B(n14868), .Z(n14870) );
  NAND U15255 ( .A(n14871), .B(n14870), .Z(n14884) );
  XNOR U15256 ( .A(n14883), .B(n14884), .Z(n14885) );
  XNOR U15257 ( .A(n14886), .B(n14885), .Z(n14878) );
  XNOR U15258 ( .A(n14877), .B(n14878), .Z(n14879) );
  XNOR U15259 ( .A(n14880), .B(n14879), .Z(n15021) );
  XNOR U15260 ( .A(n15021), .B(sreg[210]), .Z(n15023) );
  NAND U15261 ( .A(n14872), .B(sreg[209]), .Z(n14876) );
  OR U15262 ( .A(n14874), .B(n14873), .Z(n14875) );
  AND U15263 ( .A(n14876), .B(n14875), .Z(n15022) );
  XOR U15264 ( .A(n15023), .B(n15022), .Z(c[210]) );
  NANDN U15265 ( .A(n14878), .B(n14877), .Z(n14882) );
  NAND U15266 ( .A(n14880), .B(n14879), .Z(n14881) );
  NAND U15267 ( .A(n14882), .B(n14881), .Z(n15029) );
  NANDN U15268 ( .A(n14884), .B(n14883), .Z(n14888) );
  NAND U15269 ( .A(n14886), .B(n14885), .Z(n14887) );
  NAND U15270 ( .A(n14888), .B(n14887), .Z(n15027) );
  NANDN U15271 ( .A(n14890), .B(n14889), .Z(n14894) );
  NANDN U15272 ( .A(n14892), .B(n14891), .Z(n14893) );
  NAND U15273 ( .A(n14894), .B(n14893), .Z(n15163) );
  NAND U15274 ( .A(n14896), .B(n14895), .Z(n14900) );
  NAND U15275 ( .A(n14898), .B(n14897), .Z(n14899) );
  NAND U15276 ( .A(n14900), .B(n14899), .Z(n15164) );
  XNOR U15277 ( .A(n15163), .B(n15164), .Z(n15165) );
  NANDN U15278 ( .A(n14902), .B(n14901), .Z(n14906) );
  NANDN U15279 ( .A(n14904), .B(n14903), .Z(n14905) );
  NAND U15280 ( .A(n14906), .B(n14905), .Z(n15150) );
  OR U15281 ( .A(n14908), .B(n14907), .Z(n14912) );
  NAND U15282 ( .A(n14910), .B(n14909), .Z(n14911) );
  NAND U15283 ( .A(n14912), .B(n14911), .Z(n15088) );
  OR U15284 ( .A(n14914), .B(n14913), .Z(n14918) );
  NANDN U15285 ( .A(n14916), .B(n14915), .Z(n14917) );
  NAND U15286 ( .A(n14918), .B(n14917), .Z(n15087) );
  OR U15287 ( .A(n14920), .B(n14919), .Z(n14924) );
  NANDN U15288 ( .A(n14922), .B(n14921), .Z(n14923) );
  NAND U15289 ( .A(n14924), .B(n14923), .Z(n15086) );
  XOR U15290 ( .A(n15088), .B(n15089), .Z(n15147) );
  NANDN U15291 ( .A(n14926), .B(n14925), .Z(n14930) );
  NAND U15292 ( .A(n14928), .B(n14927), .Z(n14929) );
  NAND U15293 ( .A(n14930), .B(n14929), .Z(n15101) );
  NANDN U15294 ( .A(n14931), .B(n18832), .Z(n14933) );
  XOR U15295 ( .A(b[19]), .B(n17038), .Z(n15044) );
  NANDN U15296 ( .A(n15044), .B(n18834), .Z(n14932) );
  NAND U15297 ( .A(n14933), .B(n14932), .Z(n15113) );
  XNOR U15298 ( .A(b[27]), .B(a[89]), .Z(n15047) );
  NANDN U15299 ( .A(n15047), .B(n19336), .Z(n14936) );
  NANDN U15300 ( .A(n14934), .B(n19337), .Z(n14935) );
  NAND U15301 ( .A(n14936), .B(n14935), .Z(n15110) );
  XOR U15302 ( .A(a[111]), .B(b[5]), .Z(n15050) );
  NAND U15303 ( .A(n15050), .B(n17310), .Z(n14939) );
  NANDN U15304 ( .A(n14937), .B(n17311), .Z(n14938) );
  AND U15305 ( .A(n14939), .B(n14938), .Z(n15111) );
  XNOR U15306 ( .A(n15110), .B(n15111), .Z(n15112) );
  XNOR U15307 ( .A(n15113), .B(n15112), .Z(n15099) );
  XOR U15308 ( .A(b[17]), .B(a[99]), .Z(n15053) );
  NAND U15309 ( .A(n15053), .B(n18673), .Z(n14942) );
  NAND U15310 ( .A(n14940), .B(n18674), .Z(n14941) );
  NAND U15311 ( .A(n14942), .B(n14941), .Z(n15071) );
  XNOR U15312 ( .A(b[31]), .B(a[85]), .Z(n15056) );
  NANDN U15313 ( .A(n15056), .B(n19472), .Z(n14945) );
  NANDN U15314 ( .A(n14943), .B(n19473), .Z(n14944) );
  NAND U15315 ( .A(n14945), .B(n14944), .Z(n15068) );
  OR U15316 ( .A(n14946), .B(n16988), .Z(n14948) );
  XNOR U15317 ( .A(a[113]), .B(b[3]), .Z(n15059) );
  NANDN U15318 ( .A(n15059), .B(n16990), .Z(n14947) );
  AND U15319 ( .A(n14948), .B(n14947), .Z(n15069) );
  XNOR U15320 ( .A(n15068), .B(n15069), .Z(n15070) );
  XOR U15321 ( .A(n15071), .B(n15070), .Z(n15098) );
  XNOR U15322 ( .A(n15099), .B(n15098), .Z(n15100) );
  XNOR U15323 ( .A(n15101), .B(n15100), .Z(n15148) );
  XNOR U15324 ( .A(n15147), .B(n15148), .Z(n15149) );
  XNOR U15325 ( .A(n15150), .B(n15149), .Z(n15160) );
  NANDN U15326 ( .A(n14950), .B(n14949), .Z(n14954) );
  NANDN U15327 ( .A(n14952), .B(n14951), .Z(n14953) );
  NAND U15328 ( .A(n14954), .B(n14953), .Z(n15157) );
  NANDN U15329 ( .A(n14956), .B(n14955), .Z(n14960) );
  NANDN U15330 ( .A(n14958), .B(n14957), .Z(n14959) );
  NAND U15331 ( .A(n14960), .B(n14959), .Z(n15154) );
  OR U15332 ( .A(n14962), .B(n14961), .Z(n14966) );
  NAND U15333 ( .A(n14964), .B(n14963), .Z(n14965) );
  NAND U15334 ( .A(n14966), .B(n14965), .Z(n15151) );
  NANDN U15335 ( .A(n14968), .B(n14967), .Z(n14972) );
  NAND U15336 ( .A(n14970), .B(n14969), .Z(n14971) );
  NAND U15337 ( .A(n14972), .B(n14971), .Z(n15092) );
  NANDN U15338 ( .A(n14974), .B(n14973), .Z(n14978) );
  NAND U15339 ( .A(n14976), .B(n14975), .Z(n14977) );
  AND U15340 ( .A(n14978), .B(n14977), .Z(n15093) );
  XNOR U15341 ( .A(n15092), .B(n15093), .Z(n15094) );
  XNOR U15342 ( .A(b[9]), .B(a[107]), .Z(n15116) );
  NANDN U15343 ( .A(n15116), .B(n17814), .Z(n14981) );
  NANDN U15344 ( .A(n14979), .B(n17815), .Z(n14980) );
  NAND U15345 ( .A(n14981), .B(n14980), .Z(n15076) );
  NANDN U15346 ( .A(n14982), .B(n18513), .Z(n14984) );
  XOR U15347 ( .A(b[15]), .B(a[101]), .Z(n15119) );
  NANDN U15348 ( .A(n18512), .B(n15119), .Z(n14983) );
  AND U15349 ( .A(n14984), .B(n14983), .Z(n15074) );
  NANDN U15350 ( .A(n14985), .B(n19013), .Z(n14987) );
  XNOR U15351 ( .A(b[21]), .B(a[95]), .Z(n15122) );
  NANDN U15352 ( .A(n15122), .B(n19015), .Z(n14986) );
  AND U15353 ( .A(n14987), .B(n14986), .Z(n15075) );
  XOR U15354 ( .A(n15076), .B(n15077), .Z(n15065) );
  XNOR U15355 ( .A(b[11]), .B(a[105]), .Z(n15125) );
  OR U15356 ( .A(n15125), .B(n18194), .Z(n14990) );
  NANDN U15357 ( .A(n14988), .B(n18104), .Z(n14989) );
  NAND U15358 ( .A(n14990), .B(n14989), .Z(n15063) );
  XOR U15359 ( .A(n580), .B(a[103]), .Z(n15128) );
  NANDN U15360 ( .A(n15128), .B(n18336), .Z(n14993) );
  NANDN U15361 ( .A(n14991), .B(n18337), .Z(n14992) );
  AND U15362 ( .A(n14993), .B(n14992), .Z(n15062) );
  XNOR U15363 ( .A(n15063), .B(n15062), .Z(n15064) );
  XOR U15364 ( .A(n15065), .B(n15064), .Z(n15082) );
  NAND U15365 ( .A(n19406), .B(n14994), .Z(n14996) );
  XNOR U15366 ( .A(b[29]), .B(a[87]), .Z(n15135) );
  OR U15367 ( .A(n15135), .B(n576), .Z(n14995) );
  NAND U15368 ( .A(n14996), .B(n14995), .Z(n15038) );
  NANDN U15369 ( .A(n585), .B(a[83]), .Z(n15039) );
  XNOR U15370 ( .A(n15038), .B(n15039), .Z(n15041) );
  NANDN U15371 ( .A(n577), .B(a[115]), .Z(n14997) );
  XOR U15372 ( .A(n17151), .B(n14997), .Z(n14999) );
  IV U15373 ( .A(a[114]), .Z(n18751) );
  NANDN U15374 ( .A(n18751), .B(n577), .Z(n14998) );
  AND U15375 ( .A(n14999), .B(n14998), .Z(n15040) );
  XOR U15376 ( .A(n15041), .B(n15040), .Z(n15080) );
  XOR U15377 ( .A(b[23]), .B(a[93]), .Z(n15138) );
  NANDN U15378 ( .A(n19127), .B(n15138), .Z(n15002) );
  NAND U15379 ( .A(n15000), .B(n19128), .Z(n15001) );
  NAND U15380 ( .A(n15002), .B(n15001), .Z(n15107) );
  NANDN U15381 ( .A(n15003), .B(n17553), .Z(n15005) );
  XOR U15382 ( .A(a[109]), .B(b[7]), .Z(n15141) );
  NAND U15383 ( .A(n15141), .B(n17555), .Z(n15004) );
  NAND U15384 ( .A(n15005), .B(n15004), .Z(n15104) );
  XOR U15385 ( .A(b[25]), .B(a[91]), .Z(n15144) );
  NAND U15386 ( .A(n15144), .B(n19240), .Z(n15008) );
  NAND U15387 ( .A(n15006), .B(n19242), .Z(n15007) );
  AND U15388 ( .A(n15008), .B(n15007), .Z(n15105) );
  XNOR U15389 ( .A(n15104), .B(n15105), .Z(n15106) );
  XNOR U15390 ( .A(n15107), .B(n15106), .Z(n15081) );
  XOR U15391 ( .A(n15080), .B(n15081), .Z(n15083) );
  XNOR U15392 ( .A(n15082), .B(n15083), .Z(n15095) );
  XOR U15393 ( .A(n15094), .B(n15095), .Z(n15152) );
  XNOR U15394 ( .A(n15151), .B(n15152), .Z(n15153) );
  XOR U15395 ( .A(n15154), .B(n15153), .Z(n15158) );
  XNOR U15396 ( .A(n15157), .B(n15158), .Z(n15159) );
  XOR U15397 ( .A(n15160), .B(n15159), .Z(n15166) );
  XOR U15398 ( .A(n15165), .B(n15166), .Z(n15034) );
  NANDN U15399 ( .A(n15010), .B(n15009), .Z(n15014) );
  NANDN U15400 ( .A(n15012), .B(n15011), .Z(n15013) );
  NAND U15401 ( .A(n15014), .B(n15013), .Z(n15033) );
  OR U15402 ( .A(n15016), .B(n15015), .Z(n15020) );
  OR U15403 ( .A(n15018), .B(n15017), .Z(n15019) );
  AND U15404 ( .A(n15020), .B(n15019), .Z(n15032) );
  XNOR U15405 ( .A(n15033), .B(n15032), .Z(n15035) );
  XOR U15406 ( .A(n15034), .B(n15035), .Z(n15026) );
  XOR U15407 ( .A(n15027), .B(n15026), .Z(n15028) );
  XNOR U15408 ( .A(n15029), .B(n15028), .Z(n15169) );
  XNOR U15409 ( .A(n15169), .B(sreg[211]), .Z(n15171) );
  NAND U15410 ( .A(n15021), .B(sreg[210]), .Z(n15025) );
  OR U15411 ( .A(n15023), .B(n15022), .Z(n15024) );
  AND U15412 ( .A(n15025), .B(n15024), .Z(n15170) );
  XOR U15413 ( .A(n15171), .B(n15170), .Z(c[211]) );
  NAND U15414 ( .A(n15027), .B(n15026), .Z(n15031) );
  NAND U15415 ( .A(n15029), .B(n15028), .Z(n15030) );
  NAND U15416 ( .A(n15031), .B(n15030), .Z(n15177) );
  NANDN U15417 ( .A(n15033), .B(n15032), .Z(n15037) );
  NAND U15418 ( .A(n15035), .B(n15034), .Z(n15036) );
  NAND U15419 ( .A(n15037), .B(n15036), .Z(n15175) );
  NANDN U15420 ( .A(n15039), .B(n15038), .Z(n15043) );
  NAND U15421 ( .A(n15041), .B(n15040), .Z(n15042) );
  NAND U15422 ( .A(n15043), .B(n15042), .Z(n15261) );
  NANDN U15423 ( .A(n15044), .B(n18832), .Z(n15046) );
  XNOR U15424 ( .A(b[19]), .B(a[98]), .Z(n15204) );
  NANDN U15425 ( .A(n15204), .B(n18834), .Z(n15045) );
  NAND U15426 ( .A(n15046), .B(n15045), .Z(n15271) );
  XNOR U15427 ( .A(b[27]), .B(a[90]), .Z(n15207) );
  NANDN U15428 ( .A(n15207), .B(n19336), .Z(n15049) );
  NANDN U15429 ( .A(n15047), .B(n19337), .Z(n15048) );
  NAND U15430 ( .A(n15049), .B(n15048), .Z(n15268) );
  XNOR U15431 ( .A(a[112]), .B(b[5]), .Z(n15210) );
  NANDN U15432 ( .A(n15210), .B(n17310), .Z(n15052) );
  NAND U15433 ( .A(n15050), .B(n17311), .Z(n15051) );
  AND U15434 ( .A(n15052), .B(n15051), .Z(n15269) );
  XNOR U15435 ( .A(n15268), .B(n15269), .Z(n15270) );
  XNOR U15436 ( .A(n15271), .B(n15270), .Z(n15259) );
  XNOR U15437 ( .A(b[17]), .B(a[100]), .Z(n15213) );
  NANDN U15438 ( .A(n15213), .B(n18673), .Z(n15055) );
  NAND U15439 ( .A(n15053), .B(n18674), .Z(n15054) );
  NAND U15440 ( .A(n15055), .B(n15054), .Z(n15231) );
  XOR U15441 ( .A(b[31]), .B(n15429), .Z(n15216) );
  NANDN U15442 ( .A(n15216), .B(n19472), .Z(n15058) );
  NANDN U15443 ( .A(n15056), .B(n19473), .Z(n15057) );
  NAND U15444 ( .A(n15058), .B(n15057), .Z(n15228) );
  OR U15445 ( .A(n15059), .B(n16988), .Z(n15061) );
  XOR U15446 ( .A(a[114]), .B(n578), .Z(n15219) );
  NANDN U15447 ( .A(n15219), .B(n16990), .Z(n15060) );
  AND U15448 ( .A(n15061), .B(n15060), .Z(n15229) );
  XNOR U15449 ( .A(n15228), .B(n15229), .Z(n15230) );
  XOR U15450 ( .A(n15231), .B(n15230), .Z(n15258) );
  XNOR U15451 ( .A(n15259), .B(n15258), .Z(n15260) );
  XNOR U15452 ( .A(n15261), .B(n15260), .Z(n15304) );
  NANDN U15453 ( .A(n15063), .B(n15062), .Z(n15067) );
  NAND U15454 ( .A(n15065), .B(n15064), .Z(n15066) );
  NAND U15455 ( .A(n15067), .B(n15066), .Z(n15249) );
  NANDN U15456 ( .A(n15069), .B(n15068), .Z(n15073) );
  NAND U15457 ( .A(n15071), .B(n15070), .Z(n15072) );
  NAND U15458 ( .A(n15073), .B(n15072), .Z(n15247) );
  OR U15459 ( .A(n15075), .B(n15074), .Z(n15079) );
  NANDN U15460 ( .A(n15077), .B(n15076), .Z(n15078) );
  NAND U15461 ( .A(n15079), .B(n15078), .Z(n15246) );
  XNOR U15462 ( .A(n15249), .B(n15248), .Z(n15305) );
  XOR U15463 ( .A(n15304), .B(n15305), .Z(n15307) );
  NANDN U15464 ( .A(n15081), .B(n15080), .Z(n15085) );
  OR U15465 ( .A(n15083), .B(n15082), .Z(n15084) );
  NAND U15466 ( .A(n15085), .B(n15084), .Z(n15306) );
  XOR U15467 ( .A(n15307), .B(n15306), .Z(n15194) );
  OR U15468 ( .A(n15087), .B(n15086), .Z(n15091) );
  NANDN U15469 ( .A(n15089), .B(n15088), .Z(n15090) );
  NAND U15470 ( .A(n15091), .B(n15090), .Z(n15193) );
  NANDN U15471 ( .A(n15093), .B(n15092), .Z(n15097) );
  NANDN U15472 ( .A(n15095), .B(n15094), .Z(n15096) );
  NAND U15473 ( .A(n15097), .B(n15096), .Z(n15312) );
  NANDN U15474 ( .A(n15099), .B(n15098), .Z(n15103) );
  NAND U15475 ( .A(n15101), .B(n15100), .Z(n15102) );
  NAND U15476 ( .A(n15103), .B(n15102), .Z(n15311) );
  NANDN U15477 ( .A(n15105), .B(n15104), .Z(n15109) );
  NAND U15478 ( .A(n15107), .B(n15106), .Z(n15108) );
  NAND U15479 ( .A(n15109), .B(n15108), .Z(n15252) );
  NANDN U15480 ( .A(n15111), .B(n15110), .Z(n15115) );
  NAND U15481 ( .A(n15113), .B(n15112), .Z(n15114) );
  AND U15482 ( .A(n15115), .B(n15114), .Z(n15253) );
  XNOR U15483 ( .A(n15252), .B(n15253), .Z(n15254) );
  XOR U15484 ( .A(a[108]), .B(n579), .Z(n15274) );
  NANDN U15485 ( .A(n15274), .B(n17814), .Z(n15118) );
  NANDN U15486 ( .A(n15116), .B(n17815), .Z(n15117) );
  NAND U15487 ( .A(n15118), .B(n15117), .Z(n15236) );
  NAND U15488 ( .A(n15119), .B(n18513), .Z(n15121) );
  XNOR U15489 ( .A(b[15]), .B(a[102]), .Z(n15277) );
  OR U15490 ( .A(n15277), .B(n18512), .Z(n15120) );
  AND U15491 ( .A(n15121), .B(n15120), .Z(n15234) );
  NANDN U15492 ( .A(n15122), .B(n19013), .Z(n15124) );
  XNOR U15493 ( .A(b[21]), .B(a[96]), .Z(n15280) );
  NANDN U15494 ( .A(n15280), .B(n19015), .Z(n15123) );
  AND U15495 ( .A(n15124), .B(n15123), .Z(n15235) );
  XOR U15496 ( .A(n15236), .B(n15237), .Z(n15225) );
  XOR U15497 ( .A(b[11]), .B(n17690), .Z(n15283) );
  OR U15498 ( .A(n15283), .B(n18194), .Z(n15127) );
  NANDN U15499 ( .A(n15125), .B(n18104), .Z(n15126) );
  NAND U15500 ( .A(n15127), .B(n15126), .Z(n15223) );
  XOR U15501 ( .A(n580), .B(a[104]), .Z(n15286) );
  NANDN U15502 ( .A(n15286), .B(n18336), .Z(n15130) );
  NANDN U15503 ( .A(n15128), .B(n18337), .Z(n15129) );
  AND U15504 ( .A(n15130), .B(n15129), .Z(n15222) );
  XNOR U15505 ( .A(n15223), .B(n15222), .Z(n15224) );
  XOR U15506 ( .A(n15225), .B(n15224), .Z(n15242) );
  NANDN U15507 ( .A(n577), .B(a[116]), .Z(n15131) );
  XOR U15508 ( .A(n17151), .B(n15131), .Z(n15133) );
  IV U15509 ( .A(a[115]), .Z(n19022) );
  NANDN U15510 ( .A(n19022), .B(n577), .Z(n15132) );
  AND U15511 ( .A(n15133), .B(n15132), .Z(n15201) );
  ANDN U15512 ( .B(b[31]), .A(n15134), .Z(n15198) );
  NANDN U15513 ( .A(n15135), .B(n19406), .Z(n15137) );
  XNOR U15514 ( .A(n584), .B(a[88]), .Z(n15292) );
  NANDN U15515 ( .A(n576), .B(n15292), .Z(n15136) );
  NAND U15516 ( .A(n15137), .B(n15136), .Z(n15199) );
  XOR U15517 ( .A(n15198), .B(n15199), .Z(n15200) );
  XNOR U15518 ( .A(n15201), .B(n15200), .Z(n15240) );
  XNOR U15519 ( .A(b[23]), .B(a[94]), .Z(n15295) );
  OR U15520 ( .A(n15295), .B(n19127), .Z(n15140) );
  NAND U15521 ( .A(n15138), .B(n19128), .Z(n15139) );
  NAND U15522 ( .A(n15140), .B(n15139), .Z(n15265) );
  NAND U15523 ( .A(n15141), .B(n17553), .Z(n15143) );
  XNOR U15524 ( .A(a[110]), .B(b[7]), .Z(n15298) );
  NANDN U15525 ( .A(n15298), .B(n17555), .Z(n15142) );
  NAND U15526 ( .A(n15143), .B(n15142), .Z(n15262) );
  XOR U15527 ( .A(b[25]), .B(a[92]), .Z(n15301) );
  NAND U15528 ( .A(n15301), .B(n19240), .Z(n15146) );
  NAND U15529 ( .A(n15144), .B(n19242), .Z(n15145) );
  AND U15530 ( .A(n15146), .B(n15145), .Z(n15263) );
  XNOR U15531 ( .A(n15262), .B(n15263), .Z(n15264) );
  XNOR U15532 ( .A(n15265), .B(n15264), .Z(n15241) );
  XNOR U15533 ( .A(n15240), .B(n15241), .Z(n15243) );
  XNOR U15534 ( .A(n15242), .B(n15243), .Z(n15255) );
  XNOR U15535 ( .A(n15254), .B(n15255), .Z(n15310) );
  XNOR U15536 ( .A(n15311), .B(n15310), .Z(n15313) );
  XNOR U15537 ( .A(n15312), .B(n15313), .Z(n15192) );
  XOR U15538 ( .A(n15193), .B(n15192), .Z(n15195) );
  NANDN U15539 ( .A(n15152), .B(n15151), .Z(n15156) );
  NAND U15540 ( .A(n15154), .B(n15153), .Z(n15155) );
  AND U15541 ( .A(n15156), .B(n15155), .Z(n15186) );
  XNOR U15542 ( .A(n15187), .B(n15186), .Z(n15188) );
  XOR U15543 ( .A(n15189), .B(n15188), .Z(n15182) );
  NANDN U15544 ( .A(n15158), .B(n15157), .Z(n15162) );
  NAND U15545 ( .A(n15160), .B(n15159), .Z(n15161) );
  NAND U15546 ( .A(n15162), .B(n15161), .Z(n15180) );
  NANDN U15547 ( .A(n15164), .B(n15163), .Z(n15168) );
  NAND U15548 ( .A(n15166), .B(n15165), .Z(n15167) );
  AND U15549 ( .A(n15168), .B(n15167), .Z(n15181) );
  XNOR U15550 ( .A(n15180), .B(n15181), .Z(n15183) );
  XOR U15551 ( .A(n15182), .B(n15183), .Z(n15174) );
  XOR U15552 ( .A(n15175), .B(n15174), .Z(n15176) );
  XNOR U15553 ( .A(n15177), .B(n15176), .Z(n15316) );
  XNOR U15554 ( .A(n15316), .B(sreg[212]), .Z(n15318) );
  NAND U15555 ( .A(n15169), .B(sreg[211]), .Z(n15173) );
  OR U15556 ( .A(n15171), .B(n15170), .Z(n15172) );
  AND U15557 ( .A(n15173), .B(n15172), .Z(n15317) );
  XOR U15558 ( .A(n15318), .B(n15317), .Z(c[212]) );
  NAND U15559 ( .A(n15175), .B(n15174), .Z(n15179) );
  NAND U15560 ( .A(n15177), .B(n15176), .Z(n15178) );
  NAND U15561 ( .A(n15179), .B(n15178), .Z(n15324) );
  NANDN U15562 ( .A(n15181), .B(n15180), .Z(n15185) );
  NAND U15563 ( .A(n15183), .B(n15182), .Z(n15184) );
  NAND U15564 ( .A(n15185), .B(n15184), .Z(n15322) );
  NANDN U15565 ( .A(n15187), .B(n15186), .Z(n15191) );
  NAND U15566 ( .A(n15189), .B(n15188), .Z(n15190) );
  NAND U15567 ( .A(n15191), .B(n15190), .Z(n15327) );
  NANDN U15568 ( .A(n15193), .B(n15192), .Z(n15197) );
  OR U15569 ( .A(n15195), .B(n15194), .Z(n15196) );
  NAND U15570 ( .A(n15197), .B(n15196), .Z(n15328) );
  XNOR U15571 ( .A(n15327), .B(n15328), .Z(n15329) );
  OR U15572 ( .A(n15199), .B(n15198), .Z(n15203) );
  NANDN U15573 ( .A(n15201), .B(n15200), .Z(n15202) );
  NAND U15574 ( .A(n15203), .B(n15202), .Z(n15395) );
  NANDN U15575 ( .A(n15204), .B(n18832), .Z(n15206) );
  XNOR U15576 ( .A(b[19]), .B(a[99]), .Z(n15339) );
  NANDN U15577 ( .A(n15339), .B(n18834), .Z(n15205) );
  NAND U15578 ( .A(n15206), .B(n15205), .Z(n15408) );
  XNOR U15579 ( .A(b[27]), .B(a[91]), .Z(n15342) );
  NANDN U15580 ( .A(n15342), .B(n19336), .Z(n15209) );
  NANDN U15581 ( .A(n15207), .B(n19337), .Z(n15208) );
  NAND U15582 ( .A(n15209), .B(n15208), .Z(n15405) );
  XOR U15583 ( .A(a[113]), .B(b[5]), .Z(n15345) );
  NAND U15584 ( .A(n15345), .B(n17310), .Z(n15212) );
  NANDN U15585 ( .A(n15210), .B(n17311), .Z(n15211) );
  AND U15586 ( .A(n15212), .B(n15211), .Z(n15406) );
  XNOR U15587 ( .A(n15405), .B(n15406), .Z(n15407) );
  XNOR U15588 ( .A(n15408), .B(n15407), .Z(n15394) );
  XOR U15589 ( .A(b[17]), .B(a[101]), .Z(n15348) );
  NAND U15590 ( .A(n15348), .B(n18673), .Z(n15215) );
  NANDN U15591 ( .A(n15213), .B(n18674), .Z(n15214) );
  NAND U15592 ( .A(n15215), .B(n15214), .Z(n15366) );
  XNOR U15593 ( .A(b[31]), .B(a[87]), .Z(n15351) );
  NANDN U15594 ( .A(n15351), .B(n19472), .Z(n15218) );
  NANDN U15595 ( .A(n15216), .B(n19473), .Z(n15217) );
  NAND U15596 ( .A(n15218), .B(n15217), .Z(n15363) );
  OR U15597 ( .A(n15219), .B(n16988), .Z(n15221) );
  XOR U15598 ( .A(a[115]), .B(n578), .Z(n15354) );
  NANDN U15599 ( .A(n15354), .B(n16990), .Z(n15220) );
  AND U15600 ( .A(n15221), .B(n15220), .Z(n15364) );
  XNOR U15601 ( .A(n15363), .B(n15364), .Z(n15365) );
  XOR U15602 ( .A(n15366), .B(n15365), .Z(n15393) );
  XOR U15603 ( .A(n15394), .B(n15393), .Z(n15396) );
  XNOR U15604 ( .A(n15395), .B(n15396), .Z(n15442) );
  NANDN U15605 ( .A(n15223), .B(n15222), .Z(n15227) );
  NAND U15606 ( .A(n15225), .B(n15224), .Z(n15226) );
  NAND U15607 ( .A(n15227), .B(n15226), .Z(n15384) );
  NANDN U15608 ( .A(n15229), .B(n15228), .Z(n15233) );
  NAND U15609 ( .A(n15231), .B(n15230), .Z(n15232) );
  NAND U15610 ( .A(n15233), .B(n15232), .Z(n15382) );
  OR U15611 ( .A(n15235), .B(n15234), .Z(n15239) );
  NANDN U15612 ( .A(n15237), .B(n15236), .Z(n15238) );
  NAND U15613 ( .A(n15239), .B(n15238), .Z(n15381) );
  XNOR U15614 ( .A(n15384), .B(n15383), .Z(n15443) );
  XNOR U15615 ( .A(n15442), .B(n15443), .Z(n15444) );
  OR U15616 ( .A(n15241), .B(n15240), .Z(n15245) );
  OR U15617 ( .A(n15243), .B(n15242), .Z(n15244) );
  NAND U15618 ( .A(n15245), .B(n15244), .Z(n15445) );
  XNOR U15619 ( .A(n15444), .B(n15445), .Z(n15462) );
  OR U15620 ( .A(n15247), .B(n15246), .Z(n15251) );
  NAND U15621 ( .A(n15249), .B(n15248), .Z(n15250) );
  NAND U15622 ( .A(n15251), .B(n15250), .Z(n15461) );
  NANDN U15623 ( .A(n15253), .B(n15252), .Z(n15257) );
  NANDN U15624 ( .A(n15255), .B(n15254), .Z(n15256) );
  NAND U15625 ( .A(n15257), .B(n15256), .Z(n15450) );
  NANDN U15626 ( .A(n15263), .B(n15262), .Z(n15267) );
  NAND U15627 ( .A(n15265), .B(n15264), .Z(n15266) );
  NAND U15628 ( .A(n15267), .B(n15266), .Z(n15387) );
  NANDN U15629 ( .A(n15269), .B(n15268), .Z(n15273) );
  NAND U15630 ( .A(n15271), .B(n15270), .Z(n15272) );
  AND U15631 ( .A(n15273), .B(n15272), .Z(n15388) );
  XNOR U15632 ( .A(n15387), .B(n15388), .Z(n15389) );
  XNOR U15633 ( .A(a[109]), .B(b[9]), .Z(n15411) );
  NANDN U15634 ( .A(n15411), .B(n17814), .Z(n15276) );
  NANDN U15635 ( .A(n15274), .B(n17815), .Z(n15275) );
  NAND U15636 ( .A(n15276), .B(n15275), .Z(n15371) );
  NANDN U15637 ( .A(n15277), .B(n18513), .Z(n15279) );
  XOR U15638 ( .A(b[15]), .B(a[103]), .Z(n15414) );
  NANDN U15639 ( .A(n18512), .B(n15414), .Z(n15278) );
  AND U15640 ( .A(n15279), .B(n15278), .Z(n15369) );
  NANDN U15641 ( .A(n15280), .B(n19013), .Z(n15282) );
  XOR U15642 ( .A(b[21]), .B(n17038), .Z(n15417) );
  NANDN U15643 ( .A(n15417), .B(n19015), .Z(n15281) );
  AND U15644 ( .A(n15282), .B(n15281), .Z(n15370) );
  XOR U15645 ( .A(n15371), .B(n15372), .Z(n15360) );
  XNOR U15646 ( .A(b[11]), .B(a[107]), .Z(n15420) );
  OR U15647 ( .A(n15420), .B(n18194), .Z(n15285) );
  NANDN U15648 ( .A(n15283), .B(n18104), .Z(n15284) );
  NAND U15649 ( .A(n15285), .B(n15284), .Z(n15358) );
  XOR U15650 ( .A(n580), .B(a[105]), .Z(n15423) );
  NANDN U15651 ( .A(n15423), .B(n18336), .Z(n15288) );
  NANDN U15652 ( .A(n15286), .B(n18337), .Z(n15287) );
  AND U15653 ( .A(n15288), .B(n15287), .Z(n15357) );
  XNOR U15654 ( .A(n15358), .B(n15357), .Z(n15359) );
  XOR U15655 ( .A(n15360), .B(n15359), .Z(n15377) );
  NANDN U15656 ( .A(n577), .B(a[117]), .Z(n15289) );
  XOR U15657 ( .A(n17151), .B(n15289), .Z(n15291) );
  IV U15658 ( .A(a[116]), .Z(n18950) );
  NANDN U15659 ( .A(n18950), .B(n577), .Z(n15290) );
  AND U15660 ( .A(n15291), .B(n15290), .Z(n15335) );
  NAND U15661 ( .A(n15292), .B(n19406), .Z(n15294) );
  XNOR U15662 ( .A(b[29]), .B(a[89]), .Z(n15430) );
  OR U15663 ( .A(n15430), .B(n576), .Z(n15293) );
  NAND U15664 ( .A(n15294), .B(n15293), .Z(n15333) );
  NANDN U15665 ( .A(n585), .B(a[85]), .Z(n15334) );
  XNOR U15666 ( .A(n15333), .B(n15334), .Z(n15336) );
  XOR U15667 ( .A(n15335), .B(n15336), .Z(n15375) );
  XOR U15668 ( .A(b[23]), .B(a[95]), .Z(n15433) );
  NANDN U15669 ( .A(n19127), .B(n15433), .Z(n15297) );
  NANDN U15670 ( .A(n15295), .B(n19128), .Z(n15296) );
  NAND U15671 ( .A(n15297), .B(n15296), .Z(n15402) );
  NANDN U15672 ( .A(n15298), .B(n17553), .Z(n15300) );
  XOR U15673 ( .A(a[111]), .B(b[7]), .Z(n15436) );
  NAND U15674 ( .A(n15436), .B(n17555), .Z(n15299) );
  NAND U15675 ( .A(n15300), .B(n15299), .Z(n15399) );
  XOR U15676 ( .A(b[25]), .B(a[93]), .Z(n15439) );
  NAND U15677 ( .A(n15439), .B(n19240), .Z(n15303) );
  NAND U15678 ( .A(n15301), .B(n19242), .Z(n15302) );
  AND U15679 ( .A(n15303), .B(n15302), .Z(n15400) );
  XNOR U15680 ( .A(n15399), .B(n15400), .Z(n15401) );
  XNOR U15681 ( .A(n15402), .B(n15401), .Z(n15376) );
  XOR U15682 ( .A(n15375), .B(n15376), .Z(n15378) );
  XNOR U15683 ( .A(n15377), .B(n15378), .Z(n15390) );
  XNOR U15684 ( .A(n15389), .B(n15390), .Z(n15448) );
  XNOR U15685 ( .A(n15449), .B(n15448), .Z(n15451) );
  XNOR U15686 ( .A(n15450), .B(n15451), .Z(n15460) );
  XOR U15687 ( .A(n15461), .B(n15460), .Z(n15463) );
  NANDN U15688 ( .A(n15305), .B(n15304), .Z(n15309) );
  OR U15689 ( .A(n15307), .B(n15306), .Z(n15308) );
  NAND U15690 ( .A(n15309), .B(n15308), .Z(n15454) );
  NAND U15691 ( .A(n15311), .B(n15310), .Z(n15315) );
  NANDN U15692 ( .A(n15313), .B(n15312), .Z(n15314) );
  NAND U15693 ( .A(n15315), .B(n15314), .Z(n15455) );
  XNOR U15694 ( .A(n15454), .B(n15455), .Z(n15456) );
  XOR U15695 ( .A(n15457), .B(n15456), .Z(n15330) );
  XOR U15696 ( .A(n15329), .B(n15330), .Z(n15321) );
  XOR U15697 ( .A(n15322), .B(n15321), .Z(n15323) );
  XNOR U15698 ( .A(n15324), .B(n15323), .Z(n15466) );
  XNOR U15699 ( .A(n15466), .B(sreg[213]), .Z(n15468) );
  NAND U15700 ( .A(n15316), .B(sreg[212]), .Z(n15320) );
  OR U15701 ( .A(n15318), .B(n15317), .Z(n15319) );
  AND U15702 ( .A(n15320), .B(n15319), .Z(n15467) );
  XOR U15703 ( .A(n15468), .B(n15467), .Z(c[213]) );
  NAND U15704 ( .A(n15322), .B(n15321), .Z(n15326) );
  NAND U15705 ( .A(n15324), .B(n15323), .Z(n15325) );
  NAND U15706 ( .A(n15326), .B(n15325), .Z(n15474) );
  NANDN U15707 ( .A(n15328), .B(n15327), .Z(n15332) );
  NAND U15708 ( .A(n15330), .B(n15329), .Z(n15331) );
  NAND U15709 ( .A(n15332), .B(n15331), .Z(n15472) );
  NANDN U15710 ( .A(n15334), .B(n15333), .Z(n15338) );
  NAND U15711 ( .A(n15336), .B(n15335), .Z(n15337) );
  NAND U15712 ( .A(n15338), .B(n15337), .Z(n15546) );
  NANDN U15713 ( .A(n15339), .B(n18832), .Z(n15341) );
  XOR U15714 ( .A(b[19]), .B(n17447), .Z(n15513) );
  NANDN U15715 ( .A(n15513), .B(n18834), .Z(n15340) );
  NAND U15716 ( .A(n15341), .B(n15340), .Z(n15558) );
  XNOR U15717 ( .A(b[27]), .B(a[92]), .Z(n15516) );
  NANDN U15718 ( .A(n15516), .B(n19336), .Z(n15344) );
  NANDN U15719 ( .A(n15342), .B(n19337), .Z(n15343) );
  NAND U15720 ( .A(n15344), .B(n15343), .Z(n15555) );
  XNOR U15721 ( .A(a[114]), .B(b[5]), .Z(n15519) );
  NANDN U15722 ( .A(n15519), .B(n17310), .Z(n15347) );
  NAND U15723 ( .A(n15345), .B(n17311), .Z(n15346) );
  AND U15724 ( .A(n15347), .B(n15346), .Z(n15556) );
  XNOR U15725 ( .A(n15555), .B(n15556), .Z(n15557) );
  XNOR U15726 ( .A(n15558), .B(n15557), .Z(n15543) );
  XNOR U15727 ( .A(b[17]), .B(a[102]), .Z(n15522) );
  NANDN U15728 ( .A(n15522), .B(n18673), .Z(n15350) );
  NAND U15729 ( .A(n15348), .B(n18674), .Z(n15349) );
  NAND U15730 ( .A(n15350), .B(n15349), .Z(n15497) );
  XNOR U15731 ( .A(b[31]), .B(a[88]), .Z(n15525) );
  NANDN U15732 ( .A(n15525), .B(n19472), .Z(n15353) );
  NANDN U15733 ( .A(n15351), .B(n19473), .Z(n15352) );
  AND U15734 ( .A(n15353), .B(n15352), .Z(n15495) );
  OR U15735 ( .A(n15354), .B(n16988), .Z(n15356) );
  XOR U15736 ( .A(a[116]), .B(n578), .Z(n15528) );
  NANDN U15737 ( .A(n15528), .B(n16990), .Z(n15355) );
  AND U15738 ( .A(n15356), .B(n15355), .Z(n15496) );
  XOR U15739 ( .A(n15497), .B(n15498), .Z(n15544) );
  XOR U15740 ( .A(n15543), .B(n15544), .Z(n15545) );
  XNOR U15741 ( .A(n15546), .B(n15545), .Z(n15591) );
  NANDN U15742 ( .A(n15358), .B(n15357), .Z(n15362) );
  NAND U15743 ( .A(n15360), .B(n15359), .Z(n15361) );
  NAND U15744 ( .A(n15362), .B(n15361), .Z(n15534) );
  NANDN U15745 ( .A(n15364), .B(n15363), .Z(n15368) );
  NAND U15746 ( .A(n15366), .B(n15365), .Z(n15367) );
  NAND U15747 ( .A(n15368), .B(n15367), .Z(n15532) );
  OR U15748 ( .A(n15370), .B(n15369), .Z(n15374) );
  NANDN U15749 ( .A(n15372), .B(n15371), .Z(n15373) );
  NAND U15750 ( .A(n15374), .B(n15373), .Z(n15531) );
  XNOR U15751 ( .A(n15534), .B(n15533), .Z(n15592) );
  XOR U15752 ( .A(n15591), .B(n15592), .Z(n15594) );
  NANDN U15753 ( .A(n15376), .B(n15375), .Z(n15380) );
  OR U15754 ( .A(n15378), .B(n15377), .Z(n15379) );
  NAND U15755 ( .A(n15380), .B(n15379), .Z(n15593) );
  XOR U15756 ( .A(n15594), .B(n15593), .Z(n15611) );
  OR U15757 ( .A(n15382), .B(n15381), .Z(n15386) );
  NAND U15758 ( .A(n15384), .B(n15383), .Z(n15385) );
  NAND U15759 ( .A(n15386), .B(n15385), .Z(n15610) );
  NANDN U15760 ( .A(n15388), .B(n15387), .Z(n15392) );
  NANDN U15761 ( .A(n15390), .B(n15389), .Z(n15391) );
  NAND U15762 ( .A(n15392), .B(n15391), .Z(n15599) );
  NANDN U15763 ( .A(n15394), .B(n15393), .Z(n15398) );
  OR U15764 ( .A(n15396), .B(n15395), .Z(n15397) );
  NAND U15765 ( .A(n15398), .B(n15397), .Z(n15598) );
  NANDN U15766 ( .A(n15400), .B(n15399), .Z(n15404) );
  NAND U15767 ( .A(n15402), .B(n15401), .Z(n15403) );
  NAND U15768 ( .A(n15404), .B(n15403), .Z(n15537) );
  NANDN U15769 ( .A(n15406), .B(n15405), .Z(n15410) );
  NAND U15770 ( .A(n15408), .B(n15407), .Z(n15409) );
  AND U15771 ( .A(n15410), .B(n15409), .Z(n15538) );
  XNOR U15772 ( .A(n15537), .B(n15538), .Z(n15539) );
  XOR U15773 ( .A(a[110]), .B(n579), .Z(n15561) );
  NANDN U15774 ( .A(n15561), .B(n17814), .Z(n15413) );
  NANDN U15775 ( .A(n15411), .B(n17815), .Z(n15412) );
  NAND U15776 ( .A(n15413), .B(n15412), .Z(n15503) );
  NAND U15777 ( .A(n15414), .B(n18513), .Z(n15416) );
  XNOR U15778 ( .A(b[15]), .B(a[104]), .Z(n15564) );
  OR U15779 ( .A(n15564), .B(n18512), .Z(n15415) );
  AND U15780 ( .A(n15416), .B(n15415), .Z(n15501) );
  NANDN U15781 ( .A(n15417), .B(n19013), .Z(n15419) );
  XNOR U15782 ( .A(b[21]), .B(a[98]), .Z(n15567) );
  NANDN U15783 ( .A(n15567), .B(n19015), .Z(n15418) );
  AND U15784 ( .A(n15419), .B(n15418), .Z(n15502) );
  XOR U15785 ( .A(n15503), .B(n15504), .Z(n15492) );
  XOR U15786 ( .A(b[11]), .B(n18198), .Z(n15570) );
  OR U15787 ( .A(n15570), .B(n18194), .Z(n15422) );
  NANDN U15788 ( .A(n15420), .B(n18104), .Z(n15421) );
  NAND U15789 ( .A(n15422), .B(n15421), .Z(n15490) );
  XOR U15790 ( .A(n580), .B(a[106]), .Z(n15573) );
  NANDN U15791 ( .A(n15573), .B(n18336), .Z(n15425) );
  NANDN U15792 ( .A(n15423), .B(n18337), .Z(n15424) );
  NAND U15793 ( .A(n15425), .B(n15424), .Z(n15489) );
  XOR U15794 ( .A(n15492), .B(n15491), .Z(n15486) );
  NANDN U15795 ( .A(n577), .B(a[118]), .Z(n15426) );
  XOR U15796 ( .A(n17151), .B(n15426), .Z(n15428) );
  IV U15797 ( .A(a[117]), .Z(n19136) );
  NANDN U15798 ( .A(n19136), .B(n577), .Z(n15427) );
  AND U15799 ( .A(n15428), .B(n15427), .Z(n15510) );
  ANDN U15800 ( .B(b[31]), .A(n15429), .Z(n15507) );
  NANDN U15801 ( .A(n15430), .B(n19406), .Z(n15432) );
  XNOR U15802 ( .A(n584), .B(a[90]), .Z(n15579) );
  NANDN U15803 ( .A(n576), .B(n15579), .Z(n15431) );
  NAND U15804 ( .A(n15432), .B(n15431), .Z(n15508) );
  XOR U15805 ( .A(n15507), .B(n15508), .Z(n15509) );
  XNOR U15806 ( .A(n15510), .B(n15509), .Z(n15483) );
  XOR U15807 ( .A(b[23]), .B(a[96]), .Z(n15582) );
  NANDN U15808 ( .A(n19127), .B(n15582), .Z(n15435) );
  NAND U15809 ( .A(n15433), .B(n19128), .Z(n15434) );
  NAND U15810 ( .A(n15435), .B(n15434), .Z(n15552) );
  NAND U15811 ( .A(n15436), .B(n17553), .Z(n15438) );
  XNOR U15812 ( .A(a[112]), .B(b[7]), .Z(n15585) );
  NANDN U15813 ( .A(n15585), .B(n17555), .Z(n15437) );
  NAND U15814 ( .A(n15438), .B(n15437), .Z(n15549) );
  XNOR U15815 ( .A(b[25]), .B(a[94]), .Z(n15588) );
  NANDN U15816 ( .A(n15588), .B(n19240), .Z(n15441) );
  NAND U15817 ( .A(n15439), .B(n19242), .Z(n15440) );
  AND U15818 ( .A(n15441), .B(n15440), .Z(n15550) );
  XNOR U15819 ( .A(n15549), .B(n15550), .Z(n15551) );
  XNOR U15820 ( .A(n15552), .B(n15551), .Z(n15484) );
  XOR U15821 ( .A(n15486), .B(n15485), .Z(n15540) );
  XNOR U15822 ( .A(n15539), .B(n15540), .Z(n15597) );
  XNOR U15823 ( .A(n15598), .B(n15597), .Z(n15600) );
  XNOR U15824 ( .A(n15599), .B(n15600), .Z(n15609) );
  XOR U15825 ( .A(n15610), .B(n15609), .Z(n15612) );
  NANDN U15826 ( .A(n15443), .B(n15442), .Z(n15447) );
  NANDN U15827 ( .A(n15445), .B(n15444), .Z(n15446) );
  NAND U15828 ( .A(n15447), .B(n15446), .Z(n15603) );
  NAND U15829 ( .A(n15449), .B(n15448), .Z(n15453) );
  NANDN U15830 ( .A(n15451), .B(n15450), .Z(n15452) );
  NAND U15831 ( .A(n15453), .B(n15452), .Z(n15604) );
  XNOR U15832 ( .A(n15603), .B(n15604), .Z(n15605) );
  XOR U15833 ( .A(n15606), .B(n15605), .Z(n15479) );
  NANDN U15834 ( .A(n15455), .B(n15454), .Z(n15459) );
  NAND U15835 ( .A(n15457), .B(n15456), .Z(n15458) );
  NAND U15836 ( .A(n15459), .B(n15458), .Z(n15477) );
  NANDN U15837 ( .A(n15461), .B(n15460), .Z(n15465) );
  OR U15838 ( .A(n15463), .B(n15462), .Z(n15464) );
  NAND U15839 ( .A(n15465), .B(n15464), .Z(n15478) );
  XNOR U15840 ( .A(n15477), .B(n15478), .Z(n15480) );
  XOR U15841 ( .A(n15479), .B(n15480), .Z(n15471) );
  XOR U15842 ( .A(n15472), .B(n15471), .Z(n15473) );
  XNOR U15843 ( .A(n15474), .B(n15473), .Z(n15615) );
  XNOR U15844 ( .A(n15615), .B(sreg[214]), .Z(n15617) );
  NAND U15845 ( .A(n15466), .B(sreg[213]), .Z(n15470) );
  OR U15846 ( .A(n15468), .B(n15467), .Z(n15469) );
  AND U15847 ( .A(n15470), .B(n15469), .Z(n15616) );
  XOR U15848 ( .A(n15617), .B(n15616), .Z(c[214]) );
  NAND U15849 ( .A(n15472), .B(n15471), .Z(n15476) );
  NAND U15850 ( .A(n15474), .B(n15473), .Z(n15475) );
  NAND U15851 ( .A(n15476), .B(n15475), .Z(n15623) );
  NANDN U15852 ( .A(n15478), .B(n15477), .Z(n15482) );
  NAND U15853 ( .A(n15480), .B(n15479), .Z(n15481) );
  NAND U15854 ( .A(n15482), .B(n15481), .Z(n15621) );
  OR U15855 ( .A(n15484), .B(n15483), .Z(n15488) );
  NANDN U15856 ( .A(n15486), .B(n15485), .Z(n15487) );
  NAND U15857 ( .A(n15488), .B(n15487), .Z(n15753) );
  OR U15858 ( .A(n15490), .B(n15489), .Z(n15494) );
  NAND U15859 ( .A(n15492), .B(n15491), .Z(n15493) );
  NAND U15860 ( .A(n15494), .B(n15493), .Z(n15692) );
  OR U15861 ( .A(n15496), .B(n15495), .Z(n15500) );
  NANDN U15862 ( .A(n15498), .B(n15497), .Z(n15499) );
  NAND U15863 ( .A(n15500), .B(n15499), .Z(n15691) );
  OR U15864 ( .A(n15502), .B(n15501), .Z(n15506) );
  NANDN U15865 ( .A(n15504), .B(n15503), .Z(n15505) );
  NAND U15866 ( .A(n15506), .B(n15505), .Z(n15690) );
  XOR U15867 ( .A(n15692), .B(n15693), .Z(n15751) );
  OR U15868 ( .A(n15508), .B(n15507), .Z(n15512) );
  NANDN U15869 ( .A(n15510), .B(n15509), .Z(n15511) );
  NAND U15870 ( .A(n15512), .B(n15511), .Z(n15704) );
  NANDN U15871 ( .A(n15513), .B(n18832), .Z(n15515) );
  XNOR U15872 ( .A(b[19]), .B(a[101]), .Z(n15648) );
  NANDN U15873 ( .A(n15648), .B(n18834), .Z(n15514) );
  NAND U15874 ( .A(n15515), .B(n15514), .Z(n15717) );
  XNOR U15875 ( .A(b[27]), .B(a[93]), .Z(n15651) );
  NANDN U15876 ( .A(n15651), .B(n19336), .Z(n15518) );
  NANDN U15877 ( .A(n15516), .B(n19337), .Z(n15517) );
  NAND U15878 ( .A(n15518), .B(n15517), .Z(n15714) );
  XNOR U15879 ( .A(a[115]), .B(b[5]), .Z(n15654) );
  NANDN U15880 ( .A(n15654), .B(n17310), .Z(n15521) );
  NANDN U15881 ( .A(n15519), .B(n17311), .Z(n15520) );
  AND U15882 ( .A(n15521), .B(n15520), .Z(n15715) );
  XNOR U15883 ( .A(n15714), .B(n15715), .Z(n15716) );
  XNOR U15884 ( .A(n15717), .B(n15716), .Z(n15703) );
  XOR U15885 ( .A(b[17]), .B(a[103]), .Z(n15657) );
  NAND U15886 ( .A(n15657), .B(n18673), .Z(n15524) );
  NANDN U15887 ( .A(n15522), .B(n18674), .Z(n15523) );
  NAND U15888 ( .A(n15524), .B(n15523), .Z(n15675) );
  XNOR U15889 ( .A(b[31]), .B(a[89]), .Z(n15660) );
  NANDN U15890 ( .A(n15660), .B(n19472), .Z(n15527) );
  NANDN U15891 ( .A(n15525), .B(n19473), .Z(n15526) );
  NAND U15892 ( .A(n15527), .B(n15526), .Z(n15672) );
  OR U15893 ( .A(n15528), .B(n16988), .Z(n15530) );
  XOR U15894 ( .A(a[117]), .B(n578), .Z(n15663) );
  NANDN U15895 ( .A(n15663), .B(n16990), .Z(n15529) );
  AND U15896 ( .A(n15530), .B(n15529), .Z(n15673) );
  XNOR U15897 ( .A(n15672), .B(n15673), .Z(n15674) );
  XOR U15898 ( .A(n15675), .B(n15674), .Z(n15702) );
  XOR U15899 ( .A(n15703), .B(n15702), .Z(n15705) );
  XOR U15900 ( .A(n15704), .B(n15705), .Z(n15750) );
  XOR U15901 ( .A(n15751), .B(n15750), .Z(n15752) );
  XNOR U15902 ( .A(n15753), .B(n15752), .Z(n15639) );
  OR U15903 ( .A(n15532), .B(n15531), .Z(n15536) );
  NAND U15904 ( .A(n15534), .B(n15533), .Z(n15535) );
  NAND U15905 ( .A(n15536), .B(n15535), .Z(n15637) );
  NANDN U15906 ( .A(n15538), .B(n15537), .Z(n15542) );
  NANDN U15907 ( .A(n15540), .B(n15539), .Z(n15541) );
  NAND U15908 ( .A(n15542), .B(n15541), .Z(n15758) );
  OR U15909 ( .A(n15544), .B(n15543), .Z(n15548) );
  NAND U15910 ( .A(n15546), .B(n15545), .Z(n15547) );
  NAND U15911 ( .A(n15548), .B(n15547), .Z(n15757) );
  NANDN U15912 ( .A(n15550), .B(n15549), .Z(n15554) );
  NAND U15913 ( .A(n15552), .B(n15551), .Z(n15553) );
  NAND U15914 ( .A(n15554), .B(n15553), .Z(n15696) );
  NANDN U15915 ( .A(n15556), .B(n15555), .Z(n15560) );
  NAND U15916 ( .A(n15558), .B(n15557), .Z(n15559) );
  AND U15917 ( .A(n15560), .B(n15559), .Z(n15697) );
  XNOR U15918 ( .A(n15696), .B(n15697), .Z(n15698) );
  XNOR U15919 ( .A(a[111]), .B(b[9]), .Z(n15720) );
  NANDN U15920 ( .A(n15720), .B(n17814), .Z(n15563) );
  NANDN U15921 ( .A(n15561), .B(n17815), .Z(n15562) );
  NAND U15922 ( .A(n15563), .B(n15562), .Z(n15680) );
  NANDN U15923 ( .A(n15564), .B(n18513), .Z(n15566) );
  XOR U15924 ( .A(b[15]), .B(a[105]), .Z(n15723) );
  NANDN U15925 ( .A(n18512), .B(n15723), .Z(n15565) );
  AND U15926 ( .A(n15566), .B(n15565), .Z(n15678) );
  NANDN U15927 ( .A(n15567), .B(n19013), .Z(n15569) );
  XNOR U15928 ( .A(b[21]), .B(a[99]), .Z(n15726) );
  NANDN U15929 ( .A(n15726), .B(n19015), .Z(n15568) );
  AND U15930 ( .A(n15569), .B(n15568), .Z(n15679) );
  XOR U15931 ( .A(n15680), .B(n15681), .Z(n15669) );
  XNOR U15932 ( .A(b[11]), .B(a[109]), .Z(n15729) );
  OR U15933 ( .A(n15729), .B(n18194), .Z(n15572) );
  NANDN U15934 ( .A(n15570), .B(n18104), .Z(n15571) );
  NAND U15935 ( .A(n15572), .B(n15571), .Z(n15667) );
  XOR U15936 ( .A(n580), .B(a[107]), .Z(n15732) );
  NANDN U15937 ( .A(n15732), .B(n18336), .Z(n15575) );
  NANDN U15938 ( .A(n15573), .B(n18337), .Z(n15574) );
  AND U15939 ( .A(n15575), .B(n15574), .Z(n15666) );
  XNOR U15940 ( .A(n15667), .B(n15666), .Z(n15668) );
  XOR U15941 ( .A(n15669), .B(n15668), .Z(n15686) );
  NANDN U15942 ( .A(n577), .B(a[119]), .Z(n15576) );
  XOR U15943 ( .A(n17151), .B(n15576), .Z(n15578) );
  IV U15944 ( .A(a[118]), .Z(n19077) );
  NANDN U15945 ( .A(n19077), .B(n577), .Z(n15577) );
  AND U15946 ( .A(n15578), .B(n15577), .Z(n15644) );
  NAND U15947 ( .A(n15579), .B(n19406), .Z(n15581) );
  XNOR U15948 ( .A(n584), .B(a[91]), .Z(n15738) );
  NANDN U15949 ( .A(n576), .B(n15738), .Z(n15580) );
  NAND U15950 ( .A(n15581), .B(n15580), .Z(n15642) );
  NANDN U15951 ( .A(n585), .B(a[87]), .Z(n15643) );
  XNOR U15952 ( .A(n15642), .B(n15643), .Z(n15645) );
  XOR U15953 ( .A(n15644), .B(n15645), .Z(n15684) );
  XNOR U15954 ( .A(b[23]), .B(a[97]), .Z(n15741) );
  OR U15955 ( .A(n15741), .B(n19127), .Z(n15584) );
  NAND U15956 ( .A(n15582), .B(n19128), .Z(n15583) );
  NAND U15957 ( .A(n15584), .B(n15583), .Z(n15711) );
  NANDN U15958 ( .A(n15585), .B(n17553), .Z(n15587) );
  XOR U15959 ( .A(a[113]), .B(b[7]), .Z(n15744) );
  NAND U15960 ( .A(n15744), .B(n17555), .Z(n15586) );
  NAND U15961 ( .A(n15587), .B(n15586), .Z(n15708) );
  XOR U15962 ( .A(b[25]), .B(a[95]), .Z(n15747) );
  NAND U15963 ( .A(n15747), .B(n19240), .Z(n15590) );
  NANDN U15964 ( .A(n15588), .B(n19242), .Z(n15589) );
  AND U15965 ( .A(n15590), .B(n15589), .Z(n15709) );
  XNOR U15966 ( .A(n15708), .B(n15709), .Z(n15710) );
  XNOR U15967 ( .A(n15711), .B(n15710), .Z(n15685) );
  XOR U15968 ( .A(n15684), .B(n15685), .Z(n15687) );
  XNOR U15969 ( .A(n15686), .B(n15687), .Z(n15699) );
  XNOR U15970 ( .A(n15698), .B(n15699), .Z(n15756) );
  XNOR U15971 ( .A(n15757), .B(n15756), .Z(n15759) );
  XNOR U15972 ( .A(n15758), .B(n15759), .Z(n15636) );
  XNOR U15973 ( .A(n15637), .B(n15636), .Z(n15638) );
  XOR U15974 ( .A(n15639), .B(n15638), .Z(n15633) );
  NANDN U15975 ( .A(n15592), .B(n15591), .Z(n15596) );
  OR U15976 ( .A(n15594), .B(n15593), .Z(n15595) );
  NAND U15977 ( .A(n15596), .B(n15595), .Z(n15630) );
  NAND U15978 ( .A(n15598), .B(n15597), .Z(n15602) );
  NANDN U15979 ( .A(n15600), .B(n15599), .Z(n15601) );
  NAND U15980 ( .A(n15602), .B(n15601), .Z(n15631) );
  XNOR U15981 ( .A(n15630), .B(n15631), .Z(n15632) );
  XNOR U15982 ( .A(n15633), .B(n15632), .Z(n15627) );
  NANDN U15983 ( .A(n15604), .B(n15603), .Z(n15608) );
  NAND U15984 ( .A(n15606), .B(n15605), .Z(n15607) );
  NAND U15985 ( .A(n15608), .B(n15607), .Z(n15624) );
  NANDN U15986 ( .A(n15610), .B(n15609), .Z(n15614) );
  OR U15987 ( .A(n15612), .B(n15611), .Z(n15613) );
  NAND U15988 ( .A(n15614), .B(n15613), .Z(n15625) );
  XNOR U15989 ( .A(n15624), .B(n15625), .Z(n15626) );
  XNOR U15990 ( .A(n15627), .B(n15626), .Z(n15620) );
  XOR U15991 ( .A(n15621), .B(n15620), .Z(n15622) );
  XNOR U15992 ( .A(n15623), .B(n15622), .Z(n15762) );
  XNOR U15993 ( .A(n15762), .B(sreg[215]), .Z(n15764) );
  NAND U15994 ( .A(n15615), .B(sreg[214]), .Z(n15619) );
  OR U15995 ( .A(n15617), .B(n15616), .Z(n15618) );
  AND U15996 ( .A(n15619), .B(n15618), .Z(n15763) );
  XOR U15997 ( .A(n15764), .B(n15763), .Z(c[215]) );
  NANDN U15998 ( .A(n15625), .B(n15624), .Z(n15629) );
  NANDN U15999 ( .A(n15627), .B(n15626), .Z(n15628) );
  NAND U16000 ( .A(n15629), .B(n15628), .Z(n15768) );
  NANDN U16001 ( .A(n15631), .B(n15630), .Z(n15635) );
  NAND U16002 ( .A(n15633), .B(n15632), .Z(n15634) );
  NAND U16003 ( .A(n15635), .B(n15634), .Z(n15773) );
  NANDN U16004 ( .A(n15637), .B(n15636), .Z(n15641) );
  NANDN U16005 ( .A(n15639), .B(n15638), .Z(n15640) );
  NAND U16006 ( .A(n15641), .B(n15640), .Z(n15774) );
  XNOR U16007 ( .A(n15773), .B(n15774), .Z(n15775) );
  NANDN U16008 ( .A(n15643), .B(n15642), .Z(n15647) );
  NAND U16009 ( .A(n15645), .B(n15644), .Z(n15646) );
  NAND U16010 ( .A(n15647), .B(n15646), .Z(n15854) );
  NANDN U16011 ( .A(n15648), .B(n18832), .Z(n15650) );
  XOR U16012 ( .A(b[19]), .B(n17208), .Z(n15797) );
  NANDN U16013 ( .A(n15797), .B(n18834), .Z(n15649) );
  NAND U16014 ( .A(n15650), .B(n15649), .Z(n15864) );
  XOR U16015 ( .A(b[27]), .B(n16590), .Z(n15800) );
  NANDN U16016 ( .A(n15800), .B(n19336), .Z(n15653) );
  NANDN U16017 ( .A(n15651), .B(n19337), .Z(n15652) );
  NAND U16018 ( .A(n15653), .B(n15652), .Z(n15861) );
  XNOR U16019 ( .A(a[116]), .B(b[5]), .Z(n15803) );
  NANDN U16020 ( .A(n15803), .B(n17310), .Z(n15656) );
  NANDN U16021 ( .A(n15654), .B(n17311), .Z(n15655) );
  AND U16022 ( .A(n15656), .B(n15655), .Z(n15862) );
  XNOR U16023 ( .A(n15861), .B(n15862), .Z(n15863) );
  XNOR U16024 ( .A(n15864), .B(n15863), .Z(n15852) );
  XNOR U16025 ( .A(b[17]), .B(a[104]), .Z(n15806) );
  NANDN U16026 ( .A(n15806), .B(n18673), .Z(n15659) );
  NAND U16027 ( .A(n15657), .B(n18674), .Z(n15658) );
  NAND U16028 ( .A(n15659), .B(n15658), .Z(n15824) );
  XNOR U16029 ( .A(b[31]), .B(a[90]), .Z(n15809) );
  NANDN U16030 ( .A(n15809), .B(n19472), .Z(n15662) );
  NANDN U16031 ( .A(n15660), .B(n19473), .Z(n15661) );
  NAND U16032 ( .A(n15662), .B(n15661), .Z(n15821) );
  OR U16033 ( .A(n15663), .B(n16988), .Z(n15665) );
  XOR U16034 ( .A(a[118]), .B(n578), .Z(n15812) );
  NANDN U16035 ( .A(n15812), .B(n16990), .Z(n15664) );
  AND U16036 ( .A(n15665), .B(n15664), .Z(n15822) );
  XNOR U16037 ( .A(n15821), .B(n15822), .Z(n15823) );
  XOR U16038 ( .A(n15824), .B(n15823), .Z(n15851) );
  XNOR U16039 ( .A(n15852), .B(n15851), .Z(n15853) );
  XNOR U16040 ( .A(n15854), .B(n15853), .Z(n15897) );
  NANDN U16041 ( .A(n15667), .B(n15666), .Z(n15671) );
  NAND U16042 ( .A(n15669), .B(n15668), .Z(n15670) );
  NAND U16043 ( .A(n15671), .B(n15670), .Z(n15842) );
  NANDN U16044 ( .A(n15673), .B(n15672), .Z(n15677) );
  NAND U16045 ( .A(n15675), .B(n15674), .Z(n15676) );
  NAND U16046 ( .A(n15677), .B(n15676), .Z(n15840) );
  OR U16047 ( .A(n15679), .B(n15678), .Z(n15683) );
  NANDN U16048 ( .A(n15681), .B(n15680), .Z(n15682) );
  NAND U16049 ( .A(n15683), .B(n15682), .Z(n15839) );
  XNOR U16050 ( .A(n15842), .B(n15841), .Z(n15898) );
  XOR U16051 ( .A(n15897), .B(n15898), .Z(n15900) );
  NANDN U16052 ( .A(n15685), .B(n15684), .Z(n15689) );
  OR U16053 ( .A(n15687), .B(n15686), .Z(n15688) );
  NAND U16054 ( .A(n15689), .B(n15688), .Z(n15899) );
  XOR U16055 ( .A(n15900), .B(n15899), .Z(n15787) );
  OR U16056 ( .A(n15691), .B(n15690), .Z(n15695) );
  NANDN U16057 ( .A(n15693), .B(n15692), .Z(n15694) );
  NAND U16058 ( .A(n15695), .B(n15694), .Z(n15786) );
  NANDN U16059 ( .A(n15697), .B(n15696), .Z(n15701) );
  NANDN U16060 ( .A(n15699), .B(n15698), .Z(n15700) );
  NAND U16061 ( .A(n15701), .B(n15700), .Z(n15905) );
  NANDN U16062 ( .A(n15703), .B(n15702), .Z(n15707) );
  OR U16063 ( .A(n15705), .B(n15704), .Z(n15706) );
  NAND U16064 ( .A(n15707), .B(n15706), .Z(n15904) );
  NANDN U16065 ( .A(n15709), .B(n15708), .Z(n15713) );
  NAND U16066 ( .A(n15711), .B(n15710), .Z(n15712) );
  NAND U16067 ( .A(n15713), .B(n15712), .Z(n15845) );
  NANDN U16068 ( .A(n15715), .B(n15714), .Z(n15719) );
  NAND U16069 ( .A(n15717), .B(n15716), .Z(n15718) );
  AND U16070 ( .A(n15719), .B(n15718), .Z(n15846) );
  XNOR U16071 ( .A(n15845), .B(n15846), .Z(n15847) );
  XOR U16072 ( .A(a[112]), .B(n579), .Z(n15867) );
  NANDN U16073 ( .A(n15867), .B(n17814), .Z(n15722) );
  NANDN U16074 ( .A(n15720), .B(n17815), .Z(n15721) );
  NAND U16075 ( .A(n15722), .B(n15721), .Z(n15829) );
  NAND U16076 ( .A(n15723), .B(n18513), .Z(n15725) );
  XNOR U16077 ( .A(b[15]), .B(a[106]), .Z(n15870) );
  OR U16078 ( .A(n15870), .B(n18512), .Z(n15724) );
  AND U16079 ( .A(n15725), .B(n15724), .Z(n15827) );
  NANDN U16080 ( .A(n15726), .B(n19013), .Z(n15728) );
  XOR U16081 ( .A(b[21]), .B(n17447), .Z(n15873) );
  NANDN U16082 ( .A(n15873), .B(n19015), .Z(n15727) );
  AND U16083 ( .A(n15728), .B(n15727), .Z(n15828) );
  XOR U16084 ( .A(n15829), .B(n15830), .Z(n15818) );
  XOR U16085 ( .A(n18415), .B(b[11]), .Z(n15876) );
  OR U16086 ( .A(n15876), .B(n18194), .Z(n15731) );
  NANDN U16087 ( .A(n15729), .B(n18104), .Z(n15730) );
  NAND U16088 ( .A(n15731), .B(n15730), .Z(n15816) );
  XOR U16089 ( .A(n580), .B(a[108]), .Z(n15879) );
  NANDN U16090 ( .A(n15879), .B(n18336), .Z(n15734) );
  NANDN U16091 ( .A(n15732), .B(n18337), .Z(n15733) );
  AND U16092 ( .A(n15734), .B(n15733), .Z(n15815) );
  XNOR U16093 ( .A(n15816), .B(n15815), .Z(n15817) );
  XOR U16094 ( .A(n15818), .B(n15817), .Z(n15835) );
  NANDN U16095 ( .A(n577), .B(a[120]), .Z(n15735) );
  XOR U16096 ( .A(n17151), .B(n15735), .Z(n15737) );
  IV U16097 ( .A(a[119]), .Z(n19239) );
  NANDN U16098 ( .A(n19239), .B(n577), .Z(n15736) );
  AND U16099 ( .A(n15737), .B(n15736), .Z(n15793) );
  NAND U16100 ( .A(n19406), .B(n15738), .Z(n15740) );
  XNOR U16101 ( .A(n584), .B(a[92]), .Z(n15885) );
  NANDN U16102 ( .A(n576), .B(n15885), .Z(n15739) );
  NAND U16103 ( .A(n15740), .B(n15739), .Z(n15791) );
  NANDN U16104 ( .A(n585), .B(a[88]), .Z(n15792) );
  XNOR U16105 ( .A(n15791), .B(n15792), .Z(n15794) );
  XOR U16106 ( .A(n15793), .B(n15794), .Z(n15833) );
  XOR U16107 ( .A(b[23]), .B(a[98]), .Z(n15888) );
  NANDN U16108 ( .A(n19127), .B(n15888), .Z(n15743) );
  NANDN U16109 ( .A(n15741), .B(n19128), .Z(n15742) );
  NAND U16110 ( .A(n15743), .B(n15742), .Z(n15858) );
  NAND U16111 ( .A(n15744), .B(n17553), .Z(n15746) );
  XNOR U16112 ( .A(a[114]), .B(b[7]), .Z(n15891) );
  NANDN U16113 ( .A(n15891), .B(n17555), .Z(n15745) );
  NAND U16114 ( .A(n15746), .B(n15745), .Z(n15855) );
  XOR U16115 ( .A(b[25]), .B(a[96]), .Z(n15894) );
  NAND U16116 ( .A(n15894), .B(n19240), .Z(n15749) );
  NAND U16117 ( .A(n15747), .B(n19242), .Z(n15748) );
  AND U16118 ( .A(n15749), .B(n15748), .Z(n15856) );
  XNOR U16119 ( .A(n15855), .B(n15856), .Z(n15857) );
  XNOR U16120 ( .A(n15858), .B(n15857), .Z(n15834) );
  XOR U16121 ( .A(n15833), .B(n15834), .Z(n15836) );
  XNOR U16122 ( .A(n15835), .B(n15836), .Z(n15848) );
  XNOR U16123 ( .A(n15847), .B(n15848), .Z(n15903) );
  XNOR U16124 ( .A(n15904), .B(n15903), .Z(n15906) );
  XNOR U16125 ( .A(n15905), .B(n15906), .Z(n15785) );
  XOR U16126 ( .A(n15786), .B(n15785), .Z(n15788) );
  NAND U16127 ( .A(n15751), .B(n15750), .Z(n15755) );
  NAND U16128 ( .A(n15753), .B(n15752), .Z(n15754) );
  NAND U16129 ( .A(n15755), .B(n15754), .Z(n15780) );
  NAND U16130 ( .A(n15757), .B(n15756), .Z(n15761) );
  NANDN U16131 ( .A(n15759), .B(n15758), .Z(n15760) );
  AND U16132 ( .A(n15761), .B(n15760), .Z(n15779) );
  XNOR U16133 ( .A(n15780), .B(n15779), .Z(n15781) );
  XOR U16134 ( .A(n15782), .B(n15781), .Z(n15776) );
  XOR U16135 ( .A(n15775), .B(n15776), .Z(n15767) );
  XOR U16136 ( .A(n15768), .B(n15767), .Z(n15769) );
  XNOR U16137 ( .A(n15770), .B(n15769), .Z(n15909) );
  XNOR U16138 ( .A(n15909), .B(sreg[216]), .Z(n15911) );
  NAND U16139 ( .A(n15762), .B(sreg[215]), .Z(n15766) );
  OR U16140 ( .A(n15764), .B(n15763), .Z(n15765) );
  AND U16141 ( .A(n15766), .B(n15765), .Z(n15910) );
  XOR U16142 ( .A(n15911), .B(n15910), .Z(c[216]) );
  NAND U16143 ( .A(n15768), .B(n15767), .Z(n15772) );
  NAND U16144 ( .A(n15770), .B(n15769), .Z(n15771) );
  NAND U16145 ( .A(n15772), .B(n15771), .Z(n15917) );
  NANDN U16146 ( .A(n15774), .B(n15773), .Z(n15778) );
  NAND U16147 ( .A(n15776), .B(n15775), .Z(n15777) );
  NAND U16148 ( .A(n15778), .B(n15777), .Z(n15915) );
  NANDN U16149 ( .A(n15780), .B(n15779), .Z(n15784) );
  NAND U16150 ( .A(n15782), .B(n15781), .Z(n15783) );
  NAND U16151 ( .A(n15784), .B(n15783), .Z(n15920) );
  NANDN U16152 ( .A(n15786), .B(n15785), .Z(n15790) );
  OR U16153 ( .A(n15788), .B(n15787), .Z(n15789) );
  NAND U16154 ( .A(n15790), .B(n15789), .Z(n15921) );
  XNOR U16155 ( .A(n15920), .B(n15921), .Z(n15922) );
  NANDN U16156 ( .A(n15792), .B(n15791), .Z(n15796) );
  NAND U16157 ( .A(n15794), .B(n15793), .Z(n15795) );
  NAND U16158 ( .A(n15796), .B(n15795), .Z(n16001) );
  NANDN U16159 ( .A(n15797), .B(n18832), .Z(n15799) );
  XNOR U16160 ( .A(b[19]), .B(a[103]), .Z(n15968) );
  NANDN U16161 ( .A(n15968), .B(n18834), .Z(n15798) );
  NAND U16162 ( .A(n15799), .B(n15798), .Z(n16013) );
  XNOR U16163 ( .A(b[27]), .B(a[95]), .Z(n15971) );
  NANDN U16164 ( .A(n15971), .B(n19336), .Z(n15802) );
  NANDN U16165 ( .A(n15800), .B(n19337), .Z(n15801) );
  NAND U16166 ( .A(n15802), .B(n15801), .Z(n16010) );
  XNOR U16167 ( .A(a[117]), .B(b[5]), .Z(n15974) );
  NANDN U16168 ( .A(n15974), .B(n17310), .Z(n15805) );
  NANDN U16169 ( .A(n15803), .B(n17311), .Z(n15804) );
  AND U16170 ( .A(n15805), .B(n15804), .Z(n16011) );
  XNOR U16171 ( .A(n16010), .B(n16011), .Z(n16012) );
  XNOR U16172 ( .A(n16013), .B(n16012), .Z(n15998) );
  XOR U16173 ( .A(b[17]), .B(a[105]), .Z(n15977) );
  NAND U16174 ( .A(n15977), .B(n18673), .Z(n15808) );
  NANDN U16175 ( .A(n15806), .B(n18674), .Z(n15807) );
  NAND U16176 ( .A(n15808), .B(n15807), .Z(n15952) );
  XNOR U16177 ( .A(b[31]), .B(a[91]), .Z(n15980) );
  NANDN U16178 ( .A(n15980), .B(n19472), .Z(n15811) );
  NANDN U16179 ( .A(n15809), .B(n19473), .Z(n15810) );
  AND U16180 ( .A(n15811), .B(n15810), .Z(n15950) );
  OR U16181 ( .A(n15812), .B(n16988), .Z(n15814) );
  XOR U16182 ( .A(a[119]), .B(n578), .Z(n15983) );
  NANDN U16183 ( .A(n15983), .B(n16990), .Z(n15813) );
  AND U16184 ( .A(n15814), .B(n15813), .Z(n15951) );
  XOR U16185 ( .A(n15952), .B(n15953), .Z(n15999) );
  XOR U16186 ( .A(n15998), .B(n15999), .Z(n16000) );
  XNOR U16187 ( .A(n16001), .B(n16000), .Z(n16046) );
  NANDN U16188 ( .A(n15816), .B(n15815), .Z(n15820) );
  NAND U16189 ( .A(n15818), .B(n15817), .Z(n15819) );
  NAND U16190 ( .A(n15820), .B(n15819), .Z(n15989) );
  NANDN U16191 ( .A(n15822), .B(n15821), .Z(n15826) );
  NAND U16192 ( .A(n15824), .B(n15823), .Z(n15825) );
  NAND U16193 ( .A(n15826), .B(n15825), .Z(n15987) );
  OR U16194 ( .A(n15828), .B(n15827), .Z(n15832) );
  NANDN U16195 ( .A(n15830), .B(n15829), .Z(n15831) );
  NAND U16196 ( .A(n15832), .B(n15831), .Z(n15986) );
  XNOR U16197 ( .A(n15989), .B(n15988), .Z(n16047) );
  XOR U16198 ( .A(n16046), .B(n16047), .Z(n16049) );
  NANDN U16199 ( .A(n15834), .B(n15833), .Z(n15838) );
  OR U16200 ( .A(n15836), .B(n15835), .Z(n15837) );
  NAND U16201 ( .A(n15838), .B(n15837), .Z(n16048) );
  XOR U16202 ( .A(n16049), .B(n16048), .Z(n15934) );
  OR U16203 ( .A(n15840), .B(n15839), .Z(n15844) );
  NAND U16204 ( .A(n15842), .B(n15841), .Z(n15843) );
  NAND U16205 ( .A(n15844), .B(n15843), .Z(n15933) );
  NANDN U16206 ( .A(n15846), .B(n15845), .Z(n15850) );
  NANDN U16207 ( .A(n15848), .B(n15847), .Z(n15849) );
  NAND U16208 ( .A(n15850), .B(n15849), .Z(n16054) );
  NANDN U16209 ( .A(n15856), .B(n15855), .Z(n15860) );
  NAND U16210 ( .A(n15858), .B(n15857), .Z(n15859) );
  NAND U16211 ( .A(n15860), .B(n15859), .Z(n15992) );
  NANDN U16212 ( .A(n15862), .B(n15861), .Z(n15866) );
  NAND U16213 ( .A(n15864), .B(n15863), .Z(n15865) );
  AND U16214 ( .A(n15866), .B(n15865), .Z(n15993) );
  XNOR U16215 ( .A(n15992), .B(n15993), .Z(n15994) );
  XNOR U16216 ( .A(a[113]), .B(b[9]), .Z(n16016) );
  NANDN U16217 ( .A(n16016), .B(n17814), .Z(n15869) );
  NANDN U16218 ( .A(n15867), .B(n17815), .Z(n15868) );
  NAND U16219 ( .A(n15869), .B(n15868), .Z(n15958) );
  NANDN U16220 ( .A(n15870), .B(n18513), .Z(n15872) );
  XOR U16221 ( .A(b[15]), .B(a[107]), .Z(n16019) );
  NANDN U16222 ( .A(n18512), .B(n16019), .Z(n15871) );
  AND U16223 ( .A(n15872), .B(n15871), .Z(n15956) );
  NANDN U16224 ( .A(n15873), .B(n19013), .Z(n15875) );
  XNOR U16225 ( .A(b[21]), .B(a[101]), .Z(n16022) );
  NANDN U16226 ( .A(n16022), .B(n19015), .Z(n15874) );
  AND U16227 ( .A(n15875), .B(n15874), .Z(n15957) );
  XOR U16228 ( .A(n15958), .B(n15959), .Z(n15947) );
  XNOR U16229 ( .A(a[111]), .B(b[11]), .Z(n16025) );
  OR U16230 ( .A(n16025), .B(n18194), .Z(n15878) );
  NANDN U16231 ( .A(n15876), .B(n18104), .Z(n15877) );
  NAND U16232 ( .A(n15878), .B(n15877), .Z(n15945) );
  XOR U16233 ( .A(n580), .B(a[109]), .Z(n16028) );
  NANDN U16234 ( .A(n16028), .B(n18336), .Z(n15881) );
  NANDN U16235 ( .A(n15879), .B(n18337), .Z(n15880) );
  NAND U16236 ( .A(n15881), .B(n15880), .Z(n15944) );
  XOR U16237 ( .A(n15947), .B(n15946), .Z(n15941) );
  NANDN U16238 ( .A(n577), .B(a[121]), .Z(n15882) );
  XOR U16239 ( .A(n17151), .B(n15882), .Z(n15884) );
  IV U16240 ( .A(a[120]), .Z(n19188) );
  NANDN U16241 ( .A(n19188), .B(n577), .Z(n15883) );
  AND U16242 ( .A(n15884), .B(n15883), .Z(n15964) );
  NAND U16243 ( .A(n19406), .B(n15885), .Z(n15887) );
  XNOR U16244 ( .A(n584), .B(a[93]), .Z(n16034) );
  NANDN U16245 ( .A(n576), .B(n16034), .Z(n15886) );
  NAND U16246 ( .A(n15887), .B(n15886), .Z(n15962) );
  NANDN U16247 ( .A(n585), .B(a[89]), .Z(n15963) );
  XNOR U16248 ( .A(n15962), .B(n15963), .Z(n15965) );
  XNOR U16249 ( .A(n15964), .B(n15965), .Z(n15939) );
  XOR U16250 ( .A(b[23]), .B(a[99]), .Z(n16037) );
  NANDN U16251 ( .A(n19127), .B(n16037), .Z(n15890) );
  NAND U16252 ( .A(n15888), .B(n19128), .Z(n15889) );
  NAND U16253 ( .A(n15890), .B(n15889), .Z(n16007) );
  NANDN U16254 ( .A(n15891), .B(n17553), .Z(n15893) );
  XNOR U16255 ( .A(a[115]), .B(b[7]), .Z(n16040) );
  NANDN U16256 ( .A(n16040), .B(n17555), .Z(n15892) );
  NAND U16257 ( .A(n15893), .B(n15892), .Z(n16004) );
  XNOR U16258 ( .A(b[25]), .B(a[97]), .Z(n16043) );
  NANDN U16259 ( .A(n16043), .B(n19240), .Z(n15896) );
  NAND U16260 ( .A(n15894), .B(n19242), .Z(n15895) );
  AND U16261 ( .A(n15896), .B(n15895), .Z(n16005) );
  XNOR U16262 ( .A(n16004), .B(n16005), .Z(n16006) );
  XOR U16263 ( .A(n16007), .B(n16006), .Z(n15938) );
  XOR U16264 ( .A(n15941), .B(n15940), .Z(n15995) );
  XNOR U16265 ( .A(n15994), .B(n15995), .Z(n16052) );
  XNOR U16266 ( .A(n16053), .B(n16052), .Z(n16055) );
  XNOR U16267 ( .A(n16054), .B(n16055), .Z(n15932) );
  XOR U16268 ( .A(n15933), .B(n15932), .Z(n15935) );
  NANDN U16269 ( .A(n15898), .B(n15897), .Z(n15902) );
  OR U16270 ( .A(n15900), .B(n15899), .Z(n15901) );
  NAND U16271 ( .A(n15902), .B(n15901), .Z(n15926) );
  NAND U16272 ( .A(n15904), .B(n15903), .Z(n15908) );
  NANDN U16273 ( .A(n15906), .B(n15905), .Z(n15907) );
  NAND U16274 ( .A(n15908), .B(n15907), .Z(n15927) );
  XNOR U16275 ( .A(n15926), .B(n15927), .Z(n15928) );
  XOR U16276 ( .A(n15929), .B(n15928), .Z(n15923) );
  XOR U16277 ( .A(n15922), .B(n15923), .Z(n15914) );
  XOR U16278 ( .A(n15915), .B(n15914), .Z(n15916) );
  XNOR U16279 ( .A(n15917), .B(n15916), .Z(n16058) );
  XNOR U16280 ( .A(n16058), .B(sreg[217]), .Z(n16060) );
  NAND U16281 ( .A(n15909), .B(sreg[216]), .Z(n15913) );
  OR U16282 ( .A(n15911), .B(n15910), .Z(n15912) );
  AND U16283 ( .A(n15913), .B(n15912), .Z(n16059) );
  XOR U16284 ( .A(n16060), .B(n16059), .Z(c[217]) );
  NAND U16285 ( .A(n15915), .B(n15914), .Z(n15919) );
  NAND U16286 ( .A(n15917), .B(n15916), .Z(n15918) );
  NAND U16287 ( .A(n15919), .B(n15918), .Z(n16066) );
  NANDN U16288 ( .A(n15921), .B(n15920), .Z(n15925) );
  NAND U16289 ( .A(n15923), .B(n15922), .Z(n15924) );
  NAND U16290 ( .A(n15925), .B(n15924), .Z(n16064) );
  NANDN U16291 ( .A(n15927), .B(n15926), .Z(n15931) );
  NAND U16292 ( .A(n15929), .B(n15928), .Z(n15930) );
  NAND U16293 ( .A(n15931), .B(n15930), .Z(n16069) );
  NANDN U16294 ( .A(n15933), .B(n15932), .Z(n15937) );
  OR U16295 ( .A(n15935), .B(n15934), .Z(n15936) );
  NAND U16296 ( .A(n15937), .B(n15936), .Z(n16070) );
  XNOR U16297 ( .A(n16069), .B(n16070), .Z(n16071) );
  NANDN U16298 ( .A(n15939), .B(n15938), .Z(n15943) );
  NANDN U16299 ( .A(n15941), .B(n15940), .Z(n15942) );
  NAND U16300 ( .A(n15943), .B(n15942), .Z(n16186) );
  OR U16301 ( .A(n15945), .B(n15944), .Z(n15949) );
  NAND U16302 ( .A(n15947), .B(n15946), .Z(n15948) );
  NAND U16303 ( .A(n15949), .B(n15948), .Z(n16125) );
  OR U16304 ( .A(n15951), .B(n15950), .Z(n15955) );
  NANDN U16305 ( .A(n15953), .B(n15952), .Z(n15954) );
  NAND U16306 ( .A(n15955), .B(n15954), .Z(n16124) );
  OR U16307 ( .A(n15957), .B(n15956), .Z(n15961) );
  NANDN U16308 ( .A(n15959), .B(n15958), .Z(n15960) );
  NAND U16309 ( .A(n15961), .B(n15960), .Z(n16123) );
  XOR U16310 ( .A(n16125), .B(n16126), .Z(n16183) );
  NANDN U16311 ( .A(n15963), .B(n15962), .Z(n15967) );
  NAND U16312 ( .A(n15965), .B(n15964), .Z(n15966) );
  NAND U16313 ( .A(n15967), .B(n15966), .Z(n16138) );
  NANDN U16314 ( .A(n15968), .B(n18832), .Z(n15970) );
  XOR U16315 ( .A(b[19]), .B(n17716), .Z(n16081) );
  NANDN U16316 ( .A(n16081), .B(n18834), .Z(n15969) );
  NAND U16317 ( .A(n15970), .B(n15969), .Z(n16150) );
  XNOR U16318 ( .A(b[27]), .B(a[96]), .Z(n16084) );
  NANDN U16319 ( .A(n16084), .B(n19336), .Z(n15973) );
  NANDN U16320 ( .A(n15971), .B(n19337), .Z(n15972) );
  NAND U16321 ( .A(n15973), .B(n15972), .Z(n16147) );
  XNOR U16322 ( .A(a[118]), .B(b[5]), .Z(n16087) );
  NANDN U16323 ( .A(n16087), .B(n17310), .Z(n15976) );
  NANDN U16324 ( .A(n15974), .B(n17311), .Z(n15975) );
  AND U16325 ( .A(n15976), .B(n15975), .Z(n16148) );
  XNOR U16326 ( .A(n16147), .B(n16148), .Z(n16149) );
  XNOR U16327 ( .A(n16150), .B(n16149), .Z(n16136) );
  XNOR U16328 ( .A(b[17]), .B(a[106]), .Z(n16090) );
  NANDN U16329 ( .A(n16090), .B(n18673), .Z(n15979) );
  NAND U16330 ( .A(n15977), .B(n18674), .Z(n15978) );
  NAND U16331 ( .A(n15979), .B(n15978), .Z(n16108) );
  XNOR U16332 ( .A(b[31]), .B(a[92]), .Z(n16093) );
  NANDN U16333 ( .A(n16093), .B(n19472), .Z(n15982) );
  NANDN U16334 ( .A(n15980), .B(n19473), .Z(n15981) );
  NAND U16335 ( .A(n15982), .B(n15981), .Z(n16105) );
  OR U16336 ( .A(n15983), .B(n16988), .Z(n15985) );
  XOR U16337 ( .A(a[120]), .B(n578), .Z(n16096) );
  NANDN U16338 ( .A(n16096), .B(n16990), .Z(n15984) );
  AND U16339 ( .A(n15985), .B(n15984), .Z(n16106) );
  XNOR U16340 ( .A(n16105), .B(n16106), .Z(n16107) );
  XOR U16341 ( .A(n16108), .B(n16107), .Z(n16135) );
  XNOR U16342 ( .A(n16136), .B(n16135), .Z(n16137) );
  XNOR U16343 ( .A(n16138), .B(n16137), .Z(n16184) );
  XNOR U16344 ( .A(n16183), .B(n16184), .Z(n16185) );
  XNOR U16345 ( .A(n16186), .B(n16185), .Z(n16204) );
  OR U16346 ( .A(n15987), .B(n15986), .Z(n15991) );
  NAND U16347 ( .A(n15989), .B(n15988), .Z(n15990) );
  NAND U16348 ( .A(n15991), .B(n15990), .Z(n16202) );
  NANDN U16349 ( .A(n15993), .B(n15992), .Z(n15997) );
  NANDN U16350 ( .A(n15995), .B(n15994), .Z(n15996) );
  NAND U16351 ( .A(n15997), .B(n15996), .Z(n16191) );
  OR U16352 ( .A(n15999), .B(n15998), .Z(n16003) );
  NAND U16353 ( .A(n16001), .B(n16000), .Z(n16002) );
  NAND U16354 ( .A(n16003), .B(n16002), .Z(n16190) );
  NANDN U16355 ( .A(n16005), .B(n16004), .Z(n16009) );
  NAND U16356 ( .A(n16007), .B(n16006), .Z(n16008) );
  NAND U16357 ( .A(n16009), .B(n16008), .Z(n16129) );
  NANDN U16358 ( .A(n16011), .B(n16010), .Z(n16015) );
  NAND U16359 ( .A(n16013), .B(n16012), .Z(n16014) );
  AND U16360 ( .A(n16015), .B(n16014), .Z(n16130) );
  XNOR U16361 ( .A(n16129), .B(n16130), .Z(n16131) );
  XOR U16362 ( .A(n18751), .B(n579), .Z(n16153) );
  NAND U16363 ( .A(n17814), .B(n16153), .Z(n16018) );
  NANDN U16364 ( .A(n16016), .B(n17815), .Z(n16017) );
  NAND U16365 ( .A(n16018), .B(n16017), .Z(n16113) );
  NAND U16366 ( .A(n16019), .B(n18513), .Z(n16021) );
  XNOR U16367 ( .A(b[15]), .B(a[108]), .Z(n16156) );
  OR U16368 ( .A(n16156), .B(n18512), .Z(n16020) );
  AND U16369 ( .A(n16021), .B(n16020), .Z(n16111) );
  NANDN U16370 ( .A(n16022), .B(n19013), .Z(n16024) );
  XOR U16371 ( .A(n582), .B(n17208), .Z(n16159) );
  NAND U16372 ( .A(n16159), .B(n19015), .Z(n16023) );
  AND U16373 ( .A(n16024), .B(n16023), .Z(n16112) );
  XOR U16374 ( .A(n16113), .B(n16114), .Z(n16102) );
  XOR U16375 ( .A(n18582), .B(b[11]), .Z(n16162) );
  OR U16376 ( .A(n16162), .B(n18194), .Z(n16027) );
  NANDN U16377 ( .A(n16025), .B(n18104), .Z(n16026) );
  NAND U16378 ( .A(n16027), .B(n16026), .Z(n16100) );
  XOR U16379 ( .A(n580), .B(a[110]), .Z(n16165) );
  NANDN U16380 ( .A(n16165), .B(n18336), .Z(n16030) );
  NANDN U16381 ( .A(n16028), .B(n18337), .Z(n16029) );
  AND U16382 ( .A(n16030), .B(n16029), .Z(n16099) );
  XNOR U16383 ( .A(n16100), .B(n16099), .Z(n16101) );
  XOR U16384 ( .A(n16102), .B(n16101), .Z(n16119) );
  NANDN U16385 ( .A(n577), .B(a[122]), .Z(n16031) );
  XOR U16386 ( .A(n17151), .B(n16031), .Z(n16033) );
  IV U16387 ( .A(a[121]), .Z(n19347) );
  NANDN U16388 ( .A(n19347), .B(n577), .Z(n16032) );
  AND U16389 ( .A(n16033), .B(n16032), .Z(n16077) );
  NAND U16390 ( .A(n19406), .B(n16034), .Z(n16036) );
  XOR U16391 ( .A(n584), .B(n16590), .Z(n16168) );
  NANDN U16392 ( .A(n576), .B(n16168), .Z(n16035) );
  NAND U16393 ( .A(n16036), .B(n16035), .Z(n16075) );
  NANDN U16394 ( .A(n585), .B(a[90]), .Z(n16076) );
  XNOR U16395 ( .A(n16075), .B(n16076), .Z(n16078) );
  XOR U16396 ( .A(n16077), .B(n16078), .Z(n16117) );
  XNOR U16397 ( .A(b[23]), .B(a[100]), .Z(n16174) );
  OR U16398 ( .A(n16174), .B(n19127), .Z(n16039) );
  NAND U16399 ( .A(n16037), .B(n19128), .Z(n16038) );
  NAND U16400 ( .A(n16039), .B(n16038), .Z(n16144) );
  NANDN U16401 ( .A(n16040), .B(n17553), .Z(n16042) );
  XNOR U16402 ( .A(a[116]), .B(b[7]), .Z(n16177) );
  NANDN U16403 ( .A(n16177), .B(n17555), .Z(n16041) );
  NAND U16404 ( .A(n16042), .B(n16041), .Z(n16141) );
  XOR U16405 ( .A(b[25]), .B(a[98]), .Z(n16180) );
  NAND U16406 ( .A(n16180), .B(n19240), .Z(n16045) );
  NANDN U16407 ( .A(n16043), .B(n19242), .Z(n16044) );
  AND U16408 ( .A(n16045), .B(n16044), .Z(n16142) );
  XNOR U16409 ( .A(n16141), .B(n16142), .Z(n16143) );
  XNOR U16410 ( .A(n16144), .B(n16143), .Z(n16118) );
  XOR U16411 ( .A(n16117), .B(n16118), .Z(n16120) );
  XNOR U16412 ( .A(n16119), .B(n16120), .Z(n16132) );
  XNOR U16413 ( .A(n16131), .B(n16132), .Z(n16189) );
  XNOR U16414 ( .A(n16190), .B(n16189), .Z(n16192) );
  XNOR U16415 ( .A(n16191), .B(n16192), .Z(n16201) );
  XNOR U16416 ( .A(n16202), .B(n16201), .Z(n16203) );
  XOR U16417 ( .A(n16204), .B(n16203), .Z(n16198) );
  NANDN U16418 ( .A(n16047), .B(n16046), .Z(n16051) );
  OR U16419 ( .A(n16049), .B(n16048), .Z(n16050) );
  NAND U16420 ( .A(n16051), .B(n16050), .Z(n16195) );
  NAND U16421 ( .A(n16053), .B(n16052), .Z(n16057) );
  NANDN U16422 ( .A(n16055), .B(n16054), .Z(n16056) );
  NAND U16423 ( .A(n16057), .B(n16056), .Z(n16196) );
  XNOR U16424 ( .A(n16195), .B(n16196), .Z(n16197) );
  XOR U16425 ( .A(n16198), .B(n16197), .Z(n16072) );
  XOR U16426 ( .A(n16071), .B(n16072), .Z(n16063) );
  XOR U16427 ( .A(n16064), .B(n16063), .Z(n16065) );
  XNOR U16428 ( .A(n16066), .B(n16065), .Z(n16207) );
  XNOR U16429 ( .A(n16207), .B(sreg[218]), .Z(n16209) );
  NAND U16430 ( .A(n16058), .B(sreg[217]), .Z(n16062) );
  OR U16431 ( .A(n16060), .B(n16059), .Z(n16061) );
  AND U16432 ( .A(n16062), .B(n16061), .Z(n16208) );
  XOR U16433 ( .A(n16209), .B(n16208), .Z(c[218]) );
  NAND U16434 ( .A(n16064), .B(n16063), .Z(n16068) );
  NAND U16435 ( .A(n16066), .B(n16065), .Z(n16067) );
  NAND U16436 ( .A(n16068), .B(n16067), .Z(n16215) );
  NANDN U16437 ( .A(n16070), .B(n16069), .Z(n16074) );
  NAND U16438 ( .A(n16072), .B(n16071), .Z(n16073) );
  NAND U16439 ( .A(n16074), .B(n16073), .Z(n16213) );
  NANDN U16440 ( .A(n16076), .B(n16075), .Z(n16080) );
  NAND U16441 ( .A(n16078), .B(n16077), .Z(n16079) );
  NAND U16442 ( .A(n16080), .B(n16079), .Z(n16297) );
  NANDN U16443 ( .A(n16081), .B(n18832), .Z(n16083) );
  XNOR U16444 ( .A(n581), .B(a[105]), .Z(n16242) );
  NAND U16445 ( .A(n16242), .B(n18834), .Z(n16082) );
  NAND U16446 ( .A(n16083), .B(n16082), .Z(n16337) );
  XOR U16447 ( .A(n583), .B(n17038), .Z(n16248) );
  NAND U16448 ( .A(n19336), .B(n16248), .Z(n16086) );
  NANDN U16449 ( .A(n16084), .B(n19337), .Z(n16085) );
  NAND U16450 ( .A(n16086), .B(n16085), .Z(n16334) );
  XNOR U16451 ( .A(n19239), .B(b[5]), .Z(n16245) );
  NAND U16452 ( .A(n16245), .B(n17310), .Z(n16089) );
  NANDN U16453 ( .A(n16087), .B(n17311), .Z(n16088) );
  AND U16454 ( .A(n16089), .B(n16088), .Z(n16335) );
  XNOR U16455 ( .A(n16334), .B(n16335), .Z(n16336) );
  XNOR U16456 ( .A(n16337), .B(n16336), .Z(n16295) );
  XOR U16457 ( .A(b[17]), .B(a[107]), .Z(n16251) );
  NAND U16458 ( .A(n16251), .B(n18673), .Z(n16092) );
  NANDN U16459 ( .A(n16090), .B(n18674), .Z(n16091) );
  NAND U16460 ( .A(n16092), .B(n16091), .Z(n16269) );
  XNOR U16461 ( .A(b[31]), .B(a[93]), .Z(n16254) );
  NANDN U16462 ( .A(n16254), .B(n19472), .Z(n16095) );
  NANDN U16463 ( .A(n16093), .B(n19473), .Z(n16094) );
  NAND U16464 ( .A(n16095), .B(n16094), .Z(n16266) );
  OR U16465 ( .A(n16096), .B(n16988), .Z(n16098) );
  XOR U16466 ( .A(a[121]), .B(n578), .Z(n16257) );
  NANDN U16467 ( .A(n16257), .B(n16990), .Z(n16097) );
  AND U16468 ( .A(n16098), .B(n16097), .Z(n16267) );
  XNOR U16469 ( .A(n16266), .B(n16267), .Z(n16268) );
  XOR U16470 ( .A(n16269), .B(n16268), .Z(n16294) );
  XNOR U16471 ( .A(n16295), .B(n16294), .Z(n16296) );
  XNOR U16472 ( .A(n16297), .B(n16296), .Z(n16340) );
  NANDN U16473 ( .A(n16100), .B(n16099), .Z(n16104) );
  NAND U16474 ( .A(n16102), .B(n16101), .Z(n16103) );
  NAND U16475 ( .A(n16104), .B(n16103), .Z(n16285) );
  NANDN U16476 ( .A(n16106), .B(n16105), .Z(n16110) );
  NAND U16477 ( .A(n16108), .B(n16107), .Z(n16109) );
  NAND U16478 ( .A(n16110), .B(n16109), .Z(n16283) );
  OR U16479 ( .A(n16112), .B(n16111), .Z(n16116) );
  NANDN U16480 ( .A(n16114), .B(n16113), .Z(n16115) );
  NAND U16481 ( .A(n16116), .B(n16115), .Z(n16282) );
  XNOR U16482 ( .A(n16285), .B(n16284), .Z(n16341) );
  XOR U16483 ( .A(n16340), .B(n16341), .Z(n16343) );
  NANDN U16484 ( .A(n16118), .B(n16117), .Z(n16122) );
  OR U16485 ( .A(n16120), .B(n16119), .Z(n16121) );
  NAND U16486 ( .A(n16122), .B(n16121), .Z(n16342) );
  XOR U16487 ( .A(n16343), .B(n16342), .Z(n16232) );
  OR U16488 ( .A(n16124), .B(n16123), .Z(n16128) );
  NANDN U16489 ( .A(n16126), .B(n16125), .Z(n16127) );
  NAND U16490 ( .A(n16128), .B(n16127), .Z(n16231) );
  NANDN U16491 ( .A(n16130), .B(n16129), .Z(n16134) );
  NANDN U16492 ( .A(n16132), .B(n16131), .Z(n16133) );
  NAND U16493 ( .A(n16134), .B(n16133), .Z(n16348) );
  NANDN U16494 ( .A(n16136), .B(n16135), .Z(n16140) );
  NAND U16495 ( .A(n16138), .B(n16137), .Z(n16139) );
  NAND U16496 ( .A(n16140), .B(n16139), .Z(n16347) );
  NANDN U16497 ( .A(n16142), .B(n16141), .Z(n16146) );
  NAND U16498 ( .A(n16144), .B(n16143), .Z(n16145) );
  NAND U16499 ( .A(n16146), .B(n16145), .Z(n16288) );
  NANDN U16500 ( .A(n16148), .B(n16147), .Z(n16152) );
  NAND U16501 ( .A(n16150), .B(n16149), .Z(n16151) );
  AND U16502 ( .A(n16152), .B(n16151), .Z(n16289) );
  XNOR U16503 ( .A(n16288), .B(n16289), .Z(n16290) );
  XOR U16504 ( .A(a[115]), .B(n579), .Z(n16298) );
  NANDN U16505 ( .A(n16298), .B(n17814), .Z(n16155) );
  NAND U16506 ( .A(n17815), .B(n16153), .Z(n16154) );
  NAND U16507 ( .A(n16155), .B(n16154), .Z(n16274) );
  XNOR U16508 ( .A(b[15]), .B(a[109]), .Z(n16301) );
  OR U16509 ( .A(n16301), .B(n18512), .Z(n16158) );
  NANDN U16510 ( .A(n16156), .B(n18513), .Z(n16157) );
  NAND U16511 ( .A(n16158), .B(n16157), .Z(n16272) );
  XNOR U16512 ( .A(b[21]), .B(a[103]), .Z(n16304) );
  NANDN U16513 ( .A(n16304), .B(n19015), .Z(n16161) );
  NAND U16514 ( .A(n19013), .B(n16159), .Z(n16160) );
  NAND U16515 ( .A(n16161), .B(n16160), .Z(n16273) );
  XNOR U16516 ( .A(n16272), .B(n16273), .Z(n16275) );
  XOR U16517 ( .A(n16274), .B(n16275), .Z(n16263) );
  XNOR U16518 ( .A(a[113]), .B(b[11]), .Z(n16307) );
  OR U16519 ( .A(n16307), .B(n18194), .Z(n16164) );
  NANDN U16520 ( .A(n16162), .B(n18104), .Z(n16163) );
  NAND U16521 ( .A(n16164), .B(n16163), .Z(n16261) );
  XOR U16522 ( .A(n580), .B(a[111]), .Z(n16310) );
  NANDN U16523 ( .A(n16310), .B(n18336), .Z(n16167) );
  NANDN U16524 ( .A(n16165), .B(n18337), .Z(n16166) );
  AND U16525 ( .A(n16167), .B(n16166), .Z(n16260) );
  XNOR U16526 ( .A(n16261), .B(n16260), .Z(n16262) );
  XNOR U16527 ( .A(n16263), .B(n16262), .Z(n16279) );
  NAND U16528 ( .A(n19406), .B(n16168), .Z(n16170) );
  XNOR U16529 ( .A(n584), .B(a[95]), .Z(n16325) );
  NANDN U16530 ( .A(n576), .B(n16325), .Z(n16169) );
  NAND U16531 ( .A(n16170), .B(n16169), .Z(n16236) );
  NANDN U16532 ( .A(n585), .B(a[91]), .Z(n16237) );
  XNOR U16533 ( .A(n16236), .B(n16237), .Z(n16239) );
  NANDN U16534 ( .A(n577), .B(a[123]), .Z(n16171) );
  XOR U16535 ( .A(n17151), .B(n16171), .Z(n16173) );
  IV U16536 ( .A(a[122]), .Z(n19276) );
  NANDN U16537 ( .A(n19276), .B(n577), .Z(n16172) );
  AND U16538 ( .A(n16173), .B(n16172), .Z(n16238) );
  XNOR U16539 ( .A(n16239), .B(n16238), .Z(n16277) );
  XOR U16540 ( .A(b[23]), .B(a[101]), .Z(n16316) );
  NANDN U16541 ( .A(n19127), .B(n16316), .Z(n16176) );
  NANDN U16542 ( .A(n16174), .B(n19128), .Z(n16175) );
  NAND U16543 ( .A(n16176), .B(n16175), .Z(n16331) );
  NANDN U16544 ( .A(n16177), .B(n17553), .Z(n16179) );
  XNOR U16545 ( .A(a[117]), .B(b[7]), .Z(n16319) );
  NANDN U16546 ( .A(n16319), .B(n17555), .Z(n16178) );
  NAND U16547 ( .A(n16179), .B(n16178), .Z(n16328) );
  XOR U16548 ( .A(b[25]), .B(a[99]), .Z(n16313) );
  NAND U16549 ( .A(n16313), .B(n19240), .Z(n16182) );
  NAND U16550 ( .A(n16180), .B(n19242), .Z(n16181) );
  AND U16551 ( .A(n16182), .B(n16181), .Z(n16329) );
  XNOR U16552 ( .A(n16328), .B(n16329), .Z(n16330) );
  XOR U16553 ( .A(n16331), .B(n16330), .Z(n16276) );
  XOR U16554 ( .A(n16279), .B(n16278), .Z(n16291) );
  XOR U16555 ( .A(n16290), .B(n16291), .Z(n16346) );
  XNOR U16556 ( .A(n16347), .B(n16346), .Z(n16349) );
  XNOR U16557 ( .A(n16348), .B(n16349), .Z(n16230) );
  XOR U16558 ( .A(n16231), .B(n16230), .Z(n16233) );
  NANDN U16559 ( .A(n16184), .B(n16183), .Z(n16188) );
  NAND U16560 ( .A(n16186), .B(n16185), .Z(n16187) );
  NAND U16561 ( .A(n16188), .B(n16187), .Z(n16225) );
  NAND U16562 ( .A(n16190), .B(n16189), .Z(n16194) );
  NANDN U16563 ( .A(n16192), .B(n16191), .Z(n16193) );
  AND U16564 ( .A(n16194), .B(n16193), .Z(n16224) );
  XNOR U16565 ( .A(n16225), .B(n16224), .Z(n16226) );
  XOR U16566 ( .A(n16227), .B(n16226), .Z(n16220) );
  NANDN U16567 ( .A(n16196), .B(n16195), .Z(n16200) );
  NAND U16568 ( .A(n16198), .B(n16197), .Z(n16199) );
  NAND U16569 ( .A(n16200), .B(n16199), .Z(n16218) );
  NANDN U16570 ( .A(n16202), .B(n16201), .Z(n16206) );
  NANDN U16571 ( .A(n16204), .B(n16203), .Z(n16205) );
  NAND U16572 ( .A(n16206), .B(n16205), .Z(n16219) );
  XNOR U16573 ( .A(n16218), .B(n16219), .Z(n16221) );
  XOR U16574 ( .A(n16220), .B(n16221), .Z(n16212) );
  XOR U16575 ( .A(n16213), .B(n16212), .Z(n16214) );
  XNOR U16576 ( .A(n16215), .B(n16214), .Z(n16352) );
  XNOR U16577 ( .A(n16352), .B(sreg[219]), .Z(n16354) );
  NAND U16578 ( .A(n16207), .B(sreg[218]), .Z(n16211) );
  OR U16579 ( .A(n16209), .B(n16208), .Z(n16210) );
  AND U16580 ( .A(n16211), .B(n16210), .Z(n16353) );
  XOR U16581 ( .A(n16354), .B(n16353), .Z(c[219]) );
  NAND U16582 ( .A(n16213), .B(n16212), .Z(n16217) );
  NAND U16583 ( .A(n16215), .B(n16214), .Z(n16216) );
  NAND U16584 ( .A(n16217), .B(n16216), .Z(n16360) );
  NANDN U16585 ( .A(n16219), .B(n16218), .Z(n16223) );
  NAND U16586 ( .A(n16221), .B(n16220), .Z(n16222) );
  NAND U16587 ( .A(n16223), .B(n16222), .Z(n16358) );
  NANDN U16588 ( .A(n16225), .B(n16224), .Z(n16229) );
  NAND U16589 ( .A(n16227), .B(n16226), .Z(n16228) );
  NAND U16590 ( .A(n16229), .B(n16228), .Z(n16363) );
  NANDN U16591 ( .A(n16231), .B(n16230), .Z(n16235) );
  OR U16592 ( .A(n16233), .B(n16232), .Z(n16234) );
  NAND U16593 ( .A(n16235), .B(n16234), .Z(n16364) );
  XNOR U16594 ( .A(n16363), .B(n16364), .Z(n16365) );
  NANDN U16595 ( .A(n16237), .B(n16236), .Z(n16241) );
  NAND U16596 ( .A(n16239), .B(n16238), .Z(n16240) );
  NAND U16597 ( .A(n16241), .B(n16240), .Z(n16440) );
  XOR U16598 ( .A(n581), .B(a[106]), .Z(n16412) );
  NANDN U16599 ( .A(n16412), .B(n18834), .Z(n16244) );
  NAND U16600 ( .A(n18832), .B(n16242), .Z(n16243) );
  NAND U16601 ( .A(n16244), .B(n16243), .Z(n16480) );
  XOR U16602 ( .A(n19188), .B(b[5]), .Z(n16415) );
  NANDN U16603 ( .A(n16415), .B(n17310), .Z(n16247) );
  NAND U16604 ( .A(n17311), .B(n16245), .Z(n16246) );
  AND U16605 ( .A(n16247), .B(n16246), .Z(n16479) );
  XNOR U16606 ( .A(n16480), .B(n16479), .Z(n16481) );
  XOR U16607 ( .A(n583), .B(a[98]), .Z(n16418) );
  NANDN U16608 ( .A(n16418), .B(n19336), .Z(n16250) );
  NAND U16609 ( .A(n19337), .B(n16248), .Z(n16249) );
  NAND U16610 ( .A(n16250), .B(n16249), .Z(n16482) );
  XOR U16611 ( .A(n16481), .B(n16482), .Z(n16437) );
  XNOR U16612 ( .A(b[17]), .B(a[108]), .Z(n16403) );
  NANDN U16613 ( .A(n16403), .B(n18673), .Z(n16253) );
  NAND U16614 ( .A(n16251), .B(n18674), .Z(n16252) );
  NAND U16615 ( .A(n16253), .B(n16252), .Z(n16394) );
  XOR U16616 ( .A(b[31]), .B(n16590), .Z(n16406) );
  NANDN U16617 ( .A(n16406), .B(n19472), .Z(n16256) );
  NANDN U16618 ( .A(n16254), .B(n19473), .Z(n16255) );
  NAND U16619 ( .A(n16256), .B(n16255), .Z(n16391) );
  OR U16620 ( .A(n16257), .B(n16988), .Z(n16259) );
  XOR U16621 ( .A(a[122]), .B(n578), .Z(n16409) );
  NANDN U16622 ( .A(n16409), .B(n16990), .Z(n16258) );
  AND U16623 ( .A(n16259), .B(n16258), .Z(n16392) );
  XNOR U16624 ( .A(n16391), .B(n16392), .Z(n16393) );
  XNOR U16625 ( .A(n16394), .B(n16393), .Z(n16438) );
  XNOR U16626 ( .A(n16437), .B(n16438), .Z(n16439) );
  XNOR U16627 ( .A(n16440), .B(n16439), .Z(n16376) );
  NANDN U16628 ( .A(n16261), .B(n16260), .Z(n16265) );
  NAND U16629 ( .A(n16263), .B(n16262), .Z(n16264) );
  NAND U16630 ( .A(n16265), .B(n16264), .Z(n16429) );
  NANDN U16631 ( .A(n16267), .B(n16266), .Z(n16271) );
  NAND U16632 ( .A(n16269), .B(n16268), .Z(n16270) );
  NAND U16633 ( .A(n16271), .B(n16270), .Z(n16428) );
  XNOR U16634 ( .A(n16428), .B(n16427), .Z(n16430) );
  XOR U16635 ( .A(n16429), .B(n16430), .Z(n16375) );
  XOR U16636 ( .A(n16376), .B(n16375), .Z(n16377) );
  NANDN U16637 ( .A(n16277), .B(n16276), .Z(n16281) );
  NAND U16638 ( .A(n16279), .B(n16278), .Z(n16280) );
  NAND U16639 ( .A(n16281), .B(n16280), .Z(n16378) );
  XNOR U16640 ( .A(n16377), .B(n16378), .Z(n16493) );
  OR U16641 ( .A(n16283), .B(n16282), .Z(n16287) );
  NAND U16642 ( .A(n16285), .B(n16284), .Z(n16286) );
  NAND U16643 ( .A(n16287), .B(n16286), .Z(n16492) );
  NANDN U16644 ( .A(n16289), .B(n16288), .Z(n16293) );
  NAND U16645 ( .A(n16291), .B(n16290), .Z(n16292) );
  NAND U16646 ( .A(n16293), .B(n16292), .Z(n16372) );
  XOR U16647 ( .A(a[116]), .B(n579), .Z(n16458) );
  NANDN U16648 ( .A(n16458), .B(n17814), .Z(n16300) );
  NANDN U16649 ( .A(n16298), .B(n17815), .Z(n16299) );
  NAND U16650 ( .A(n16300), .B(n16299), .Z(n16400) );
  NANDN U16651 ( .A(n16301), .B(n18513), .Z(n16303) );
  XNOR U16652 ( .A(b[15]), .B(a[110]), .Z(n16461) );
  OR U16653 ( .A(n16461), .B(n18512), .Z(n16302) );
  NAND U16654 ( .A(n16303), .B(n16302), .Z(n16397) );
  NANDN U16655 ( .A(n16304), .B(n19013), .Z(n16306) );
  XOR U16656 ( .A(b[21]), .B(n17716), .Z(n16464) );
  NANDN U16657 ( .A(n16464), .B(n19015), .Z(n16305) );
  AND U16658 ( .A(n16306), .B(n16305), .Z(n16398) );
  XNOR U16659 ( .A(n16397), .B(n16398), .Z(n16399) );
  XNOR U16660 ( .A(n16400), .B(n16399), .Z(n16388) );
  XOR U16661 ( .A(n18751), .B(b[11]), .Z(n16470) );
  OR U16662 ( .A(n16470), .B(n18194), .Z(n16309) );
  NANDN U16663 ( .A(n16307), .B(n18104), .Z(n16308) );
  NAND U16664 ( .A(n16309), .B(n16308), .Z(n16386) );
  XOR U16665 ( .A(n18582), .B(b[13]), .Z(n16467) );
  NANDN U16666 ( .A(n16467), .B(n18336), .Z(n16312) );
  NANDN U16667 ( .A(n16310), .B(n18337), .Z(n16311) );
  AND U16668 ( .A(n16312), .B(n16311), .Z(n16385) );
  XNOR U16669 ( .A(n16386), .B(n16385), .Z(n16387) );
  XNOR U16670 ( .A(n16388), .B(n16387), .Z(n16382) );
  XNOR U16671 ( .A(b[25]), .B(a[100]), .Z(n16455) );
  NANDN U16672 ( .A(n16455), .B(n19240), .Z(n16315) );
  NAND U16673 ( .A(n16313), .B(n19242), .Z(n16314) );
  NAND U16674 ( .A(n16315), .B(n16314), .Z(n16476) );
  XNOR U16675 ( .A(b[23]), .B(a[102]), .Z(n16449) );
  OR U16676 ( .A(n16449), .B(n19127), .Z(n16318) );
  NAND U16677 ( .A(n16316), .B(n19128), .Z(n16317) );
  NAND U16678 ( .A(n16318), .B(n16317), .Z(n16473) );
  NANDN U16679 ( .A(n16319), .B(n17553), .Z(n16321) );
  XNOR U16680 ( .A(a[118]), .B(b[7]), .Z(n16452) );
  NANDN U16681 ( .A(n16452), .B(n17555), .Z(n16320) );
  AND U16682 ( .A(n16321), .B(n16320), .Z(n16474) );
  XNOR U16683 ( .A(n16473), .B(n16474), .Z(n16475) );
  XNOR U16684 ( .A(n16476), .B(n16475), .Z(n16379) );
  NANDN U16685 ( .A(n577), .B(a[124]), .Z(n16322) );
  XOR U16686 ( .A(n17151), .B(n16322), .Z(n16324) );
  NANDN U16687 ( .A(b[0]), .B(a[123]), .Z(n16323) );
  AND U16688 ( .A(n16324), .B(n16323), .Z(n16423) );
  NAND U16689 ( .A(n19406), .B(n16325), .Z(n16327) );
  XNOR U16690 ( .A(n584), .B(a[96]), .Z(n16446) );
  NANDN U16691 ( .A(n576), .B(n16446), .Z(n16326) );
  NAND U16692 ( .A(n16327), .B(n16326), .Z(n16421) );
  NANDN U16693 ( .A(n585), .B(a[92]), .Z(n16422) );
  XNOR U16694 ( .A(n16421), .B(n16422), .Z(n16424) );
  XOR U16695 ( .A(n16423), .B(n16424), .Z(n16380) );
  XNOR U16696 ( .A(n16379), .B(n16380), .Z(n16381) );
  XOR U16697 ( .A(n16382), .B(n16381), .Z(n16434) );
  NANDN U16698 ( .A(n16329), .B(n16328), .Z(n16333) );
  NAND U16699 ( .A(n16331), .B(n16330), .Z(n16332) );
  NAND U16700 ( .A(n16333), .B(n16332), .Z(n16431) );
  NANDN U16701 ( .A(n16335), .B(n16334), .Z(n16339) );
  NAND U16702 ( .A(n16337), .B(n16336), .Z(n16338) );
  AND U16703 ( .A(n16339), .B(n16338), .Z(n16432) );
  XNOR U16704 ( .A(n16431), .B(n16432), .Z(n16433) );
  XNOR U16705 ( .A(n16434), .B(n16433), .Z(n16370) );
  XNOR U16706 ( .A(n16369), .B(n16370), .Z(n16371) );
  XOR U16707 ( .A(n16372), .B(n16371), .Z(n16491) );
  XOR U16708 ( .A(n16492), .B(n16491), .Z(n16494) );
  NANDN U16709 ( .A(n16341), .B(n16340), .Z(n16345) );
  OR U16710 ( .A(n16343), .B(n16342), .Z(n16344) );
  NAND U16711 ( .A(n16345), .B(n16344), .Z(n16485) );
  NAND U16712 ( .A(n16347), .B(n16346), .Z(n16351) );
  NANDN U16713 ( .A(n16349), .B(n16348), .Z(n16350) );
  NAND U16714 ( .A(n16351), .B(n16350), .Z(n16486) );
  XNOR U16715 ( .A(n16485), .B(n16486), .Z(n16487) );
  XOR U16716 ( .A(n16488), .B(n16487), .Z(n16366) );
  XOR U16717 ( .A(n16365), .B(n16366), .Z(n16357) );
  XOR U16718 ( .A(n16358), .B(n16357), .Z(n16359) );
  XNOR U16719 ( .A(n16360), .B(n16359), .Z(n16497) );
  XNOR U16720 ( .A(n16497), .B(sreg[220]), .Z(n16499) );
  NAND U16721 ( .A(n16352), .B(sreg[219]), .Z(n16356) );
  OR U16722 ( .A(n16354), .B(n16353), .Z(n16355) );
  AND U16723 ( .A(n16356), .B(n16355), .Z(n16498) );
  XOR U16724 ( .A(n16499), .B(n16498), .Z(c[220]) );
  NAND U16725 ( .A(n16358), .B(n16357), .Z(n16362) );
  NAND U16726 ( .A(n16360), .B(n16359), .Z(n16361) );
  NAND U16727 ( .A(n16362), .B(n16361), .Z(n16505) );
  NANDN U16728 ( .A(n16364), .B(n16363), .Z(n16368) );
  NAND U16729 ( .A(n16366), .B(n16365), .Z(n16367) );
  NAND U16730 ( .A(n16368), .B(n16367), .Z(n16502) );
  NANDN U16731 ( .A(n16370), .B(n16369), .Z(n16374) );
  NAND U16732 ( .A(n16372), .B(n16371), .Z(n16373) );
  NAND U16733 ( .A(n16374), .B(n16373), .Z(n16633) );
  XNOR U16734 ( .A(n16633), .B(n16634), .Z(n16635) );
  NANDN U16735 ( .A(n16380), .B(n16379), .Z(n16384) );
  NANDN U16736 ( .A(n16382), .B(n16381), .Z(n16383) );
  NAND U16737 ( .A(n16384), .B(n16383), .Z(n16523) );
  NANDN U16738 ( .A(n16386), .B(n16385), .Z(n16390) );
  NAND U16739 ( .A(n16388), .B(n16387), .Z(n16389) );
  NAND U16740 ( .A(n16390), .B(n16389), .Z(n16577) );
  NANDN U16741 ( .A(n16392), .B(n16391), .Z(n16396) );
  NAND U16742 ( .A(n16394), .B(n16393), .Z(n16395) );
  NAND U16743 ( .A(n16396), .B(n16395), .Z(n16575) );
  NANDN U16744 ( .A(n16398), .B(n16397), .Z(n16402) );
  NAND U16745 ( .A(n16400), .B(n16399), .Z(n16401) );
  AND U16746 ( .A(n16402), .B(n16401), .Z(n16574) );
  XNOR U16747 ( .A(n16575), .B(n16574), .Z(n16576) );
  XNOR U16748 ( .A(n16577), .B(n16576), .Z(n16520) );
  XOR U16749 ( .A(b[17]), .B(a[109]), .Z(n16532) );
  NAND U16750 ( .A(n16532), .B(n18673), .Z(n16405) );
  NANDN U16751 ( .A(n16403), .B(n18674), .Z(n16404) );
  NAND U16752 ( .A(n16405), .B(n16404), .Z(n16565) );
  XNOR U16753 ( .A(b[31]), .B(a[95]), .Z(n16535) );
  NANDN U16754 ( .A(n16535), .B(n19472), .Z(n16408) );
  NANDN U16755 ( .A(n16406), .B(n19473), .Z(n16407) );
  NAND U16756 ( .A(n16408), .B(n16407), .Z(n16562) );
  OR U16757 ( .A(n16409), .B(n16988), .Z(n16411) );
  XNOR U16758 ( .A(a[123]), .B(b[3]), .Z(n16538) );
  NANDN U16759 ( .A(n16538), .B(n16990), .Z(n16410) );
  AND U16760 ( .A(n16411), .B(n16410), .Z(n16563) );
  XNOR U16761 ( .A(n16562), .B(n16563), .Z(n16564) );
  XNOR U16762 ( .A(n16565), .B(n16564), .Z(n16586) );
  XNOR U16763 ( .A(b[19]), .B(a[107]), .Z(n16547) );
  NANDN U16764 ( .A(n16547), .B(n18834), .Z(n16414) );
  NANDN U16765 ( .A(n16412), .B(n18832), .Z(n16413) );
  NAND U16766 ( .A(n16414), .B(n16413), .Z(n16628) );
  XNOR U16767 ( .A(a[121]), .B(b[5]), .Z(n16544) );
  NANDN U16768 ( .A(n16544), .B(n17310), .Z(n16417) );
  NANDN U16769 ( .A(n16415), .B(n17311), .Z(n16416) );
  AND U16770 ( .A(n16417), .B(n16416), .Z(n16627) );
  XNOR U16771 ( .A(n16628), .B(n16627), .Z(n16629) );
  XNOR U16772 ( .A(b[27]), .B(a[99]), .Z(n16541) );
  NANDN U16773 ( .A(n16541), .B(n19336), .Z(n16420) );
  NANDN U16774 ( .A(n16418), .B(n19337), .Z(n16419) );
  AND U16775 ( .A(n16420), .B(n16419), .Z(n16630) );
  XNOR U16776 ( .A(n16629), .B(n16630), .Z(n16587) );
  XNOR U16777 ( .A(n16586), .B(n16587), .Z(n16588) );
  NANDN U16778 ( .A(n16422), .B(n16421), .Z(n16426) );
  NAND U16779 ( .A(n16424), .B(n16423), .Z(n16425) );
  AND U16780 ( .A(n16426), .B(n16425), .Z(n16589) );
  XNOR U16781 ( .A(n16588), .B(n16589), .Z(n16521) );
  XOR U16782 ( .A(n16520), .B(n16521), .Z(n16522) );
  XOR U16783 ( .A(n16523), .B(n16522), .Z(n16641) );
  NANDN U16784 ( .A(n16432), .B(n16431), .Z(n16436) );
  NAND U16785 ( .A(n16434), .B(n16433), .Z(n16435) );
  NAND U16786 ( .A(n16436), .B(n16435), .Z(n16517) );
  NANDN U16787 ( .A(n16438), .B(n16437), .Z(n16442) );
  NAND U16788 ( .A(n16440), .B(n16439), .Z(n16441) );
  NAND U16789 ( .A(n16442), .B(n16441), .Z(n16514) );
  IV U16790 ( .A(a[125]), .Z(n19402) );
  NANDN U16791 ( .A(n19402), .B(b[0]), .Z(n16443) );
  XOR U16792 ( .A(n17151), .B(n16443), .Z(n16445) );
  IV U16793 ( .A(a[124]), .Z(n19373) );
  NANDN U16794 ( .A(n19373), .B(n577), .Z(n16444) );
  AND U16795 ( .A(n16445), .B(n16444), .Z(n16552) );
  NAND U16796 ( .A(n19406), .B(n16446), .Z(n16448) );
  XOR U16797 ( .A(b[29]), .B(n17038), .Z(n16594) );
  OR U16798 ( .A(n16594), .B(n576), .Z(n16447) );
  NAND U16799 ( .A(n16448), .B(n16447), .Z(n16550) );
  NANDN U16800 ( .A(n585), .B(a[93]), .Z(n16551) );
  XNOR U16801 ( .A(n16550), .B(n16551), .Z(n16553) );
  XOR U16802 ( .A(n16552), .B(n16553), .Z(n16529) );
  XOR U16803 ( .A(b[23]), .B(a[103]), .Z(n16600) );
  NANDN U16804 ( .A(n19127), .B(n16600), .Z(n16451) );
  NANDN U16805 ( .A(n16449), .B(n19128), .Z(n16450) );
  NAND U16806 ( .A(n16451), .B(n16450), .Z(n16624) );
  NANDN U16807 ( .A(n16452), .B(n17553), .Z(n16454) );
  XNOR U16808 ( .A(a[119]), .B(b[7]), .Z(n16603) );
  NANDN U16809 ( .A(n16603), .B(n17555), .Z(n16453) );
  NAND U16810 ( .A(n16454), .B(n16453), .Z(n16621) );
  XOR U16811 ( .A(b[25]), .B(a[101]), .Z(n16597) );
  NAND U16812 ( .A(n16597), .B(n19240), .Z(n16457) );
  NANDN U16813 ( .A(n16455), .B(n19242), .Z(n16456) );
  AND U16814 ( .A(n16457), .B(n16456), .Z(n16622) );
  XNOR U16815 ( .A(n16621), .B(n16622), .Z(n16623) );
  XNOR U16816 ( .A(n16624), .B(n16623), .Z(n16526) );
  XOR U16817 ( .A(a[117]), .B(n579), .Z(n16615) );
  NANDN U16818 ( .A(n16615), .B(n17814), .Z(n16460) );
  NANDN U16819 ( .A(n16458), .B(n17815), .Z(n16459) );
  NAND U16820 ( .A(n16460), .B(n16459), .Z(n16571) );
  NANDN U16821 ( .A(n16461), .B(n18513), .Z(n16463) );
  XOR U16822 ( .A(b[15]), .B(a[111]), .Z(n16618) );
  NANDN U16823 ( .A(n18512), .B(n16618), .Z(n16462) );
  NAND U16824 ( .A(n16463), .B(n16462), .Z(n16568) );
  NANDN U16825 ( .A(n16464), .B(n19013), .Z(n16466) );
  XNOR U16826 ( .A(b[21]), .B(a[105]), .Z(n16612) );
  NANDN U16827 ( .A(n16612), .B(n19015), .Z(n16465) );
  AND U16828 ( .A(n16466), .B(n16465), .Z(n16569) );
  XNOR U16829 ( .A(n16568), .B(n16569), .Z(n16570) );
  XNOR U16830 ( .A(n16571), .B(n16570), .Z(n16559) );
  XNOR U16831 ( .A(a[113]), .B(b[13]), .Z(n16609) );
  NANDN U16832 ( .A(n16609), .B(n18336), .Z(n16469) );
  NANDN U16833 ( .A(n16467), .B(n18337), .Z(n16468) );
  NAND U16834 ( .A(n16469), .B(n16468), .Z(n16557) );
  XNOR U16835 ( .A(a[115]), .B(b[11]), .Z(n16606) );
  OR U16836 ( .A(n16606), .B(n18194), .Z(n16472) );
  NANDN U16837 ( .A(n16470), .B(n18104), .Z(n16471) );
  AND U16838 ( .A(n16472), .B(n16471), .Z(n16556) );
  XNOR U16839 ( .A(n16557), .B(n16556), .Z(n16558) );
  XNOR U16840 ( .A(n16559), .B(n16558), .Z(n16527) );
  XNOR U16841 ( .A(n16529), .B(n16528), .Z(n16583) );
  NANDN U16842 ( .A(n16474), .B(n16473), .Z(n16478) );
  NAND U16843 ( .A(n16476), .B(n16475), .Z(n16477) );
  NAND U16844 ( .A(n16478), .B(n16477), .Z(n16580) );
  NANDN U16845 ( .A(n16480), .B(n16479), .Z(n16484) );
  NANDN U16846 ( .A(n16482), .B(n16481), .Z(n16483) );
  NAND U16847 ( .A(n16484), .B(n16483), .Z(n16581) );
  XNOR U16848 ( .A(n16580), .B(n16581), .Z(n16582) );
  XOR U16849 ( .A(n16583), .B(n16582), .Z(n16515) );
  XNOR U16850 ( .A(n16514), .B(n16515), .Z(n16516) );
  XNOR U16851 ( .A(n16517), .B(n16516), .Z(n16639) );
  XNOR U16852 ( .A(n16640), .B(n16639), .Z(n16642) );
  XNOR U16853 ( .A(n16641), .B(n16642), .Z(n16636) );
  XOR U16854 ( .A(n16635), .B(n16636), .Z(n16511) );
  NANDN U16855 ( .A(n16486), .B(n16485), .Z(n16490) );
  NAND U16856 ( .A(n16488), .B(n16487), .Z(n16489) );
  NAND U16857 ( .A(n16490), .B(n16489), .Z(n16508) );
  NANDN U16858 ( .A(n16492), .B(n16491), .Z(n16496) );
  OR U16859 ( .A(n16494), .B(n16493), .Z(n16495) );
  NAND U16860 ( .A(n16496), .B(n16495), .Z(n16509) );
  XNOR U16861 ( .A(n16508), .B(n16509), .Z(n16510) );
  XNOR U16862 ( .A(n16511), .B(n16510), .Z(n16503) );
  XNOR U16863 ( .A(n16502), .B(n16503), .Z(n16504) );
  XNOR U16864 ( .A(n16505), .B(n16504), .Z(n16645) );
  XNOR U16865 ( .A(n16645), .B(sreg[221]), .Z(n16647) );
  NAND U16866 ( .A(n16497), .B(sreg[220]), .Z(n16501) );
  OR U16867 ( .A(n16499), .B(n16498), .Z(n16500) );
  AND U16868 ( .A(n16501), .B(n16500), .Z(n16646) );
  XOR U16869 ( .A(n16647), .B(n16646), .Z(c[221]) );
  NANDN U16870 ( .A(n16503), .B(n16502), .Z(n16507) );
  NAND U16871 ( .A(n16505), .B(n16504), .Z(n16506) );
  NAND U16872 ( .A(n16507), .B(n16506), .Z(n16653) );
  NANDN U16873 ( .A(n16509), .B(n16508), .Z(n16513) );
  NAND U16874 ( .A(n16511), .B(n16510), .Z(n16512) );
  NAND U16875 ( .A(n16513), .B(n16512), .Z(n16650) );
  NANDN U16876 ( .A(n16515), .B(n16514), .Z(n16519) );
  NAND U16877 ( .A(n16517), .B(n16516), .Z(n16518) );
  NAND U16878 ( .A(n16519), .B(n16518), .Z(n16666) );
  OR U16879 ( .A(n16521), .B(n16520), .Z(n16525) );
  NAND U16880 ( .A(n16523), .B(n16522), .Z(n16524) );
  NAND U16881 ( .A(n16525), .B(n16524), .Z(n16667) );
  XNOR U16882 ( .A(n16666), .B(n16667), .Z(n16668) );
  NANDN U16883 ( .A(n16527), .B(n16526), .Z(n16531) );
  NANDN U16884 ( .A(n16529), .B(n16528), .Z(n16530) );
  NAND U16885 ( .A(n16531), .B(n16530), .Z(n16789) );
  XNOR U16886 ( .A(b[17]), .B(a[110]), .Z(n16741) );
  NANDN U16887 ( .A(n16741), .B(n18673), .Z(n16534) );
  NAND U16888 ( .A(n16532), .B(n18674), .Z(n16533) );
  NAND U16889 ( .A(n16534), .B(n16533), .Z(n16764) );
  XNOR U16890 ( .A(b[31]), .B(a[96]), .Z(n16744) );
  NANDN U16891 ( .A(n16744), .B(n19472), .Z(n16537) );
  NANDN U16892 ( .A(n16535), .B(n19473), .Z(n16536) );
  AND U16893 ( .A(n16537), .B(n16536), .Z(n16762) );
  OR U16894 ( .A(n16538), .B(n16988), .Z(n16540) );
  XOR U16895 ( .A(a[124]), .B(n578), .Z(n16747) );
  NANDN U16896 ( .A(n16747), .B(n16990), .Z(n16539) );
  AND U16897 ( .A(n16540), .B(n16539), .Z(n16763) );
  XOR U16898 ( .A(n16764), .B(n16765), .Z(n16678) );
  XOR U16899 ( .A(n583), .B(n17447), .Z(n16738) );
  NAND U16900 ( .A(n19336), .B(n16738), .Z(n16543) );
  NANDN U16901 ( .A(n16541), .B(n19337), .Z(n16542) );
  NAND U16902 ( .A(n16543), .B(n16542), .Z(n16723) );
  XNOR U16903 ( .A(n19276), .B(b[5]), .Z(n16735) );
  NAND U16904 ( .A(n16735), .B(n17310), .Z(n16546) );
  NANDN U16905 ( .A(n16544), .B(n17311), .Z(n16545) );
  NAND U16906 ( .A(n16546), .B(n16545), .Z(n16720) );
  NANDN U16907 ( .A(n16547), .B(n18832), .Z(n16549) );
  XOR U16908 ( .A(n581), .B(n18198), .Z(n16732) );
  NAND U16909 ( .A(n16732), .B(n18834), .Z(n16548) );
  AND U16910 ( .A(n16549), .B(n16548), .Z(n16721) );
  XNOR U16911 ( .A(n16720), .B(n16721), .Z(n16722) );
  XOR U16912 ( .A(n16723), .B(n16722), .Z(n16679) );
  XNOR U16913 ( .A(n16678), .B(n16679), .Z(n16680) );
  NANDN U16914 ( .A(n16551), .B(n16550), .Z(n16555) );
  NAND U16915 ( .A(n16553), .B(n16552), .Z(n16554) );
  AND U16916 ( .A(n16555), .B(n16554), .Z(n16681) );
  XNOR U16917 ( .A(n16680), .B(n16681), .Z(n16787) );
  NANDN U16918 ( .A(n16557), .B(n16556), .Z(n16561) );
  NAND U16919 ( .A(n16559), .B(n16558), .Z(n16560) );
  NAND U16920 ( .A(n16561), .B(n16560), .Z(n16729) );
  NANDN U16921 ( .A(n16563), .B(n16562), .Z(n16567) );
  NAND U16922 ( .A(n16565), .B(n16564), .Z(n16566) );
  NAND U16923 ( .A(n16567), .B(n16566), .Z(n16727) );
  NANDN U16924 ( .A(n16569), .B(n16568), .Z(n16573) );
  NAND U16925 ( .A(n16571), .B(n16570), .Z(n16572) );
  AND U16926 ( .A(n16573), .B(n16572), .Z(n16726) );
  XNOR U16927 ( .A(n16727), .B(n16726), .Z(n16728) );
  XOR U16928 ( .A(n16729), .B(n16728), .Z(n16786) );
  XNOR U16929 ( .A(n16787), .B(n16786), .Z(n16788) );
  XNOR U16930 ( .A(n16789), .B(n16788), .Z(n16665) );
  NANDN U16931 ( .A(n16575), .B(n16574), .Z(n16579) );
  NAND U16932 ( .A(n16577), .B(n16576), .Z(n16578) );
  NAND U16933 ( .A(n16579), .B(n16578), .Z(n16663) );
  NANDN U16934 ( .A(n16581), .B(n16580), .Z(n16585) );
  NANDN U16935 ( .A(n16583), .B(n16582), .Z(n16584) );
  NAND U16936 ( .A(n16585), .B(n16584), .Z(n16780) );
  XNOR U16937 ( .A(n16780), .B(n16781), .Z(n16782) );
  ANDN U16938 ( .B(b[31]), .A(n16590), .Z(n16753) );
  IV U16939 ( .A(a[126]), .Z(n19295) );
  NANDN U16940 ( .A(n19295), .B(b[0]), .Z(n16591) );
  XOR U16941 ( .A(n17151), .B(n16591), .Z(n16593) );
  NANDN U16942 ( .A(n19402), .B(n577), .Z(n16592) );
  AND U16943 ( .A(n16593), .B(n16592), .Z(n16751) );
  NANDN U16944 ( .A(n16594), .B(n19406), .Z(n16596) );
  XNOR U16945 ( .A(n584), .B(a[98]), .Z(n16696) );
  NANDN U16946 ( .A(n576), .B(n16696), .Z(n16595) );
  AND U16947 ( .A(n16596), .B(n16595), .Z(n16750) );
  XNOR U16948 ( .A(n16751), .B(n16750), .Z(n16752) );
  XOR U16949 ( .A(n16753), .B(n16752), .Z(n16774) );
  XNOR U16950 ( .A(b[25]), .B(a[102]), .Z(n16684) );
  NANDN U16951 ( .A(n16684), .B(n19240), .Z(n16599) );
  NAND U16952 ( .A(n16597), .B(n19242), .Z(n16598) );
  NAND U16953 ( .A(n16599), .B(n16598), .Z(n16717) );
  XNOR U16954 ( .A(b[23]), .B(a[104]), .Z(n16687) );
  OR U16955 ( .A(n16687), .B(n19127), .Z(n16602) );
  NAND U16956 ( .A(n16600), .B(n19128), .Z(n16601) );
  NAND U16957 ( .A(n16602), .B(n16601), .Z(n16714) );
  NANDN U16958 ( .A(n16603), .B(n17553), .Z(n16605) );
  XNOR U16959 ( .A(a[120]), .B(b[7]), .Z(n16690) );
  NANDN U16960 ( .A(n16690), .B(n17555), .Z(n16604) );
  AND U16961 ( .A(n16605), .B(n16604), .Z(n16715) );
  XNOR U16962 ( .A(n16714), .B(n16715), .Z(n16716) );
  XNOR U16963 ( .A(n16717), .B(n16716), .Z(n16775) );
  XOR U16964 ( .A(n16774), .B(n16775), .Z(n16777) );
  XNOR U16965 ( .A(n18950), .B(b[11]), .Z(n16711) );
  NANDN U16966 ( .A(n18194), .B(n16711), .Z(n16608) );
  NANDN U16967 ( .A(n16606), .B(n18104), .Z(n16607) );
  AND U16968 ( .A(n16608), .B(n16607), .Z(n16759) );
  XOR U16969 ( .A(n18751), .B(n580), .Z(n16708) );
  NAND U16970 ( .A(n16708), .B(n18336), .Z(n16611) );
  NANDN U16971 ( .A(n16609), .B(n18337), .Z(n16610) );
  AND U16972 ( .A(n16611), .B(n16610), .Z(n16756) );
  NANDN U16973 ( .A(n16612), .B(n19013), .Z(n16614) );
  XOR U16974 ( .A(b[21]), .B(n17690), .Z(n16705) );
  NANDN U16975 ( .A(n16705), .B(n19015), .Z(n16613) );
  AND U16976 ( .A(n16614), .B(n16613), .Z(n16768) );
  XOR U16977 ( .A(a[118]), .B(n579), .Z(n16702) );
  NANDN U16978 ( .A(n16702), .B(n17814), .Z(n16617) );
  NANDN U16979 ( .A(n16615), .B(n17815), .Z(n16616) );
  AND U16980 ( .A(n16617), .B(n16616), .Z(n16769) );
  NAND U16981 ( .A(n16618), .B(n18513), .Z(n16620) );
  XNOR U16982 ( .A(b[15]), .B(a[112]), .Z(n16699) );
  OR U16983 ( .A(n16699), .B(n18512), .Z(n16619) );
  NAND U16984 ( .A(n16620), .B(n16619), .Z(n16771) );
  XNOR U16985 ( .A(n16770), .B(n16771), .Z(n16757) );
  XOR U16986 ( .A(n16759), .B(n16758), .Z(n16776) );
  XNOR U16987 ( .A(n16777), .B(n16776), .Z(n16674) );
  NANDN U16988 ( .A(n16622), .B(n16621), .Z(n16626) );
  NAND U16989 ( .A(n16624), .B(n16623), .Z(n16625) );
  NAND U16990 ( .A(n16626), .B(n16625), .Z(n16672) );
  NANDN U16991 ( .A(n16628), .B(n16627), .Z(n16632) );
  NAND U16992 ( .A(n16630), .B(n16629), .Z(n16631) );
  NAND U16993 ( .A(n16632), .B(n16631), .Z(n16673) );
  XNOR U16994 ( .A(n16672), .B(n16673), .Z(n16675) );
  XOR U16995 ( .A(n16674), .B(n16675), .Z(n16783) );
  XOR U16996 ( .A(n16782), .B(n16783), .Z(n16662) );
  XNOR U16997 ( .A(n16663), .B(n16662), .Z(n16664) );
  XOR U16998 ( .A(n16665), .B(n16664), .Z(n16669) );
  XNOR U16999 ( .A(n16668), .B(n16669), .Z(n16659) );
  NANDN U17000 ( .A(n16634), .B(n16633), .Z(n16638) );
  NANDN U17001 ( .A(n16636), .B(n16635), .Z(n16637) );
  NAND U17002 ( .A(n16638), .B(n16637), .Z(n16657) );
  OR U17003 ( .A(n16640), .B(n16639), .Z(n16644) );
  OR U17004 ( .A(n16642), .B(n16641), .Z(n16643) );
  AND U17005 ( .A(n16644), .B(n16643), .Z(n16656) );
  XNOR U17006 ( .A(n16657), .B(n16656), .Z(n16658) );
  XNOR U17007 ( .A(n16659), .B(n16658), .Z(n16651) );
  XNOR U17008 ( .A(n16650), .B(n16651), .Z(n16652) );
  XNOR U17009 ( .A(n16653), .B(n16652), .Z(n16790) );
  XNOR U17010 ( .A(n16790), .B(sreg[222]), .Z(n16792) );
  NAND U17011 ( .A(n16645), .B(sreg[221]), .Z(n16649) );
  OR U17012 ( .A(n16647), .B(n16646), .Z(n16648) );
  AND U17013 ( .A(n16649), .B(n16648), .Z(n16791) );
  XOR U17014 ( .A(n16792), .B(n16791), .Z(c[222]) );
  NANDN U17015 ( .A(n16651), .B(n16650), .Z(n16655) );
  NAND U17016 ( .A(n16653), .B(n16652), .Z(n16654) );
  NAND U17017 ( .A(n16655), .B(n16654), .Z(n16798) );
  NANDN U17018 ( .A(n16657), .B(n16656), .Z(n16661) );
  NAND U17019 ( .A(n16659), .B(n16658), .Z(n16660) );
  NAND U17020 ( .A(n16661), .B(n16660), .Z(n16795) );
  NANDN U17021 ( .A(n16667), .B(n16666), .Z(n16671) );
  NAND U17022 ( .A(n16669), .B(n16668), .Z(n16670) );
  AND U17023 ( .A(n16671), .B(n16670), .Z(n16933) );
  XNOR U17024 ( .A(n16932), .B(n16933), .Z(n16934) );
  NANDN U17025 ( .A(n16673), .B(n16672), .Z(n16677) );
  NAND U17026 ( .A(n16675), .B(n16674), .Z(n16676) );
  NAND U17027 ( .A(n16677), .B(n16676), .Z(n16917) );
  NANDN U17028 ( .A(n16679), .B(n16678), .Z(n16683) );
  NAND U17029 ( .A(n16681), .B(n16680), .Z(n16682) );
  NAND U17030 ( .A(n16683), .B(n16682), .Z(n16914) );
  XOR U17031 ( .A(b[25]), .B(a[103]), .Z(n16837) );
  NAND U17032 ( .A(n16837), .B(n19240), .Z(n16686) );
  NANDN U17033 ( .A(n16684), .B(n19242), .Z(n16685) );
  NAND U17034 ( .A(n16686), .B(n16685), .Z(n16828) );
  XOR U17035 ( .A(b[23]), .B(a[105]), .Z(n16831) );
  NANDN U17036 ( .A(n19127), .B(n16831), .Z(n16689) );
  NANDN U17037 ( .A(n16687), .B(n19128), .Z(n16688) );
  NAND U17038 ( .A(n16689), .B(n16688), .Z(n16825) );
  NANDN U17039 ( .A(n16690), .B(n17553), .Z(n16692) );
  XNOR U17040 ( .A(a[121]), .B(b[7]), .Z(n16834) );
  NANDN U17041 ( .A(n16834), .B(n17555), .Z(n16691) );
  AND U17042 ( .A(n16692), .B(n16691), .Z(n16826) );
  XNOR U17043 ( .A(n16825), .B(n16826), .Z(n16827) );
  XOR U17044 ( .A(n16828), .B(n16827), .Z(n16866) );
  NANDN U17045 ( .A(n577), .B(a[127]), .Z(n16693) );
  XOR U17046 ( .A(n17151), .B(n16693), .Z(n16695) );
  NANDN U17047 ( .A(n19295), .B(n577), .Z(n16694) );
  AND U17048 ( .A(n16695), .B(n16694), .Z(n16874) );
  NAND U17049 ( .A(n16696), .B(n19406), .Z(n16698) );
  XNOR U17050 ( .A(n584), .B(a[99]), .Z(n16842) );
  NANDN U17051 ( .A(n576), .B(n16842), .Z(n16697) );
  NAND U17052 ( .A(n16698), .B(n16697), .Z(n16872) );
  NANDN U17053 ( .A(n585), .B(a[95]), .Z(n16873) );
  XNOR U17054 ( .A(n16872), .B(n16873), .Z(n16875) );
  XOR U17055 ( .A(n16874), .B(n16875), .Z(n16867) );
  XNOR U17056 ( .A(n16866), .B(n16867), .Z(n16869) );
  NANDN U17057 ( .A(n16699), .B(n18513), .Z(n16701) );
  XOR U17058 ( .A(b[15]), .B(a[113]), .Z(n16845) );
  NANDN U17059 ( .A(n18512), .B(n16845), .Z(n16700) );
  NAND U17060 ( .A(n16701), .B(n16700), .Z(n16910) );
  XOR U17061 ( .A(a[119]), .B(n579), .Z(n16851) );
  NANDN U17062 ( .A(n16851), .B(n17814), .Z(n16704) );
  NANDN U17063 ( .A(n16702), .B(n17815), .Z(n16703) );
  AND U17064 ( .A(n16704), .B(n16703), .Z(n16908) );
  NANDN U17065 ( .A(n16705), .B(n19013), .Z(n16707) );
  XNOR U17066 ( .A(b[21]), .B(a[107]), .Z(n16848) );
  NANDN U17067 ( .A(n16848), .B(n19015), .Z(n16706) );
  AND U17068 ( .A(n16707), .B(n16706), .Z(n16909) );
  XOR U17069 ( .A(n16910), .B(n16911), .Z(n16905) );
  XOR U17070 ( .A(n19022), .B(b[13]), .Z(n16854) );
  NANDN U17071 ( .A(n16854), .B(n18336), .Z(n16710) );
  NAND U17072 ( .A(n18337), .B(n16708), .Z(n16709) );
  NAND U17073 ( .A(n16710), .B(n16709), .Z(n16903) );
  XOR U17074 ( .A(n19136), .B(b[11]), .Z(n16857) );
  OR U17075 ( .A(n16857), .B(n18194), .Z(n16713) );
  NAND U17076 ( .A(n18104), .B(n16711), .Z(n16712) );
  AND U17077 ( .A(n16713), .B(n16712), .Z(n16902) );
  XNOR U17078 ( .A(n16903), .B(n16902), .Z(n16904) );
  XOR U17079 ( .A(n16905), .B(n16904), .Z(n16868) );
  XNOR U17080 ( .A(n16869), .B(n16868), .Z(n16816) );
  NANDN U17081 ( .A(n16715), .B(n16714), .Z(n16719) );
  NAND U17082 ( .A(n16717), .B(n16716), .Z(n16718) );
  NAND U17083 ( .A(n16719), .B(n16718), .Z(n16813) );
  NANDN U17084 ( .A(n16721), .B(n16720), .Z(n16725) );
  NAND U17085 ( .A(n16723), .B(n16722), .Z(n16724) );
  AND U17086 ( .A(n16725), .B(n16724), .Z(n16814) );
  XNOR U17087 ( .A(n16813), .B(n16814), .Z(n16815) );
  XOR U17088 ( .A(n16816), .B(n16815), .Z(n16915) );
  XOR U17089 ( .A(n16914), .B(n16915), .Z(n16916) );
  XNOR U17090 ( .A(n16917), .B(n16916), .Z(n16929) );
  NANDN U17091 ( .A(n16727), .B(n16726), .Z(n16731) );
  NAND U17092 ( .A(n16729), .B(n16728), .Z(n16730) );
  NAND U17093 ( .A(n16731), .B(n16730), .Z(n16927) );
  XNOR U17094 ( .A(b[19]), .B(a[109]), .Z(n16887) );
  NANDN U17095 ( .A(n16887), .B(n18834), .Z(n16734) );
  NAND U17096 ( .A(n18832), .B(n16732), .Z(n16733) );
  NAND U17097 ( .A(n16734), .B(n16733), .Z(n16820) );
  XOR U17098 ( .A(a[123]), .B(b[5]), .Z(n16893) );
  NAND U17099 ( .A(n17310), .B(n16893), .Z(n16737) );
  NAND U17100 ( .A(n17311), .B(n16735), .Z(n16736) );
  AND U17101 ( .A(n16737), .B(n16736), .Z(n16819) );
  XNOR U17102 ( .A(n16820), .B(n16819), .Z(n16821) );
  XNOR U17103 ( .A(b[27]), .B(a[101]), .Z(n16890) );
  NANDN U17104 ( .A(n16890), .B(n19336), .Z(n16740) );
  NAND U17105 ( .A(n19337), .B(n16738), .Z(n16739) );
  NAND U17106 ( .A(n16740), .B(n16739), .Z(n16822) );
  XOR U17107 ( .A(n16821), .B(n16822), .Z(n16860) );
  XOR U17108 ( .A(b[17]), .B(a[111]), .Z(n16878) );
  NAND U17109 ( .A(n16878), .B(n18673), .Z(n16743) );
  NANDN U17110 ( .A(n16741), .B(n18674), .Z(n16742) );
  NAND U17111 ( .A(n16743), .B(n16742), .Z(n16899) );
  XOR U17112 ( .A(b[31]), .B(n17038), .Z(n16881) );
  NANDN U17113 ( .A(n16881), .B(n19472), .Z(n16746) );
  NANDN U17114 ( .A(n16744), .B(n19473), .Z(n16745) );
  NAND U17115 ( .A(n16746), .B(n16745), .Z(n16896) );
  OR U17116 ( .A(n16747), .B(n16988), .Z(n16749) );
  XOR U17117 ( .A(a[125]), .B(n578), .Z(n16884) );
  NANDN U17118 ( .A(n16884), .B(n16990), .Z(n16748) );
  AND U17119 ( .A(n16749), .B(n16748), .Z(n16897) );
  XNOR U17120 ( .A(n16896), .B(n16897), .Z(n16898) );
  XNOR U17121 ( .A(n16899), .B(n16898), .Z(n16861) );
  XNOR U17122 ( .A(n16860), .B(n16861), .Z(n16862) );
  NANDN U17123 ( .A(n16751), .B(n16750), .Z(n16755) );
  NANDN U17124 ( .A(n16753), .B(n16752), .Z(n16754) );
  NAND U17125 ( .A(n16755), .B(n16754), .Z(n16863) );
  XOR U17126 ( .A(n16862), .B(n16863), .Z(n16921) );
  OR U17127 ( .A(n16757), .B(n16756), .Z(n16761) );
  OR U17128 ( .A(n16759), .B(n16758), .Z(n16760) );
  NAND U17129 ( .A(n16761), .B(n16760), .Z(n16810) );
  OR U17130 ( .A(n16763), .B(n16762), .Z(n16767) );
  NANDN U17131 ( .A(n16765), .B(n16764), .Z(n16766) );
  NAND U17132 ( .A(n16767), .B(n16766), .Z(n16808) );
  OR U17133 ( .A(n16769), .B(n16768), .Z(n16773) );
  NAND U17134 ( .A(n16771), .B(n16770), .Z(n16772) );
  NAND U17135 ( .A(n16773), .B(n16772), .Z(n16807) );
  XNOR U17136 ( .A(n16810), .B(n16809), .Z(n16920) );
  XNOR U17137 ( .A(n16921), .B(n16920), .Z(n16923) );
  NANDN U17138 ( .A(n16775), .B(n16774), .Z(n16779) );
  NANDN U17139 ( .A(n16777), .B(n16776), .Z(n16778) );
  AND U17140 ( .A(n16779), .B(n16778), .Z(n16922) );
  XNOR U17141 ( .A(n16923), .B(n16922), .Z(n16926) );
  XOR U17142 ( .A(n16927), .B(n16926), .Z(n16928) );
  XOR U17143 ( .A(n16929), .B(n16928), .Z(n16804) );
  NANDN U17144 ( .A(n16781), .B(n16780), .Z(n16785) );
  NAND U17145 ( .A(n16783), .B(n16782), .Z(n16784) );
  NAND U17146 ( .A(n16785), .B(n16784), .Z(n16801) );
  XNOR U17147 ( .A(n16801), .B(n16802), .Z(n16803) );
  XOR U17148 ( .A(n16804), .B(n16803), .Z(n16935) );
  XNOR U17149 ( .A(n16934), .B(n16935), .Z(n16796) );
  XNOR U17150 ( .A(n16795), .B(n16796), .Z(n16797) );
  XNOR U17151 ( .A(n16798), .B(n16797), .Z(n16938) );
  XNOR U17152 ( .A(n16938), .B(sreg[223]), .Z(n16940) );
  NAND U17153 ( .A(n16790), .B(sreg[222]), .Z(n16794) );
  OR U17154 ( .A(n16792), .B(n16791), .Z(n16793) );
  AND U17155 ( .A(n16794), .B(n16793), .Z(n16939) );
  XOR U17156 ( .A(n16940), .B(n16939), .Z(c[223]) );
  NANDN U17157 ( .A(n16796), .B(n16795), .Z(n16800) );
  NAND U17158 ( .A(n16798), .B(n16797), .Z(n16799) );
  NAND U17159 ( .A(n16800), .B(n16799), .Z(n16948) );
  NANDN U17160 ( .A(n16802), .B(n16801), .Z(n16806) );
  NANDN U17161 ( .A(n16804), .B(n16803), .Z(n16805) );
  NAND U17162 ( .A(n16806), .B(n16805), .Z(n17084) );
  OR U17163 ( .A(n16808), .B(n16807), .Z(n16812) );
  NANDN U17164 ( .A(n16810), .B(n16809), .Z(n16811) );
  AND U17165 ( .A(n16812), .B(n16811), .Z(n17075) );
  NANDN U17166 ( .A(n16814), .B(n16813), .Z(n16818) );
  NANDN U17167 ( .A(n16816), .B(n16815), .Z(n16817) );
  NAND U17168 ( .A(n16818), .B(n16817), .Z(n16960) );
  NANDN U17169 ( .A(n16820), .B(n16819), .Z(n16824) );
  NANDN U17170 ( .A(n16822), .B(n16821), .Z(n16823) );
  NAND U17171 ( .A(n16824), .B(n16823), .Z(n17057) );
  NANDN U17172 ( .A(n16826), .B(n16825), .Z(n16830) );
  NAND U17173 ( .A(n16828), .B(n16827), .Z(n16829) );
  NAND U17174 ( .A(n16830), .B(n16829), .Z(n17058) );
  XNOR U17175 ( .A(n17057), .B(n17058), .Z(n17059) );
  XNOR U17176 ( .A(b[23]), .B(a[106]), .Z(n17029) );
  OR U17177 ( .A(n17029), .B(n19127), .Z(n16833) );
  NAND U17178 ( .A(n16831), .B(n19128), .Z(n16832) );
  NAND U17179 ( .A(n16833), .B(n16832), .Z(n17054) );
  NANDN U17180 ( .A(n16834), .B(n17553), .Z(n16836) );
  XNOR U17181 ( .A(a[122]), .B(b[7]), .Z(n17020) );
  NANDN U17182 ( .A(n17020), .B(n17555), .Z(n16835) );
  NAND U17183 ( .A(n16836), .B(n16835), .Z(n17051) );
  XNOR U17184 ( .A(b[25]), .B(a[104]), .Z(n16985) );
  NANDN U17185 ( .A(n16985), .B(n19240), .Z(n16839) );
  NAND U17186 ( .A(n16837), .B(n19242), .Z(n16838) );
  AND U17187 ( .A(n16839), .B(n16838), .Z(n17052) );
  XNOR U17188 ( .A(n17051), .B(n17052), .Z(n17053) );
  XNOR U17189 ( .A(n17054), .B(n17053), .Z(n16967) );
  NANDN U17190 ( .A(n577), .B(b[1]), .Z(n16841) );
  IV U17191 ( .A(a[127]), .Z(n19502) );
  NANDN U17192 ( .A(n17151), .B(n19502), .Z(n16840) );
  NAND U17193 ( .A(n16841), .B(n16840), .Z(n16976) );
  NAND U17194 ( .A(n19406), .B(n16842), .Z(n16844) );
  XOR U17195 ( .A(b[29]), .B(n17447), .Z(n17039) );
  OR U17196 ( .A(n17039), .B(n576), .Z(n16843) );
  NAND U17197 ( .A(n16844), .B(n16843), .Z(n16973) );
  NANDN U17198 ( .A(n585), .B(a[96]), .Z(n16974) );
  XNOR U17199 ( .A(n16973), .B(n16974), .Z(n16975) );
  XOR U17200 ( .A(n16976), .B(n16975), .Z(n16968) );
  XOR U17201 ( .A(n16967), .B(n16968), .Z(n16970) );
  NAND U17202 ( .A(n16845), .B(n18513), .Z(n16847) );
  XNOR U17203 ( .A(a[114]), .B(b[15]), .Z(n16982) );
  OR U17204 ( .A(n16982), .B(n18512), .Z(n16846) );
  NAND U17205 ( .A(n16847), .B(n16846), .Z(n17011) );
  NANDN U17206 ( .A(n16848), .B(n19013), .Z(n16850) );
  XOR U17207 ( .A(b[21]), .B(n18198), .Z(n17032) );
  NANDN U17208 ( .A(n17032), .B(n19015), .Z(n16849) );
  NAND U17209 ( .A(n16850), .B(n16849), .Z(n17008) );
  XOR U17210 ( .A(a[120]), .B(n579), .Z(n17014) );
  NANDN U17211 ( .A(n17014), .B(n17814), .Z(n16853) );
  NANDN U17212 ( .A(n16851), .B(n17815), .Z(n16852) );
  AND U17213 ( .A(n16853), .B(n16852), .Z(n17009) );
  XNOR U17214 ( .A(n17008), .B(n17009), .Z(n17010) );
  XNOR U17215 ( .A(n17011), .B(n17010), .Z(n16999) );
  XOR U17216 ( .A(a[116]), .B(n580), .Z(n17023) );
  NANDN U17217 ( .A(n17023), .B(n18336), .Z(n16856) );
  NANDN U17218 ( .A(n16854), .B(n18337), .Z(n16855) );
  NAND U17219 ( .A(n16856), .B(n16855), .Z(n16997) );
  XNOR U17220 ( .A(a[118]), .B(b[11]), .Z(n17017) );
  OR U17221 ( .A(n17017), .B(n18194), .Z(n16859) );
  NANDN U17222 ( .A(n16857), .B(n18104), .Z(n16858) );
  AND U17223 ( .A(n16859), .B(n16858), .Z(n16996) );
  XNOR U17224 ( .A(n16997), .B(n16996), .Z(n16998) );
  XOR U17225 ( .A(n16999), .B(n16998), .Z(n16969) );
  XNOR U17226 ( .A(n16970), .B(n16969), .Z(n17060) );
  XNOR U17227 ( .A(n17059), .B(n17060), .Z(n16957) );
  NANDN U17228 ( .A(n16861), .B(n16860), .Z(n16865) );
  NANDN U17229 ( .A(n16863), .B(n16862), .Z(n16864) );
  AND U17230 ( .A(n16865), .B(n16864), .Z(n16958) );
  XNOR U17231 ( .A(n16957), .B(n16958), .Z(n16959) );
  XOR U17232 ( .A(n16960), .B(n16959), .Z(n17076) );
  OR U17233 ( .A(n16867), .B(n16866), .Z(n16871) );
  NANDN U17234 ( .A(n16869), .B(n16868), .Z(n16870) );
  NAND U17235 ( .A(n16871), .B(n16870), .Z(n16952) );
  NANDN U17236 ( .A(n16873), .B(n16872), .Z(n16877) );
  NAND U17237 ( .A(n16875), .B(n16874), .Z(n16876) );
  NAND U17238 ( .A(n16877), .B(n16876), .Z(n17065) );
  XNOR U17239 ( .A(b[17]), .B(a[112]), .Z(n16993) );
  NANDN U17240 ( .A(n16993), .B(n18673), .Z(n16880) );
  NAND U17241 ( .A(n16878), .B(n18674), .Z(n16879) );
  NAND U17242 ( .A(n16880), .B(n16879), .Z(n17005) );
  XNOR U17243 ( .A(n585), .B(a[98]), .Z(n17042) );
  NAND U17244 ( .A(n17042), .B(n19472), .Z(n16883) );
  NANDN U17245 ( .A(n16881), .B(n19473), .Z(n16882) );
  NAND U17246 ( .A(n16883), .B(n16882), .Z(n17002) );
  OR U17247 ( .A(n16884), .B(n16988), .Z(n16886) );
  XOR U17248 ( .A(a[126]), .B(n578), .Z(n16989) );
  NANDN U17249 ( .A(n16989), .B(n16990), .Z(n16885) );
  AND U17250 ( .A(n16886), .B(n16885), .Z(n17003) );
  XNOR U17251 ( .A(n17002), .B(n17003), .Z(n17004) );
  XNOR U17252 ( .A(n17005), .B(n17004), .Z(n17063) );
  NANDN U17253 ( .A(n16887), .B(n18832), .Z(n16889) );
  XOR U17254 ( .A(b[19]), .B(n18415), .Z(n17026) );
  NANDN U17255 ( .A(n17026), .B(n18834), .Z(n16888) );
  NAND U17256 ( .A(n16889), .B(n16888), .Z(n17048) );
  XOR U17257 ( .A(b[27]), .B(n17208), .Z(n16979) );
  NANDN U17258 ( .A(n16979), .B(n19336), .Z(n16892) );
  NANDN U17259 ( .A(n16890), .B(n19337), .Z(n16891) );
  NAND U17260 ( .A(n16892), .B(n16891), .Z(n17045) );
  XNOR U17261 ( .A(a[124]), .B(b[5]), .Z(n17035) );
  NANDN U17262 ( .A(n17035), .B(n17310), .Z(n16895) );
  NAND U17263 ( .A(n16893), .B(n17311), .Z(n16894) );
  AND U17264 ( .A(n16895), .B(n16894), .Z(n17046) );
  XNOR U17265 ( .A(n17045), .B(n17046), .Z(n17047) );
  XOR U17266 ( .A(n17048), .B(n17047), .Z(n17064) );
  XOR U17267 ( .A(n17063), .B(n17064), .Z(n17066) );
  XOR U17268 ( .A(n17065), .B(n17066), .Z(n16951) );
  XNOR U17269 ( .A(n16952), .B(n16951), .Z(n16953) );
  NANDN U17270 ( .A(n16897), .B(n16896), .Z(n16901) );
  NAND U17271 ( .A(n16899), .B(n16898), .Z(n16900) );
  NAND U17272 ( .A(n16901), .B(n16900), .Z(n16964) );
  NANDN U17273 ( .A(n16903), .B(n16902), .Z(n16907) );
  NAND U17274 ( .A(n16905), .B(n16904), .Z(n16906) );
  NAND U17275 ( .A(n16907), .B(n16906), .Z(n16961) );
  OR U17276 ( .A(n16909), .B(n16908), .Z(n16913) );
  NANDN U17277 ( .A(n16911), .B(n16910), .Z(n16912) );
  NAND U17278 ( .A(n16913), .B(n16912), .Z(n16962) );
  XNOR U17279 ( .A(n16961), .B(n16962), .Z(n16963) );
  XOR U17280 ( .A(n16964), .B(n16963), .Z(n16954) );
  XOR U17281 ( .A(n16953), .B(n16954), .Z(n17077) );
  XOR U17282 ( .A(n17078), .B(n17077), .Z(n17072) );
  OR U17283 ( .A(n16915), .B(n16914), .Z(n16919) );
  NAND U17284 ( .A(n16917), .B(n16916), .Z(n16918) );
  NAND U17285 ( .A(n16919), .B(n16918), .Z(n17069) );
  NAND U17286 ( .A(n16921), .B(n16920), .Z(n16925) );
  NANDN U17287 ( .A(n16923), .B(n16922), .Z(n16924) );
  NAND U17288 ( .A(n16925), .B(n16924), .Z(n17070) );
  XNOR U17289 ( .A(n17069), .B(n17070), .Z(n17071) );
  XNOR U17290 ( .A(n17072), .B(n17071), .Z(n17082) );
  NAND U17291 ( .A(n16927), .B(n16926), .Z(n16931) );
  NAND U17292 ( .A(n16929), .B(n16928), .Z(n16930) );
  AND U17293 ( .A(n16931), .B(n16930), .Z(n17081) );
  XNOR U17294 ( .A(n17082), .B(n17081), .Z(n17083) );
  XNOR U17295 ( .A(n17084), .B(n17083), .Z(n16945) );
  NANDN U17296 ( .A(n16933), .B(n16932), .Z(n16937) );
  NANDN U17297 ( .A(n16935), .B(n16934), .Z(n16936) );
  NAND U17298 ( .A(n16937), .B(n16936), .Z(n16946) );
  XNOR U17299 ( .A(n16945), .B(n16946), .Z(n16947) );
  XOR U17300 ( .A(n16948), .B(n16947), .Z(n16944) );
  NAND U17301 ( .A(n16938), .B(sreg[223]), .Z(n16942) );
  OR U17302 ( .A(n16940), .B(n16939), .Z(n16941) );
  AND U17303 ( .A(n16942), .B(n16941), .Z(n16943) );
  XOR U17304 ( .A(n16944), .B(n16943), .Z(c[224]) );
  OR U17305 ( .A(n16944), .B(n16943), .Z(n17227) );
  NANDN U17306 ( .A(n16946), .B(n16945), .Z(n16950) );
  NAND U17307 ( .A(n16948), .B(n16947), .Z(n16949) );
  NAND U17308 ( .A(n16950), .B(n16949), .Z(n17090) );
  NAND U17309 ( .A(n16952), .B(n16951), .Z(n16956) );
  OR U17310 ( .A(n16954), .B(n16953), .Z(n16955) );
  NAND U17311 ( .A(n16956), .B(n16955), .Z(n17097) );
  XNOR U17312 ( .A(n17097), .B(n17098), .Z(n17099) );
  NANDN U17313 ( .A(n16962), .B(n16961), .Z(n16966) );
  NANDN U17314 ( .A(n16964), .B(n16963), .Z(n16965) );
  NAND U17315 ( .A(n16966), .B(n16965), .Z(n17220) );
  NANDN U17316 ( .A(n16968), .B(n16967), .Z(n16972) );
  NANDN U17317 ( .A(n16970), .B(n16969), .Z(n16971) );
  NAND U17318 ( .A(n16972), .B(n16971), .Z(n17175) );
  NANDN U17319 ( .A(n16974), .B(n16973), .Z(n16978) );
  NAND U17320 ( .A(n16976), .B(n16975), .Z(n16977) );
  NAND U17321 ( .A(n16978), .B(n16977), .Z(n17170) );
  XNOR U17322 ( .A(b[27]), .B(a[103]), .Z(n17145) );
  NANDN U17323 ( .A(n17145), .B(n19336), .Z(n16981) );
  NANDN U17324 ( .A(n16979), .B(n19337), .Z(n16980) );
  NAND U17325 ( .A(n16981), .B(n16980), .Z(n17141) );
  NANDN U17326 ( .A(n16982), .B(n18513), .Z(n16984) );
  XNOR U17327 ( .A(a[115]), .B(b[15]), .Z(n17204) );
  OR U17328 ( .A(n17204), .B(n18512), .Z(n16983) );
  AND U17329 ( .A(n16984), .B(n16983), .Z(n17139) );
  XOR U17330 ( .A(b[1]), .B(n17139), .Z(n17140) );
  XNOR U17331 ( .A(n17141), .B(n17140), .Z(n17168) );
  XOR U17332 ( .A(b[25]), .B(a[105]), .Z(n17136) );
  NAND U17333 ( .A(n17136), .B(n19240), .Z(n16987) );
  NANDN U17334 ( .A(n16985), .B(n19242), .Z(n16986) );
  NAND U17335 ( .A(n16987), .B(n16986), .Z(n17112) );
  OR U17336 ( .A(n16989), .B(n16988), .Z(n16992) );
  XNOR U17337 ( .A(n19502), .B(b[3]), .Z(n17153) );
  NAND U17338 ( .A(n17153), .B(n16990), .Z(n16991) );
  NAND U17339 ( .A(n16992), .B(n16991), .Z(n17109) );
  XOR U17340 ( .A(b[17]), .B(a[113]), .Z(n17148) );
  NAND U17341 ( .A(n17148), .B(n18673), .Z(n16995) );
  NANDN U17342 ( .A(n16993), .B(n18674), .Z(n16994) );
  AND U17343 ( .A(n16995), .B(n16994), .Z(n17110) );
  XNOR U17344 ( .A(n17109), .B(n17110), .Z(n17111) );
  XOR U17345 ( .A(n17112), .B(n17111), .Z(n17169) );
  XOR U17346 ( .A(n17168), .B(n17169), .Z(n17171) );
  XOR U17347 ( .A(n17170), .B(n17171), .Z(n17174) );
  XNOR U17348 ( .A(n17175), .B(n17174), .Z(n17177) );
  NANDN U17349 ( .A(n16997), .B(n16996), .Z(n17001) );
  NAND U17350 ( .A(n16999), .B(n16998), .Z(n17000) );
  NAND U17351 ( .A(n17001), .B(n17000), .Z(n17195) );
  NANDN U17352 ( .A(n17003), .B(n17002), .Z(n17007) );
  NAND U17353 ( .A(n17005), .B(n17004), .Z(n17006) );
  NAND U17354 ( .A(n17007), .B(n17006), .Z(n17193) );
  NANDN U17355 ( .A(n17009), .B(n17008), .Z(n17013) );
  NAND U17356 ( .A(n17011), .B(n17010), .Z(n17012) );
  AND U17357 ( .A(n17013), .B(n17012), .Z(n17192) );
  XNOR U17358 ( .A(n17193), .B(n17192), .Z(n17194) );
  XOR U17359 ( .A(n17195), .B(n17194), .Z(n17176) );
  XNOR U17360 ( .A(n17177), .B(n17176), .Z(n17219) );
  XNOR U17361 ( .A(n17220), .B(n17219), .Z(n17221) );
  XOR U17362 ( .A(a[121]), .B(n579), .Z(n17121) );
  NANDN U17363 ( .A(n17121), .B(n17814), .Z(n17016) );
  NANDN U17364 ( .A(n17014), .B(n17815), .Z(n17015) );
  NAND U17365 ( .A(n17016), .B(n17015), .Z(n17106) );
  XNOR U17366 ( .A(a[119]), .B(b[11]), .Z(n17133) );
  OR U17367 ( .A(n17133), .B(n18194), .Z(n17019) );
  NANDN U17368 ( .A(n17017), .B(n18104), .Z(n17018) );
  NAND U17369 ( .A(n17019), .B(n17018), .Z(n17103) );
  NANDN U17370 ( .A(n17020), .B(n17553), .Z(n17022) );
  XOR U17371 ( .A(a[123]), .B(b[7]), .Z(n17124) );
  NAND U17372 ( .A(n17124), .B(n17555), .Z(n17021) );
  NAND U17373 ( .A(n17022), .B(n17021), .Z(n17118) );
  XOR U17374 ( .A(a[117]), .B(n580), .Z(n17130) );
  NANDN U17375 ( .A(n17130), .B(n18336), .Z(n17025) );
  NANDN U17376 ( .A(n17023), .B(n18337), .Z(n17024) );
  NAND U17377 ( .A(n17025), .B(n17024), .Z(n17115) );
  NANDN U17378 ( .A(n17026), .B(n18832), .Z(n17028) );
  XNOR U17379 ( .A(n581), .B(a[111]), .Z(n17156) );
  NAND U17380 ( .A(n17156), .B(n18834), .Z(n17027) );
  AND U17381 ( .A(n17028), .B(n17027), .Z(n17116) );
  XNOR U17382 ( .A(n17115), .B(n17116), .Z(n17117) );
  XNOR U17383 ( .A(n17118), .B(n17117), .Z(n17104) );
  XNOR U17384 ( .A(n17103), .B(n17104), .Z(n17105) );
  XOR U17385 ( .A(n17106), .B(n17105), .Z(n17165) );
  XOR U17386 ( .A(b[23]), .B(a[107]), .Z(n17142) );
  NANDN U17387 ( .A(n19127), .B(n17142), .Z(n17031) );
  NANDN U17388 ( .A(n17029), .B(n19128), .Z(n17030) );
  NAND U17389 ( .A(n17031), .B(n17030), .Z(n17201) );
  NANDN U17390 ( .A(n17032), .B(n19013), .Z(n17034) );
  XNOR U17391 ( .A(b[21]), .B(a[109]), .Z(n17127) );
  NANDN U17392 ( .A(n17127), .B(n19015), .Z(n17033) );
  NAND U17393 ( .A(n17034), .B(n17033), .Z(n17198) );
  XNOR U17394 ( .A(n19402), .B(b[5]), .Z(n17159) );
  NAND U17395 ( .A(n17159), .B(n17310), .Z(n17037) );
  NANDN U17396 ( .A(n17035), .B(n17311), .Z(n17036) );
  AND U17397 ( .A(n17037), .B(n17036), .Z(n17199) );
  XNOR U17398 ( .A(n17198), .B(n17199), .Z(n17200) );
  XOR U17399 ( .A(n17201), .B(n17200), .Z(n17163) );
  ANDN U17400 ( .B(b[31]), .A(n17038), .Z(n17269) );
  IV U17401 ( .A(n17269), .Z(n17406) );
  NANDN U17402 ( .A(n17039), .B(n19406), .Z(n17041) );
  XNOR U17403 ( .A(n584), .B(a[101]), .Z(n17207) );
  NANDN U17404 ( .A(n576), .B(n17207), .Z(n17040) );
  AND U17405 ( .A(n17041), .B(n17040), .Z(n17214) );
  XOR U17406 ( .A(n17406), .B(n17214), .Z(n17216) );
  XNOR U17407 ( .A(b[31]), .B(a[99]), .Z(n17211) );
  NANDN U17408 ( .A(n17211), .B(n19472), .Z(n17044) );
  NAND U17409 ( .A(n19473), .B(n17042), .Z(n17043) );
  NAND U17410 ( .A(n17044), .B(n17043), .Z(n17215) );
  XOR U17411 ( .A(n17216), .B(n17215), .Z(n17162) );
  XOR U17412 ( .A(n17163), .B(n17162), .Z(n17164) );
  XOR U17413 ( .A(n17165), .B(n17164), .Z(n17189) );
  NANDN U17414 ( .A(n17046), .B(n17045), .Z(n17050) );
  NAND U17415 ( .A(n17048), .B(n17047), .Z(n17049) );
  NAND U17416 ( .A(n17050), .B(n17049), .Z(n17186) );
  NANDN U17417 ( .A(n17052), .B(n17051), .Z(n17056) );
  NAND U17418 ( .A(n17054), .B(n17053), .Z(n17055) );
  AND U17419 ( .A(n17056), .B(n17055), .Z(n17187) );
  XNOR U17420 ( .A(n17186), .B(n17187), .Z(n17188) );
  XNOR U17421 ( .A(n17189), .B(n17188), .Z(n17183) );
  NANDN U17422 ( .A(n17058), .B(n17057), .Z(n17062) );
  NAND U17423 ( .A(n17060), .B(n17059), .Z(n17061) );
  NAND U17424 ( .A(n17062), .B(n17061), .Z(n17180) );
  NANDN U17425 ( .A(n17064), .B(n17063), .Z(n17068) );
  OR U17426 ( .A(n17066), .B(n17065), .Z(n17067) );
  AND U17427 ( .A(n17068), .B(n17067), .Z(n17181) );
  XNOR U17428 ( .A(n17180), .B(n17181), .Z(n17182) );
  XOR U17429 ( .A(n17183), .B(n17182), .Z(n17222) );
  XOR U17430 ( .A(n17221), .B(n17222), .Z(n17100) );
  XNOR U17431 ( .A(n17099), .B(n17100), .Z(n17095) );
  NANDN U17432 ( .A(n17070), .B(n17069), .Z(n17074) );
  NAND U17433 ( .A(n17072), .B(n17071), .Z(n17073) );
  NAND U17434 ( .A(n17074), .B(n17073), .Z(n17093) );
  OR U17435 ( .A(n17076), .B(n17075), .Z(n17080) );
  NANDN U17436 ( .A(n17078), .B(n17077), .Z(n17079) );
  NAND U17437 ( .A(n17080), .B(n17079), .Z(n17094) );
  XNOR U17438 ( .A(n17093), .B(n17094), .Z(n17096) );
  XNOR U17439 ( .A(n17095), .B(n17096), .Z(n17087) );
  NANDN U17440 ( .A(n17082), .B(n17081), .Z(n17086) );
  NAND U17441 ( .A(n17084), .B(n17083), .Z(n17085) );
  NAND U17442 ( .A(n17086), .B(n17085), .Z(n17088) );
  XNOR U17443 ( .A(n17087), .B(n17088), .Z(n17089) );
  XOR U17444 ( .A(n17090), .B(n17089), .Z(n17226) );
  XOR U17445 ( .A(n17227), .B(n17226), .Z(c[225]) );
  NANDN U17446 ( .A(n17088), .B(n17087), .Z(n17092) );
  NAND U17447 ( .A(n17090), .B(n17089), .Z(n17091) );
  AND U17448 ( .A(n17092), .B(n17091), .Z(n17232) );
  NANDN U17449 ( .A(n17098), .B(n17097), .Z(n17102) );
  NAND U17450 ( .A(n17100), .B(n17099), .Z(n17101) );
  NAND U17451 ( .A(n17102), .B(n17101), .Z(n17360) );
  NANDN U17452 ( .A(n17104), .B(n17103), .Z(n17108) );
  NAND U17453 ( .A(n17106), .B(n17105), .Z(n17107) );
  NAND U17454 ( .A(n17108), .B(n17107), .Z(n17344) );
  NANDN U17455 ( .A(n17110), .B(n17109), .Z(n17114) );
  NAND U17456 ( .A(n17112), .B(n17111), .Z(n17113) );
  NAND U17457 ( .A(n17114), .B(n17113), .Z(n17343) );
  NANDN U17458 ( .A(n17116), .B(n17115), .Z(n17120) );
  NAND U17459 ( .A(n17118), .B(n17117), .Z(n17119) );
  NAND U17460 ( .A(n17120), .B(n17119), .Z(n17253) );
  XOR U17461 ( .A(a[122]), .B(n579), .Z(n17306) );
  NANDN U17462 ( .A(n17306), .B(n17814), .Z(n17123) );
  NANDN U17463 ( .A(n17121), .B(n17815), .Z(n17122) );
  NAND U17464 ( .A(n17123), .B(n17122), .Z(n17287) );
  NAND U17465 ( .A(n17124), .B(n17553), .Z(n17126) );
  XNOR U17466 ( .A(a[124]), .B(b[7]), .Z(n17333) );
  NANDN U17467 ( .A(n17333), .B(n17555), .Z(n17125) );
  NAND U17468 ( .A(n17126), .B(n17125), .Z(n17284) );
  NANDN U17469 ( .A(n17127), .B(n19013), .Z(n17129) );
  XOR U17470 ( .A(b[21]), .B(n18415), .Z(n17339) );
  NANDN U17471 ( .A(n17339), .B(n19015), .Z(n17128) );
  AND U17472 ( .A(n17129), .B(n17128), .Z(n17285) );
  XNOR U17473 ( .A(n17284), .B(n17285), .Z(n17286) );
  XNOR U17474 ( .A(n17287), .B(n17286), .Z(n17251) );
  XOR U17475 ( .A(a[118]), .B(n580), .Z(n17257) );
  NANDN U17476 ( .A(n17257), .B(n18336), .Z(n17132) );
  NANDN U17477 ( .A(n17130), .B(n18337), .Z(n17131) );
  NAND U17478 ( .A(n17132), .B(n17131), .Z(n17297) );
  XNOR U17479 ( .A(a[120]), .B(b[11]), .Z(n17324) );
  OR U17480 ( .A(n17324), .B(n18194), .Z(n17135) );
  NANDN U17481 ( .A(n17133), .B(n18104), .Z(n17134) );
  NAND U17482 ( .A(n17135), .B(n17134), .Z(n17294) );
  XNOR U17483 ( .A(b[25]), .B(a[106]), .Z(n17327) );
  NANDN U17484 ( .A(n17327), .B(n19240), .Z(n17138) );
  NAND U17485 ( .A(n17136), .B(n19242), .Z(n17137) );
  AND U17486 ( .A(n17138), .B(n17137), .Z(n17295) );
  XNOR U17487 ( .A(n17294), .B(n17295), .Z(n17296) );
  XOR U17488 ( .A(n17297), .B(n17296), .Z(n17252) );
  XOR U17489 ( .A(n17251), .B(n17252), .Z(n17254) );
  XOR U17490 ( .A(n17253), .B(n17254), .Z(n17342) );
  XOR U17491 ( .A(n17343), .B(n17342), .Z(n17345) );
  XOR U17492 ( .A(n17344), .B(n17345), .Z(n17352) );
  XNOR U17493 ( .A(b[23]), .B(a[108]), .Z(n17300) );
  OR U17494 ( .A(n17300), .B(n19127), .Z(n17144) );
  NAND U17495 ( .A(n17142), .B(n19128), .Z(n17143) );
  NAND U17496 ( .A(n17144), .B(n17143), .Z(n17275) );
  XOR U17497 ( .A(b[27]), .B(n17716), .Z(n17330) );
  NANDN U17498 ( .A(n17330), .B(n19336), .Z(n17147) );
  NANDN U17499 ( .A(n17145), .B(n19337), .Z(n17146) );
  NAND U17500 ( .A(n17147), .B(n17146), .Z(n17272) );
  XNOR U17501 ( .A(b[17]), .B(a[114]), .Z(n17263) );
  NANDN U17502 ( .A(n17263), .B(n18673), .Z(n17150) );
  NAND U17503 ( .A(n17148), .B(n18674), .Z(n17149) );
  AND U17504 ( .A(n17150), .B(n17149), .Z(n17273) );
  XNOR U17505 ( .A(n17272), .B(n17273), .Z(n17274) );
  XNOR U17506 ( .A(n17275), .B(n17274), .Z(n17291) );
  NANDN U17507 ( .A(n17151), .B(b[2]), .Z(n17309) );
  XOR U17508 ( .A(n578), .B(n17309), .Z(n17155) );
  XOR U17509 ( .A(b[2]), .B(n17151), .Z(n17152) );
  NANDN U17510 ( .A(n17153), .B(n17152), .Z(n17154) );
  AND U17511 ( .A(n17155), .B(n17154), .Z(n17266) );
  NANDN U17512 ( .A(n585), .B(a[98]), .Z(n17267) );
  XNOR U17513 ( .A(n17266), .B(n17267), .Z(n17268) );
  XOR U17514 ( .A(n17406), .B(n17268), .Z(n17281) );
  XOR U17515 ( .A(n581), .B(a[112]), .Z(n17315) );
  NANDN U17516 ( .A(n17315), .B(n18834), .Z(n17158) );
  NAND U17517 ( .A(n18832), .B(n17156), .Z(n17157) );
  NAND U17518 ( .A(n17158), .B(n17157), .Z(n17279) );
  XOR U17519 ( .A(n19295), .B(b[5]), .Z(n17312) );
  NANDN U17520 ( .A(n17312), .B(n17310), .Z(n17161) );
  NAND U17521 ( .A(n17311), .B(n17159), .Z(n17160) );
  AND U17522 ( .A(n17161), .B(n17160), .Z(n17278) );
  XNOR U17523 ( .A(n17279), .B(n17278), .Z(n17280) );
  XNOR U17524 ( .A(n17281), .B(n17280), .Z(n17290) );
  XOR U17525 ( .A(n17291), .B(n17290), .Z(n17292) );
  XOR U17526 ( .A(n17293), .B(n17292), .Z(n17236) );
  NANDN U17527 ( .A(n17163), .B(n17162), .Z(n17167) );
  OR U17528 ( .A(n17165), .B(n17164), .Z(n17166) );
  NAND U17529 ( .A(n17167), .B(n17166), .Z(n17234) );
  NANDN U17530 ( .A(n17169), .B(n17168), .Z(n17173) );
  OR U17531 ( .A(n17171), .B(n17170), .Z(n17172) );
  AND U17532 ( .A(n17173), .B(n17172), .Z(n17233) );
  XNOR U17533 ( .A(n17234), .B(n17233), .Z(n17235) );
  XNOR U17534 ( .A(n17236), .B(n17235), .Z(n17353) );
  NAND U17535 ( .A(n17175), .B(n17174), .Z(n17179) );
  NANDN U17536 ( .A(n17177), .B(n17176), .Z(n17178) );
  NAND U17537 ( .A(n17179), .B(n17178), .Z(n17355) );
  XOR U17538 ( .A(n17354), .B(n17355), .Z(n17351) );
  NANDN U17539 ( .A(n17181), .B(n17180), .Z(n17185) );
  NANDN U17540 ( .A(n17183), .B(n17182), .Z(n17184) );
  NAND U17541 ( .A(n17185), .B(n17184), .Z(n17349) );
  NANDN U17542 ( .A(n17187), .B(n17186), .Z(n17191) );
  NANDN U17543 ( .A(n17189), .B(n17188), .Z(n17190) );
  NAND U17544 ( .A(n17191), .B(n17190), .Z(n17242) );
  NANDN U17545 ( .A(n17193), .B(n17192), .Z(n17197) );
  NAND U17546 ( .A(n17195), .B(n17194), .Z(n17196) );
  NAND U17547 ( .A(n17197), .B(n17196), .Z(n17240) );
  NANDN U17548 ( .A(n17199), .B(n17198), .Z(n17203) );
  NAND U17549 ( .A(n17201), .B(n17200), .Z(n17202) );
  NAND U17550 ( .A(n17203), .B(n17202), .Z(n17247) );
  NANDN U17551 ( .A(n17204), .B(n18513), .Z(n17206) );
  XNOR U17552 ( .A(a[116]), .B(b[15]), .Z(n17260) );
  OR U17553 ( .A(n17260), .B(n18512), .Z(n17205) );
  NAND U17554 ( .A(n17206), .B(n17205), .Z(n17321) );
  NAND U17555 ( .A(n17207), .B(n19406), .Z(n17210) );
  XOR U17556 ( .A(n584), .B(n17208), .Z(n17303) );
  NANDN U17557 ( .A(n576), .B(n17303), .Z(n17209) );
  NAND U17558 ( .A(n17210), .B(n17209), .Z(n17318) );
  XOR U17559 ( .A(b[31]), .B(n17447), .Z(n17336) );
  NANDN U17560 ( .A(n17336), .B(n19472), .Z(n17213) );
  NANDN U17561 ( .A(n17211), .B(n19473), .Z(n17212) );
  AND U17562 ( .A(n17213), .B(n17212), .Z(n17319) );
  XNOR U17563 ( .A(n17318), .B(n17319), .Z(n17320) );
  XNOR U17564 ( .A(n17321), .B(n17320), .Z(n17245) );
  NANDN U17565 ( .A(n17406), .B(n17214), .Z(n17218) );
  OR U17566 ( .A(n17216), .B(n17215), .Z(n17217) );
  AND U17567 ( .A(n17218), .B(n17217), .Z(n17246) );
  XOR U17568 ( .A(n17245), .B(n17246), .Z(n17248) );
  XOR U17569 ( .A(n17247), .B(n17248), .Z(n17239) );
  XOR U17570 ( .A(n17240), .B(n17239), .Z(n17241) );
  XNOR U17571 ( .A(n17242), .B(n17241), .Z(n17348) );
  XOR U17572 ( .A(n17349), .B(n17348), .Z(n17350) );
  XNOR U17573 ( .A(n17351), .B(n17350), .Z(n17358) );
  NAND U17574 ( .A(n17220), .B(n17219), .Z(n17224) );
  OR U17575 ( .A(n17222), .B(n17221), .Z(n17223) );
  NAND U17576 ( .A(n17224), .B(n17223), .Z(n17359) );
  XOR U17577 ( .A(n17358), .B(n17359), .Z(n17361) );
  XOR U17578 ( .A(n17360), .B(n17361), .Z(n17230) );
  XNOR U17579 ( .A(n17231), .B(n17230), .Z(n17225) );
  XOR U17580 ( .A(n17232), .B(n17225), .Z(n17228) );
  OR U17581 ( .A(n17227), .B(n17226), .Z(n17229) );
  XNOR U17582 ( .A(n17228), .B(n17229), .Z(c[226]) );
  NANDN U17583 ( .A(n17229), .B(n17228), .Z(n17365) );
  NANDN U17584 ( .A(n17234), .B(n17233), .Z(n17238) );
  NAND U17585 ( .A(n17236), .B(n17235), .Z(n17237) );
  NAND U17586 ( .A(n17238), .B(n17237), .Z(n17378) );
  NAND U17587 ( .A(n17240), .B(n17239), .Z(n17244) );
  NANDN U17588 ( .A(n17242), .B(n17241), .Z(n17243) );
  NAND U17589 ( .A(n17244), .B(n17243), .Z(n17379) );
  XNOR U17590 ( .A(n17378), .B(n17379), .Z(n17380) );
  NANDN U17591 ( .A(n17246), .B(n17245), .Z(n17250) );
  OR U17592 ( .A(n17248), .B(n17247), .Z(n17249) );
  NAND U17593 ( .A(n17250), .B(n17249), .Z(n17484) );
  NANDN U17594 ( .A(n17252), .B(n17251), .Z(n17256) );
  OR U17595 ( .A(n17254), .B(n17253), .Z(n17255) );
  NAND U17596 ( .A(n17256), .B(n17255), .Z(n17482) );
  XOR U17597 ( .A(a[119]), .B(n580), .Z(n17418) );
  NANDN U17598 ( .A(n17418), .B(n18336), .Z(n17259) );
  NANDN U17599 ( .A(n17257), .B(n18337), .Z(n17258) );
  NAND U17600 ( .A(n17259), .B(n17258), .Z(n17424) );
  NANDN U17601 ( .A(n17260), .B(n18513), .Z(n17262) );
  XNOR U17602 ( .A(a[117]), .B(b[15]), .Z(n17412) );
  OR U17603 ( .A(n17412), .B(n18512), .Z(n17261) );
  NAND U17604 ( .A(n17262), .B(n17261), .Z(n17421) );
  XNOR U17605 ( .A(b[17]), .B(a[115]), .Z(n17415) );
  NANDN U17606 ( .A(n17415), .B(n18673), .Z(n17265) );
  NANDN U17607 ( .A(n17263), .B(n18674), .Z(n17264) );
  AND U17608 ( .A(n17265), .B(n17264), .Z(n17422) );
  XNOR U17609 ( .A(n17421), .B(n17422), .Z(n17423) );
  XNOR U17610 ( .A(n17424), .B(n17423), .Z(n17478) );
  NANDN U17611 ( .A(n17267), .B(n17266), .Z(n17271) );
  NANDN U17612 ( .A(n17269), .B(n17268), .Z(n17270) );
  NAND U17613 ( .A(n17271), .B(n17270), .Z(n17476) );
  NANDN U17614 ( .A(n17273), .B(n17272), .Z(n17277) );
  NAND U17615 ( .A(n17275), .B(n17274), .Z(n17276) );
  AND U17616 ( .A(n17277), .B(n17276), .Z(n17475) );
  XNOR U17617 ( .A(n17476), .B(n17475), .Z(n17477) );
  XOR U17618 ( .A(n17478), .B(n17477), .Z(n17489) );
  NANDN U17619 ( .A(n17279), .B(n17278), .Z(n17283) );
  NANDN U17620 ( .A(n17281), .B(n17280), .Z(n17282) );
  NAND U17621 ( .A(n17283), .B(n17282), .Z(n17487) );
  NANDN U17622 ( .A(n17285), .B(n17284), .Z(n17289) );
  NAND U17623 ( .A(n17287), .B(n17286), .Z(n17288) );
  NAND U17624 ( .A(n17289), .B(n17288), .Z(n17488) );
  XNOR U17625 ( .A(n17487), .B(n17488), .Z(n17490) );
  XOR U17626 ( .A(n17489), .B(n17490), .Z(n17481) );
  XOR U17627 ( .A(n17482), .B(n17481), .Z(n17483) );
  XNOR U17628 ( .A(n17484), .B(n17483), .Z(n17387) );
  NANDN U17629 ( .A(n17295), .B(n17294), .Z(n17299) );
  NAND U17630 ( .A(n17297), .B(n17296), .Z(n17298) );
  NAND U17631 ( .A(n17299), .B(n17298), .Z(n17501) );
  XOR U17632 ( .A(b[23]), .B(a[109]), .Z(n17457) );
  NANDN U17633 ( .A(n19127), .B(n17457), .Z(n17302) );
  NANDN U17634 ( .A(n17300), .B(n19128), .Z(n17301) );
  NAND U17635 ( .A(n17302), .B(n17301), .Z(n17430) );
  NAND U17636 ( .A(n19406), .B(n17303), .Z(n17305) );
  XNOR U17637 ( .A(n584), .B(a[103]), .Z(n17469) );
  NANDN U17638 ( .A(n576), .B(n17469), .Z(n17304) );
  NAND U17639 ( .A(n17305), .B(n17304), .Z(n17427) );
  XNOR U17640 ( .A(a[123]), .B(b[9]), .Z(n17439) );
  NANDN U17641 ( .A(n17439), .B(n17814), .Z(n17308) );
  NANDN U17642 ( .A(n17306), .B(n17815), .Z(n17307) );
  AND U17643 ( .A(n17308), .B(n17307), .Z(n17428) );
  XNOR U17644 ( .A(n17427), .B(n17428), .Z(n17429) );
  XNOR U17645 ( .A(n17430), .B(n17429), .Z(n17499) );
  NANDN U17646 ( .A(n585), .B(a[99]), .Z(n17409) );
  ANDN U17647 ( .B(n17309), .A(n578), .Z(n17407) );
  XNOR U17648 ( .A(n17406), .B(n17407), .Z(n17408) );
  XNOR U17649 ( .A(n17409), .B(n17408), .Z(n17400) );
  XNOR U17650 ( .A(a[127]), .B(b[5]), .Z(n17443) );
  NANDN U17651 ( .A(n17443), .B(n17310), .Z(n17314) );
  NANDN U17652 ( .A(n17312), .B(n17311), .Z(n17313) );
  NAND U17653 ( .A(n17314), .B(n17313), .Z(n17401) );
  XNOR U17654 ( .A(n17400), .B(n17401), .Z(n17402) );
  XNOR U17655 ( .A(b[19]), .B(a[113]), .Z(n17472) );
  NANDN U17656 ( .A(n17472), .B(n18834), .Z(n17317) );
  NANDN U17657 ( .A(n17315), .B(n18832), .Z(n17316) );
  AND U17658 ( .A(n17317), .B(n17316), .Z(n17403) );
  XNOR U17659 ( .A(n17402), .B(n17403), .Z(n17500) );
  XOR U17660 ( .A(n17499), .B(n17500), .Z(n17502) );
  XOR U17661 ( .A(n17501), .B(n17502), .Z(n17388) );
  NANDN U17662 ( .A(n17319), .B(n17318), .Z(n17323) );
  NAND U17663 ( .A(n17321), .B(n17320), .Z(n17322) );
  NAND U17664 ( .A(n17323), .B(n17322), .Z(n17495) );
  XNOR U17665 ( .A(a[121]), .B(b[11]), .Z(n17463) );
  OR U17666 ( .A(n17463), .B(n18194), .Z(n17326) );
  NANDN U17667 ( .A(n17324), .B(n18104), .Z(n17325) );
  NAND U17668 ( .A(n17326), .B(n17325), .Z(n17454) );
  XOR U17669 ( .A(b[25]), .B(a[107]), .Z(n17460) );
  NAND U17670 ( .A(n17460), .B(n19240), .Z(n17329) );
  NANDN U17671 ( .A(n17327), .B(n19242), .Z(n17328) );
  NAND U17672 ( .A(n17329), .B(n17328), .Z(n17451) );
  XNOR U17673 ( .A(b[27]), .B(a[105]), .Z(n17436) );
  NANDN U17674 ( .A(n17436), .B(n19336), .Z(n17332) );
  NANDN U17675 ( .A(n17330), .B(n19337), .Z(n17331) );
  AND U17676 ( .A(n17332), .B(n17331), .Z(n17452) );
  XNOR U17677 ( .A(n17451), .B(n17452), .Z(n17453) );
  XNOR U17678 ( .A(n17454), .B(n17453), .Z(n17493) );
  NANDN U17679 ( .A(n17333), .B(n17553), .Z(n17335) );
  XNOR U17680 ( .A(a[125]), .B(b[7]), .Z(n17466) );
  NANDN U17681 ( .A(n17466), .B(n17555), .Z(n17334) );
  NAND U17682 ( .A(n17335), .B(n17334), .Z(n17397) );
  XNOR U17683 ( .A(n585), .B(a[101]), .Z(n17448) );
  NAND U17684 ( .A(n17448), .B(n19472), .Z(n17338) );
  NANDN U17685 ( .A(n17336), .B(n19473), .Z(n17337) );
  NAND U17686 ( .A(n17338), .B(n17337), .Z(n17394) );
  NANDN U17687 ( .A(n17339), .B(n19013), .Z(n17341) );
  XNOR U17688 ( .A(b[21]), .B(a[111]), .Z(n17433) );
  NANDN U17689 ( .A(n17433), .B(n19015), .Z(n17340) );
  AND U17690 ( .A(n17341), .B(n17340), .Z(n17395) );
  XNOR U17691 ( .A(n17394), .B(n17395), .Z(n17396) );
  XOR U17692 ( .A(n17397), .B(n17396), .Z(n17494) );
  XOR U17693 ( .A(n17493), .B(n17494), .Z(n17496) );
  XOR U17694 ( .A(n17495), .B(n17496), .Z(n17389) );
  XOR U17695 ( .A(n17388), .B(n17389), .Z(n17390) );
  XNOR U17696 ( .A(n17391), .B(n17390), .Z(n17384) );
  NANDN U17697 ( .A(n17343), .B(n17342), .Z(n17347) );
  OR U17698 ( .A(n17345), .B(n17344), .Z(n17346) );
  NAND U17699 ( .A(n17347), .B(n17346), .Z(n17385) );
  XNOR U17700 ( .A(n17384), .B(n17385), .Z(n17386) );
  XOR U17701 ( .A(n17387), .B(n17386), .Z(n17381) );
  XNOR U17702 ( .A(n17380), .B(n17381), .Z(n17375) );
  OR U17703 ( .A(n17353), .B(n17352), .Z(n17357) );
  NANDN U17704 ( .A(n17355), .B(n17354), .Z(n17356) );
  NAND U17705 ( .A(n17357), .B(n17356), .Z(n17373) );
  XNOR U17706 ( .A(n17372), .B(n17373), .Z(n17374) );
  XNOR U17707 ( .A(n17375), .B(n17374), .Z(n17367) );
  NANDN U17708 ( .A(n17359), .B(n17358), .Z(n17363) );
  OR U17709 ( .A(n17361), .B(n17360), .Z(n17362) );
  AND U17710 ( .A(n17363), .B(n17362), .Z(n17366) );
  XNOR U17711 ( .A(n17367), .B(n17366), .Z(n17368) );
  XNOR U17712 ( .A(n17369), .B(n17368), .Z(n17364) );
  XOR U17713 ( .A(n17365), .B(n17364), .Z(c[227]) );
  OR U17714 ( .A(n17365), .B(n17364), .Z(n17637) );
  NANDN U17715 ( .A(n17367), .B(n17366), .Z(n17371) );
  NANDN U17716 ( .A(n17369), .B(n17368), .Z(n17370) );
  NAND U17717 ( .A(n17371), .B(n17370), .Z(n17508) );
  NANDN U17718 ( .A(n17373), .B(n17372), .Z(n17377) );
  NAND U17719 ( .A(n17375), .B(n17374), .Z(n17376) );
  NAND U17720 ( .A(n17377), .B(n17376), .Z(n17505) );
  NANDN U17721 ( .A(n17379), .B(n17378), .Z(n17383) );
  NAND U17722 ( .A(n17381), .B(n17380), .Z(n17382) );
  NAND U17723 ( .A(n17383), .B(n17382), .Z(n17514) );
  NAND U17724 ( .A(n17389), .B(n17388), .Z(n17393) );
  NAND U17725 ( .A(n17391), .B(n17390), .Z(n17392) );
  NAND U17726 ( .A(n17393), .B(n17392), .Z(n17609) );
  NANDN U17727 ( .A(n17395), .B(n17394), .Z(n17399) );
  NAND U17728 ( .A(n17397), .B(n17396), .Z(n17398) );
  NAND U17729 ( .A(n17399), .B(n17398), .Z(n17612) );
  NANDN U17730 ( .A(n17401), .B(n17400), .Z(n17405) );
  NAND U17731 ( .A(n17403), .B(n17402), .Z(n17404) );
  NAND U17732 ( .A(n17405), .B(n17404), .Z(n17613) );
  XNOR U17733 ( .A(n17612), .B(n17613), .Z(n17614) );
  OR U17734 ( .A(n17407), .B(n17406), .Z(n17411) );
  OR U17735 ( .A(n17409), .B(n17408), .Z(n17410) );
  AND U17736 ( .A(n17411), .B(n17410), .Z(n17600) );
  NANDN U17737 ( .A(n17412), .B(n18513), .Z(n17414) );
  XNOR U17738 ( .A(a[118]), .B(b[15]), .Z(n17535) );
  OR U17739 ( .A(n17535), .B(n18512), .Z(n17413) );
  NAND U17740 ( .A(n17414), .B(n17413), .Z(n17591) );
  XNOR U17741 ( .A(a[116]), .B(b[17]), .Z(n17541) );
  NANDN U17742 ( .A(n17541), .B(n18673), .Z(n17417) );
  NANDN U17743 ( .A(n17415), .B(n18674), .Z(n17416) );
  NAND U17744 ( .A(n17417), .B(n17416), .Z(n17588) );
  XOR U17745 ( .A(a[120]), .B(n580), .Z(n17538) );
  NANDN U17746 ( .A(n17538), .B(n18336), .Z(n17420) );
  NANDN U17747 ( .A(n17418), .B(n18337), .Z(n17419) );
  AND U17748 ( .A(n17420), .B(n17419), .Z(n17589) );
  XNOR U17749 ( .A(n17588), .B(n17589), .Z(n17590) );
  XNOR U17750 ( .A(n17591), .B(n17590), .Z(n17601) );
  XNOR U17751 ( .A(n17600), .B(n17601), .Z(n17602) );
  NANDN U17752 ( .A(n17422), .B(n17421), .Z(n17426) );
  NAND U17753 ( .A(n17424), .B(n17423), .Z(n17425) );
  AND U17754 ( .A(n17426), .B(n17425), .Z(n17603) );
  XOR U17755 ( .A(n17614), .B(n17615), .Z(n17606) );
  NANDN U17756 ( .A(n17428), .B(n17427), .Z(n17432) );
  NAND U17757 ( .A(n17430), .B(n17429), .Z(n17431) );
  NAND U17758 ( .A(n17432), .B(n17431), .Z(n17626) );
  NANDN U17759 ( .A(n17433), .B(n19013), .Z(n17435) );
  XOR U17760 ( .A(b[21]), .B(n18582), .Z(n17558) );
  NANDN U17761 ( .A(n17558), .B(n19015), .Z(n17434) );
  NAND U17762 ( .A(n17435), .B(n17434), .Z(n17597) );
  XOR U17763 ( .A(b[27]), .B(n17690), .Z(n17578) );
  NANDN U17764 ( .A(n17578), .B(n19336), .Z(n17438) );
  NANDN U17765 ( .A(n17436), .B(n19337), .Z(n17437) );
  NAND U17766 ( .A(n17438), .B(n17437), .Z(n17594) );
  XOR U17767 ( .A(a[124]), .B(n579), .Z(n17575) );
  NANDN U17768 ( .A(n17575), .B(n17814), .Z(n17441) );
  NANDN U17769 ( .A(n17439), .B(n17815), .Z(n17440) );
  AND U17770 ( .A(n17441), .B(n17440), .Z(n17595) );
  XNOR U17771 ( .A(n17594), .B(n17595), .Z(n17596) );
  XNOR U17772 ( .A(n17597), .B(n17596), .Z(n17624) );
  XNOR U17773 ( .A(b[5]), .B(n17442), .Z(n17446) );
  XOR U17774 ( .A(n578), .B(b[4]), .Z(n17444) );
  NAND U17775 ( .A(n17444), .B(n17443), .Z(n17445) );
  AND U17776 ( .A(n17446), .B(n17445), .Z(n17567) );
  ANDN U17777 ( .B(b[31]), .A(n17447), .Z(n17581) );
  XNOR U17778 ( .A(n17567), .B(n17581), .Z(n17568) );
  XOR U17779 ( .A(n585), .B(a[102]), .Z(n17582) );
  NANDN U17780 ( .A(n17582), .B(n19472), .Z(n17450) );
  NAND U17781 ( .A(n19473), .B(n17448), .Z(n17449) );
  AND U17782 ( .A(n17450), .B(n17449), .Z(n17569) );
  XNOR U17783 ( .A(n17568), .B(n17569), .Z(n17625) );
  XOR U17784 ( .A(n17624), .B(n17625), .Z(n17627) );
  XNOR U17785 ( .A(n17626), .B(n17627), .Z(n17523) );
  NANDN U17786 ( .A(n17452), .B(n17451), .Z(n17456) );
  NAND U17787 ( .A(n17454), .B(n17453), .Z(n17455) );
  NAND U17788 ( .A(n17456), .B(n17455), .Z(n17620) );
  XNOR U17789 ( .A(b[23]), .B(a[110]), .Z(n17572) );
  OR U17790 ( .A(n17572), .B(n19127), .Z(n17459) );
  NAND U17791 ( .A(n17457), .B(n19128), .Z(n17458) );
  NAND U17792 ( .A(n17459), .B(n17458), .Z(n17532) );
  XNOR U17793 ( .A(b[25]), .B(a[108]), .Z(n17544) );
  NANDN U17794 ( .A(n17544), .B(n19240), .Z(n17462) );
  NAND U17795 ( .A(n17460), .B(n19242), .Z(n17461) );
  NAND U17796 ( .A(n17462), .B(n17461), .Z(n17529) );
  XNOR U17797 ( .A(a[122]), .B(b[11]), .Z(n17547) );
  OR U17798 ( .A(n17547), .B(n18194), .Z(n17465) );
  NANDN U17799 ( .A(n17463), .B(n18104), .Z(n17464) );
  AND U17800 ( .A(n17465), .B(n17464), .Z(n17530) );
  XNOR U17801 ( .A(n17529), .B(n17530), .Z(n17531) );
  XNOR U17802 ( .A(n17532), .B(n17531), .Z(n17618) );
  NANDN U17803 ( .A(n17466), .B(n17553), .Z(n17468) );
  XNOR U17804 ( .A(a[126]), .B(b[7]), .Z(n17554) );
  NANDN U17805 ( .A(n17554), .B(n17555), .Z(n17467) );
  NAND U17806 ( .A(n17468), .B(n17467), .Z(n17564) );
  NAND U17807 ( .A(n19406), .B(n17469), .Z(n17471) );
  XOR U17808 ( .A(n584), .B(n17716), .Z(n17550) );
  NANDN U17809 ( .A(n576), .B(n17550), .Z(n17470) );
  NAND U17810 ( .A(n17471), .B(n17470), .Z(n17561) );
  NANDN U17811 ( .A(n17472), .B(n18832), .Z(n17474) );
  XOR U17812 ( .A(n581), .B(n18751), .Z(n17585) );
  NAND U17813 ( .A(n17585), .B(n18834), .Z(n17473) );
  AND U17814 ( .A(n17474), .B(n17473), .Z(n17562) );
  XNOR U17815 ( .A(n17561), .B(n17562), .Z(n17563) );
  XOR U17816 ( .A(n17564), .B(n17563), .Z(n17619) );
  XOR U17817 ( .A(n17618), .B(n17619), .Z(n17621) );
  XOR U17818 ( .A(n17620), .B(n17621), .Z(n17524) );
  XNOR U17819 ( .A(n17523), .B(n17524), .Z(n17525) );
  NANDN U17820 ( .A(n17476), .B(n17475), .Z(n17480) );
  NAND U17821 ( .A(n17478), .B(n17477), .Z(n17479) );
  NAND U17822 ( .A(n17480), .B(n17479), .Z(n17526) );
  XNOR U17823 ( .A(n17525), .B(n17526), .Z(n17607) );
  XNOR U17824 ( .A(n17606), .B(n17607), .Z(n17608) );
  XNOR U17825 ( .A(n17609), .B(n17608), .Z(n17520) );
  NAND U17826 ( .A(n17482), .B(n17481), .Z(n17486) );
  NAND U17827 ( .A(n17484), .B(n17483), .Z(n17485) );
  NAND U17828 ( .A(n17486), .B(n17485), .Z(n17517) );
  NANDN U17829 ( .A(n17488), .B(n17487), .Z(n17492) );
  NAND U17830 ( .A(n17490), .B(n17489), .Z(n17491) );
  NAND U17831 ( .A(n17492), .B(n17491), .Z(n17633) );
  NANDN U17832 ( .A(n17494), .B(n17493), .Z(n17498) );
  OR U17833 ( .A(n17496), .B(n17495), .Z(n17497) );
  NAND U17834 ( .A(n17498), .B(n17497), .Z(n17630) );
  NANDN U17835 ( .A(n17500), .B(n17499), .Z(n17504) );
  OR U17836 ( .A(n17502), .B(n17501), .Z(n17503) );
  AND U17837 ( .A(n17504), .B(n17503), .Z(n17631) );
  XNOR U17838 ( .A(n17630), .B(n17631), .Z(n17632) );
  XNOR U17839 ( .A(n17633), .B(n17632), .Z(n17518) );
  XNOR U17840 ( .A(n17517), .B(n17518), .Z(n17519) );
  XNOR U17841 ( .A(n17520), .B(n17519), .Z(n17512) );
  XNOR U17842 ( .A(n17511), .B(n17512), .Z(n17513) );
  XOR U17843 ( .A(n17514), .B(n17513), .Z(n17506) );
  XNOR U17844 ( .A(n17505), .B(n17506), .Z(n17507) );
  XOR U17845 ( .A(n17508), .B(n17507), .Z(n17636) );
  XOR U17846 ( .A(n17637), .B(n17636), .Z(c[228]) );
  NANDN U17847 ( .A(n17506), .B(n17505), .Z(n17510) );
  NAND U17848 ( .A(n17508), .B(n17507), .Z(n17509) );
  NAND U17849 ( .A(n17510), .B(n17509), .Z(n17641) );
  NANDN U17850 ( .A(n17512), .B(n17511), .Z(n17516) );
  NAND U17851 ( .A(n17514), .B(n17513), .Z(n17515) );
  NAND U17852 ( .A(n17516), .B(n17515), .Z(n17638) );
  NANDN U17853 ( .A(n17518), .B(n17517), .Z(n17522) );
  NANDN U17854 ( .A(n17520), .B(n17519), .Z(n17521) );
  NAND U17855 ( .A(n17522), .B(n17521), .Z(n17762) );
  NANDN U17856 ( .A(n17524), .B(n17523), .Z(n17528) );
  NANDN U17857 ( .A(n17526), .B(n17525), .Z(n17527) );
  NAND U17858 ( .A(n17528), .B(n17527), .Z(n17653) );
  NANDN U17859 ( .A(n17530), .B(n17529), .Z(n17534) );
  NAND U17860 ( .A(n17532), .B(n17531), .Z(n17533) );
  NAND U17861 ( .A(n17534), .B(n17533), .Z(n17661) );
  NANDN U17862 ( .A(n17535), .B(n18513), .Z(n17537) );
  XNOR U17863 ( .A(a[119]), .B(b[15]), .Z(n17738) );
  OR U17864 ( .A(n17738), .B(n18512), .Z(n17536) );
  NAND U17865 ( .A(n17537), .B(n17536), .Z(n17723) );
  XOR U17866 ( .A(a[121]), .B(n580), .Z(n17741) );
  NANDN U17867 ( .A(n17741), .B(n18336), .Z(n17540) );
  NANDN U17868 ( .A(n17538), .B(n18337), .Z(n17539) );
  NAND U17869 ( .A(n17540), .B(n17539), .Z(n17720) );
  XNOR U17870 ( .A(a[117]), .B(b[17]), .Z(n17693) );
  NANDN U17871 ( .A(n17693), .B(n18673), .Z(n17543) );
  NANDN U17872 ( .A(n17541), .B(n18674), .Z(n17542) );
  NAND U17873 ( .A(n17543), .B(n17542), .Z(n17683) );
  XOR U17874 ( .A(b[25]), .B(a[109]), .Z(n17744) );
  NAND U17875 ( .A(n17744), .B(n19240), .Z(n17546) );
  NANDN U17876 ( .A(n17544), .B(n19242), .Z(n17545) );
  NAND U17877 ( .A(n17546), .B(n17545), .Z(n17680) );
  XOR U17878 ( .A(a[123]), .B(b[11]), .Z(n17705) );
  NANDN U17879 ( .A(n18194), .B(n17705), .Z(n17549) );
  NANDN U17880 ( .A(n17547), .B(n18104), .Z(n17548) );
  AND U17881 ( .A(n17549), .B(n17548), .Z(n17681) );
  XNOR U17882 ( .A(n17680), .B(n17681), .Z(n17682) );
  XNOR U17883 ( .A(n17683), .B(n17682), .Z(n17721) );
  XNOR U17884 ( .A(n17720), .B(n17721), .Z(n17722) );
  XNOR U17885 ( .A(n17723), .B(n17722), .Z(n17667) );
  NAND U17886 ( .A(n19406), .B(n17550), .Z(n17552) );
  XNOR U17887 ( .A(n584), .B(a[105]), .Z(n17689) );
  NANDN U17888 ( .A(n576), .B(n17689), .Z(n17551) );
  NAND U17889 ( .A(n17552), .B(n17551), .Z(n17750) );
  NANDN U17890 ( .A(n17554), .B(n17553), .Z(n17557) );
  XNOR U17891 ( .A(n19502), .B(b[7]), .Z(n17713) );
  NAND U17892 ( .A(n17713), .B(n17555), .Z(n17556) );
  NAND U17893 ( .A(n17557), .B(n17556), .Z(n17747) );
  NANDN U17894 ( .A(n17558), .B(n19013), .Z(n17560) );
  XNOR U17895 ( .A(b[21]), .B(a[113]), .Z(n17702) );
  NANDN U17896 ( .A(n17702), .B(n19015), .Z(n17559) );
  AND U17897 ( .A(n17560), .B(n17559), .Z(n17748) );
  XNOR U17898 ( .A(n17747), .B(n17748), .Z(n17749) );
  XNOR U17899 ( .A(n17750), .B(n17749), .Z(n17664) );
  NANDN U17900 ( .A(n17562), .B(n17561), .Z(n17566) );
  NAND U17901 ( .A(n17564), .B(n17563), .Z(n17565) );
  NAND U17902 ( .A(n17566), .B(n17565), .Z(n17665) );
  XNOR U17903 ( .A(n17664), .B(n17665), .Z(n17666) );
  XOR U17904 ( .A(n17667), .B(n17666), .Z(n17660) );
  XNOR U17905 ( .A(n17661), .B(n17660), .Z(n17662) );
  IV U17906 ( .A(n17581), .Z(n17735) );
  OR U17907 ( .A(n17567), .B(n17735), .Z(n17571) );
  NAND U17908 ( .A(n17569), .B(n17568), .Z(n17570) );
  NAND U17909 ( .A(n17571), .B(n17570), .Z(n17671) );
  XOR U17910 ( .A(b[23]), .B(a[111]), .Z(n17699) );
  NANDN U17911 ( .A(n19127), .B(n17699), .Z(n17574) );
  NANDN U17912 ( .A(n17572), .B(n19128), .Z(n17573) );
  NAND U17913 ( .A(n17574), .B(n17573), .Z(n17729) );
  XOR U17914 ( .A(a[125]), .B(n579), .Z(n17708) );
  NANDN U17915 ( .A(n17708), .B(n17814), .Z(n17577) );
  NANDN U17916 ( .A(n17575), .B(n17815), .Z(n17576) );
  NAND U17917 ( .A(n17577), .B(n17576), .Z(n17726) );
  XNOR U17918 ( .A(b[27]), .B(a[107]), .Z(n17686) );
  NANDN U17919 ( .A(n17686), .B(n19336), .Z(n17580) );
  NANDN U17920 ( .A(n17578), .B(n19337), .Z(n17579) );
  AND U17921 ( .A(n17580), .B(n17579), .Z(n17727) );
  XNOR U17922 ( .A(n17726), .B(n17727), .Z(n17728) );
  XNOR U17923 ( .A(n17729), .B(n17728), .Z(n17668) );
  NANDN U17924 ( .A(n585), .B(a[101]), .Z(n17732) );
  XOR U17925 ( .A(n17733), .B(n17732), .Z(n17734) );
  XOR U17926 ( .A(n17581), .B(n17734), .Z(n17675) );
  XOR U17927 ( .A(n585), .B(a[103]), .Z(n17717) );
  NANDN U17928 ( .A(n17717), .B(n19472), .Z(n17584) );
  NANDN U17929 ( .A(n17582), .B(n19473), .Z(n17583) );
  NAND U17930 ( .A(n17584), .B(n17583), .Z(n17674) );
  XOR U17931 ( .A(n17675), .B(n17674), .Z(n17676) );
  XOR U17932 ( .A(n581), .B(a[115]), .Z(n17696) );
  NANDN U17933 ( .A(n17696), .B(n18834), .Z(n17587) );
  NAND U17934 ( .A(n18832), .B(n17585), .Z(n17586) );
  AND U17935 ( .A(n17587), .B(n17586), .Z(n17677) );
  XNOR U17936 ( .A(n17676), .B(n17677), .Z(n17669) );
  XNOR U17937 ( .A(n17668), .B(n17669), .Z(n17670) );
  XNOR U17938 ( .A(n17671), .B(n17670), .Z(n17756) );
  NANDN U17939 ( .A(n17589), .B(n17588), .Z(n17593) );
  NAND U17940 ( .A(n17591), .B(n17590), .Z(n17592) );
  NAND U17941 ( .A(n17593), .B(n17592), .Z(n17754) );
  NANDN U17942 ( .A(n17595), .B(n17594), .Z(n17599) );
  NAND U17943 ( .A(n17597), .B(n17596), .Z(n17598) );
  AND U17944 ( .A(n17599), .B(n17598), .Z(n17753) );
  XNOR U17945 ( .A(n17754), .B(n17753), .Z(n17755) );
  XOR U17946 ( .A(n17756), .B(n17755), .Z(n17663) );
  XOR U17947 ( .A(n17662), .B(n17663), .Z(n17650) );
  OR U17948 ( .A(n17601), .B(n17600), .Z(n17605) );
  OR U17949 ( .A(n17603), .B(n17602), .Z(n17604) );
  AND U17950 ( .A(n17605), .B(n17604), .Z(n17651) );
  XNOR U17951 ( .A(n17650), .B(n17651), .Z(n17652) );
  XNOR U17952 ( .A(n17653), .B(n17652), .Z(n17759) );
  NANDN U17953 ( .A(n17607), .B(n17606), .Z(n17611) );
  NAND U17954 ( .A(n17609), .B(n17608), .Z(n17610) );
  NAND U17955 ( .A(n17611), .B(n17610), .Z(n17647) );
  NANDN U17956 ( .A(n17613), .B(n17612), .Z(n17617) );
  NANDN U17957 ( .A(n17615), .B(n17614), .Z(n17616) );
  NAND U17958 ( .A(n17617), .B(n17616), .Z(n17657) );
  NANDN U17959 ( .A(n17619), .B(n17618), .Z(n17623) );
  OR U17960 ( .A(n17621), .B(n17620), .Z(n17622) );
  NAND U17961 ( .A(n17623), .B(n17622), .Z(n17654) );
  NANDN U17962 ( .A(n17625), .B(n17624), .Z(n17629) );
  OR U17963 ( .A(n17627), .B(n17626), .Z(n17628) );
  AND U17964 ( .A(n17629), .B(n17628), .Z(n17655) );
  XNOR U17965 ( .A(n17654), .B(n17655), .Z(n17656) );
  XOR U17966 ( .A(n17657), .B(n17656), .Z(n17644) );
  NANDN U17967 ( .A(n17631), .B(n17630), .Z(n17635) );
  NAND U17968 ( .A(n17633), .B(n17632), .Z(n17634) );
  NAND U17969 ( .A(n17635), .B(n17634), .Z(n17645) );
  XNOR U17970 ( .A(n17644), .B(n17645), .Z(n17646) );
  XNOR U17971 ( .A(n17647), .B(n17646), .Z(n17760) );
  XNOR U17972 ( .A(n17759), .B(n17760), .Z(n17761) );
  XOR U17973 ( .A(n17762), .B(n17761), .Z(n17639) );
  XNOR U17974 ( .A(n17638), .B(n17639), .Z(n17640) );
  XNOR U17975 ( .A(n17641), .B(n17640), .Z(n17765) );
  OR U17976 ( .A(n17637), .B(n17636), .Z(n17766) );
  XNOR U17977 ( .A(n17765), .B(n17766), .Z(c[229]) );
  NANDN U17978 ( .A(n17639), .B(n17638), .Z(n17643) );
  NANDN U17979 ( .A(n17641), .B(n17640), .Z(n17642) );
  NAND U17980 ( .A(n17643), .B(n17642), .Z(n17769) );
  NANDN U17981 ( .A(n17645), .B(n17644), .Z(n17649) );
  NANDN U17982 ( .A(n17647), .B(n17646), .Z(n17648) );
  NAND U17983 ( .A(n17649), .B(n17648), .Z(n17775) );
  NANDN U17984 ( .A(n17655), .B(n17654), .Z(n17659) );
  NANDN U17985 ( .A(n17657), .B(n17656), .Z(n17658) );
  NAND U17986 ( .A(n17659), .B(n17658), .Z(n17781) );
  NANDN U17987 ( .A(n17669), .B(n17668), .Z(n17673) );
  NAND U17988 ( .A(n17671), .B(n17670), .Z(n17672) );
  NAND U17989 ( .A(n17673), .B(n17672), .Z(n17865) );
  OR U17990 ( .A(n17675), .B(n17674), .Z(n17679) );
  NAND U17991 ( .A(n17677), .B(n17676), .Z(n17678) );
  NAND U17992 ( .A(n17679), .B(n17678), .Z(n17870) );
  NANDN U17993 ( .A(n17681), .B(n17680), .Z(n17685) );
  NAND U17994 ( .A(n17683), .B(n17682), .Z(n17684) );
  NAND U17995 ( .A(n17685), .B(n17684), .Z(n17871) );
  XNOR U17996 ( .A(n17870), .B(n17871), .Z(n17872) );
  XOR U17997 ( .A(b[27]), .B(n18198), .Z(n17840) );
  NANDN U17998 ( .A(n17840), .B(n19336), .Z(n17688) );
  NANDN U17999 ( .A(n17686), .B(n19337), .Z(n17687) );
  NAND U18000 ( .A(n17688), .B(n17687), .Z(n17800) );
  NAND U18001 ( .A(n19406), .B(n17689), .Z(n17692) );
  XOR U18002 ( .A(n584), .B(n17690), .Z(n17822) );
  NANDN U18003 ( .A(n576), .B(n17822), .Z(n17691) );
  NAND U18004 ( .A(n17692), .B(n17691), .Z(n17797) );
  XNOR U18005 ( .A(a[118]), .B(b[17]), .Z(n17846) );
  NANDN U18006 ( .A(n17846), .B(n18673), .Z(n17695) );
  NANDN U18007 ( .A(n17693), .B(n18674), .Z(n17694) );
  AND U18008 ( .A(n17695), .B(n17694), .Z(n17798) );
  XNOR U18009 ( .A(n17797), .B(n17798), .Z(n17799) );
  XNOR U18010 ( .A(n17800), .B(n17799), .Z(n17861) );
  XOR U18011 ( .A(a[116]), .B(n581), .Z(n17849) );
  NANDN U18012 ( .A(n17849), .B(n18834), .Z(n17698) );
  NANDN U18013 ( .A(n17696), .B(n18832), .Z(n17697) );
  NAND U18014 ( .A(n17698), .B(n17697), .Z(n17859) );
  XNOR U18015 ( .A(b[23]), .B(a[112]), .Z(n17828) );
  OR U18016 ( .A(n17828), .B(n19127), .Z(n17701) );
  NAND U18017 ( .A(n19128), .B(n17699), .Z(n17700) );
  AND U18018 ( .A(n17701), .B(n17700), .Z(n17858) );
  XNOR U18019 ( .A(n17859), .B(n17858), .Z(n17860) );
  XOR U18020 ( .A(n17861), .B(n17860), .Z(n17884) );
  NANDN U18021 ( .A(n17702), .B(n19013), .Z(n17704) );
  XOR U18022 ( .A(b[21]), .B(n18751), .Z(n17819) );
  NANDN U18023 ( .A(n17819), .B(n19015), .Z(n17703) );
  NAND U18024 ( .A(n17704), .B(n17703), .Z(n17806) );
  XNOR U18025 ( .A(a[124]), .B(b[11]), .Z(n17843) );
  OR U18026 ( .A(n17843), .B(n18194), .Z(n17707) );
  NAND U18027 ( .A(n17705), .B(n18104), .Z(n17706) );
  NAND U18028 ( .A(n17707), .B(n17706), .Z(n17803) );
  XOR U18029 ( .A(a[126]), .B(n579), .Z(n17816) );
  NANDN U18030 ( .A(n17816), .B(n17814), .Z(n17710) );
  NANDN U18031 ( .A(n17708), .B(n17815), .Z(n17709) );
  AND U18032 ( .A(n17710), .B(n17709), .Z(n17804) );
  XNOR U18033 ( .A(n17803), .B(n17804), .Z(n17805) );
  XNOR U18034 ( .A(n17806), .B(n17805), .Z(n17882) );
  XNOR U18035 ( .A(b[7]), .B(n17711), .Z(n17715) );
  XNOR U18036 ( .A(b[6]), .B(b[5]), .Z(n17712) );
  NANDN U18037 ( .A(n17713), .B(n17712), .Z(n17714) );
  AND U18038 ( .A(n17715), .B(n17714), .Z(n17809) );
  AND U18039 ( .A(a[102]), .B(b[31]), .Z(n17973) );
  XNOR U18040 ( .A(n17809), .B(n17973), .Z(n17810) );
  XOR U18041 ( .A(b[31]), .B(n17716), .Z(n17825) );
  NANDN U18042 ( .A(n17825), .B(n19472), .Z(n17719) );
  NANDN U18043 ( .A(n17717), .B(n19473), .Z(n17718) );
  AND U18044 ( .A(n17719), .B(n17718), .Z(n17811) );
  XNOR U18045 ( .A(n17810), .B(n17811), .Z(n17883) );
  XOR U18046 ( .A(n17882), .B(n17883), .Z(n17885) );
  XNOR U18047 ( .A(n17884), .B(n17885), .Z(n17873) );
  XOR U18048 ( .A(n17872), .B(n17873), .Z(n17864) );
  XOR U18049 ( .A(n17865), .B(n17864), .Z(n17866) );
  XNOR U18050 ( .A(n17867), .B(n17866), .Z(n17788) );
  NANDN U18051 ( .A(n17721), .B(n17720), .Z(n17725) );
  NAND U18052 ( .A(n17723), .B(n17722), .Z(n17724) );
  NAND U18053 ( .A(n17725), .B(n17724), .Z(n17794) );
  NANDN U18054 ( .A(n17727), .B(n17726), .Z(n17731) );
  NAND U18055 ( .A(n17729), .B(n17728), .Z(n17730) );
  NAND U18056 ( .A(n17731), .B(n17730), .Z(n17876) );
  OR U18057 ( .A(n17733), .B(n17732), .Z(n17737) );
  NANDN U18058 ( .A(n17735), .B(n17734), .Z(n17736) );
  AND U18059 ( .A(n17737), .B(n17736), .Z(n17877) );
  XNOR U18060 ( .A(n17876), .B(n17877), .Z(n17878) );
  NANDN U18061 ( .A(n17738), .B(n18513), .Z(n17740) );
  XNOR U18062 ( .A(a[120]), .B(b[15]), .Z(n17855) );
  OR U18063 ( .A(n17855), .B(n18512), .Z(n17739) );
  NAND U18064 ( .A(n17740), .B(n17739), .Z(n17834) );
  XOR U18065 ( .A(a[122]), .B(n580), .Z(n17852) );
  NANDN U18066 ( .A(n17852), .B(n18336), .Z(n17743) );
  NANDN U18067 ( .A(n17741), .B(n18337), .Z(n17742) );
  NAND U18068 ( .A(n17743), .B(n17742), .Z(n17831) );
  XNOR U18069 ( .A(b[25]), .B(a[110]), .Z(n17837) );
  NANDN U18070 ( .A(n17837), .B(n19240), .Z(n17746) );
  NAND U18071 ( .A(n17744), .B(n19242), .Z(n17745) );
  AND U18072 ( .A(n17746), .B(n17745), .Z(n17832) );
  XNOR U18073 ( .A(n17831), .B(n17832), .Z(n17833) );
  XNOR U18074 ( .A(n17834), .B(n17833), .Z(n17879) );
  XOR U18075 ( .A(n17878), .B(n17879), .Z(n17791) );
  NANDN U18076 ( .A(n17748), .B(n17747), .Z(n17752) );
  NAND U18077 ( .A(n17750), .B(n17749), .Z(n17751) );
  NAND U18078 ( .A(n17752), .B(n17751), .Z(n17792) );
  XNOR U18079 ( .A(n17791), .B(n17792), .Z(n17793) );
  XOR U18080 ( .A(n17794), .B(n17793), .Z(n17785) );
  NANDN U18081 ( .A(n17754), .B(n17753), .Z(n17758) );
  NANDN U18082 ( .A(n17756), .B(n17755), .Z(n17757) );
  NAND U18083 ( .A(n17758), .B(n17757), .Z(n17786) );
  XNOR U18084 ( .A(n17785), .B(n17786), .Z(n17787) );
  XOR U18085 ( .A(n17788), .B(n17787), .Z(n17779) );
  XOR U18086 ( .A(n17780), .B(n17779), .Z(n17782) );
  XOR U18087 ( .A(n17781), .B(n17782), .Z(n17773) );
  XNOR U18088 ( .A(n17774), .B(n17773), .Z(n17776) );
  XNOR U18089 ( .A(n17775), .B(n17776), .Z(n17767) );
  NANDN U18090 ( .A(n17760), .B(n17759), .Z(n17764) );
  NAND U18091 ( .A(n17762), .B(n17761), .Z(n17763) );
  AND U18092 ( .A(n17764), .B(n17763), .Z(n17768) );
  XNOR U18093 ( .A(n17767), .B(n17768), .Z(n17770) );
  XNOR U18094 ( .A(n17769), .B(n17770), .Z(n17888) );
  NANDN U18095 ( .A(n17766), .B(n17765), .Z(n17889) );
  XNOR U18096 ( .A(n17888), .B(n17889), .Z(c[230]) );
  NAND U18097 ( .A(n17768), .B(n17767), .Z(n17772) );
  NANDN U18098 ( .A(n17770), .B(n17769), .Z(n17771) );
  NAND U18099 ( .A(n17772), .B(n17771), .Z(n17892) );
  NAND U18100 ( .A(n17774), .B(n17773), .Z(n17778) );
  NANDN U18101 ( .A(n17776), .B(n17775), .Z(n17777) );
  NAND U18102 ( .A(n17778), .B(n17777), .Z(n17891) );
  NANDN U18103 ( .A(n17780), .B(n17779), .Z(n17784) );
  OR U18104 ( .A(n17782), .B(n17781), .Z(n17783) );
  NAND U18105 ( .A(n17784), .B(n17783), .Z(n17898) );
  NANDN U18106 ( .A(n17786), .B(n17785), .Z(n17790) );
  NAND U18107 ( .A(n17788), .B(n17787), .Z(n17789) );
  NAND U18108 ( .A(n17790), .B(n17789), .Z(n17897) );
  NANDN U18109 ( .A(n17792), .B(n17791), .Z(n17796) );
  NANDN U18110 ( .A(n17794), .B(n17793), .Z(n17795) );
  NAND U18111 ( .A(n17796), .B(n17795), .Z(n18007) );
  NANDN U18112 ( .A(n17798), .B(n17797), .Z(n17802) );
  NAND U18113 ( .A(n17800), .B(n17799), .Z(n17801) );
  NAND U18114 ( .A(n17802), .B(n17801), .Z(n17914) );
  NANDN U18115 ( .A(n17804), .B(n17803), .Z(n17808) );
  NAND U18116 ( .A(n17806), .B(n17805), .Z(n17807) );
  AND U18117 ( .A(n17808), .B(n17807), .Z(n17915) );
  XNOR U18118 ( .A(n17914), .B(n17915), .Z(n17916) );
  NANDN U18119 ( .A(n17809), .B(n17973), .Z(n17813) );
  NAND U18120 ( .A(n17811), .B(n17810), .Z(n17812) );
  NAND U18121 ( .A(n17813), .B(n17812), .Z(n17923) );
  XNOR U18122 ( .A(n19502), .B(b[9]), .Z(n17965) );
  NAND U18123 ( .A(n17814), .B(n17965), .Z(n17818) );
  NANDN U18124 ( .A(n17816), .B(n17815), .Z(n17817) );
  NAND U18125 ( .A(n17818), .B(n17817), .Z(n17998) );
  NANDN U18126 ( .A(n17819), .B(n19013), .Z(n17821) );
  XOR U18127 ( .A(b[21]), .B(n19022), .Z(n17995) );
  NANDN U18128 ( .A(n17995), .B(n19015), .Z(n17820) );
  AND U18129 ( .A(n17821), .B(n17820), .Z(n17999) );
  XNOR U18130 ( .A(n17998), .B(n17999), .Z(n18000) );
  NANDN U18131 ( .A(n585), .B(a[103]), .Z(n17971) );
  XOR U18132 ( .A(n17972), .B(n17971), .Z(n17974) );
  XNOR U18133 ( .A(n17973), .B(n17974), .Z(n18001) );
  XNOR U18134 ( .A(n18000), .B(n18001), .Z(n17920) );
  NAND U18135 ( .A(n19406), .B(n17822), .Z(n17824) );
  XNOR U18136 ( .A(n584), .B(a[107]), .Z(n17992) );
  NANDN U18137 ( .A(n576), .B(n17992), .Z(n17823) );
  NAND U18138 ( .A(n17824), .B(n17823), .Z(n17980) );
  XNOR U18139 ( .A(n585), .B(a[105]), .Z(n17968) );
  NAND U18140 ( .A(n17968), .B(n19472), .Z(n17827) );
  NANDN U18141 ( .A(n17825), .B(n19473), .Z(n17826) );
  NAND U18142 ( .A(n17827), .B(n17826), .Z(n17977) );
  XOR U18143 ( .A(b[23]), .B(a[113]), .Z(n17942) );
  NANDN U18144 ( .A(n19127), .B(n17942), .Z(n17830) );
  NANDN U18145 ( .A(n17828), .B(n19128), .Z(n17829) );
  AND U18146 ( .A(n17830), .B(n17829), .Z(n17978) );
  XNOR U18147 ( .A(n17977), .B(n17978), .Z(n17979) );
  XOR U18148 ( .A(n17980), .B(n17979), .Z(n17921) );
  XOR U18149 ( .A(n17920), .B(n17921), .Z(n17922) );
  XOR U18150 ( .A(n17923), .B(n17922), .Z(n17917) );
  XOR U18151 ( .A(n17916), .B(n17917), .Z(n18004) );
  NANDN U18152 ( .A(n17832), .B(n17831), .Z(n17836) );
  NAND U18153 ( .A(n17834), .B(n17833), .Z(n17835) );
  NAND U18154 ( .A(n17836), .B(n17835), .Z(n17930) );
  XOR U18155 ( .A(b[25]), .B(a[111]), .Z(n17936) );
  NAND U18156 ( .A(n17936), .B(n19240), .Z(n17839) );
  NANDN U18157 ( .A(n17837), .B(n19242), .Z(n17838) );
  NAND U18158 ( .A(n17839), .B(n17838), .Z(n17960) );
  XNOR U18159 ( .A(b[27]), .B(a[109]), .Z(n17939) );
  NANDN U18160 ( .A(n17939), .B(n19336), .Z(n17842) );
  NANDN U18161 ( .A(n17840), .B(n19337), .Z(n17841) );
  NAND U18162 ( .A(n17842), .B(n17841), .Z(n17957) );
  XNOR U18163 ( .A(a[125]), .B(b[11]), .Z(n17989) );
  OR U18164 ( .A(n17989), .B(n18194), .Z(n17845) );
  NANDN U18165 ( .A(n17843), .B(n18104), .Z(n17844) );
  AND U18166 ( .A(n17845), .B(n17844), .Z(n17958) );
  XNOR U18167 ( .A(n17957), .B(n17958), .Z(n17959) );
  XNOR U18168 ( .A(n17960), .B(n17959), .Z(n17927) );
  XNOR U18169 ( .A(n19239), .B(b[17]), .Z(n17945) );
  NAND U18170 ( .A(n17945), .B(n18673), .Z(n17848) );
  NANDN U18171 ( .A(n17846), .B(n18674), .Z(n17847) );
  NAND U18172 ( .A(n17848), .B(n17847), .Z(n17986) );
  NANDN U18173 ( .A(n17849), .B(n18832), .Z(n17851) );
  XOR U18174 ( .A(b[19]), .B(n19136), .Z(n17951) );
  NANDN U18175 ( .A(n17951), .B(n18834), .Z(n17850) );
  NAND U18176 ( .A(n17851), .B(n17850), .Z(n17983) );
  XNOR U18177 ( .A(a[123]), .B(b[13]), .Z(n17954) );
  NANDN U18178 ( .A(n17954), .B(n18336), .Z(n17854) );
  NANDN U18179 ( .A(n17852), .B(n18337), .Z(n17853) );
  AND U18180 ( .A(n17854), .B(n17853), .Z(n17984) );
  XNOR U18181 ( .A(n17983), .B(n17984), .Z(n17985) );
  XNOR U18182 ( .A(n17986), .B(n17985), .Z(n17924) );
  XNOR U18183 ( .A(a[121]), .B(b[15]), .Z(n17948) );
  OR U18184 ( .A(n17948), .B(n18512), .Z(n17857) );
  NANDN U18185 ( .A(n17855), .B(n18513), .Z(n17856) );
  NAND U18186 ( .A(n17857), .B(n17856), .Z(n17925) );
  XNOR U18187 ( .A(n17924), .B(n17925), .Z(n17926) );
  XOR U18188 ( .A(n17927), .B(n17926), .Z(n17931) );
  XNOR U18189 ( .A(n17930), .B(n17931), .Z(n17932) );
  NANDN U18190 ( .A(n17859), .B(n17858), .Z(n17863) );
  NAND U18191 ( .A(n17861), .B(n17860), .Z(n17862) );
  NAND U18192 ( .A(n17863), .B(n17862), .Z(n17933) );
  XNOR U18193 ( .A(n17932), .B(n17933), .Z(n18005) );
  XNOR U18194 ( .A(n18004), .B(n18005), .Z(n18006) );
  XNOR U18195 ( .A(n18007), .B(n18006), .Z(n17905) );
  NAND U18196 ( .A(n17865), .B(n17864), .Z(n17869) );
  NAND U18197 ( .A(n17867), .B(n17866), .Z(n17868) );
  NAND U18198 ( .A(n17869), .B(n17868), .Z(n17902) );
  NANDN U18199 ( .A(n17871), .B(n17870), .Z(n17875) );
  NAND U18200 ( .A(n17873), .B(n17872), .Z(n17874) );
  NAND U18201 ( .A(n17875), .B(n17874), .Z(n17911) );
  NANDN U18202 ( .A(n17877), .B(n17876), .Z(n17881) );
  NANDN U18203 ( .A(n17879), .B(n17878), .Z(n17880) );
  NAND U18204 ( .A(n17881), .B(n17880), .Z(n17908) );
  NANDN U18205 ( .A(n17883), .B(n17882), .Z(n17887) );
  NANDN U18206 ( .A(n17885), .B(n17884), .Z(n17886) );
  NAND U18207 ( .A(n17887), .B(n17886), .Z(n17909) );
  XNOR U18208 ( .A(n17908), .B(n17909), .Z(n17910) );
  XOR U18209 ( .A(n17911), .B(n17910), .Z(n17903) );
  XOR U18210 ( .A(n17902), .B(n17903), .Z(n17904) );
  XOR U18211 ( .A(n17905), .B(n17904), .Z(n17896) );
  XNOR U18212 ( .A(n17897), .B(n17896), .Z(n17899) );
  XNOR U18213 ( .A(n17898), .B(n17899), .Z(n17890) );
  XNOR U18214 ( .A(n17891), .B(n17890), .Z(n17893) );
  XNOR U18215 ( .A(n17892), .B(n17893), .Z(n18010) );
  NANDN U18216 ( .A(n17889), .B(n17888), .Z(n18011) );
  XNOR U18217 ( .A(n18010), .B(n18011), .Z(c[231]) );
  NAND U18218 ( .A(n17891), .B(n17890), .Z(n17895) );
  NANDN U18219 ( .A(n17893), .B(n17892), .Z(n17894) );
  NAND U18220 ( .A(n17895), .B(n17894), .Z(n18017) );
  NAND U18221 ( .A(n17897), .B(n17896), .Z(n17901) );
  NANDN U18222 ( .A(n17899), .B(n17898), .Z(n17900) );
  NAND U18223 ( .A(n17901), .B(n17900), .Z(n18014) );
  OR U18224 ( .A(n17903), .B(n17902), .Z(n17907) );
  NAND U18225 ( .A(n17905), .B(n17904), .Z(n17906) );
  NAND U18226 ( .A(n17907), .B(n17906), .Z(n18120) );
  NANDN U18227 ( .A(n17909), .B(n17908), .Z(n17913) );
  NANDN U18228 ( .A(n17911), .B(n17910), .Z(n17912) );
  NAND U18229 ( .A(n17913), .B(n17912), .Z(n18020) );
  NANDN U18230 ( .A(n17915), .B(n17914), .Z(n17919) );
  NANDN U18231 ( .A(n17917), .B(n17916), .Z(n17918) );
  NAND U18232 ( .A(n17919), .B(n17918), .Z(n18114) );
  NANDN U18233 ( .A(n17925), .B(n17924), .Z(n17929) );
  NAND U18234 ( .A(n17927), .B(n17926), .Z(n17928) );
  NAND U18235 ( .A(n17929), .B(n17928), .Z(n18112) );
  XNOR U18236 ( .A(n18111), .B(n18112), .Z(n18113) );
  XNOR U18237 ( .A(n18114), .B(n18113), .Z(n18021) );
  XNOR U18238 ( .A(n18020), .B(n18021), .Z(n18022) );
  NANDN U18239 ( .A(n17931), .B(n17930), .Z(n17935) );
  NANDN U18240 ( .A(n17933), .B(n17932), .Z(n17934) );
  NAND U18241 ( .A(n17935), .B(n17934), .Z(n18029) );
  XNOR U18242 ( .A(b[25]), .B(a[112]), .Z(n18060) );
  NANDN U18243 ( .A(n18060), .B(n19240), .Z(n17938) );
  NAND U18244 ( .A(n17936), .B(n19242), .Z(n17937) );
  NAND U18245 ( .A(n17938), .B(n17937), .Z(n18083) );
  XOR U18246 ( .A(b[27]), .B(n18415), .Z(n18063) );
  NANDN U18247 ( .A(n18063), .B(n19336), .Z(n17941) );
  NANDN U18248 ( .A(n17939), .B(n19337), .Z(n17940) );
  NAND U18249 ( .A(n17941), .B(n17940), .Z(n18080) );
  XNOR U18250 ( .A(b[23]), .B(a[114]), .Z(n18108) );
  OR U18251 ( .A(n18108), .B(n19127), .Z(n17944) );
  NAND U18252 ( .A(n17942), .B(n19128), .Z(n17943) );
  AND U18253 ( .A(n17944), .B(n17943), .Z(n18081) );
  XNOR U18254 ( .A(n18080), .B(n18081), .Z(n18082) );
  XNOR U18255 ( .A(n18083), .B(n18082), .Z(n18045) );
  XNOR U18256 ( .A(a[120]), .B(b[17]), .Z(n18095) );
  NANDN U18257 ( .A(n18095), .B(n18673), .Z(n17947) );
  NAND U18258 ( .A(n17945), .B(n18674), .Z(n17946) );
  NAND U18259 ( .A(n17947), .B(n17946), .Z(n18042) );
  NANDN U18260 ( .A(n17948), .B(n18513), .Z(n17950) );
  XNOR U18261 ( .A(a[122]), .B(b[15]), .Z(n18098) );
  OR U18262 ( .A(n18098), .B(n18512), .Z(n17949) );
  NAND U18263 ( .A(n17950), .B(n17949), .Z(n18089) );
  NANDN U18264 ( .A(n17951), .B(n18832), .Z(n17953) );
  XOR U18265 ( .A(a[118]), .B(n581), .Z(n18066) );
  NANDN U18266 ( .A(n18066), .B(n18834), .Z(n17952) );
  NAND U18267 ( .A(n17953), .B(n17952), .Z(n18086) );
  XOR U18268 ( .A(a[124]), .B(n580), .Z(n18101) );
  NANDN U18269 ( .A(n18101), .B(n18336), .Z(n17956) );
  NANDN U18270 ( .A(n17954), .B(n18337), .Z(n17955) );
  AND U18271 ( .A(n17956), .B(n17955), .Z(n18087) );
  XNOR U18272 ( .A(n18086), .B(n18087), .Z(n18088) );
  XNOR U18273 ( .A(n18089), .B(n18088), .Z(n18043) );
  XNOR U18274 ( .A(n18042), .B(n18043), .Z(n18044) );
  XOR U18275 ( .A(n18045), .B(n18044), .Z(n18035) );
  NANDN U18276 ( .A(n17958), .B(n17957), .Z(n17962) );
  NAND U18277 ( .A(n17960), .B(n17959), .Z(n17961) );
  NAND U18278 ( .A(n17962), .B(n17961), .Z(n18051) );
  XOR U18279 ( .A(n579), .B(n17963), .Z(n17967) );
  XNOR U18280 ( .A(b[8]), .B(b[7]), .Z(n17964) );
  NANDN U18281 ( .A(n17965), .B(n17964), .Z(n17966) );
  AND U18282 ( .A(n17967), .B(n17966), .Z(n18075) );
  AND U18283 ( .A(a[104]), .B(b[31]), .Z(n18151) );
  XOR U18284 ( .A(n18075), .B(n18151), .Z(n18077) );
  XOR U18285 ( .A(n585), .B(a[106]), .Z(n18069) );
  NANDN U18286 ( .A(n18069), .B(n19472), .Z(n17970) );
  NAND U18287 ( .A(n19473), .B(n17968), .Z(n17969) );
  NAND U18288 ( .A(n17970), .B(n17969), .Z(n18076) );
  XNOR U18289 ( .A(n18077), .B(n18076), .Z(n18048) );
  OR U18290 ( .A(n17972), .B(n17971), .Z(n17976) );
  NAND U18291 ( .A(n17974), .B(n17973), .Z(n17975) );
  AND U18292 ( .A(n17976), .B(n17975), .Z(n18049) );
  XNOR U18293 ( .A(n18048), .B(n18049), .Z(n18050) );
  XNOR U18294 ( .A(n18051), .B(n18050), .Z(n18032) );
  NANDN U18295 ( .A(n17978), .B(n17977), .Z(n17982) );
  NAND U18296 ( .A(n17980), .B(n17979), .Z(n17981) );
  NAND U18297 ( .A(n17982), .B(n17981), .Z(n18033) );
  XNOR U18298 ( .A(n18032), .B(n18033), .Z(n18034) );
  XNOR U18299 ( .A(n18035), .B(n18034), .Z(n18026) );
  NANDN U18300 ( .A(n17984), .B(n17983), .Z(n17988) );
  NAND U18301 ( .A(n17986), .B(n17985), .Z(n17987) );
  NAND U18302 ( .A(n17988), .B(n17987), .Z(n18038) );
  XNOR U18303 ( .A(n19295), .B(b[11]), .Z(n18105) );
  NANDN U18304 ( .A(n18194), .B(n18105), .Z(n17991) );
  NANDN U18305 ( .A(n17989), .B(n18104), .Z(n17990) );
  NAND U18306 ( .A(n17991), .B(n17990), .Z(n18057) );
  NAND U18307 ( .A(n19406), .B(n17992), .Z(n17994) );
  XOR U18308 ( .A(b[29]), .B(n18198), .Z(n18092) );
  OR U18309 ( .A(n18092), .B(n576), .Z(n17993) );
  NAND U18310 ( .A(n17994), .B(n17993), .Z(n18054) );
  NANDN U18311 ( .A(n17995), .B(n19013), .Z(n17997) );
  XOR U18312 ( .A(n582), .B(n18950), .Z(n18072) );
  NAND U18313 ( .A(n18072), .B(n19015), .Z(n17996) );
  AND U18314 ( .A(n17997), .B(n17996), .Z(n18055) );
  XNOR U18315 ( .A(n18054), .B(n18055), .Z(n18056) );
  XNOR U18316 ( .A(n18057), .B(n18056), .Z(n18036) );
  NANDN U18317 ( .A(n17999), .B(n17998), .Z(n18003) );
  NANDN U18318 ( .A(n18001), .B(n18000), .Z(n18002) );
  NAND U18319 ( .A(n18003), .B(n18002), .Z(n18037) );
  XOR U18320 ( .A(n18036), .B(n18037), .Z(n18039) );
  XOR U18321 ( .A(n18038), .B(n18039), .Z(n18027) );
  XNOR U18322 ( .A(n18026), .B(n18027), .Z(n18028) );
  XNOR U18323 ( .A(n18029), .B(n18028), .Z(n18023) );
  XOR U18324 ( .A(n18022), .B(n18023), .Z(n18117) );
  NANDN U18325 ( .A(n18005), .B(n18004), .Z(n18009) );
  NAND U18326 ( .A(n18007), .B(n18006), .Z(n18008) );
  AND U18327 ( .A(n18009), .B(n18008), .Z(n18118) );
  XNOR U18328 ( .A(n18117), .B(n18118), .Z(n18119) );
  XNOR U18329 ( .A(n18120), .B(n18119), .Z(n18015) );
  XNOR U18330 ( .A(n18014), .B(n18015), .Z(n18016) );
  XNOR U18331 ( .A(n18017), .B(n18016), .Z(n18013) );
  NANDN U18332 ( .A(n18011), .B(n18010), .Z(n18012) );
  XOR U18333 ( .A(n18013), .B(n18012), .Z(c[232]) );
  OR U18334 ( .A(n18013), .B(n18012), .Z(n18239) );
  NANDN U18335 ( .A(n18015), .B(n18014), .Z(n18019) );
  NAND U18336 ( .A(n18017), .B(n18016), .Z(n18018) );
  AND U18337 ( .A(n18019), .B(n18018), .Z(n18128) );
  NANDN U18338 ( .A(n18021), .B(n18020), .Z(n18025) );
  NANDN U18339 ( .A(n18023), .B(n18022), .Z(n18024) );
  NAND U18340 ( .A(n18025), .B(n18024), .Z(n18235) );
  NANDN U18341 ( .A(n18027), .B(n18026), .Z(n18031) );
  NAND U18342 ( .A(n18029), .B(n18028), .Z(n18030) );
  NAND U18343 ( .A(n18031), .B(n18030), .Z(n18233) );
  NANDN U18344 ( .A(n18037), .B(n18036), .Z(n18041) );
  OR U18345 ( .A(n18039), .B(n18038), .Z(n18040) );
  NAND U18346 ( .A(n18041), .B(n18040), .Z(n18226) );
  NANDN U18347 ( .A(n18043), .B(n18042), .Z(n18047) );
  NANDN U18348 ( .A(n18045), .B(n18044), .Z(n18046) );
  NAND U18349 ( .A(n18047), .B(n18046), .Z(n18227) );
  XNOR U18350 ( .A(n18226), .B(n18227), .Z(n18228) );
  XNOR U18351 ( .A(n18229), .B(n18228), .Z(n18134) );
  NANDN U18352 ( .A(n18049), .B(n18048), .Z(n18053) );
  NAND U18353 ( .A(n18051), .B(n18050), .Z(n18052) );
  NAND U18354 ( .A(n18053), .B(n18052), .Z(n18140) );
  NANDN U18355 ( .A(n18055), .B(n18054), .Z(n18059) );
  NAND U18356 ( .A(n18057), .B(n18056), .Z(n18058) );
  NAND U18357 ( .A(n18059), .B(n18058), .Z(n18175) );
  XOR U18358 ( .A(b[25]), .B(a[113]), .Z(n18191) );
  NAND U18359 ( .A(n18191), .B(n19240), .Z(n18062) );
  NANDN U18360 ( .A(n18060), .B(n19242), .Z(n18061) );
  NAND U18361 ( .A(n18062), .B(n18061), .Z(n18205) );
  XNOR U18362 ( .A(b[27]), .B(a[111]), .Z(n18208) );
  NANDN U18363 ( .A(n18208), .B(n19336), .Z(n18065) );
  NANDN U18364 ( .A(n18063), .B(n19337), .Z(n18064) );
  NAND U18365 ( .A(n18065), .B(n18064), .Z(n18202) );
  NANDN U18366 ( .A(n18066), .B(n18832), .Z(n18068) );
  XOR U18367 ( .A(n19239), .B(n581), .Z(n18185) );
  NAND U18368 ( .A(n18185), .B(n18834), .Z(n18067) );
  AND U18369 ( .A(n18068), .B(n18067), .Z(n18203) );
  XNOR U18370 ( .A(n18202), .B(n18203), .Z(n18204) );
  XNOR U18371 ( .A(n18205), .B(n18204), .Z(n18173) );
  NANDN U18372 ( .A(n585), .B(a[105]), .Z(n18150) );
  XNOR U18373 ( .A(n18149), .B(n18150), .Z(n18152) );
  XNOR U18374 ( .A(n18151), .B(n18152), .Z(n18179) );
  XOR U18375 ( .A(n585), .B(a[107]), .Z(n18199) );
  NANDN U18376 ( .A(n18199), .B(n19472), .Z(n18071) );
  NANDN U18377 ( .A(n18069), .B(n19473), .Z(n18070) );
  NAND U18378 ( .A(n18071), .B(n18070), .Z(n18180) );
  XOR U18379 ( .A(n18179), .B(n18180), .Z(n18181) );
  XOR U18380 ( .A(n582), .B(a[117]), .Z(n18188) );
  NANDN U18381 ( .A(n18188), .B(n19015), .Z(n18074) );
  NAND U18382 ( .A(n19013), .B(n18072), .Z(n18073) );
  AND U18383 ( .A(n18074), .B(n18073), .Z(n18182) );
  XNOR U18384 ( .A(n18181), .B(n18182), .Z(n18174) );
  XOR U18385 ( .A(n18173), .B(n18174), .Z(n18176) );
  XOR U18386 ( .A(n18175), .B(n18176), .Z(n18145) );
  NANDN U18387 ( .A(n18075), .B(n18151), .Z(n18079) );
  OR U18388 ( .A(n18077), .B(n18076), .Z(n18078) );
  NAND U18389 ( .A(n18079), .B(n18078), .Z(n18143) );
  NANDN U18390 ( .A(n18081), .B(n18080), .Z(n18085) );
  NAND U18391 ( .A(n18083), .B(n18082), .Z(n18084) );
  NAND U18392 ( .A(n18085), .B(n18084), .Z(n18144) );
  XNOR U18393 ( .A(n18143), .B(n18144), .Z(n18146) );
  XOR U18394 ( .A(n18145), .B(n18146), .Z(n18137) );
  NANDN U18395 ( .A(n18087), .B(n18086), .Z(n18091) );
  NAND U18396 ( .A(n18089), .B(n18088), .Z(n18090) );
  NAND U18397 ( .A(n18091), .B(n18090), .Z(n18169) );
  NANDN U18398 ( .A(n18092), .B(n19406), .Z(n18094) );
  XNOR U18399 ( .A(n584), .B(a[109]), .Z(n18211) );
  NANDN U18400 ( .A(n576), .B(n18211), .Z(n18093) );
  NAND U18401 ( .A(n18094), .B(n18093), .Z(n18164) );
  XNOR U18402 ( .A(a[121]), .B(b[17]), .Z(n18214) );
  NANDN U18403 ( .A(n18214), .B(n18673), .Z(n18097) );
  NANDN U18404 ( .A(n18095), .B(n18674), .Z(n18096) );
  NAND U18405 ( .A(n18097), .B(n18096), .Z(n18161) );
  NANDN U18406 ( .A(n18098), .B(n18513), .Z(n18100) );
  XOR U18407 ( .A(a[123]), .B(b[15]), .Z(n18220) );
  NANDN U18408 ( .A(n18512), .B(n18220), .Z(n18099) );
  AND U18409 ( .A(n18100), .B(n18099), .Z(n18162) );
  XNOR U18410 ( .A(n18161), .B(n18162), .Z(n18163) );
  XNOR U18411 ( .A(n18164), .B(n18163), .Z(n18167) );
  XOR U18412 ( .A(a[125]), .B(n580), .Z(n18223) );
  NANDN U18413 ( .A(n18223), .B(n18336), .Z(n18103) );
  NANDN U18414 ( .A(n18101), .B(n18337), .Z(n18102) );
  NAND U18415 ( .A(n18103), .B(n18102), .Z(n18158) );
  XNOR U18416 ( .A(n19502), .B(b[11]), .Z(n18195) );
  NANDN U18417 ( .A(n18194), .B(n18195), .Z(n18107) );
  NAND U18418 ( .A(n18105), .B(n18104), .Z(n18106) );
  NAND U18419 ( .A(n18107), .B(n18106), .Z(n18155) );
  XNOR U18420 ( .A(b[23]), .B(a[115]), .Z(n18217) );
  OR U18421 ( .A(n18217), .B(n19127), .Z(n18110) );
  NANDN U18422 ( .A(n18108), .B(n19128), .Z(n18109) );
  AND U18423 ( .A(n18110), .B(n18109), .Z(n18156) );
  XNOR U18424 ( .A(n18155), .B(n18156), .Z(n18157) );
  XOR U18425 ( .A(n18158), .B(n18157), .Z(n18168) );
  XOR U18426 ( .A(n18167), .B(n18168), .Z(n18170) );
  XOR U18427 ( .A(n18169), .B(n18170), .Z(n18138) );
  XOR U18428 ( .A(n18137), .B(n18138), .Z(n18139) );
  XOR U18429 ( .A(n18140), .B(n18139), .Z(n18131) );
  NANDN U18430 ( .A(n18112), .B(n18111), .Z(n18116) );
  NAND U18431 ( .A(n18114), .B(n18113), .Z(n18115) );
  AND U18432 ( .A(n18116), .B(n18115), .Z(n18132) );
  XNOR U18433 ( .A(n18131), .B(n18132), .Z(n18133) );
  XOR U18434 ( .A(n18134), .B(n18133), .Z(n18232) );
  XOR U18435 ( .A(n18233), .B(n18232), .Z(n18234) );
  XOR U18436 ( .A(n18235), .B(n18234), .Z(n18126) );
  IV U18437 ( .A(n18126), .Z(n18124) );
  NANDN U18438 ( .A(n18118), .B(n18117), .Z(n18122) );
  NANDN U18439 ( .A(n18120), .B(n18119), .Z(n18121) );
  AND U18440 ( .A(n18122), .B(n18121), .Z(n18125) );
  XOR U18441 ( .A(n18124), .B(n18125), .Z(n18123) );
  XNOR U18442 ( .A(n18128), .B(n18123), .Z(n18238) );
  XOR U18443 ( .A(n18239), .B(n18238), .Z(c[233]) );
  NANDN U18444 ( .A(n18124), .B(n18125), .Z(n18130) );
  NOR U18445 ( .A(n18126), .B(n18125), .Z(n18127) );
  OR U18446 ( .A(n18128), .B(n18127), .Z(n18129) );
  NAND U18447 ( .A(n18130), .B(n18129), .Z(n18242) );
  NANDN U18448 ( .A(n18132), .B(n18131), .Z(n18136) );
  NAND U18449 ( .A(n18134), .B(n18133), .Z(n18135) );
  NAND U18450 ( .A(n18136), .B(n18135), .Z(n18249) );
  NAND U18451 ( .A(n18138), .B(n18137), .Z(n18142) );
  NANDN U18452 ( .A(n18140), .B(n18139), .Z(n18141) );
  NAND U18453 ( .A(n18142), .B(n18141), .Z(n18254) );
  NANDN U18454 ( .A(n18144), .B(n18143), .Z(n18148) );
  NAND U18455 ( .A(n18146), .B(n18145), .Z(n18147) );
  NAND U18456 ( .A(n18148), .B(n18147), .Z(n18253) );
  OR U18457 ( .A(n18150), .B(n18149), .Z(n18154) );
  NANDN U18458 ( .A(n18152), .B(n18151), .Z(n18153) );
  NAND U18459 ( .A(n18154), .B(n18153), .Z(n18273) );
  NANDN U18460 ( .A(n18156), .B(n18155), .Z(n18160) );
  NAND U18461 ( .A(n18158), .B(n18157), .Z(n18159) );
  NAND U18462 ( .A(n18160), .B(n18159), .Z(n18271) );
  NANDN U18463 ( .A(n18162), .B(n18161), .Z(n18166) );
  NAND U18464 ( .A(n18164), .B(n18163), .Z(n18165) );
  AND U18465 ( .A(n18166), .B(n18165), .Z(n18270) );
  XNOR U18466 ( .A(n18271), .B(n18270), .Z(n18272) );
  XOR U18467 ( .A(n18273), .B(n18272), .Z(n18258) );
  NANDN U18468 ( .A(n18168), .B(n18167), .Z(n18172) );
  OR U18469 ( .A(n18170), .B(n18169), .Z(n18171) );
  NAND U18470 ( .A(n18172), .B(n18171), .Z(n18259) );
  XNOR U18471 ( .A(n18258), .B(n18259), .Z(n18260) );
  NANDN U18472 ( .A(n18174), .B(n18173), .Z(n18178) );
  OR U18473 ( .A(n18176), .B(n18175), .Z(n18177) );
  NAND U18474 ( .A(n18178), .B(n18177), .Z(n18267) );
  OR U18475 ( .A(n18180), .B(n18179), .Z(n18184) );
  NAND U18476 ( .A(n18182), .B(n18181), .Z(n18183) );
  NAND U18477 ( .A(n18184), .B(n18183), .Z(n18282) );
  XOR U18478 ( .A(a[120]), .B(n581), .Z(n18312) );
  NANDN U18479 ( .A(n18312), .B(n18834), .Z(n18187) );
  NAND U18480 ( .A(n18832), .B(n18185), .Z(n18186) );
  NAND U18481 ( .A(n18187), .B(n18186), .Z(n18295) );
  XOR U18482 ( .A(b[21]), .B(n19077), .Z(n18341) );
  NANDN U18483 ( .A(n18341), .B(n19015), .Z(n18190) );
  NANDN U18484 ( .A(n18188), .B(n19013), .Z(n18189) );
  AND U18485 ( .A(n18190), .B(n18189), .Z(n18294) );
  XNOR U18486 ( .A(n18295), .B(n18294), .Z(n18296) );
  XOR U18487 ( .A(b[25]), .B(n18751), .Z(n18306) );
  NANDN U18488 ( .A(n18306), .B(n19240), .Z(n18193) );
  NAND U18489 ( .A(n19242), .B(n18191), .Z(n18192) );
  AND U18490 ( .A(n18193), .B(n18192), .Z(n18297) );
  XNOR U18491 ( .A(n18296), .B(n18297), .Z(n18283) );
  XOR U18492 ( .A(n18282), .B(n18283), .Z(n18285) );
  NANDN U18493 ( .A(n579), .B(b[10]), .Z(n18332) );
  XNOR U18494 ( .A(b[11]), .B(n18332), .Z(n18197) );
  NANDN U18495 ( .A(n18195), .B(n18194), .Z(n18196) );
  AND U18496 ( .A(n18197), .B(n18196), .Z(n18321) );
  AND U18497 ( .A(a[106]), .B(b[31]), .Z(n18397) );
  XNOR U18498 ( .A(n18321), .B(n18397), .Z(n18322) );
  XOR U18499 ( .A(b[31]), .B(n18198), .Z(n18329) );
  NANDN U18500 ( .A(n18329), .B(n19472), .Z(n18201) );
  NANDN U18501 ( .A(n18199), .B(n19473), .Z(n18200) );
  AND U18502 ( .A(n18201), .B(n18200), .Z(n18323) );
  XNOR U18503 ( .A(n18322), .B(n18323), .Z(n18284) );
  XNOR U18504 ( .A(n18285), .B(n18284), .Z(n18264) );
  NANDN U18505 ( .A(n18203), .B(n18202), .Z(n18207) );
  NAND U18506 ( .A(n18205), .B(n18204), .Z(n18206) );
  NAND U18507 ( .A(n18207), .B(n18206), .Z(n18279) );
  XOR U18508 ( .A(n583), .B(n18582), .Z(n18309) );
  NAND U18509 ( .A(n19336), .B(n18309), .Z(n18210) );
  NANDN U18510 ( .A(n18208), .B(n19337), .Z(n18209) );
  NAND U18511 ( .A(n18210), .B(n18209), .Z(n18291) );
  NAND U18512 ( .A(n19406), .B(n18211), .Z(n18213) );
  XOR U18513 ( .A(n584), .B(n18415), .Z(n18333) );
  NANDN U18514 ( .A(n576), .B(n18333), .Z(n18212) );
  NAND U18515 ( .A(n18213), .B(n18212), .Z(n18288) );
  XNOR U18516 ( .A(a[122]), .B(b[17]), .Z(n18300) );
  NANDN U18517 ( .A(n18300), .B(n18673), .Z(n18216) );
  NANDN U18518 ( .A(n18214), .B(n18674), .Z(n18215) );
  AND U18519 ( .A(n18216), .B(n18215), .Z(n18289) );
  XNOR U18520 ( .A(n18288), .B(n18289), .Z(n18290) );
  XNOR U18521 ( .A(n18291), .B(n18290), .Z(n18276) );
  XNOR U18522 ( .A(b[23]), .B(a[116]), .Z(n18326) );
  OR U18523 ( .A(n18326), .B(n19127), .Z(n18219) );
  NANDN U18524 ( .A(n18217), .B(n19128), .Z(n18218) );
  NAND U18525 ( .A(n18219), .B(n18218), .Z(n18318) );
  NAND U18526 ( .A(n18220), .B(n18513), .Z(n18222) );
  XNOR U18527 ( .A(a[124]), .B(b[15]), .Z(n18303) );
  OR U18528 ( .A(n18303), .B(n18512), .Z(n18221) );
  NAND U18529 ( .A(n18222), .B(n18221), .Z(n18315) );
  XOR U18530 ( .A(a[126]), .B(n580), .Z(n18338) );
  NANDN U18531 ( .A(n18338), .B(n18336), .Z(n18225) );
  NANDN U18532 ( .A(n18223), .B(n18337), .Z(n18224) );
  AND U18533 ( .A(n18225), .B(n18224), .Z(n18316) );
  XNOR U18534 ( .A(n18315), .B(n18316), .Z(n18317) );
  XOR U18535 ( .A(n18318), .B(n18317), .Z(n18277) );
  XNOR U18536 ( .A(n18276), .B(n18277), .Z(n18278) );
  XNOR U18537 ( .A(n18279), .B(n18278), .Z(n18265) );
  XNOR U18538 ( .A(n18264), .B(n18265), .Z(n18266) );
  XOR U18539 ( .A(n18267), .B(n18266), .Z(n18261) );
  XNOR U18540 ( .A(n18260), .B(n18261), .Z(n18252) );
  XOR U18541 ( .A(n18253), .B(n18252), .Z(n18255) );
  XNOR U18542 ( .A(n18254), .B(n18255), .Z(n18246) );
  NANDN U18543 ( .A(n18227), .B(n18226), .Z(n18231) );
  NAND U18544 ( .A(n18229), .B(n18228), .Z(n18230) );
  AND U18545 ( .A(n18231), .B(n18230), .Z(n18247) );
  XNOR U18546 ( .A(n18246), .B(n18247), .Z(n18248) );
  XOR U18547 ( .A(n18249), .B(n18248), .Z(n18240) );
  NAND U18548 ( .A(n18233), .B(n18232), .Z(n18237) );
  NAND U18549 ( .A(n18235), .B(n18234), .Z(n18236) );
  AND U18550 ( .A(n18237), .B(n18236), .Z(n18241) );
  XNOR U18551 ( .A(n18240), .B(n18241), .Z(n18243) );
  XOR U18552 ( .A(n18242), .B(n18243), .Z(n18345) );
  OR U18553 ( .A(n18239), .B(n18238), .Z(n18346) );
  XNOR U18554 ( .A(n18345), .B(n18346), .Z(c[234]) );
  NANDN U18555 ( .A(n18241), .B(n18240), .Z(n18245) );
  NAND U18556 ( .A(n18243), .B(n18242), .Z(n18244) );
  NAND U18557 ( .A(n18245), .B(n18244), .Z(n18350) );
  NANDN U18558 ( .A(n18247), .B(n18246), .Z(n18251) );
  NANDN U18559 ( .A(n18249), .B(n18248), .Z(n18250) );
  NAND U18560 ( .A(n18251), .B(n18250), .Z(n18348) );
  NANDN U18561 ( .A(n18253), .B(n18252), .Z(n18257) );
  OR U18562 ( .A(n18255), .B(n18254), .Z(n18256) );
  NAND U18563 ( .A(n18257), .B(n18256), .Z(n18442) );
  NANDN U18564 ( .A(n18259), .B(n18258), .Z(n18263) );
  NANDN U18565 ( .A(n18261), .B(n18260), .Z(n18262) );
  NAND U18566 ( .A(n18263), .B(n18262), .Z(n18441) );
  NANDN U18567 ( .A(n18265), .B(n18264), .Z(n18269) );
  NANDN U18568 ( .A(n18267), .B(n18266), .Z(n18268) );
  NAND U18569 ( .A(n18269), .B(n18268), .Z(n18353) );
  NANDN U18570 ( .A(n18271), .B(n18270), .Z(n18275) );
  NANDN U18571 ( .A(n18273), .B(n18272), .Z(n18274) );
  NAND U18572 ( .A(n18275), .B(n18274), .Z(n18354) );
  XNOR U18573 ( .A(n18353), .B(n18354), .Z(n18355) );
  NANDN U18574 ( .A(n18277), .B(n18276), .Z(n18281) );
  NANDN U18575 ( .A(n18279), .B(n18278), .Z(n18280) );
  NAND U18576 ( .A(n18281), .B(n18280), .Z(n18435) );
  NANDN U18577 ( .A(n18283), .B(n18282), .Z(n18287) );
  OR U18578 ( .A(n18285), .B(n18284), .Z(n18286) );
  AND U18579 ( .A(n18287), .B(n18286), .Z(n18434) );
  XNOR U18580 ( .A(n18435), .B(n18434), .Z(n18436) );
  NANDN U18581 ( .A(n18289), .B(n18288), .Z(n18293) );
  NAND U18582 ( .A(n18291), .B(n18290), .Z(n18292) );
  NAND U18583 ( .A(n18293), .B(n18292), .Z(n18425) );
  NANDN U18584 ( .A(n18295), .B(n18294), .Z(n18299) );
  NAND U18585 ( .A(n18297), .B(n18296), .Z(n18298) );
  AND U18586 ( .A(n18299), .B(n18298), .Z(n18426) );
  XOR U18587 ( .A(a[123]), .B(b[17]), .Z(n18386) );
  NAND U18588 ( .A(n18386), .B(n18673), .Z(n18302) );
  NANDN U18589 ( .A(n18300), .B(n18674), .Z(n18301) );
  NAND U18590 ( .A(n18302), .B(n18301), .Z(n18361) );
  NANDN U18591 ( .A(n18303), .B(n18513), .Z(n18305) );
  XNOR U18592 ( .A(a[125]), .B(b[15]), .Z(n18389) );
  OR U18593 ( .A(n18389), .B(n18512), .Z(n18304) );
  NAND U18594 ( .A(n18305), .B(n18304), .Z(n18360) );
  XNOR U18595 ( .A(b[25]), .B(a[115]), .Z(n18392) );
  NANDN U18596 ( .A(n18392), .B(n19240), .Z(n18308) );
  NANDN U18597 ( .A(n18306), .B(n19242), .Z(n18307) );
  AND U18598 ( .A(n18308), .B(n18307), .Z(n18404) );
  XNOR U18599 ( .A(b[27]), .B(a[113]), .Z(n18377) );
  NANDN U18600 ( .A(n18377), .B(n19336), .Z(n18311) );
  NAND U18601 ( .A(n19337), .B(n18309), .Z(n18310) );
  NAND U18602 ( .A(n18311), .B(n18310), .Z(n18401) );
  NANDN U18603 ( .A(n18312), .B(n18832), .Z(n18314) );
  XOR U18604 ( .A(a[121]), .B(n581), .Z(n18371) );
  NANDN U18605 ( .A(n18371), .B(n18834), .Z(n18313) );
  AND U18606 ( .A(n18314), .B(n18313), .Z(n18402) );
  XNOR U18607 ( .A(n18401), .B(n18402), .Z(n18403) );
  XNOR U18608 ( .A(n18404), .B(n18403), .Z(n18359) );
  XNOR U18609 ( .A(n18360), .B(n18359), .Z(n18362) );
  XNOR U18610 ( .A(n18361), .B(n18362), .Z(n18431) );
  NANDN U18611 ( .A(n18316), .B(n18315), .Z(n18320) );
  NAND U18612 ( .A(n18318), .B(n18317), .Z(n18319) );
  NAND U18613 ( .A(n18320), .B(n18319), .Z(n18429) );
  NANDN U18614 ( .A(n18321), .B(n18397), .Z(n18325) );
  NAND U18615 ( .A(n18323), .B(n18322), .Z(n18324) );
  NAND U18616 ( .A(n18325), .B(n18324), .Z(n18421) );
  XNOR U18617 ( .A(b[23]), .B(a[117]), .Z(n18383) );
  OR U18618 ( .A(n18383), .B(n19127), .Z(n18328) );
  NANDN U18619 ( .A(n18326), .B(n19128), .Z(n18327) );
  NAND U18620 ( .A(n18328), .B(n18327), .Z(n18408) );
  XNOR U18621 ( .A(b[31]), .B(a[109]), .Z(n18416) );
  NANDN U18622 ( .A(n18416), .B(n19472), .Z(n18331) );
  NANDN U18623 ( .A(n18329), .B(n19473), .Z(n18330) );
  NAND U18624 ( .A(n18331), .B(n18330), .Z(n18405) );
  AND U18625 ( .A(n18332), .B(b[11]), .Z(n18396) );
  NANDN U18626 ( .A(n585), .B(a[107]), .Z(n18395) );
  XOR U18627 ( .A(n18396), .B(n18395), .Z(n18398) );
  XNOR U18628 ( .A(n18397), .B(n18398), .Z(n18406) );
  XNOR U18629 ( .A(n18405), .B(n18406), .Z(n18407) );
  XNOR U18630 ( .A(n18408), .B(n18407), .Z(n18420) );
  NAND U18631 ( .A(n19406), .B(n18333), .Z(n18335) );
  XNOR U18632 ( .A(n584), .B(a[111]), .Z(n18380) );
  NANDN U18633 ( .A(n576), .B(n18380), .Z(n18334) );
  NAND U18634 ( .A(n18335), .B(n18334), .Z(n18368) );
  XNOR U18635 ( .A(n19502), .B(b[13]), .Z(n18412) );
  NAND U18636 ( .A(n18412), .B(n18336), .Z(n18340) );
  NANDN U18637 ( .A(n18338), .B(n18337), .Z(n18339) );
  NAND U18638 ( .A(n18340), .B(n18339), .Z(n18365) );
  NANDN U18639 ( .A(n18341), .B(n19013), .Z(n18343) );
  XOR U18640 ( .A(b[21]), .B(n19239), .Z(n18374) );
  NANDN U18641 ( .A(n18374), .B(n19015), .Z(n18342) );
  AND U18642 ( .A(n18343), .B(n18342), .Z(n18366) );
  XNOR U18643 ( .A(n18365), .B(n18366), .Z(n18367) );
  XOR U18644 ( .A(n18368), .B(n18367), .Z(n18419) );
  XOR U18645 ( .A(n18420), .B(n18419), .Z(n18422) );
  XOR U18646 ( .A(n18421), .B(n18422), .Z(n18428) );
  XNOR U18647 ( .A(n18429), .B(n18428), .Z(n18430) );
  XOR U18648 ( .A(n18431), .B(n18430), .Z(n18427) );
  XNOR U18649 ( .A(n18426), .B(n18427), .Z(n18344) );
  XNOR U18650 ( .A(n18425), .B(n18344), .Z(n18437) );
  XOR U18651 ( .A(n18436), .B(n18437), .Z(n18356) );
  XNOR U18652 ( .A(n18355), .B(n18356), .Z(n18440) );
  XNOR U18653 ( .A(n18441), .B(n18440), .Z(n18443) );
  XNOR U18654 ( .A(n18442), .B(n18443), .Z(n18347) );
  XNOR U18655 ( .A(n18348), .B(n18347), .Z(n18349) );
  XNOR U18656 ( .A(n18350), .B(n18349), .Z(n18447) );
  NANDN U18657 ( .A(n18346), .B(n18345), .Z(n18446) );
  XOR U18658 ( .A(n18447), .B(n18446), .Z(c[235]) );
  NANDN U18659 ( .A(n18348), .B(n18347), .Z(n18352) );
  NAND U18660 ( .A(n18350), .B(n18349), .Z(n18351) );
  NAND U18661 ( .A(n18352), .B(n18351), .Z(n18453) );
  NANDN U18662 ( .A(n18354), .B(n18353), .Z(n18358) );
  NANDN U18663 ( .A(n18356), .B(n18355), .Z(n18357) );
  NAND U18664 ( .A(n18358), .B(n18357), .Z(n18536) );
  NAND U18665 ( .A(n18360), .B(n18359), .Z(n18364) );
  NANDN U18666 ( .A(n18362), .B(n18361), .Z(n18363) );
  NAND U18667 ( .A(n18364), .B(n18363), .Z(n18468) );
  NANDN U18668 ( .A(n18366), .B(n18365), .Z(n18370) );
  NAND U18669 ( .A(n18368), .B(n18367), .Z(n18369) );
  NAND U18670 ( .A(n18370), .B(n18369), .Z(n18467) );
  NANDN U18671 ( .A(n18371), .B(n18832), .Z(n18373) );
  XOR U18672 ( .A(a[122]), .B(n581), .Z(n18493) );
  NANDN U18673 ( .A(n18493), .B(n18834), .Z(n18372) );
  NAND U18674 ( .A(n18373), .B(n18372), .Z(n18502) );
  NANDN U18675 ( .A(n18374), .B(n19013), .Z(n18376) );
  XOR U18676 ( .A(n19188), .B(n582), .Z(n18496) );
  NAND U18677 ( .A(n18496), .B(n19015), .Z(n18375) );
  NAND U18678 ( .A(n18376), .B(n18375), .Z(n18499) );
  XOR U18679 ( .A(b[27]), .B(n18751), .Z(n18487) );
  NANDN U18680 ( .A(n18487), .B(n19336), .Z(n18379) );
  NANDN U18681 ( .A(n18377), .B(n19337), .Z(n18378) );
  NAND U18682 ( .A(n18379), .B(n18378), .Z(n18508) );
  NAND U18683 ( .A(n19406), .B(n18380), .Z(n18382) );
  XOR U18684 ( .A(n584), .B(n18582), .Z(n18490) );
  NANDN U18685 ( .A(n576), .B(n18490), .Z(n18381) );
  AND U18686 ( .A(n18382), .B(n18381), .Z(n18505) );
  XNOR U18687 ( .A(b[23]), .B(a[118]), .Z(n18478) );
  OR U18688 ( .A(n18478), .B(n19127), .Z(n18385) );
  NANDN U18689 ( .A(n18383), .B(n19128), .Z(n18384) );
  AND U18690 ( .A(n18385), .B(n18384), .Z(n18506) );
  XNOR U18691 ( .A(n18508), .B(n18507), .Z(n18500) );
  XNOR U18692 ( .A(n18499), .B(n18500), .Z(n18501) );
  XNOR U18693 ( .A(n18502), .B(n18501), .Z(n18528) );
  XNOR U18694 ( .A(a[124]), .B(b[17]), .Z(n18481) );
  NANDN U18695 ( .A(n18481), .B(n18673), .Z(n18388) );
  NAND U18696 ( .A(n18386), .B(n18674), .Z(n18387) );
  NAND U18697 ( .A(n18388), .B(n18387), .Z(n18475) );
  NANDN U18698 ( .A(n18389), .B(n18513), .Z(n18391) );
  XNOR U18699 ( .A(a[126]), .B(b[15]), .Z(n18514) );
  OR U18700 ( .A(n18514), .B(n18512), .Z(n18390) );
  NAND U18701 ( .A(n18391), .B(n18390), .Z(n18472) );
  XNOR U18702 ( .A(b[25]), .B(n18950), .Z(n18517) );
  NAND U18703 ( .A(n18517), .B(n19240), .Z(n18394) );
  NANDN U18704 ( .A(n18392), .B(n19242), .Z(n18393) );
  AND U18705 ( .A(n18394), .B(n18393), .Z(n18473) );
  XNOR U18706 ( .A(n18472), .B(n18473), .Z(n18474) );
  XNOR U18707 ( .A(n18475), .B(n18474), .Z(n18525) );
  OR U18708 ( .A(n18396), .B(n18395), .Z(n18400) );
  NAND U18709 ( .A(n18398), .B(n18397), .Z(n18399) );
  NAND U18710 ( .A(n18400), .B(n18399), .Z(n18526) );
  XNOR U18711 ( .A(n18525), .B(n18526), .Z(n18527) );
  XOR U18712 ( .A(n18528), .B(n18527), .Z(n18466) );
  XOR U18713 ( .A(n18467), .B(n18466), .Z(n18469) );
  XOR U18714 ( .A(n18468), .B(n18469), .Z(n18531) );
  NANDN U18715 ( .A(n18406), .B(n18405), .Z(n18410) );
  NAND U18716 ( .A(n18408), .B(n18407), .Z(n18409) );
  AND U18717 ( .A(n18410), .B(n18409), .Z(n18461) );
  XNOR U18718 ( .A(n18460), .B(n18461), .Z(n18462) );
  NAND U18719 ( .A(b[11]), .B(b[12]), .Z(n18511) );
  XOR U18720 ( .A(n580), .B(n18511), .Z(n18414) );
  XNOR U18721 ( .A(b[12]), .B(b[11]), .Z(n18411) );
  NANDN U18722 ( .A(n18412), .B(n18411), .Z(n18413) );
  AND U18723 ( .A(n18414), .B(n18413), .Z(n18521) );
  AND U18724 ( .A(a[108]), .B(b[31]), .Z(n18567) );
  XOR U18725 ( .A(b[31]), .B(n18415), .Z(n18484) );
  NANDN U18726 ( .A(n18484), .B(n19472), .Z(n18418) );
  NANDN U18727 ( .A(n18416), .B(n19473), .Z(n18417) );
  AND U18728 ( .A(n18418), .B(n18417), .Z(n18520) );
  XOR U18729 ( .A(n18567), .B(n18520), .Z(n18522) );
  XOR U18730 ( .A(n18521), .B(n18522), .Z(n18463) );
  XNOR U18731 ( .A(n18462), .B(n18463), .Z(n18529) );
  NANDN U18732 ( .A(n18420), .B(n18419), .Z(n18424) );
  OR U18733 ( .A(n18422), .B(n18421), .Z(n18423) );
  NAND U18734 ( .A(n18424), .B(n18423), .Z(n18530) );
  XNOR U18735 ( .A(n18529), .B(n18530), .Z(n18532) );
  XNOR U18736 ( .A(n18531), .B(n18532), .Z(n18458) );
  OR U18737 ( .A(n18429), .B(n18428), .Z(n18433) );
  OR U18738 ( .A(n18431), .B(n18430), .Z(n18432) );
  AND U18739 ( .A(n18433), .B(n18432), .Z(n18456) );
  XNOR U18740 ( .A(n18457), .B(n18456), .Z(n18459) );
  XNOR U18741 ( .A(n18458), .B(n18459), .Z(n18533) );
  NANDN U18742 ( .A(n18435), .B(n18434), .Z(n18439) );
  NANDN U18743 ( .A(n18437), .B(n18436), .Z(n18438) );
  NAND U18744 ( .A(n18439), .B(n18438), .Z(n18534) );
  XNOR U18745 ( .A(n18533), .B(n18534), .Z(n18535) );
  XOR U18746 ( .A(n18536), .B(n18535), .Z(n18450) );
  NAND U18747 ( .A(n18441), .B(n18440), .Z(n18445) );
  NANDN U18748 ( .A(n18443), .B(n18442), .Z(n18444) );
  AND U18749 ( .A(n18445), .B(n18444), .Z(n18451) );
  XNOR U18750 ( .A(n18450), .B(n18451), .Z(n18452) );
  XNOR U18751 ( .A(n18453), .B(n18452), .Z(n18449) );
  OR U18752 ( .A(n18447), .B(n18446), .Z(n18448) );
  XOR U18753 ( .A(n18449), .B(n18448), .Z(c[236]) );
  OR U18754 ( .A(n18449), .B(n18448), .Z(n18632) );
  NANDN U18755 ( .A(n18451), .B(n18450), .Z(n18455) );
  NAND U18756 ( .A(n18453), .B(n18452), .Z(n18454) );
  NAND U18757 ( .A(n18455), .B(n18454), .Z(n18542) );
  NANDN U18758 ( .A(n18461), .B(n18460), .Z(n18465) );
  NAND U18759 ( .A(n18463), .B(n18462), .Z(n18464) );
  NAND U18760 ( .A(n18465), .B(n18464), .Z(n18543) );
  NANDN U18761 ( .A(n18467), .B(n18466), .Z(n18471) );
  OR U18762 ( .A(n18469), .B(n18468), .Z(n18470) );
  NAND U18763 ( .A(n18471), .B(n18470), .Z(n18544) );
  XNOR U18764 ( .A(n18543), .B(n18544), .Z(n18545) );
  NANDN U18765 ( .A(n18473), .B(n18472), .Z(n18477) );
  NAND U18766 ( .A(n18475), .B(n18474), .Z(n18476) );
  NAND U18767 ( .A(n18477), .B(n18476), .Z(n18556) );
  XNOR U18768 ( .A(b[23]), .B(a[119]), .Z(n18598) );
  OR U18769 ( .A(n18598), .B(n19127), .Z(n18480) );
  NANDN U18770 ( .A(n18478), .B(n19128), .Z(n18479) );
  NAND U18771 ( .A(n18480), .B(n18479), .Z(n18610) );
  XNOR U18772 ( .A(a[125]), .B(b[17]), .Z(n18601) );
  NANDN U18773 ( .A(n18601), .B(n18673), .Z(n18483) );
  NANDN U18774 ( .A(n18481), .B(n18674), .Z(n18482) );
  NAND U18775 ( .A(n18483), .B(n18482), .Z(n18607) );
  XNOR U18776 ( .A(b[31]), .B(a[111]), .Z(n18583) );
  NANDN U18777 ( .A(n18583), .B(n19472), .Z(n18486) );
  NANDN U18778 ( .A(n18484), .B(n19473), .Z(n18485) );
  AND U18779 ( .A(n18486), .B(n18485), .Z(n18608) );
  XNOR U18780 ( .A(n18607), .B(n18608), .Z(n18609) );
  XNOR U18781 ( .A(n18610), .B(n18609), .Z(n18564) );
  XOR U18782 ( .A(b[27]), .B(n19022), .Z(n18586) );
  NANDN U18783 ( .A(n18586), .B(n19336), .Z(n18489) );
  NANDN U18784 ( .A(n18487), .B(n19337), .Z(n18488) );
  NAND U18785 ( .A(n18489), .B(n18488), .Z(n18616) );
  NAND U18786 ( .A(n19406), .B(n18490), .Z(n18492) );
  XNOR U18787 ( .A(n584), .B(a[113]), .Z(n18589) );
  NANDN U18788 ( .A(n576), .B(n18589), .Z(n18491) );
  NAND U18789 ( .A(n18492), .B(n18491), .Z(n18613) );
  NANDN U18790 ( .A(n18493), .B(n18832), .Z(n18495) );
  XNOR U18791 ( .A(a[123]), .B(n581), .Z(n18604) );
  NAND U18792 ( .A(n18604), .B(n18834), .Z(n18494) );
  AND U18793 ( .A(n18495), .B(n18494), .Z(n18614) );
  XNOR U18794 ( .A(n18613), .B(n18614), .Z(n18615) );
  XNOR U18795 ( .A(n18616), .B(n18615), .Z(n18561) );
  XOR U18796 ( .A(a[121]), .B(n582), .Z(n18595) );
  NANDN U18797 ( .A(n18595), .B(n19015), .Z(n18498) );
  NAND U18798 ( .A(n19013), .B(n18496), .Z(n18497) );
  NAND U18799 ( .A(n18498), .B(n18497), .Z(n18562) );
  XNOR U18800 ( .A(n18561), .B(n18562), .Z(n18563) );
  XOR U18801 ( .A(n18564), .B(n18563), .Z(n18555) );
  XOR U18802 ( .A(n18556), .B(n18555), .Z(n18558) );
  NANDN U18803 ( .A(n18500), .B(n18499), .Z(n18504) );
  NAND U18804 ( .A(n18502), .B(n18501), .Z(n18503) );
  NAND U18805 ( .A(n18504), .B(n18503), .Z(n18557) );
  XNOR U18806 ( .A(n18558), .B(n18557), .Z(n18622) );
  OR U18807 ( .A(n18506), .B(n18505), .Z(n18510) );
  NAND U18808 ( .A(n18508), .B(n18507), .Z(n18509) );
  NAND U18809 ( .A(n18510), .B(n18509), .Z(n18550) );
  NAND U18810 ( .A(b[13]), .B(n18511), .Z(n18565) );
  NANDN U18811 ( .A(n585), .B(a[109]), .Z(n18566) );
  XOR U18812 ( .A(n18565), .B(n18566), .Z(n18568) );
  XNOR U18813 ( .A(n18567), .B(n18568), .Z(n18571) );
  XNOR U18814 ( .A(a[127]), .B(b[15]), .Z(n18578) );
  OR U18815 ( .A(n18578), .B(n18512), .Z(n18516) );
  NANDN U18816 ( .A(n18514), .B(n18513), .Z(n18515) );
  NAND U18817 ( .A(n18516), .B(n18515), .Z(n18572) );
  XOR U18818 ( .A(n18571), .B(n18572), .Z(n18573) );
  XNOR U18819 ( .A(b[25]), .B(a[117]), .Z(n18592) );
  NANDN U18820 ( .A(n18592), .B(n19240), .Z(n18519) );
  NAND U18821 ( .A(n19242), .B(n18517), .Z(n18518) );
  AND U18822 ( .A(n18519), .B(n18518), .Z(n18574) );
  XOR U18823 ( .A(n18573), .B(n18574), .Z(n18549) );
  XOR U18824 ( .A(n18550), .B(n18549), .Z(n18552) );
  OR U18825 ( .A(n18567), .B(n18520), .Z(n18524) );
  NAND U18826 ( .A(n18522), .B(n18521), .Z(n18523) );
  NAND U18827 ( .A(n18524), .B(n18523), .Z(n18551) );
  XNOR U18828 ( .A(n18552), .B(n18551), .Z(n18619) );
  XNOR U18829 ( .A(n18619), .B(n18620), .Z(n18621) );
  XNOR U18830 ( .A(n18622), .B(n18621), .Z(n18546) );
  XOR U18831 ( .A(n18545), .B(n18546), .Z(n18625) );
  XNOR U18832 ( .A(n18625), .B(n18626), .Z(n18627) );
  XOR U18833 ( .A(n18628), .B(n18627), .Z(n18540) );
  NANDN U18834 ( .A(n18534), .B(n18533), .Z(n18538) );
  NANDN U18835 ( .A(n18536), .B(n18535), .Z(n18537) );
  AND U18836 ( .A(n18538), .B(n18537), .Z(n18541) );
  XOR U18837 ( .A(n18540), .B(n18541), .Z(n18539) );
  XOR U18838 ( .A(n18542), .B(n18539), .Z(n18631) );
  XNOR U18839 ( .A(n18632), .B(n18631), .Z(c[237]) );
  NANDN U18840 ( .A(n18544), .B(n18543), .Z(n18548) );
  NANDN U18841 ( .A(n18546), .B(n18545), .Z(n18547) );
  NAND U18842 ( .A(n18548), .B(n18547), .Z(n18713) );
  NANDN U18843 ( .A(n18550), .B(n18549), .Z(n18554) );
  OR U18844 ( .A(n18552), .B(n18551), .Z(n18553) );
  NAND U18845 ( .A(n18554), .B(n18553), .Z(n18640) );
  NANDN U18846 ( .A(n18556), .B(n18555), .Z(n18560) );
  OR U18847 ( .A(n18558), .B(n18557), .Z(n18559) );
  AND U18848 ( .A(n18560), .B(n18559), .Z(n18639) );
  XNOR U18849 ( .A(n18640), .B(n18639), .Z(n18641) );
  NANDN U18850 ( .A(n18566), .B(n18565), .Z(n18570) );
  NANDN U18851 ( .A(n18568), .B(n18567), .Z(n18569) );
  NAND U18852 ( .A(n18570), .B(n18569), .Z(n18649) );
  OR U18853 ( .A(n18572), .B(n18571), .Z(n18576) );
  NAND U18854 ( .A(n18574), .B(n18573), .Z(n18575) );
  NAND U18855 ( .A(n18576), .B(n18575), .Z(n18650) );
  XNOR U18856 ( .A(n18649), .B(n18650), .Z(n18651) );
  XNOR U18857 ( .A(b[15]), .B(n18577), .Z(n18581) );
  XOR U18858 ( .A(b[14]), .B(n580), .Z(n18579) );
  NAND U18859 ( .A(n18579), .B(n18578), .Z(n18580) );
  AND U18860 ( .A(n18581), .B(n18580), .Z(n18700) );
  AND U18861 ( .A(a[110]), .B(b[31]), .Z(n18769) );
  XOR U18862 ( .A(b[31]), .B(n18582), .Z(n18684) );
  NANDN U18863 ( .A(n18684), .B(n19472), .Z(n18585) );
  NANDN U18864 ( .A(n18583), .B(n19473), .Z(n18584) );
  AND U18865 ( .A(n18585), .B(n18584), .Z(n18699) );
  XOR U18866 ( .A(n18769), .B(n18699), .Z(n18701) );
  XOR U18867 ( .A(n18700), .B(n18701), .Z(n18652) );
  XOR U18868 ( .A(n18651), .B(n18652), .Z(n18645) );
  XNOR U18869 ( .A(n18646), .B(n18645), .Z(n18647) );
  XOR U18870 ( .A(b[27]), .B(n18950), .Z(n18690) );
  NANDN U18871 ( .A(n18690), .B(n19336), .Z(n18588) );
  NANDN U18872 ( .A(n18586), .B(n19337), .Z(n18587) );
  NAND U18873 ( .A(n18588), .B(n18587), .Z(n18681) );
  NAND U18874 ( .A(n19406), .B(n18589), .Z(n18591) );
  XOR U18875 ( .A(n584), .B(n18751), .Z(n18693) );
  NANDN U18876 ( .A(n576), .B(n18693), .Z(n18590) );
  NAND U18877 ( .A(n18591), .B(n18590), .Z(n18678) );
  XNOR U18878 ( .A(b[25]), .B(a[118]), .Z(n18687) );
  NANDN U18879 ( .A(n18687), .B(n19240), .Z(n18594) );
  NANDN U18880 ( .A(n18592), .B(n19242), .Z(n18593) );
  AND U18881 ( .A(n18594), .B(n18593), .Z(n18679) );
  XNOR U18882 ( .A(n18678), .B(n18679), .Z(n18680) );
  XNOR U18883 ( .A(n18681), .B(n18680), .Z(n18707) );
  NANDN U18884 ( .A(n18595), .B(n19013), .Z(n18597) );
  XOR U18885 ( .A(a[122]), .B(n582), .Z(n18696) );
  NANDN U18886 ( .A(n18696), .B(n19015), .Z(n18596) );
  NAND U18887 ( .A(n18597), .B(n18596), .Z(n18664) );
  XNOR U18888 ( .A(b[23]), .B(a[120]), .Z(n18667) );
  OR U18889 ( .A(n18667), .B(n19127), .Z(n18600) );
  NANDN U18890 ( .A(n18598), .B(n19128), .Z(n18599) );
  NAND U18891 ( .A(n18600), .B(n18599), .Z(n18661) );
  XNOR U18892 ( .A(a[126]), .B(b[17]), .Z(n18675) );
  NANDN U18893 ( .A(n18675), .B(n18673), .Z(n18603) );
  NANDN U18894 ( .A(n18601), .B(n18674), .Z(n18602) );
  AND U18895 ( .A(n18603), .B(n18602), .Z(n18662) );
  XNOR U18896 ( .A(n18661), .B(n18662), .Z(n18663) );
  XNOR U18897 ( .A(n18664), .B(n18663), .Z(n18704) );
  XOR U18898 ( .A(a[124]), .B(n581), .Z(n18670) );
  NANDN U18899 ( .A(n18670), .B(n18834), .Z(n18606) );
  NAND U18900 ( .A(n18832), .B(n18604), .Z(n18605) );
  NAND U18901 ( .A(n18606), .B(n18605), .Z(n18705) );
  XNOR U18902 ( .A(n18704), .B(n18705), .Z(n18706) );
  XOR U18903 ( .A(n18707), .B(n18706), .Z(n18658) );
  NANDN U18904 ( .A(n18608), .B(n18607), .Z(n18612) );
  NAND U18905 ( .A(n18610), .B(n18609), .Z(n18611) );
  NAND U18906 ( .A(n18612), .B(n18611), .Z(n18655) );
  NANDN U18907 ( .A(n18614), .B(n18613), .Z(n18618) );
  NAND U18908 ( .A(n18616), .B(n18615), .Z(n18617) );
  AND U18909 ( .A(n18618), .B(n18617), .Z(n18656) );
  XNOR U18910 ( .A(n18655), .B(n18656), .Z(n18657) );
  XOR U18911 ( .A(n18658), .B(n18657), .Z(n18648) );
  XNOR U18912 ( .A(n18647), .B(n18648), .Z(n18642) );
  XNOR U18913 ( .A(n18641), .B(n18642), .Z(n18710) );
  NANDN U18914 ( .A(n18620), .B(n18619), .Z(n18624) );
  NAND U18915 ( .A(n18622), .B(n18621), .Z(n18623) );
  NAND U18916 ( .A(n18624), .B(n18623), .Z(n18711) );
  XNOR U18917 ( .A(n18710), .B(n18711), .Z(n18712) );
  XOR U18918 ( .A(n18713), .B(n18712), .Z(n18633) );
  NANDN U18919 ( .A(n18626), .B(n18625), .Z(n18630) );
  NANDN U18920 ( .A(n18628), .B(n18627), .Z(n18629) );
  NAND U18921 ( .A(n18630), .B(n18629), .Z(n18634) );
  XNOR U18922 ( .A(n18633), .B(n18634), .Z(n18636) );
  XOR U18923 ( .A(n18635), .B(n18636), .Z(n18714) );
  NANDN U18924 ( .A(n18632), .B(n18631), .Z(n18715) );
  XNOR U18925 ( .A(n18714), .B(n18715), .Z(c[238]) );
  NANDN U18926 ( .A(n18634), .B(n18633), .Z(n18638) );
  NAND U18927 ( .A(n18636), .B(n18635), .Z(n18637) );
  NAND U18928 ( .A(n18638), .B(n18637), .Z(n18718) );
  NANDN U18929 ( .A(n18640), .B(n18639), .Z(n18644) );
  NAND U18930 ( .A(n18642), .B(n18641), .Z(n18643) );
  NAND U18931 ( .A(n18644), .B(n18643), .Z(n18794) );
  NANDN U18932 ( .A(n18650), .B(n18649), .Z(n18654) );
  NAND U18933 ( .A(n18652), .B(n18651), .Z(n18653) );
  NAND U18934 ( .A(n18654), .B(n18653), .Z(n18722) );
  NANDN U18935 ( .A(n18656), .B(n18655), .Z(n18660) );
  NANDN U18936 ( .A(n18658), .B(n18657), .Z(n18659) );
  AND U18937 ( .A(n18660), .B(n18659), .Z(n18723) );
  XNOR U18938 ( .A(n18722), .B(n18723), .Z(n18724) );
  NANDN U18939 ( .A(n18662), .B(n18661), .Z(n18666) );
  NAND U18940 ( .A(n18664), .B(n18663), .Z(n18665) );
  NAND U18941 ( .A(n18666), .B(n18665), .Z(n18788) );
  XNOR U18942 ( .A(b[23]), .B(a[121]), .Z(n18779) );
  OR U18943 ( .A(n18779), .B(n19127), .Z(n18669) );
  NANDN U18944 ( .A(n18667), .B(n19128), .Z(n18668) );
  NAND U18945 ( .A(n18669), .B(n18668), .Z(n18735) );
  NANDN U18946 ( .A(n18670), .B(n18832), .Z(n18672) );
  XOR U18947 ( .A(a[125]), .B(n581), .Z(n18741) );
  NANDN U18948 ( .A(n18741), .B(n18834), .Z(n18671) );
  NAND U18949 ( .A(n18672), .B(n18671), .Z(n18732) );
  XNOR U18950 ( .A(n19502), .B(b[17]), .Z(n18748) );
  NAND U18951 ( .A(n18748), .B(n18673), .Z(n18677) );
  NANDN U18952 ( .A(n18675), .B(n18674), .Z(n18676) );
  AND U18953 ( .A(n18677), .B(n18676), .Z(n18733) );
  XNOR U18954 ( .A(n18732), .B(n18733), .Z(n18734) );
  XNOR U18955 ( .A(n18735), .B(n18734), .Z(n18786) );
  NANDN U18956 ( .A(n18679), .B(n18678), .Z(n18683) );
  NAND U18957 ( .A(n18681), .B(n18680), .Z(n18682) );
  NAND U18958 ( .A(n18683), .B(n18682), .Z(n18787) );
  XOR U18959 ( .A(n18786), .B(n18787), .Z(n18789) );
  XNOR U18960 ( .A(n18788), .B(n18789), .Z(n18731) );
  XNOR U18961 ( .A(b[31]), .B(a[113]), .Z(n18752) );
  NANDN U18962 ( .A(n18752), .B(n19472), .Z(n18686) );
  NANDN U18963 ( .A(n18684), .B(n19473), .Z(n18685) );
  NAND U18964 ( .A(n18686), .B(n18685), .Z(n18755) );
  XNOR U18965 ( .A(b[25]), .B(a[119]), .Z(n18773) );
  NANDN U18966 ( .A(n18773), .B(n19240), .Z(n18689) );
  NANDN U18967 ( .A(n18687), .B(n19242), .Z(n18688) );
  AND U18968 ( .A(n18689), .B(n18688), .Z(n18756) );
  XNOR U18969 ( .A(n18755), .B(n18756), .Z(n18757) );
  NANDN U18970 ( .A(n585), .B(a[111]), .Z(n18767) );
  XOR U18971 ( .A(n18768), .B(n18767), .Z(n18770) );
  XNOR U18972 ( .A(n18769), .B(n18770), .Z(n18758) );
  XOR U18973 ( .A(n18757), .B(n18758), .Z(n18785) );
  XOR U18974 ( .A(b[27]), .B(n19136), .Z(n18744) );
  NANDN U18975 ( .A(n18744), .B(n19336), .Z(n18692) );
  NANDN U18976 ( .A(n18690), .B(n19337), .Z(n18691) );
  NAND U18977 ( .A(n18692), .B(n18691), .Z(n18764) );
  NAND U18978 ( .A(n19406), .B(n18693), .Z(n18695) );
  XOR U18979 ( .A(n584), .B(n19022), .Z(n18776) );
  NANDN U18980 ( .A(n576), .B(n18776), .Z(n18694) );
  NAND U18981 ( .A(n18695), .B(n18694), .Z(n18761) );
  NANDN U18982 ( .A(n18696), .B(n19013), .Z(n18698) );
  XNOR U18983 ( .A(a[123]), .B(b[21]), .Z(n18738) );
  NANDN U18984 ( .A(n18738), .B(n19015), .Z(n18697) );
  AND U18985 ( .A(n18698), .B(n18697), .Z(n18762) );
  XNOR U18986 ( .A(n18761), .B(n18762), .Z(n18763) );
  XNOR U18987 ( .A(n18764), .B(n18763), .Z(n18782) );
  OR U18988 ( .A(n18769), .B(n18699), .Z(n18703) );
  NAND U18989 ( .A(n18701), .B(n18700), .Z(n18702) );
  NAND U18990 ( .A(n18703), .B(n18702), .Z(n18783) );
  XNOR U18991 ( .A(n18782), .B(n18783), .Z(n18784) );
  XNOR U18992 ( .A(n18785), .B(n18784), .Z(n18728) );
  NANDN U18993 ( .A(n18705), .B(n18704), .Z(n18709) );
  NAND U18994 ( .A(n18707), .B(n18706), .Z(n18708) );
  NAND U18995 ( .A(n18709), .B(n18708), .Z(n18729) );
  XNOR U18996 ( .A(n18728), .B(n18729), .Z(n18730) );
  XNOR U18997 ( .A(n18731), .B(n18730), .Z(n18725) );
  XNOR U18998 ( .A(n18724), .B(n18725), .Z(n18792) );
  XNOR U18999 ( .A(n18793), .B(n18792), .Z(n18795) );
  XNOR U19000 ( .A(n18794), .B(n18795), .Z(n18716) );
  XNOR U19001 ( .A(n18716), .B(n18717), .Z(n18719) );
  XNOR U19002 ( .A(n18718), .B(n18719), .Z(n18798) );
  NANDN U19003 ( .A(n18715), .B(n18714), .Z(n18799) );
  XNOR U19004 ( .A(n18798), .B(n18799), .Z(c[239]) );
  NAND U19005 ( .A(n18717), .B(n18716), .Z(n18721) );
  NANDN U19006 ( .A(n18719), .B(n18718), .Z(n18720) );
  NAND U19007 ( .A(n18721), .B(n18720), .Z(n18805) );
  NANDN U19008 ( .A(n18723), .B(n18722), .Z(n18727) );
  NANDN U19009 ( .A(n18725), .B(n18724), .Z(n18726) );
  NAND U19010 ( .A(n18727), .B(n18726), .Z(n18810) );
  NANDN U19011 ( .A(n18733), .B(n18732), .Z(n18737) );
  NAND U19012 ( .A(n18735), .B(n18734), .Z(n18736) );
  NAND U19013 ( .A(n18737), .B(n18736), .Z(n18858) );
  NANDN U19014 ( .A(n18738), .B(n19013), .Z(n18740) );
  XOR U19015 ( .A(a[124]), .B(n582), .Z(n18847) );
  NANDN U19016 ( .A(n18847), .B(n19015), .Z(n18739) );
  NAND U19017 ( .A(n18740), .B(n18739), .Z(n18871) );
  NANDN U19018 ( .A(n18741), .B(n18832), .Z(n18743) );
  XOR U19019 ( .A(a[126]), .B(n581), .Z(n18833) );
  NANDN U19020 ( .A(n18833), .B(n18834), .Z(n18742) );
  NAND U19021 ( .A(n18743), .B(n18742), .Z(n18868) );
  XOR U19022 ( .A(b[27]), .B(n19077), .Z(n18837) );
  NANDN U19023 ( .A(n18837), .B(n19336), .Z(n18746) );
  NANDN U19024 ( .A(n18744), .B(n19337), .Z(n18745) );
  AND U19025 ( .A(n18746), .B(n18745), .Z(n18869) );
  XNOR U19026 ( .A(n18868), .B(n18869), .Z(n18870) );
  XNOR U19027 ( .A(n18871), .B(n18870), .Z(n18856) );
  NAND U19028 ( .A(b[15]), .B(b[16]), .Z(n18840) );
  XNOR U19029 ( .A(b[17]), .B(n18840), .Z(n18750) );
  XNOR U19030 ( .A(b[16]), .B(b[15]), .Z(n18747) );
  NANDN U19031 ( .A(n18748), .B(n18747), .Z(n18749) );
  AND U19032 ( .A(n18750), .B(n18749), .Z(n18875) );
  AND U19033 ( .A(a[112]), .B(b[31]), .Z(n18942) );
  XOR U19034 ( .A(b[31]), .B(n18751), .Z(n18850) );
  NANDN U19035 ( .A(n18850), .B(n19472), .Z(n18754) );
  NANDN U19036 ( .A(n18752), .B(n19473), .Z(n18753) );
  AND U19037 ( .A(n18754), .B(n18753), .Z(n18874) );
  XOR U19038 ( .A(n18942), .B(n18874), .Z(n18876) );
  XOR U19039 ( .A(n18875), .B(n18876), .Z(n18857) );
  XOR U19040 ( .A(n18856), .B(n18857), .Z(n18859) );
  XNOR U19041 ( .A(n18858), .B(n18859), .Z(n18820) );
  NANDN U19042 ( .A(n18756), .B(n18755), .Z(n18760) );
  NANDN U19043 ( .A(n18758), .B(n18757), .Z(n18759) );
  AND U19044 ( .A(n18760), .B(n18759), .Z(n18821) );
  XNOR U19045 ( .A(n18820), .B(n18821), .Z(n18822) );
  NANDN U19046 ( .A(n18762), .B(n18761), .Z(n18766) );
  NAND U19047 ( .A(n18764), .B(n18763), .Z(n18765) );
  NAND U19048 ( .A(n18766), .B(n18765), .Z(n18865) );
  OR U19049 ( .A(n18768), .B(n18767), .Z(n18772) );
  NAND U19050 ( .A(n18770), .B(n18769), .Z(n18771) );
  NAND U19051 ( .A(n18772), .B(n18771), .Z(n18862) );
  XNOR U19052 ( .A(b[25]), .B(a[120]), .Z(n18853) );
  NANDN U19053 ( .A(n18853), .B(n19240), .Z(n18775) );
  NANDN U19054 ( .A(n18773), .B(n19242), .Z(n18774) );
  NAND U19055 ( .A(n18775), .B(n18774), .Z(n18829) );
  NAND U19056 ( .A(n19406), .B(n18776), .Z(n18778) );
  XOR U19057 ( .A(n584), .B(n18950), .Z(n18841) );
  NANDN U19058 ( .A(n576), .B(n18841), .Z(n18777) );
  NAND U19059 ( .A(n18778), .B(n18777), .Z(n18826) );
  XNOR U19060 ( .A(a[122]), .B(b[23]), .Z(n18844) );
  OR U19061 ( .A(n18844), .B(n19127), .Z(n18781) );
  NANDN U19062 ( .A(n18779), .B(n19128), .Z(n18780) );
  AND U19063 ( .A(n18781), .B(n18780), .Z(n18827) );
  XNOR U19064 ( .A(n18826), .B(n18827), .Z(n18828) );
  XNOR U19065 ( .A(n18829), .B(n18828), .Z(n18863) );
  XNOR U19066 ( .A(n18862), .B(n18863), .Z(n18864) );
  XNOR U19067 ( .A(n18865), .B(n18864), .Z(n18823) );
  XOR U19068 ( .A(n18822), .B(n18823), .Z(n18817) );
  NANDN U19069 ( .A(n18787), .B(n18786), .Z(n18791) );
  OR U19070 ( .A(n18789), .B(n18788), .Z(n18790) );
  AND U19071 ( .A(n18791), .B(n18790), .Z(n18815) );
  XNOR U19072 ( .A(n18814), .B(n18815), .Z(n18816) );
  XOR U19073 ( .A(n18817), .B(n18816), .Z(n18808) );
  XOR U19074 ( .A(n18809), .B(n18808), .Z(n18811) );
  XNOR U19075 ( .A(n18810), .B(n18811), .Z(n18802) );
  NAND U19076 ( .A(n18793), .B(n18792), .Z(n18797) );
  NANDN U19077 ( .A(n18795), .B(n18794), .Z(n18796) );
  AND U19078 ( .A(n18797), .B(n18796), .Z(n18803) );
  XNOR U19079 ( .A(n18802), .B(n18803), .Z(n18804) );
  XNOR U19080 ( .A(n18805), .B(n18804), .Z(n18801) );
  NANDN U19081 ( .A(n18799), .B(n18798), .Z(n18800) );
  XOR U19082 ( .A(n18801), .B(n18800), .Z(c[240]) );
  OR U19083 ( .A(n18801), .B(n18800), .Z(n18955) );
  NANDN U19084 ( .A(n18803), .B(n18802), .Z(n18807) );
  NAND U19085 ( .A(n18805), .B(n18804), .Z(n18806) );
  AND U19086 ( .A(n18807), .B(n18806), .Z(n18882) );
  NANDN U19087 ( .A(n18809), .B(n18808), .Z(n18813) );
  OR U19088 ( .A(n18811), .B(n18810), .Z(n18812) );
  AND U19089 ( .A(n18813), .B(n18812), .Z(n18881) );
  NANDN U19090 ( .A(n18815), .B(n18814), .Z(n18819) );
  NAND U19091 ( .A(n18817), .B(n18816), .Z(n18818) );
  NAND U19092 ( .A(n18819), .B(n18818), .Z(n18886) );
  NANDN U19093 ( .A(n18821), .B(n18820), .Z(n18825) );
  NANDN U19094 ( .A(n18823), .B(n18822), .Z(n18824) );
  NAND U19095 ( .A(n18825), .B(n18824), .Z(n18884) );
  NANDN U19096 ( .A(n18827), .B(n18826), .Z(n18831) );
  NAND U19097 ( .A(n18829), .B(n18828), .Z(n18830) );
  NAND U19098 ( .A(n18831), .B(n18830), .Z(n18904) );
  NANDN U19099 ( .A(n18833), .B(n18832), .Z(n18836) );
  XNOR U19100 ( .A(n19502), .B(b[19]), .Z(n18947) );
  NAND U19101 ( .A(n18947), .B(n18834), .Z(n18835) );
  NAND U19102 ( .A(n18836), .B(n18835), .Z(n18934) );
  XOR U19103 ( .A(b[27]), .B(n19239), .Z(n18925) );
  NANDN U19104 ( .A(n18925), .B(n19336), .Z(n18839) );
  NANDN U19105 ( .A(n18837), .B(n19337), .Z(n18838) );
  AND U19106 ( .A(n18839), .B(n18838), .Z(n18935) );
  XNOR U19107 ( .A(n18934), .B(n18935), .Z(n18936) );
  AND U19108 ( .A(n18840), .B(b[17]), .Z(n18941) );
  NANDN U19109 ( .A(n585), .B(a[113]), .Z(n18940) );
  XOR U19110 ( .A(n18941), .B(n18940), .Z(n18943) );
  XNOR U19111 ( .A(n18942), .B(n18943), .Z(n18937) );
  XOR U19112 ( .A(n18936), .B(n18937), .Z(n18901) );
  NAND U19113 ( .A(n19406), .B(n18841), .Z(n18843) );
  XOR U19114 ( .A(n584), .B(n19136), .Z(n18922) );
  NANDN U19115 ( .A(n576), .B(n18922), .Z(n18842) );
  NAND U19116 ( .A(n18843), .B(n18842), .Z(n18910) );
  XOR U19117 ( .A(a[123]), .B(b[23]), .Z(n18931) );
  NANDN U19118 ( .A(n19127), .B(n18931), .Z(n18846) );
  NANDN U19119 ( .A(n18844), .B(n19128), .Z(n18845) );
  NAND U19120 ( .A(n18846), .B(n18845), .Z(n18907) );
  NANDN U19121 ( .A(n18847), .B(n19013), .Z(n18849) );
  XOR U19122 ( .A(a[125]), .B(n582), .Z(n18928) );
  NANDN U19123 ( .A(n18928), .B(n19015), .Z(n18848) );
  NAND U19124 ( .A(n18849), .B(n18848), .Z(n18916) );
  XOR U19125 ( .A(b[31]), .B(n19022), .Z(n18951) );
  NANDN U19126 ( .A(n18951), .B(n19472), .Z(n18852) );
  NANDN U19127 ( .A(n18850), .B(n19473), .Z(n18851) );
  NAND U19128 ( .A(n18852), .B(n18851), .Z(n18913) );
  XNOR U19129 ( .A(b[25]), .B(a[121]), .Z(n18919) );
  NANDN U19130 ( .A(n18919), .B(n19240), .Z(n18855) );
  NANDN U19131 ( .A(n18853), .B(n19242), .Z(n18854) );
  AND U19132 ( .A(n18855), .B(n18854), .Z(n18914) );
  XNOR U19133 ( .A(n18913), .B(n18914), .Z(n18915) );
  XNOR U19134 ( .A(n18916), .B(n18915), .Z(n18908) );
  XNOR U19135 ( .A(n18907), .B(n18908), .Z(n18909) );
  XOR U19136 ( .A(n18910), .B(n18909), .Z(n18902) );
  XNOR U19137 ( .A(n18901), .B(n18902), .Z(n18903) );
  XOR U19138 ( .A(n18904), .B(n18903), .Z(n18889) );
  NANDN U19139 ( .A(n18857), .B(n18856), .Z(n18861) );
  OR U19140 ( .A(n18859), .B(n18858), .Z(n18860) );
  NAND U19141 ( .A(n18861), .B(n18860), .Z(n18890) );
  XNOR U19142 ( .A(n18889), .B(n18890), .Z(n18891) );
  NANDN U19143 ( .A(n18863), .B(n18862), .Z(n18867) );
  NAND U19144 ( .A(n18865), .B(n18864), .Z(n18866) );
  NAND U19145 ( .A(n18867), .B(n18866), .Z(n18898) );
  NANDN U19146 ( .A(n18869), .B(n18868), .Z(n18873) );
  NAND U19147 ( .A(n18871), .B(n18870), .Z(n18872) );
  NAND U19148 ( .A(n18873), .B(n18872), .Z(n18895) );
  OR U19149 ( .A(n18942), .B(n18874), .Z(n18878) );
  NAND U19150 ( .A(n18876), .B(n18875), .Z(n18877) );
  AND U19151 ( .A(n18878), .B(n18877), .Z(n18896) );
  XNOR U19152 ( .A(n18895), .B(n18896), .Z(n18897) );
  XOR U19153 ( .A(n18898), .B(n18897), .Z(n18892) );
  XOR U19154 ( .A(n18891), .B(n18892), .Z(n18883) );
  XNOR U19155 ( .A(n18884), .B(n18883), .Z(n18885) );
  XOR U19156 ( .A(n18886), .B(n18885), .Z(n18880) );
  XNOR U19157 ( .A(n18881), .B(n18880), .Z(n18879) );
  XNOR U19158 ( .A(n18882), .B(n18879), .Z(n18954) );
  XOR U19159 ( .A(n18955), .B(n18954), .Z(c[241]) );
  NAND U19160 ( .A(n18884), .B(n18883), .Z(n18888) );
  OR U19161 ( .A(n18886), .B(n18885), .Z(n18887) );
  NAND U19162 ( .A(n18888), .B(n18887), .Z(n18957) );
  NANDN U19163 ( .A(n18890), .B(n18889), .Z(n18894) );
  NAND U19164 ( .A(n18892), .B(n18891), .Z(n18893) );
  NAND U19165 ( .A(n18894), .B(n18893), .Z(n18964) );
  NANDN U19166 ( .A(n18896), .B(n18895), .Z(n18900) );
  NAND U19167 ( .A(n18898), .B(n18897), .Z(n18899) );
  NAND U19168 ( .A(n18900), .B(n18899), .Z(n18963) );
  NANDN U19169 ( .A(n18902), .B(n18901), .Z(n18906) );
  NANDN U19170 ( .A(n18904), .B(n18903), .Z(n18905) );
  NAND U19171 ( .A(n18906), .B(n18905), .Z(n18970) );
  NANDN U19172 ( .A(n18908), .B(n18907), .Z(n18912) );
  NAND U19173 ( .A(n18910), .B(n18909), .Z(n18911) );
  NAND U19174 ( .A(n18912), .B(n18911), .Z(n18969) );
  NANDN U19175 ( .A(n18914), .B(n18913), .Z(n18918) );
  NAND U19176 ( .A(n18916), .B(n18915), .Z(n18917) );
  NAND U19177 ( .A(n18918), .B(n18917), .Z(n18973) );
  XNOR U19178 ( .A(b[25]), .B(n19276), .Z(n19004) );
  NAND U19179 ( .A(n19004), .B(n19240), .Z(n18921) );
  NANDN U19180 ( .A(n18919), .B(n19242), .Z(n18920) );
  NAND U19181 ( .A(n18921), .B(n18920), .Z(n18998) );
  NAND U19182 ( .A(n19406), .B(n18922), .Z(n18924) );
  XOR U19183 ( .A(b[29]), .B(n19077), .Z(n19001) );
  OR U19184 ( .A(n19001), .B(n576), .Z(n18923) );
  NAND U19185 ( .A(n18924), .B(n18923), .Z(n18995) );
  XOR U19186 ( .A(n583), .B(n19188), .Z(n19018) );
  NAND U19187 ( .A(n19336), .B(n19018), .Z(n18927) );
  NANDN U19188 ( .A(n18925), .B(n19337), .Z(n18926) );
  AND U19189 ( .A(n18927), .B(n18926), .Z(n18996) );
  XNOR U19190 ( .A(n18995), .B(n18996), .Z(n18997) );
  XNOR U19191 ( .A(n18998), .B(n18997), .Z(n18981) );
  NANDN U19192 ( .A(n18928), .B(n19013), .Z(n18930) );
  XOR U19193 ( .A(a[126]), .B(n582), .Z(n19014) );
  NANDN U19194 ( .A(n19014), .B(n19015), .Z(n18929) );
  NAND U19195 ( .A(n18930), .B(n18929), .Z(n18978) );
  XNOR U19196 ( .A(a[124]), .B(b[23]), .Z(n19007) );
  OR U19197 ( .A(n19007), .B(n19127), .Z(n18933) );
  NAND U19198 ( .A(n18931), .B(n19128), .Z(n18932) );
  AND U19199 ( .A(n18933), .B(n18932), .Z(n18979) );
  XNOR U19200 ( .A(n18978), .B(n18979), .Z(n18980) );
  XNOR U19201 ( .A(n18981), .B(n18980), .Z(n18972) );
  XNOR U19202 ( .A(n18973), .B(n18972), .Z(n18975) );
  NANDN U19203 ( .A(n18935), .B(n18934), .Z(n18939) );
  NANDN U19204 ( .A(n18937), .B(n18936), .Z(n18938) );
  NAND U19205 ( .A(n18939), .B(n18938), .Z(n18986) );
  OR U19206 ( .A(n18941), .B(n18940), .Z(n18945) );
  NAND U19207 ( .A(n18943), .B(n18942), .Z(n18944) );
  NAND U19208 ( .A(n18945), .B(n18944), .Z(n18985) );
  NAND U19209 ( .A(b[17]), .B(b[18]), .Z(n19021) );
  XOR U19210 ( .A(n581), .B(n19021), .Z(n18949) );
  XNOR U19211 ( .A(b[18]), .B(b[17]), .Z(n18946) );
  NANDN U19212 ( .A(n18947), .B(n18946), .Z(n18948) );
  AND U19213 ( .A(n18949), .B(n18948), .Z(n18991) );
  AND U19214 ( .A(a[114]), .B(b[31]), .Z(n19055) );
  XOR U19215 ( .A(n585), .B(n18950), .Z(n19010) );
  NAND U19216 ( .A(n19010), .B(n19472), .Z(n18953) );
  NANDN U19217 ( .A(n18951), .B(n19473), .Z(n18952) );
  AND U19218 ( .A(n18953), .B(n18952), .Z(n18990) );
  XOR U19219 ( .A(n19055), .B(n18990), .Z(n18992) );
  XOR U19220 ( .A(n18991), .B(n18992), .Z(n18984) );
  XNOR U19221 ( .A(n18985), .B(n18984), .Z(n18987) );
  XNOR U19222 ( .A(n18986), .B(n18987), .Z(n18974) );
  XNOR U19223 ( .A(n18975), .B(n18974), .Z(n18968) );
  XNOR U19224 ( .A(n18969), .B(n18968), .Z(n18971) );
  XOR U19225 ( .A(n18970), .B(n18971), .Z(n18962) );
  XNOR U19226 ( .A(n18963), .B(n18962), .Z(n18965) );
  XNOR U19227 ( .A(n18964), .B(n18965), .Z(n18956) );
  XNOR U19228 ( .A(n18957), .B(n18956), .Z(n18959) );
  XNOR U19229 ( .A(n18958), .B(n18959), .Z(n19023) );
  OR U19230 ( .A(n18955), .B(n18954), .Z(n19024) );
  XNOR U19231 ( .A(n19023), .B(n19024), .Z(c[242]) );
  NAND U19232 ( .A(n18957), .B(n18956), .Z(n18961) );
  NANDN U19233 ( .A(n18959), .B(n18958), .Z(n18960) );
  NAND U19234 ( .A(n18961), .B(n18960), .Z(n19027) );
  NAND U19235 ( .A(n18963), .B(n18962), .Z(n18967) );
  NANDN U19236 ( .A(n18965), .B(n18964), .Z(n18966) );
  NAND U19237 ( .A(n18967), .B(n18966), .Z(n19026) );
  NAND U19238 ( .A(n18973), .B(n18972), .Z(n18977) );
  NANDN U19239 ( .A(n18975), .B(n18974), .Z(n18976) );
  NAND U19240 ( .A(n18977), .B(n18976), .Z(n19032) );
  NANDN U19241 ( .A(n18979), .B(n18978), .Z(n18983) );
  NANDN U19242 ( .A(n18981), .B(n18980), .Z(n18982) );
  NAND U19243 ( .A(n18983), .B(n18982), .Z(n19037) );
  NAND U19244 ( .A(n18985), .B(n18984), .Z(n18989) );
  NANDN U19245 ( .A(n18987), .B(n18986), .Z(n18988) );
  AND U19246 ( .A(n18989), .B(n18988), .Z(n19038) );
  XNOR U19247 ( .A(n19037), .B(n19038), .Z(n19039) );
  OR U19248 ( .A(n19055), .B(n18990), .Z(n18994) );
  NAND U19249 ( .A(n18992), .B(n18991), .Z(n18993) );
  NAND U19250 ( .A(n18994), .B(n18993), .Z(n19043) );
  NANDN U19251 ( .A(n18996), .B(n18995), .Z(n19000) );
  NAND U19252 ( .A(n18998), .B(n18997), .Z(n18999) );
  AND U19253 ( .A(n19000), .B(n18999), .Z(n19044) );
  XNOR U19254 ( .A(n19043), .B(n19044), .Z(n19045) );
  NANDN U19255 ( .A(n19001), .B(n19406), .Z(n19003) );
  XOR U19256 ( .A(b[29]), .B(n19239), .Z(n19090) );
  OR U19257 ( .A(n19090), .B(n576), .Z(n19002) );
  AND U19258 ( .A(n19003), .B(n19002), .Z(n19067) );
  XOR U19259 ( .A(b[25]), .B(a[123]), .Z(n19081) );
  NAND U19260 ( .A(n19081), .B(n19240), .Z(n19006) );
  NAND U19261 ( .A(n19004), .B(n19242), .Z(n19005) );
  NAND U19262 ( .A(n19006), .B(n19005), .Z(n19052) );
  XNOR U19263 ( .A(a[125]), .B(b[23]), .Z(n19084) );
  OR U19264 ( .A(n19084), .B(n19127), .Z(n19009) );
  NANDN U19265 ( .A(n19007), .B(n19128), .Z(n19008) );
  AND U19266 ( .A(n19009), .B(n19008), .Z(n19049) );
  XOR U19267 ( .A(n585), .B(n19136), .Z(n19078) );
  NAND U19268 ( .A(n19078), .B(n19472), .Z(n19012) );
  NAND U19269 ( .A(n19010), .B(n19473), .Z(n19011) );
  AND U19270 ( .A(n19012), .B(n19011), .Z(n19050) );
  XNOR U19271 ( .A(n19052), .B(n19051), .Z(n19068) );
  NANDN U19272 ( .A(n19014), .B(n19013), .Z(n19017) );
  XNOR U19273 ( .A(n19502), .B(b[21]), .Z(n19074) );
  NAND U19274 ( .A(n19074), .B(n19015), .Z(n19016) );
  AND U19275 ( .A(n19017), .B(n19016), .Z(n19061) );
  XOR U19276 ( .A(b[27]), .B(n19347), .Z(n19087) );
  NANDN U19277 ( .A(n19087), .B(n19336), .Z(n19020) );
  NAND U19278 ( .A(n19018), .B(n19337), .Z(n19019) );
  AND U19279 ( .A(n19020), .B(n19019), .Z(n19062) );
  ANDN U19280 ( .B(n19021), .A(n581), .Z(n19056) );
  XOR U19281 ( .A(n19056), .B(n19055), .Z(n19058) );
  NANDN U19282 ( .A(n19022), .B(b[31]), .Z(n19057) );
  XOR U19283 ( .A(n19058), .B(n19057), .Z(n19063) );
  XOR U19284 ( .A(n19045), .B(n19046), .Z(n19040) );
  XOR U19285 ( .A(n19039), .B(n19040), .Z(n19031) );
  XNOR U19286 ( .A(n19032), .B(n19031), .Z(n19034) );
  XNOR U19287 ( .A(n19033), .B(n19034), .Z(n19025) );
  XNOR U19288 ( .A(n19026), .B(n19025), .Z(n19028) );
  XNOR U19289 ( .A(n19027), .B(n19028), .Z(n19093) );
  NANDN U19290 ( .A(n19024), .B(n19023), .Z(n19094) );
  XNOR U19291 ( .A(n19093), .B(n19094), .Z(c[243]) );
  NAND U19292 ( .A(n19026), .B(n19025), .Z(n19030) );
  NANDN U19293 ( .A(n19028), .B(n19027), .Z(n19029) );
  NAND U19294 ( .A(n19030), .B(n19029), .Z(n19100) );
  NAND U19295 ( .A(n19032), .B(n19031), .Z(n19036) );
  NANDN U19296 ( .A(n19034), .B(n19033), .Z(n19035) );
  NAND U19297 ( .A(n19036), .B(n19035), .Z(n19097) );
  NANDN U19298 ( .A(n19038), .B(n19037), .Z(n19042) );
  NAND U19299 ( .A(n19040), .B(n19039), .Z(n19041) );
  NAND U19300 ( .A(n19042), .B(n19041), .Z(n19106) );
  NANDN U19301 ( .A(n19044), .B(n19043), .Z(n19048) );
  NAND U19302 ( .A(n19046), .B(n19045), .Z(n19047) );
  NAND U19303 ( .A(n19048), .B(n19047), .Z(n19103) );
  OR U19304 ( .A(n19050), .B(n19049), .Z(n19054) );
  NAND U19305 ( .A(n19052), .B(n19051), .Z(n19053) );
  NAND U19306 ( .A(n19054), .B(n19053), .Z(n19154) );
  NANDN U19307 ( .A(n19056), .B(n19055), .Z(n19060) );
  OR U19308 ( .A(n19058), .B(n19057), .Z(n19059) );
  NAND U19309 ( .A(n19060), .B(n19059), .Z(n19152) );
  OR U19310 ( .A(n19062), .B(n19061), .Z(n19066) );
  NANDN U19311 ( .A(n19064), .B(n19063), .Z(n19065) );
  NAND U19312 ( .A(n19066), .B(n19065), .Z(n19151) );
  XOR U19313 ( .A(n19154), .B(n19153), .Z(n19112) );
  OR U19314 ( .A(n19068), .B(n19067), .Z(n19072) );
  NANDN U19315 ( .A(n19070), .B(n19069), .Z(n19071) );
  AND U19316 ( .A(n19072), .B(n19071), .Z(n19109) );
  NANDN U19317 ( .A(n581), .B(b[20]), .Z(n19135) );
  XOR U19318 ( .A(n582), .B(n19135), .Z(n19076) );
  XOR U19319 ( .A(b[20]), .B(n581), .Z(n19073) );
  NANDN U19320 ( .A(n19074), .B(n19073), .Z(n19075) );
  AND U19321 ( .A(n19076), .B(n19075), .Z(n19146) );
  AND U19322 ( .A(a[116]), .B(b[31]), .Z(n19200) );
  XNOR U19323 ( .A(n19146), .B(n19200), .Z(n19147) );
  XOR U19324 ( .A(b[31]), .B(n19077), .Z(n19143) );
  NANDN U19325 ( .A(n19143), .B(n19472), .Z(n19080) );
  NAND U19326 ( .A(n19473), .B(n19078), .Z(n19079) );
  AND U19327 ( .A(n19080), .B(n19079), .Z(n19148) );
  XNOR U19328 ( .A(n19147), .B(n19148), .Z(n19117) );
  XNOR U19329 ( .A(a[124]), .B(b[25]), .Z(n19137) );
  NANDN U19330 ( .A(n19137), .B(n19240), .Z(n19083) );
  NAND U19331 ( .A(n19081), .B(n19242), .Z(n19082) );
  NAND U19332 ( .A(n19083), .B(n19082), .Z(n19124) );
  XNOR U19333 ( .A(a[126]), .B(b[23]), .Z(n19129) );
  OR U19334 ( .A(n19129), .B(n19127), .Z(n19086) );
  NANDN U19335 ( .A(n19084), .B(n19128), .Z(n19085) );
  NAND U19336 ( .A(n19086), .B(n19085), .Z(n19121) );
  XOR U19337 ( .A(b[27]), .B(n19276), .Z(n19132) );
  NANDN U19338 ( .A(n19132), .B(n19336), .Z(n19089) );
  NANDN U19339 ( .A(n19087), .B(n19337), .Z(n19088) );
  AND U19340 ( .A(n19089), .B(n19088), .Z(n19122) );
  XNOR U19341 ( .A(n19121), .B(n19122), .Z(n19123) );
  XNOR U19342 ( .A(n19124), .B(n19123), .Z(n19115) );
  NANDN U19343 ( .A(n19090), .B(n19406), .Z(n19092) );
  XNOR U19344 ( .A(n584), .B(a[120]), .Z(n19140) );
  NANDN U19345 ( .A(n576), .B(n19140), .Z(n19091) );
  NAND U19346 ( .A(n19092), .B(n19091), .Z(n19116) );
  XOR U19347 ( .A(n19115), .B(n19116), .Z(n19118) );
  XOR U19348 ( .A(n19117), .B(n19118), .Z(n19110) );
  XNOR U19349 ( .A(n19112), .B(n19111), .Z(n19104) );
  XNOR U19350 ( .A(n19103), .B(n19104), .Z(n19105) );
  XNOR U19351 ( .A(n19106), .B(n19105), .Z(n19098) );
  XNOR U19352 ( .A(n19097), .B(n19098), .Z(n19099) );
  XNOR U19353 ( .A(n19100), .B(n19099), .Z(n19096) );
  NANDN U19354 ( .A(n19094), .B(n19093), .Z(n19095) );
  XOR U19355 ( .A(n19096), .B(n19095), .Z(c[244]) );
  OR U19356 ( .A(n19096), .B(n19095), .Z(n19159) );
  NANDN U19357 ( .A(n19098), .B(n19097), .Z(n19102) );
  NAND U19358 ( .A(n19100), .B(n19099), .Z(n19101) );
  NAND U19359 ( .A(n19102), .B(n19101), .Z(n19206) );
  NANDN U19360 ( .A(n19104), .B(n19103), .Z(n19108) );
  NAND U19361 ( .A(n19106), .B(n19105), .Z(n19107) );
  AND U19362 ( .A(n19108), .B(n19107), .Z(n19205) );
  OR U19363 ( .A(n19110), .B(n19109), .Z(n19114) );
  NAND U19364 ( .A(n19112), .B(n19111), .Z(n19113) );
  AND U19365 ( .A(n19114), .B(n19113), .Z(n19209) );
  NANDN U19366 ( .A(n19116), .B(n19115), .Z(n19120) );
  OR U19367 ( .A(n19118), .B(n19117), .Z(n19119) );
  NAND U19368 ( .A(n19120), .B(n19119), .Z(n19163) );
  NANDN U19369 ( .A(n19122), .B(n19121), .Z(n19126) );
  NAND U19370 ( .A(n19124), .B(n19123), .Z(n19125) );
  NAND U19371 ( .A(n19126), .B(n19125), .Z(n19167) );
  XNOR U19372 ( .A(n19502), .B(b[23]), .Z(n19185) );
  NANDN U19373 ( .A(n19127), .B(n19185), .Z(n19131) );
  NANDN U19374 ( .A(n19129), .B(n19128), .Z(n19130) );
  NAND U19375 ( .A(n19131), .B(n19130), .Z(n19192) );
  XNOR U19376 ( .A(b[27]), .B(a[123]), .Z(n19174) );
  NANDN U19377 ( .A(n19174), .B(n19336), .Z(n19134) );
  NANDN U19378 ( .A(n19132), .B(n19337), .Z(n19133) );
  AND U19379 ( .A(n19134), .B(n19133), .Z(n19193) );
  XNOR U19380 ( .A(n19192), .B(n19193), .Z(n19194) );
  NANDN U19381 ( .A(n582), .B(n19135), .Z(n19199) );
  ANDN U19382 ( .B(b[31]), .A(n19136), .Z(n19198) );
  XNOR U19383 ( .A(n19199), .B(n19198), .Z(n19201) );
  XOR U19384 ( .A(n19200), .B(n19201), .Z(n19195) );
  XNOR U19385 ( .A(n19194), .B(n19195), .Z(n19164) );
  XNOR U19386 ( .A(a[125]), .B(b[25]), .Z(n19177) );
  NANDN U19387 ( .A(n19177), .B(n19240), .Z(n19139) );
  NANDN U19388 ( .A(n19137), .B(n19242), .Z(n19138) );
  NAND U19389 ( .A(n19139), .B(n19138), .Z(n19171) );
  NAND U19390 ( .A(n19140), .B(n19406), .Z(n19142) );
  XOR U19391 ( .A(n584), .B(n19347), .Z(n19180) );
  NANDN U19392 ( .A(n576), .B(n19180), .Z(n19141) );
  NAND U19393 ( .A(n19142), .B(n19141), .Z(n19168) );
  XOR U19394 ( .A(n585), .B(n19239), .Z(n19189) );
  NAND U19395 ( .A(n19189), .B(n19472), .Z(n19145) );
  NANDN U19396 ( .A(n19143), .B(n19473), .Z(n19144) );
  AND U19397 ( .A(n19145), .B(n19144), .Z(n19169) );
  XNOR U19398 ( .A(n19168), .B(n19169), .Z(n19170) );
  XOR U19399 ( .A(n19171), .B(n19170), .Z(n19165) );
  XOR U19400 ( .A(n19164), .B(n19165), .Z(n19166) );
  XNOR U19401 ( .A(n19167), .B(n19166), .Z(n19160) );
  NANDN U19402 ( .A(n19146), .B(n19200), .Z(n19150) );
  NAND U19403 ( .A(n19148), .B(n19147), .Z(n19149) );
  AND U19404 ( .A(n19150), .B(n19149), .Z(n19161) );
  XNOR U19405 ( .A(n19160), .B(n19161), .Z(n19162) );
  XNOR U19406 ( .A(n19163), .B(n19162), .Z(n19207) );
  OR U19407 ( .A(n19152), .B(n19151), .Z(n19156) );
  NANDN U19408 ( .A(n19154), .B(n19153), .Z(n19155) );
  NAND U19409 ( .A(n19156), .B(n19155), .Z(n19208) );
  XOR U19410 ( .A(n19207), .B(n19208), .Z(n19210) );
  XOR U19411 ( .A(n19205), .B(n19204), .Z(n19157) );
  XOR U19412 ( .A(n19206), .B(n19157), .Z(n19158) );
  XNOR U19413 ( .A(n19159), .B(n19158), .Z(c[245]) );
  NANDN U19414 ( .A(n19159), .B(n19158), .Z(n19215) );
  NANDN U19415 ( .A(n19169), .B(n19168), .Z(n19173) );
  NAND U19416 ( .A(n19171), .B(n19170), .Z(n19172) );
  NAND U19417 ( .A(n19173), .B(n19172), .Z(n19250) );
  XOR U19418 ( .A(b[27]), .B(n19373), .Z(n19236) );
  NANDN U19419 ( .A(n19236), .B(n19336), .Z(n19176) );
  NANDN U19420 ( .A(n19174), .B(n19337), .Z(n19175) );
  NAND U19421 ( .A(n19176), .B(n19175), .Z(n19225) );
  XNOR U19422 ( .A(n19295), .B(b[25]), .Z(n19241) );
  NAND U19423 ( .A(n19241), .B(n19240), .Z(n19179) );
  NANDN U19424 ( .A(n19177), .B(n19242), .Z(n19178) );
  NAND U19425 ( .A(n19179), .B(n19178), .Z(n19222) );
  NAND U19426 ( .A(n19406), .B(n19180), .Z(n19182) );
  XOR U19427 ( .A(b[29]), .B(n19276), .Z(n19245) );
  OR U19428 ( .A(n19245), .B(n576), .Z(n19181) );
  AND U19429 ( .A(n19182), .B(n19181), .Z(n19223) );
  XNOR U19430 ( .A(n19222), .B(n19223), .Z(n19224) );
  XNOR U19431 ( .A(n19225), .B(n19224), .Z(n19248) );
  XNOR U19432 ( .A(b[23]), .B(n19183), .Z(n19187) );
  XOR U19433 ( .A(b[22]), .B(n582), .Z(n19184) );
  NANDN U19434 ( .A(n19185), .B(n19184), .Z(n19186) );
  AND U19435 ( .A(n19187), .B(n19186), .Z(n19228) );
  AND U19436 ( .A(a[118]), .B(b[31]), .Z(n19288) );
  XNOR U19437 ( .A(n19228), .B(n19288), .Z(n19229) );
  XOR U19438 ( .A(b[31]), .B(n19188), .Z(n19233) );
  NANDN U19439 ( .A(n19233), .B(n19472), .Z(n19191) );
  NAND U19440 ( .A(n19473), .B(n19189), .Z(n19190) );
  AND U19441 ( .A(n19191), .B(n19190), .Z(n19230) );
  XNOR U19442 ( .A(n19229), .B(n19230), .Z(n19249) );
  XOR U19443 ( .A(n19248), .B(n19249), .Z(n19251) );
  XNOR U19444 ( .A(n19250), .B(n19251), .Z(n19219) );
  NANDN U19445 ( .A(n19193), .B(n19192), .Z(n19197) );
  NANDN U19446 ( .A(n19195), .B(n19194), .Z(n19196) );
  NAND U19447 ( .A(n19197), .B(n19196), .Z(n19216) );
  NAND U19448 ( .A(n19199), .B(n19198), .Z(n19203) );
  NANDN U19449 ( .A(n19201), .B(n19200), .Z(n19202) );
  AND U19450 ( .A(n19203), .B(n19202), .Z(n19217) );
  XNOR U19451 ( .A(n19216), .B(n19217), .Z(n19218) );
  XNOR U19452 ( .A(n19219), .B(n19218), .Z(n19255) );
  XNOR U19453 ( .A(n19254), .B(n19255), .Z(n19256) );
  XOR U19454 ( .A(n19257), .B(n19256), .Z(n19261) );
  NANDN U19455 ( .A(n19208), .B(n19207), .Z(n19212) );
  OR U19456 ( .A(n19210), .B(n19209), .Z(n19211) );
  NAND U19457 ( .A(n19212), .B(n19211), .Z(n19260) );
  XOR U19458 ( .A(n19262), .B(n19260), .Z(n19213) );
  XNOR U19459 ( .A(n19261), .B(n19213), .Z(n19214) );
  XNOR U19460 ( .A(n19215), .B(n19214), .Z(c[246]) );
  NANDN U19461 ( .A(n19215), .B(n19214), .Z(n19312) );
  NANDN U19462 ( .A(n19217), .B(n19216), .Z(n19221) );
  NAND U19463 ( .A(n19219), .B(n19218), .Z(n19220) );
  NAND U19464 ( .A(n19221), .B(n19220), .Z(n19307) );
  NANDN U19465 ( .A(n19223), .B(n19222), .Z(n19227) );
  NAND U19466 ( .A(n19225), .B(n19224), .Z(n19226) );
  NAND U19467 ( .A(n19227), .B(n19226), .Z(n19270) );
  NANDN U19468 ( .A(n19228), .B(n19288), .Z(n19232) );
  NAND U19469 ( .A(n19230), .B(n19229), .Z(n19231) );
  NAND U19470 ( .A(n19232), .B(n19231), .Z(n19268) );
  XOR U19471 ( .A(n585), .B(n19347), .Z(n19277) );
  NAND U19472 ( .A(n19277), .B(n19472), .Z(n19235) );
  NANDN U19473 ( .A(n19233), .B(n19473), .Z(n19234) );
  NAND U19474 ( .A(n19235), .B(n19234), .Z(n19301) );
  XOR U19475 ( .A(b[27]), .B(n19402), .Z(n19296) );
  NANDN U19476 ( .A(n19296), .B(n19336), .Z(n19238) );
  NANDN U19477 ( .A(n19236), .B(n19337), .Z(n19237) );
  NAND U19478 ( .A(n19238), .B(n19237), .Z(n19300) );
  NANDN U19479 ( .A(n19239), .B(b[31]), .Z(n19286) );
  XOR U19480 ( .A(n19287), .B(n19286), .Z(n19289) );
  XNOR U19481 ( .A(n19288), .B(n19289), .Z(n19283) );
  XNOR U19482 ( .A(a[127]), .B(b[25]), .Z(n19272) );
  NANDN U19483 ( .A(n19272), .B(n19240), .Z(n19244) );
  NAND U19484 ( .A(n19242), .B(n19241), .Z(n19243) );
  NAND U19485 ( .A(n19244), .B(n19243), .Z(n19280) );
  NANDN U19486 ( .A(n19245), .B(n19406), .Z(n19247) );
  XNOR U19487 ( .A(b[29]), .B(a[123]), .Z(n19292) );
  OR U19488 ( .A(n19292), .B(n576), .Z(n19246) );
  NAND U19489 ( .A(n19247), .B(n19246), .Z(n19281) );
  XOR U19490 ( .A(n19280), .B(n19281), .Z(n19282) );
  XNOR U19491 ( .A(n19283), .B(n19282), .Z(n19299) );
  XNOR U19492 ( .A(n19300), .B(n19299), .Z(n19302) );
  XNOR U19493 ( .A(n19301), .B(n19302), .Z(n19267) );
  XNOR U19494 ( .A(n19268), .B(n19267), .Z(n19269) );
  XNOR U19495 ( .A(n19270), .B(n19269), .Z(n19305) );
  NANDN U19496 ( .A(n19249), .B(n19248), .Z(n19253) );
  OR U19497 ( .A(n19251), .B(n19250), .Z(n19252) );
  AND U19498 ( .A(n19253), .B(n19252), .Z(n19306) );
  XOR U19499 ( .A(n19305), .B(n19306), .Z(n19308) );
  XNOR U19500 ( .A(n19307), .B(n19308), .Z(n19265) );
  NANDN U19501 ( .A(n19255), .B(n19254), .Z(n19259) );
  NANDN U19502 ( .A(n19257), .B(n19256), .Z(n19258) );
  NAND U19503 ( .A(n19259), .B(n19258), .Z(n19264) );
  XNOR U19504 ( .A(n19264), .B(n19266), .Z(n19263) );
  XOR U19505 ( .A(n19265), .B(n19263), .Z(n19311) );
  XOR U19506 ( .A(n19312), .B(n19311), .Z(c[247]) );
  XNOR U19507 ( .A(b[25]), .B(n19271), .Z(n19275) );
  XNOR U19508 ( .A(b[24]), .B(b[23]), .Z(n19273) );
  NAND U19509 ( .A(n19273), .B(n19272), .Z(n19274) );
  AND U19510 ( .A(n19275), .B(n19274), .Z(n19333) );
  AND U19511 ( .A(a[120]), .B(b[31]), .Z(n19382) );
  XNOR U19512 ( .A(n19333), .B(n19382), .Z(n19334) );
  XOR U19513 ( .A(b[31]), .B(n19276), .Z(n19344) );
  NANDN U19514 ( .A(n19344), .B(n19472), .Z(n19279) );
  NAND U19515 ( .A(n19473), .B(n19277), .Z(n19278) );
  AND U19516 ( .A(n19279), .B(n19278), .Z(n19335) );
  XNOR U19517 ( .A(n19334), .B(n19335), .Z(n19323) );
  NAND U19518 ( .A(n19281), .B(n19280), .Z(n19285) );
  NANDN U19519 ( .A(n19283), .B(n19282), .Z(n19284) );
  AND U19520 ( .A(n19285), .B(n19284), .Z(n19324) );
  XNOR U19521 ( .A(n19323), .B(n19324), .Z(n19325) );
  OR U19522 ( .A(n19287), .B(n19286), .Z(n19291) );
  NAND U19523 ( .A(n19289), .B(n19288), .Z(n19290) );
  NAND U19524 ( .A(n19291), .B(n19290), .Z(n19332) );
  NANDN U19525 ( .A(n19292), .B(n19406), .Z(n19294) );
  XNOR U19526 ( .A(n584), .B(a[124]), .Z(n19341) );
  NANDN U19527 ( .A(n576), .B(n19341), .Z(n19293) );
  NAND U19528 ( .A(n19294), .B(n19293), .Z(n19329) );
  XOR U19529 ( .A(b[27]), .B(n19295), .Z(n19338) );
  NANDN U19530 ( .A(n19338), .B(n19336), .Z(n19298) );
  NANDN U19531 ( .A(n19296), .B(n19337), .Z(n19297) );
  AND U19532 ( .A(n19298), .B(n19297), .Z(n19330) );
  XNOR U19533 ( .A(n19329), .B(n19330), .Z(n19331) );
  XOR U19534 ( .A(n19332), .B(n19331), .Z(n19326) );
  XNOR U19535 ( .A(n19325), .B(n19326), .Z(n19319) );
  NAND U19536 ( .A(n19300), .B(n19299), .Z(n19304) );
  NANDN U19537 ( .A(n19302), .B(n19301), .Z(n19303) );
  NAND U19538 ( .A(n19304), .B(n19303), .Z(n19320) );
  XNOR U19539 ( .A(n19319), .B(n19320), .Z(n19321) );
  XOR U19540 ( .A(n19322), .B(n19321), .Z(n19313) );
  NANDN U19541 ( .A(n19306), .B(n19305), .Z(n19310) );
  OR U19542 ( .A(n19308), .B(n19307), .Z(n19309) );
  NAND U19543 ( .A(n19310), .B(n19309), .Z(n19314) );
  XNOR U19544 ( .A(n19313), .B(n19314), .Z(n19316) );
  XOR U19545 ( .A(n19315), .B(n19316), .Z(n19348) );
  OR U19546 ( .A(n19312), .B(n19311), .Z(n19349) );
  XNOR U19547 ( .A(n19348), .B(n19349), .Z(c[248]) );
  NANDN U19548 ( .A(n19314), .B(n19313), .Z(n19318) );
  NAND U19549 ( .A(n19316), .B(n19315), .Z(n19317) );
  NAND U19550 ( .A(n19318), .B(n19317), .Z(n19355) );
  NANDN U19551 ( .A(n19324), .B(n19323), .Z(n19328) );
  NAND U19552 ( .A(n19326), .B(n19325), .Z(n19327) );
  NAND U19553 ( .A(n19328), .B(n19327), .Z(n19361) );
  XNOR U19554 ( .A(n19502), .B(b[27]), .Z(n19370) );
  NAND U19555 ( .A(n19336), .B(n19370), .Z(n19340) );
  NANDN U19556 ( .A(n19338), .B(n19337), .Z(n19339) );
  NAND U19557 ( .A(n19340), .B(n19339), .Z(n19365) );
  NAND U19558 ( .A(n19341), .B(n19406), .Z(n19343) );
  XOR U19559 ( .A(b[29]), .B(n19402), .Z(n19377) );
  OR U19560 ( .A(n19377), .B(n576), .Z(n19342) );
  NAND U19561 ( .A(n19343), .B(n19342), .Z(n19386) );
  XNOR U19562 ( .A(b[31]), .B(a[123]), .Z(n19374) );
  NANDN U19563 ( .A(n19374), .B(n19472), .Z(n19346) );
  NANDN U19564 ( .A(n19344), .B(n19473), .Z(n19345) );
  AND U19565 ( .A(n19346), .B(n19345), .Z(n19387) );
  XNOR U19566 ( .A(n19386), .B(n19387), .Z(n19388) );
  NANDN U19567 ( .A(n19347), .B(b[31]), .Z(n19380) );
  XOR U19568 ( .A(n19381), .B(n19380), .Z(n19383) );
  XNOR U19569 ( .A(n19382), .B(n19383), .Z(n19389) );
  XNOR U19570 ( .A(n19388), .B(n19389), .Z(n19364) );
  XNOR U19571 ( .A(n19365), .B(n19364), .Z(n19367) );
  XOR U19572 ( .A(n19366), .B(n19367), .Z(n19358) );
  XOR U19573 ( .A(n19359), .B(n19358), .Z(n19360) );
  XOR U19574 ( .A(n19361), .B(n19360), .Z(n19352) );
  XNOR U19575 ( .A(n19353), .B(n19352), .Z(n19354) );
  XNOR U19576 ( .A(n19355), .B(n19354), .Z(n19351) );
  NANDN U19577 ( .A(n19349), .B(n19348), .Z(n19350) );
  XOR U19578 ( .A(n19351), .B(n19350), .Z(c[249]) );
  OR U19579 ( .A(n19351), .B(n19350), .Z(n19420) );
  NANDN U19580 ( .A(n19353), .B(n19352), .Z(n19357) );
  NAND U19581 ( .A(n19355), .B(n19354), .Z(n19356) );
  AND U19582 ( .A(n19357), .B(n19356), .Z(n19395) );
  NAND U19583 ( .A(n19359), .B(n19358), .Z(n19363) );
  NAND U19584 ( .A(n19361), .B(n19360), .Z(n19362) );
  NAND U19585 ( .A(n19363), .B(n19362), .Z(n19393) );
  XOR U19586 ( .A(n583), .B(n19368), .Z(n19372) );
  XNOR U19587 ( .A(b[26]), .B(b[25]), .Z(n19369) );
  NANDN U19588 ( .A(n19370), .B(n19369), .Z(n19371) );
  AND U19589 ( .A(n19372), .B(n19371), .Z(n19410) );
  AND U19590 ( .A(a[122]), .B(b[31]), .Z(n19451) );
  XNOR U19591 ( .A(n19410), .B(n19451), .Z(n19411) );
  XOR U19592 ( .A(b[31]), .B(n19373), .Z(n19403) );
  NANDN U19593 ( .A(n19403), .B(n19472), .Z(n19376) );
  NANDN U19594 ( .A(n19374), .B(n19473), .Z(n19375) );
  AND U19595 ( .A(n19376), .B(n19375), .Z(n19412) );
  XOR U19596 ( .A(n19411), .B(n19412), .Z(n19399) );
  NANDN U19597 ( .A(n19377), .B(n19406), .Z(n19379) );
  XNOR U19598 ( .A(n584), .B(a[126]), .Z(n19407) );
  NANDN U19599 ( .A(n576), .B(n19407), .Z(n19378) );
  NAND U19600 ( .A(n19379), .B(n19378), .Z(n19396) );
  OR U19601 ( .A(n19381), .B(n19380), .Z(n19385) );
  NAND U19602 ( .A(n19383), .B(n19382), .Z(n19384) );
  NAND U19603 ( .A(n19385), .B(n19384), .Z(n19397) );
  XOR U19604 ( .A(n19396), .B(n19397), .Z(n19398) );
  XOR U19605 ( .A(n19399), .B(n19398), .Z(n19413) );
  NANDN U19606 ( .A(n19387), .B(n19386), .Z(n19391) );
  NANDN U19607 ( .A(n19389), .B(n19388), .Z(n19390) );
  NAND U19608 ( .A(n19391), .B(n19390), .Z(n19414) );
  XOR U19609 ( .A(n19413), .B(n19414), .Z(n19416) );
  XOR U19610 ( .A(n19415), .B(n19416), .Z(n19394) );
  XOR U19611 ( .A(n19393), .B(n19394), .Z(n19392) );
  XNOR U19612 ( .A(n19395), .B(n19392), .Z(n19419) );
  XOR U19613 ( .A(n19420), .B(n19419), .Z(c[250]) );
  NAND U19614 ( .A(n19397), .B(n19396), .Z(n19401) );
  NANDN U19615 ( .A(n19399), .B(n19398), .Z(n19400) );
  NAND U19616 ( .A(n19401), .B(n19400), .Z(n19432) );
  XOR U19617 ( .A(n585), .B(n19402), .Z(n19446) );
  NAND U19618 ( .A(n19446), .B(n19472), .Z(n19405) );
  NANDN U19619 ( .A(n19403), .B(n19473), .Z(n19404) );
  NAND U19620 ( .A(n19405), .B(n19404), .Z(n19435) );
  NAND U19621 ( .A(n19407), .B(n19406), .Z(n19409) );
  XOR U19622 ( .A(b[29]), .B(n19502), .Z(n19443) );
  OR U19623 ( .A(n19443), .B(n576), .Z(n19408) );
  AND U19624 ( .A(n19409), .B(n19408), .Z(n19436) );
  XNOR U19625 ( .A(n19435), .B(n19436), .Z(n19437) );
  NANDN U19626 ( .A(n585), .B(a[123]), .Z(n19449) );
  XOR U19627 ( .A(n19450), .B(n19449), .Z(n19452) );
  XNOR U19628 ( .A(n19451), .B(n19452), .Z(n19438) );
  XOR U19629 ( .A(n19437), .B(n19438), .Z(n19429) );
  XNOR U19630 ( .A(n19429), .B(n19430), .Z(n19431) );
  XOR U19631 ( .A(n19432), .B(n19431), .Z(n19423) );
  NANDN U19632 ( .A(n19414), .B(n19413), .Z(n19418) );
  OR U19633 ( .A(n19416), .B(n19415), .Z(n19417) );
  NAND U19634 ( .A(n19418), .B(n19417), .Z(n19424) );
  XNOR U19635 ( .A(n19423), .B(n19424), .Z(n19426) );
  XOR U19636 ( .A(n19425), .B(n19426), .Z(n19421) );
  OR U19637 ( .A(n19420), .B(n19419), .Z(n19422) );
  XNOR U19638 ( .A(n19421), .B(n19422), .Z(c[251]) );
  NANDN U19639 ( .A(n19422), .B(n19421), .Z(n19457) );
  NANDN U19640 ( .A(n19424), .B(n19423), .Z(n19428) );
  NAND U19641 ( .A(n19426), .B(n19425), .Z(n19427) );
  NAND U19642 ( .A(n19428), .B(n19427), .Z(n19460) );
  NANDN U19643 ( .A(n19430), .B(n19429), .Z(n19434) );
  NANDN U19644 ( .A(n19432), .B(n19431), .Z(n19433) );
  AND U19645 ( .A(n19434), .B(n19433), .Z(n19459) );
  NANDN U19646 ( .A(n19436), .B(n19435), .Z(n19440) );
  NANDN U19647 ( .A(n19438), .B(n19437), .Z(n19439) );
  NAND U19648 ( .A(n19440), .B(n19439), .Z(n19464) );
  NANDN U19649 ( .A(n19441), .B(n576), .Z(n19442) );
  XOR U19650 ( .A(n584), .B(n19442), .Z(n19445) );
  NANDN U19651 ( .A(n575), .B(n19443), .Z(n19444) );
  AND U19652 ( .A(n19445), .B(n19444), .Z(n19467) );
  AND U19653 ( .A(a[124]), .B(b[31]), .Z(n19485) );
  XNOR U19654 ( .A(n19467), .B(n19485), .Z(n19468) );
  XOR U19655 ( .A(n585), .B(a[126]), .Z(n19474) );
  NANDN U19656 ( .A(n19474), .B(n19472), .Z(n19448) );
  NAND U19657 ( .A(n19473), .B(n19446), .Z(n19447) );
  NAND U19658 ( .A(n19448), .B(n19447), .Z(n19469) );
  XOR U19659 ( .A(n19468), .B(n19469), .Z(n19461) );
  OR U19660 ( .A(n19450), .B(n19449), .Z(n19454) );
  NAND U19661 ( .A(n19452), .B(n19451), .Z(n19453) );
  AND U19662 ( .A(n19454), .B(n19453), .Z(n19462) );
  XNOR U19663 ( .A(n19461), .B(n19462), .Z(n19463) );
  XOR U19664 ( .A(n19464), .B(n19463), .Z(n19458) );
  XOR U19665 ( .A(n19459), .B(n19458), .Z(n19455) );
  XOR U19666 ( .A(n19460), .B(n19455), .Z(n19456) );
  XNOR U19667 ( .A(n19457), .B(n19456), .Z(c[252]) );
  NANDN U19668 ( .A(n19457), .B(n19456), .Z(n19501) );
  NANDN U19669 ( .A(n19462), .B(n19461), .Z(n19466) );
  NAND U19670 ( .A(n19464), .B(n19463), .Z(n19465) );
  AND U19671 ( .A(n19466), .B(n19465), .Z(n19491) );
  NANDN U19672 ( .A(n585), .B(a[125]), .Z(n19484) );
  XNOR U19673 ( .A(n19483), .B(n19484), .Z(n19486) );
  XOR U19674 ( .A(n19485), .B(n19486), .Z(n19496) );
  NANDN U19675 ( .A(n19467), .B(n19485), .Z(n19471) );
  NANDN U19676 ( .A(n19469), .B(n19468), .Z(n19470) );
  NAND U19677 ( .A(n19471), .B(n19470), .Z(n19494) );
  XNOR U19678 ( .A(b[31]), .B(a[127]), .Z(n19479) );
  NANDN U19679 ( .A(n19479), .B(n19472), .Z(n19476) );
  NANDN U19680 ( .A(n19474), .B(n19473), .Z(n19475) );
  NAND U19681 ( .A(n19476), .B(n19475), .Z(n19493) );
  XNOR U19682 ( .A(n19494), .B(n19493), .Z(n19495) );
  XNOR U19683 ( .A(n19496), .B(n19495), .Z(n19490) );
  XNOR U19684 ( .A(n19491), .B(n19490), .Z(n19477) );
  XOR U19685 ( .A(n19492), .B(n19477), .Z(n19500) );
  XNOR U19686 ( .A(n19501), .B(n19500), .Z(c[253]) );
  NANDN U19687 ( .A(n584), .B(b[30]), .Z(n19478) );
  XOR U19688 ( .A(n585), .B(n19478), .Z(n19482) );
  XOR U19689 ( .A(b[30]), .B(n584), .Z(n19480) );
  NAND U19690 ( .A(n19480), .B(n19479), .Z(n19481) );
  AND U19691 ( .A(n19482), .B(n19481), .Z(n19508) );
  IV U19692 ( .A(n19508), .Z(n19506) );
  OR U19693 ( .A(n19484), .B(n19483), .Z(n19488) );
  NANDN U19694 ( .A(n19486), .B(n19485), .Z(n19487) );
  NAND U19695 ( .A(n19488), .B(n19487), .Z(n19509) );
  AND U19696 ( .A(b[31]), .B(a[126]), .Z(n19507) );
  XNOR U19697 ( .A(n19509), .B(n19507), .Z(n19489) );
  XOR U19698 ( .A(n19506), .B(n19489), .Z(n19505) );
  NANDN U19699 ( .A(n19494), .B(n19493), .Z(n19498) );
  NANDN U19700 ( .A(n19496), .B(n19495), .Z(n19497) );
  NAND U19701 ( .A(n19498), .B(n19497), .Z(n19503) );
  XOR U19702 ( .A(n19504), .B(n19503), .Z(n19499) );
  XNOR U19703 ( .A(n19505), .B(n19499), .Z(n19511) );
  NANDN U19704 ( .A(n19501), .B(n19500), .Z(n19510) );
  XNOR U19705 ( .A(n19511), .B(n19510), .Z(c[254]) );
endmodule

