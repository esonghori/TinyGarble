
module sum_N128_CC4 ( clk, rst, a, b, c );
  input [31:0] a;
  input [31:0] b;
  output [31:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, \ADD_/c[31] , \ADD_/c[30] , \ADD_/c[29] ,
         \ADD_/c[28] , \ADD_/c[27] , \ADD_/c[26] , \ADD_/c[25] , \ADD_/c[24] ,
         \ADD_/c[23] , \ADD_/c[22] , \ADD_/c[21] , \ADD_/c[20] , \ADD_/c[19] ,
         \ADD_/c[18] , \ADD_/c[17] , \ADD_/c[16] , \ADD_/c[15] , \ADD_/c[14] ,
         \ADD_/c[13] , \ADD_/c[12] , \ADD_/c[11] , \ADD_/c[10] , \ADD_/c[9] ,
         \ADD_/c[8] , \ADD_/c[7] , \ADD_/c[6] , \ADD_/c[5] , \ADD_/c[4] ,
         \ADD_/c[3] , \ADD_/c[2] , \ADD_/c[1] , \ADD_/FAINST[0].FA_/n3 ,
         \ADD_/FAINST[0].FA_/n2 , \ADD_/FAINST[0].FA_/n1 ,
         \ADD_/FAINST[31].FA_/n3 , \ADD_/FAINST[31].FA_/n2 ,
         \ADD_/FAINST[31].FA_/n1 , \ADD_/FAINST[30].FA_/n3 ,
         \ADD_/FAINST[30].FA_/n2 , \ADD_/FAINST[30].FA_/n1 ,
         \ADD_/FAINST[29].FA_/n3 , \ADD_/FAINST[29].FA_/n2 ,
         \ADD_/FAINST[29].FA_/n1 , \ADD_/FAINST[28].FA_/n3 ,
         \ADD_/FAINST[28].FA_/n2 , \ADD_/FAINST[28].FA_/n1 ,
         \ADD_/FAINST[27].FA_/n3 , \ADD_/FAINST[27].FA_/n2 ,
         \ADD_/FAINST[27].FA_/n1 , \ADD_/FAINST[26].FA_/n3 ,
         \ADD_/FAINST[26].FA_/n2 , \ADD_/FAINST[26].FA_/n1 ,
         \ADD_/FAINST[25].FA_/n3 , \ADD_/FAINST[25].FA_/n2 ,
         \ADD_/FAINST[25].FA_/n1 , \ADD_/FAINST[24].FA_/n3 ,
         \ADD_/FAINST[24].FA_/n2 , \ADD_/FAINST[24].FA_/n1 ,
         \ADD_/FAINST[23].FA_/n3 , \ADD_/FAINST[23].FA_/n2 ,
         \ADD_/FAINST[23].FA_/n1 , \ADD_/FAINST[22].FA_/n3 ,
         \ADD_/FAINST[22].FA_/n2 , \ADD_/FAINST[22].FA_/n1 ,
         \ADD_/FAINST[21].FA_/n3 , \ADD_/FAINST[21].FA_/n2 ,
         \ADD_/FAINST[21].FA_/n1 , \ADD_/FAINST[20].FA_/n3 ,
         \ADD_/FAINST[20].FA_/n2 , \ADD_/FAINST[20].FA_/n1 ,
         \ADD_/FAINST[19].FA_/n3 , \ADD_/FAINST[19].FA_/n2 ,
         \ADD_/FAINST[19].FA_/n1 , \ADD_/FAINST[18].FA_/n3 ,
         \ADD_/FAINST[18].FA_/n2 , \ADD_/FAINST[18].FA_/n1 ,
         \ADD_/FAINST[17].FA_/n3 , \ADD_/FAINST[17].FA_/n2 ,
         \ADD_/FAINST[17].FA_/n1 , \ADD_/FAINST[16].FA_/n3 ,
         \ADD_/FAINST[16].FA_/n2 , \ADD_/FAINST[16].FA_/n1 ,
         \ADD_/FAINST[15].FA_/n3 , \ADD_/FAINST[15].FA_/n2 ,
         \ADD_/FAINST[15].FA_/n1 , \ADD_/FAINST[14].FA_/n3 ,
         \ADD_/FAINST[14].FA_/n2 , \ADD_/FAINST[14].FA_/n1 ,
         \ADD_/FAINST[13].FA_/n3 , \ADD_/FAINST[13].FA_/n2 ,
         \ADD_/FAINST[13].FA_/n1 , \ADD_/FAINST[12].FA_/n3 ,
         \ADD_/FAINST[12].FA_/n2 , \ADD_/FAINST[12].FA_/n1 ,
         \ADD_/FAINST[11].FA_/n3 , \ADD_/FAINST[11].FA_/n2 ,
         \ADD_/FAINST[11].FA_/n1 , \ADD_/FAINST[10].FA_/n3 ,
         \ADD_/FAINST[10].FA_/n2 , \ADD_/FAINST[10].FA_/n1 ,
         \ADD_/FAINST[9].FA_/n3 , \ADD_/FAINST[9].FA_/n2 ,
         \ADD_/FAINST[9].FA_/n1 , \ADD_/FAINST[8].FA_/n3 ,
         \ADD_/FAINST[8].FA_/n2 , \ADD_/FAINST[8].FA_/n1 ,
         \ADD_/FAINST[7].FA_/n3 , \ADD_/FAINST[7].FA_/n2 ,
         \ADD_/FAINST[7].FA_/n1 , \ADD_/FAINST[6].FA_/n3 ,
         \ADD_/FAINST[6].FA_/n2 , \ADD_/FAINST[6].FA_/n1 ,
         \ADD_/FAINST[5].FA_/n3 , \ADD_/FAINST[5].FA_/n2 ,
         \ADD_/FAINST[5].FA_/n1 , \ADD_/FAINST[4].FA_/n3 ,
         \ADD_/FAINST[4].FA_/n2 , \ADD_/FAINST[4].FA_/n1 ,
         \ADD_/FAINST[3].FA_/n3 , \ADD_/FAINST[3].FA_/n2 ,
         \ADD_/FAINST[3].FA_/n1 , \ADD_/FAINST[2].FA_/n3 ,
         \ADD_/FAINST[2].FA_/n2 , \ADD_/FAINST[2].FA_/n1 ,
         \ADD_/FAINST[1].FA_/n3 , \ADD_/FAINST[1].FA_/n2 ,
         \ADD_/FAINST[1].FA_/n1 ;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR \ADD_/FAINST[0].FA_/U5  ( .A(\ADD_/FAINST[0].FA_/n3 ), .B(carry_on), .Z(
        \ADD_/c[1] ) );
  XOR \ADD_/FAINST[0].FA_/U4  ( .A(\ADD_/FAINST[0].FA_/n1 ), .B(b[0]), .Z(c[0]) );
  AND \ADD_/FAINST[0].FA_/U3  ( .A(\ADD_/FAINST[0].FA_/n1 ), .B(
        \ADD_/FAINST[0].FA_/n2 ), .Z(\ADD_/FAINST[0].FA_/n3 ) );
  XOR \ADD_/FAINST[0].FA_/U2  ( .A(b[0]), .B(carry_on), .Z(
        \ADD_/FAINST[0].FA_/n2 ) );
  XOR \ADD_/FAINST[0].FA_/U1  ( .A(a[0]), .B(carry_on), .Z(
        \ADD_/FAINST[0].FA_/n1 ) );
  XOR \ADD_/FAINST[31].FA_/U5  ( .A(\ADD_/FAINST[31].FA_/n3 ), .B(\ADD_/c[31] ), .Z(carry_on_d) );
  XOR \ADD_/FAINST[31].FA_/U4  ( .A(\ADD_/FAINST[31].FA_/n1 ), .B(b[31]), .Z(
        c[31]) );
  AND \ADD_/FAINST[31].FA_/U3  ( .A(\ADD_/FAINST[31].FA_/n1 ), .B(
        \ADD_/FAINST[31].FA_/n2 ), .Z(\ADD_/FAINST[31].FA_/n3 ) );
  XOR \ADD_/FAINST[31].FA_/U2  ( .A(b[31]), .B(\ADD_/c[31] ), .Z(
        \ADD_/FAINST[31].FA_/n2 ) );
  XOR \ADD_/FAINST[31].FA_/U1  ( .A(a[31]), .B(\ADD_/c[31] ), .Z(
        \ADD_/FAINST[31].FA_/n1 ) );
  XOR \ADD_/FAINST[30].FA_/U5  ( .A(\ADD_/FAINST[30].FA_/n3 ), .B(\ADD_/c[30] ), .Z(\ADD_/c[31] ) );
  XOR \ADD_/FAINST[30].FA_/U4  ( .A(\ADD_/FAINST[30].FA_/n1 ), .B(b[30]), .Z(
        c[30]) );
  AND \ADD_/FAINST[30].FA_/U3  ( .A(\ADD_/FAINST[30].FA_/n1 ), .B(
        \ADD_/FAINST[30].FA_/n2 ), .Z(\ADD_/FAINST[30].FA_/n3 ) );
  XOR \ADD_/FAINST[30].FA_/U2  ( .A(b[30]), .B(\ADD_/c[30] ), .Z(
        \ADD_/FAINST[30].FA_/n2 ) );
  XOR \ADD_/FAINST[30].FA_/U1  ( .A(a[30]), .B(\ADD_/c[30] ), .Z(
        \ADD_/FAINST[30].FA_/n1 ) );
  XOR \ADD_/FAINST[29].FA_/U5  ( .A(\ADD_/FAINST[29].FA_/n3 ), .B(\ADD_/c[29] ), .Z(\ADD_/c[30] ) );
  XOR \ADD_/FAINST[29].FA_/U4  ( .A(\ADD_/FAINST[29].FA_/n1 ), .B(b[29]), .Z(
        c[29]) );
  AND \ADD_/FAINST[29].FA_/U3  ( .A(\ADD_/FAINST[29].FA_/n1 ), .B(
        \ADD_/FAINST[29].FA_/n2 ), .Z(\ADD_/FAINST[29].FA_/n3 ) );
  XOR \ADD_/FAINST[29].FA_/U2  ( .A(b[29]), .B(\ADD_/c[29] ), .Z(
        \ADD_/FAINST[29].FA_/n2 ) );
  XOR \ADD_/FAINST[29].FA_/U1  ( .A(a[29]), .B(\ADD_/c[29] ), .Z(
        \ADD_/FAINST[29].FA_/n1 ) );
  XOR \ADD_/FAINST[28].FA_/U5  ( .A(\ADD_/FAINST[28].FA_/n3 ), .B(\ADD_/c[28] ), .Z(\ADD_/c[29] ) );
  XOR \ADD_/FAINST[28].FA_/U4  ( .A(\ADD_/FAINST[28].FA_/n1 ), .B(b[28]), .Z(
        c[28]) );
  AND \ADD_/FAINST[28].FA_/U3  ( .A(\ADD_/FAINST[28].FA_/n1 ), .B(
        \ADD_/FAINST[28].FA_/n2 ), .Z(\ADD_/FAINST[28].FA_/n3 ) );
  XOR \ADD_/FAINST[28].FA_/U2  ( .A(b[28]), .B(\ADD_/c[28] ), .Z(
        \ADD_/FAINST[28].FA_/n2 ) );
  XOR \ADD_/FAINST[28].FA_/U1  ( .A(a[28]), .B(\ADD_/c[28] ), .Z(
        \ADD_/FAINST[28].FA_/n1 ) );
  XOR \ADD_/FAINST[27].FA_/U5  ( .A(\ADD_/FAINST[27].FA_/n3 ), .B(\ADD_/c[27] ), .Z(\ADD_/c[28] ) );
  XOR \ADD_/FAINST[27].FA_/U4  ( .A(\ADD_/FAINST[27].FA_/n1 ), .B(b[27]), .Z(
        c[27]) );
  AND \ADD_/FAINST[27].FA_/U3  ( .A(\ADD_/FAINST[27].FA_/n1 ), .B(
        \ADD_/FAINST[27].FA_/n2 ), .Z(\ADD_/FAINST[27].FA_/n3 ) );
  XOR \ADD_/FAINST[27].FA_/U2  ( .A(b[27]), .B(\ADD_/c[27] ), .Z(
        \ADD_/FAINST[27].FA_/n2 ) );
  XOR \ADD_/FAINST[27].FA_/U1  ( .A(a[27]), .B(\ADD_/c[27] ), .Z(
        \ADD_/FAINST[27].FA_/n1 ) );
  XOR \ADD_/FAINST[26].FA_/U5  ( .A(\ADD_/FAINST[26].FA_/n3 ), .B(\ADD_/c[26] ), .Z(\ADD_/c[27] ) );
  XOR \ADD_/FAINST[26].FA_/U4  ( .A(\ADD_/FAINST[26].FA_/n1 ), .B(b[26]), .Z(
        c[26]) );
  AND \ADD_/FAINST[26].FA_/U3  ( .A(\ADD_/FAINST[26].FA_/n1 ), .B(
        \ADD_/FAINST[26].FA_/n2 ), .Z(\ADD_/FAINST[26].FA_/n3 ) );
  XOR \ADD_/FAINST[26].FA_/U2  ( .A(b[26]), .B(\ADD_/c[26] ), .Z(
        \ADD_/FAINST[26].FA_/n2 ) );
  XOR \ADD_/FAINST[26].FA_/U1  ( .A(a[26]), .B(\ADD_/c[26] ), .Z(
        \ADD_/FAINST[26].FA_/n1 ) );
  XOR \ADD_/FAINST[25].FA_/U5  ( .A(\ADD_/FAINST[25].FA_/n3 ), .B(\ADD_/c[25] ), .Z(\ADD_/c[26] ) );
  XOR \ADD_/FAINST[25].FA_/U4  ( .A(\ADD_/FAINST[25].FA_/n1 ), .B(b[25]), .Z(
        c[25]) );
  AND \ADD_/FAINST[25].FA_/U3  ( .A(\ADD_/FAINST[25].FA_/n1 ), .B(
        \ADD_/FAINST[25].FA_/n2 ), .Z(\ADD_/FAINST[25].FA_/n3 ) );
  XOR \ADD_/FAINST[25].FA_/U2  ( .A(b[25]), .B(\ADD_/c[25] ), .Z(
        \ADD_/FAINST[25].FA_/n2 ) );
  XOR \ADD_/FAINST[25].FA_/U1  ( .A(a[25]), .B(\ADD_/c[25] ), .Z(
        \ADD_/FAINST[25].FA_/n1 ) );
  XOR \ADD_/FAINST[24].FA_/U5  ( .A(\ADD_/FAINST[24].FA_/n3 ), .B(\ADD_/c[24] ), .Z(\ADD_/c[25] ) );
  XOR \ADD_/FAINST[24].FA_/U4  ( .A(\ADD_/FAINST[24].FA_/n1 ), .B(b[24]), .Z(
        c[24]) );
  AND \ADD_/FAINST[24].FA_/U3  ( .A(\ADD_/FAINST[24].FA_/n1 ), .B(
        \ADD_/FAINST[24].FA_/n2 ), .Z(\ADD_/FAINST[24].FA_/n3 ) );
  XOR \ADD_/FAINST[24].FA_/U2  ( .A(b[24]), .B(\ADD_/c[24] ), .Z(
        \ADD_/FAINST[24].FA_/n2 ) );
  XOR \ADD_/FAINST[24].FA_/U1  ( .A(a[24]), .B(\ADD_/c[24] ), .Z(
        \ADD_/FAINST[24].FA_/n1 ) );
  XOR \ADD_/FAINST[23].FA_/U5  ( .A(\ADD_/FAINST[23].FA_/n3 ), .B(\ADD_/c[23] ), .Z(\ADD_/c[24] ) );
  XOR \ADD_/FAINST[23].FA_/U4  ( .A(\ADD_/FAINST[23].FA_/n1 ), .B(b[23]), .Z(
        c[23]) );
  AND \ADD_/FAINST[23].FA_/U3  ( .A(\ADD_/FAINST[23].FA_/n1 ), .B(
        \ADD_/FAINST[23].FA_/n2 ), .Z(\ADD_/FAINST[23].FA_/n3 ) );
  XOR \ADD_/FAINST[23].FA_/U2  ( .A(b[23]), .B(\ADD_/c[23] ), .Z(
        \ADD_/FAINST[23].FA_/n2 ) );
  XOR \ADD_/FAINST[23].FA_/U1  ( .A(a[23]), .B(\ADD_/c[23] ), .Z(
        \ADD_/FAINST[23].FA_/n1 ) );
  XOR \ADD_/FAINST[22].FA_/U5  ( .A(\ADD_/FAINST[22].FA_/n3 ), .B(\ADD_/c[22] ), .Z(\ADD_/c[23] ) );
  XOR \ADD_/FAINST[22].FA_/U4  ( .A(\ADD_/FAINST[22].FA_/n1 ), .B(b[22]), .Z(
        c[22]) );
  AND \ADD_/FAINST[22].FA_/U3  ( .A(\ADD_/FAINST[22].FA_/n1 ), .B(
        \ADD_/FAINST[22].FA_/n2 ), .Z(\ADD_/FAINST[22].FA_/n3 ) );
  XOR \ADD_/FAINST[22].FA_/U2  ( .A(b[22]), .B(\ADD_/c[22] ), .Z(
        \ADD_/FAINST[22].FA_/n2 ) );
  XOR \ADD_/FAINST[22].FA_/U1  ( .A(a[22]), .B(\ADD_/c[22] ), .Z(
        \ADD_/FAINST[22].FA_/n1 ) );
  XOR \ADD_/FAINST[21].FA_/U5  ( .A(\ADD_/FAINST[21].FA_/n3 ), .B(\ADD_/c[21] ), .Z(\ADD_/c[22] ) );
  XOR \ADD_/FAINST[21].FA_/U4  ( .A(\ADD_/FAINST[21].FA_/n1 ), .B(b[21]), .Z(
        c[21]) );
  AND \ADD_/FAINST[21].FA_/U3  ( .A(\ADD_/FAINST[21].FA_/n1 ), .B(
        \ADD_/FAINST[21].FA_/n2 ), .Z(\ADD_/FAINST[21].FA_/n3 ) );
  XOR \ADD_/FAINST[21].FA_/U2  ( .A(b[21]), .B(\ADD_/c[21] ), .Z(
        \ADD_/FAINST[21].FA_/n2 ) );
  XOR \ADD_/FAINST[21].FA_/U1  ( .A(a[21]), .B(\ADD_/c[21] ), .Z(
        \ADD_/FAINST[21].FA_/n1 ) );
  XOR \ADD_/FAINST[20].FA_/U5  ( .A(\ADD_/FAINST[20].FA_/n3 ), .B(\ADD_/c[20] ), .Z(\ADD_/c[21] ) );
  XOR \ADD_/FAINST[20].FA_/U4  ( .A(\ADD_/FAINST[20].FA_/n1 ), .B(b[20]), .Z(
        c[20]) );
  AND \ADD_/FAINST[20].FA_/U3  ( .A(\ADD_/FAINST[20].FA_/n1 ), .B(
        \ADD_/FAINST[20].FA_/n2 ), .Z(\ADD_/FAINST[20].FA_/n3 ) );
  XOR \ADD_/FAINST[20].FA_/U2  ( .A(b[20]), .B(\ADD_/c[20] ), .Z(
        \ADD_/FAINST[20].FA_/n2 ) );
  XOR \ADD_/FAINST[20].FA_/U1  ( .A(a[20]), .B(\ADD_/c[20] ), .Z(
        \ADD_/FAINST[20].FA_/n1 ) );
  XOR \ADD_/FAINST[19].FA_/U5  ( .A(\ADD_/FAINST[19].FA_/n3 ), .B(\ADD_/c[19] ), .Z(\ADD_/c[20] ) );
  XOR \ADD_/FAINST[19].FA_/U4  ( .A(\ADD_/FAINST[19].FA_/n1 ), .B(b[19]), .Z(
        c[19]) );
  AND \ADD_/FAINST[19].FA_/U3  ( .A(\ADD_/FAINST[19].FA_/n1 ), .B(
        \ADD_/FAINST[19].FA_/n2 ), .Z(\ADD_/FAINST[19].FA_/n3 ) );
  XOR \ADD_/FAINST[19].FA_/U2  ( .A(b[19]), .B(\ADD_/c[19] ), .Z(
        \ADD_/FAINST[19].FA_/n2 ) );
  XOR \ADD_/FAINST[19].FA_/U1  ( .A(a[19]), .B(\ADD_/c[19] ), .Z(
        \ADD_/FAINST[19].FA_/n1 ) );
  XOR \ADD_/FAINST[18].FA_/U5  ( .A(\ADD_/FAINST[18].FA_/n3 ), .B(\ADD_/c[18] ), .Z(\ADD_/c[19] ) );
  XOR \ADD_/FAINST[18].FA_/U4  ( .A(\ADD_/FAINST[18].FA_/n1 ), .B(b[18]), .Z(
        c[18]) );
  AND \ADD_/FAINST[18].FA_/U3  ( .A(\ADD_/FAINST[18].FA_/n1 ), .B(
        \ADD_/FAINST[18].FA_/n2 ), .Z(\ADD_/FAINST[18].FA_/n3 ) );
  XOR \ADD_/FAINST[18].FA_/U2  ( .A(b[18]), .B(\ADD_/c[18] ), .Z(
        \ADD_/FAINST[18].FA_/n2 ) );
  XOR \ADD_/FAINST[18].FA_/U1  ( .A(a[18]), .B(\ADD_/c[18] ), .Z(
        \ADD_/FAINST[18].FA_/n1 ) );
  XOR \ADD_/FAINST[17].FA_/U5  ( .A(\ADD_/FAINST[17].FA_/n3 ), .B(\ADD_/c[17] ), .Z(\ADD_/c[18] ) );
  XOR \ADD_/FAINST[17].FA_/U4  ( .A(\ADD_/FAINST[17].FA_/n1 ), .B(b[17]), .Z(
        c[17]) );
  AND \ADD_/FAINST[17].FA_/U3  ( .A(\ADD_/FAINST[17].FA_/n1 ), .B(
        \ADD_/FAINST[17].FA_/n2 ), .Z(\ADD_/FAINST[17].FA_/n3 ) );
  XOR \ADD_/FAINST[17].FA_/U2  ( .A(b[17]), .B(\ADD_/c[17] ), .Z(
        \ADD_/FAINST[17].FA_/n2 ) );
  XOR \ADD_/FAINST[17].FA_/U1  ( .A(a[17]), .B(\ADD_/c[17] ), .Z(
        \ADD_/FAINST[17].FA_/n1 ) );
  XOR \ADD_/FAINST[16].FA_/U5  ( .A(\ADD_/FAINST[16].FA_/n3 ), .B(\ADD_/c[16] ), .Z(\ADD_/c[17] ) );
  XOR \ADD_/FAINST[16].FA_/U4  ( .A(\ADD_/FAINST[16].FA_/n1 ), .B(b[16]), .Z(
        c[16]) );
  AND \ADD_/FAINST[16].FA_/U3  ( .A(\ADD_/FAINST[16].FA_/n1 ), .B(
        \ADD_/FAINST[16].FA_/n2 ), .Z(\ADD_/FAINST[16].FA_/n3 ) );
  XOR \ADD_/FAINST[16].FA_/U2  ( .A(b[16]), .B(\ADD_/c[16] ), .Z(
        \ADD_/FAINST[16].FA_/n2 ) );
  XOR \ADD_/FAINST[16].FA_/U1  ( .A(a[16]), .B(\ADD_/c[16] ), .Z(
        \ADD_/FAINST[16].FA_/n1 ) );
  XOR \ADD_/FAINST[15].FA_/U5  ( .A(\ADD_/FAINST[15].FA_/n3 ), .B(\ADD_/c[15] ), .Z(\ADD_/c[16] ) );
  XOR \ADD_/FAINST[15].FA_/U4  ( .A(\ADD_/FAINST[15].FA_/n1 ), .B(b[15]), .Z(
        c[15]) );
  AND \ADD_/FAINST[15].FA_/U3  ( .A(\ADD_/FAINST[15].FA_/n1 ), .B(
        \ADD_/FAINST[15].FA_/n2 ), .Z(\ADD_/FAINST[15].FA_/n3 ) );
  XOR \ADD_/FAINST[15].FA_/U2  ( .A(b[15]), .B(\ADD_/c[15] ), .Z(
        \ADD_/FAINST[15].FA_/n2 ) );
  XOR \ADD_/FAINST[15].FA_/U1  ( .A(a[15]), .B(\ADD_/c[15] ), .Z(
        \ADD_/FAINST[15].FA_/n1 ) );
  XOR \ADD_/FAINST[14].FA_/U5  ( .A(\ADD_/FAINST[14].FA_/n3 ), .B(\ADD_/c[14] ), .Z(\ADD_/c[15] ) );
  XOR \ADD_/FAINST[14].FA_/U4  ( .A(\ADD_/FAINST[14].FA_/n1 ), .B(b[14]), .Z(
        c[14]) );
  AND \ADD_/FAINST[14].FA_/U3  ( .A(\ADD_/FAINST[14].FA_/n1 ), .B(
        \ADD_/FAINST[14].FA_/n2 ), .Z(\ADD_/FAINST[14].FA_/n3 ) );
  XOR \ADD_/FAINST[14].FA_/U2  ( .A(b[14]), .B(\ADD_/c[14] ), .Z(
        \ADD_/FAINST[14].FA_/n2 ) );
  XOR \ADD_/FAINST[14].FA_/U1  ( .A(a[14]), .B(\ADD_/c[14] ), .Z(
        \ADD_/FAINST[14].FA_/n1 ) );
  XOR \ADD_/FAINST[13].FA_/U5  ( .A(\ADD_/FAINST[13].FA_/n3 ), .B(\ADD_/c[13] ), .Z(\ADD_/c[14] ) );
  XOR \ADD_/FAINST[13].FA_/U4  ( .A(\ADD_/FAINST[13].FA_/n1 ), .B(b[13]), .Z(
        c[13]) );
  AND \ADD_/FAINST[13].FA_/U3  ( .A(\ADD_/FAINST[13].FA_/n1 ), .B(
        \ADD_/FAINST[13].FA_/n2 ), .Z(\ADD_/FAINST[13].FA_/n3 ) );
  XOR \ADD_/FAINST[13].FA_/U2  ( .A(b[13]), .B(\ADD_/c[13] ), .Z(
        \ADD_/FAINST[13].FA_/n2 ) );
  XOR \ADD_/FAINST[13].FA_/U1  ( .A(a[13]), .B(\ADD_/c[13] ), .Z(
        \ADD_/FAINST[13].FA_/n1 ) );
  XOR \ADD_/FAINST[12].FA_/U5  ( .A(\ADD_/FAINST[12].FA_/n3 ), .B(\ADD_/c[12] ), .Z(\ADD_/c[13] ) );
  XOR \ADD_/FAINST[12].FA_/U4  ( .A(\ADD_/FAINST[12].FA_/n1 ), .B(b[12]), .Z(
        c[12]) );
  AND \ADD_/FAINST[12].FA_/U3  ( .A(\ADD_/FAINST[12].FA_/n1 ), .B(
        \ADD_/FAINST[12].FA_/n2 ), .Z(\ADD_/FAINST[12].FA_/n3 ) );
  XOR \ADD_/FAINST[12].FA_/U2  ( .A(b[12]), .B(\ADD_/c[12] ), .Z(
        \ADD_/FAINST[12].FA_/n2 ) );
  XOR \ADD_/FAINST[12].FA_/U1  ( .A(a[12]), .B(\ADD_/c[12] ), .Z(
        \ADD_/FAINST[12].FA_/n1 ) );
  XOR \ADD_/FAINST[11].FA_/U5  ( .A(\ADD_/FAINST[11].FA_/n3 ), .B(\ADD_/c[11] ), .Z(\ADD_/c[12] ) );
  XOR \ADD_/FAINST[11].FA_/U4  ( .A(\ADD_/FAINST[11].FA_/n1 ), .B(b[11]), .Z(
        c[11]) );
  AND \ADD_/FAINST[11].FA_/U3  ( .A(\ADD_/FAINST[11].FA_/n1 ), .B(
        \ADD_/FAINST[11].FA_/n2 ), .Z(\ADD_/FAINST[11].FA_/n3 ) );
  XOR \ADD_/FAINST[11].FA_/U2  ( .A(b[11]), .B(\ADD_/c[11] ), .Z(
        \ADD_/FAINST[11].FA_/n2 ) );
  XOR \ADD_/FAINST[11].FA_/U1  ( .A(a[11]), .B(\ADD_/c[11] ), .Z(
        \ADD_/FAINST[11].FA_/n1 ) );
  XOR \ADD_/FAINST[10].FA_/U5  ( .A(\ADD_/FAINST[10].FA_/n3 ), .B(\ADD_/c[10] ), .Z(\ADD_/c[11] ) );
  XOR \ADD_/FAINST[10].FA_/U4  ( .A(\ADD_/FAINST[10].FA_/n1 ), .B(b[10]), .Z(
        c[10]) );
  AND \ADD_/FAINST[10].FA_/U3  ( .A(\ADD_/FAINST[10].FA_/n1 ), .B(
        \ADD_/FAINST[10].FA_/n2 ), .Z(\ADD_/FAINST[10].FA_/n3 ) );
  XOR \ADD_/FAINST[10].FA_/U2  ( .A(b[10]), .B(\ADD_/c[10] ), .Z(
        \ADD_/FAINST[10].FA_/n2 ) );
  XOR \ADD_/FAINST[10].FA_/U1  ( .A(a[10]), .B(\ADD_/c[10] ), .Z(
        \ADD_/FAINST[10].FA_/n1 ) );
  XOR \ADD_/FAINST[9].FA_/U5  ( .A(\ADD_/FAINST[9].FA_/n3 ), .B(\ADD_/c[9] ), 
        .Z(\ADD_/c[10] ) );
  XOR \ADD_/FAINST[9].FA_/U4  ( .A(\ADD_/FAINST[9].FA_/n1 ), .B(b[9]), .Z(c[9]) );
  AND \ADD_/FAINST[9].FA_/U3  ( .A(\ADD_/FAINST[9].FA_/n1 ), .B(
        \ADD_/FAINST[9].FA_/n2 ), .Z(\ADD_/FAINST[9].FA_/n3 ) );
  XOR \ADD_/FAINST[9].FA_/U2  ( .A(b[9]), .B(\ADD_/c[9] ), .Z(
        \ADD_/FAINST[9].FA_/n2 ) );
  XOR \ADD_/FAINST[9].FA_/U1  ( .A(a[9]), .B(\ADD_/c[9] ), .Z(
        \ADD_/FAINST[9].FA_/n1 ) );
  XOR \ADD_/FAINST[8].FA_/U5  ( .A(\ADD_/FAINST[8].FA_/n3 ), .B(\ADD_/c[8] ), 
        .Z(\ADD_/c[9] ) );
  XOR \ADD_/FAINST[8].FA_/U4  ( .A(\ADD_/FAINST[8].FA_/n1 ), .B(b[8]), .Z(c[8]) );
  AND \ADD_/FAINST[8].FA_/U3  ( .A(\ADD_/FAINST[8].FA_/n1 ), .B(
        \ADD_/FAINST[8].FA_/n2 ), .Z(\ADD_/FAINST[8].FA_/n3 ) );
  XOR \ADD_/FAINST[8].FA_/U2  ( .A(b[8]), .B(\ADD_/c[8] ), .Z(
        \ADD_/FAINST[8].FA_/n2 ) );
  XOR \ADD_/FAINST[8].FA_/U1  ( .A(a[8]), .B(\ADD_/c[8] ), .Z(
        \ADD_/FAINST[8].FA_/n1 ) );
  XOR \ADD_/FAINST[7].FA_/U5  ( .A(\ADD_/FAINST[7].FA_/n3 ), .B(\ADD_/c[7] ), 
        .Z(\ADD_/c[8] ) );
  XOR \ADD_/FAINST[7].FA_/U4  ( .A(\ADD_/FAINST[7].FA_/n1 ), .B(b[7]), .Z(c[7]) );
  AND \ADD_/FAINST[7].FA_/U3  ( .A(\ADD_/FAINST[7].FA_/n1 ), .B(
        \ADD_/FAINST[7].FA_/n2 ), .Z(\ADD_/FAINST[7].FA_/n3 ) );
  XOR \ADD_/FAINST[7].FA_/U2  ( .A(b[7]), .B(\ADD_/c[7] ), .Z(
        \ADD_/FAINST[7].FA_/n2 ) );
  XOR \ADD_/FAINST[7].FA_/U1  ( .A(a[7]), .B(\ADD_/c[7] ), .Z(
        \ADD_/FAINST[7].FA_/n1 ) );
  XOR \ADD_/FAINST[6].FA_/U5  ( .A(\ADD_/FAINST[6].FA_/n3 ), .B(\ADD_/c[6] ), 
        .Z(\ADD_/c[7] ) );
  XOR \ADD_/FAINST[6].FA_/U4  ( .A(\ADD_/FAINST[6].FA_/n1 ), .B(b[6]), .Z(c[6]) );
  AND \ADD_/FAINST[6].FA_/U3  ( .A(\ADD_/FAINST[6].FA_/n1 ), .B(
        \ADD_/FAINST[6].FA_/n2 ), .Z(\ADD_/FAINST[6].FA_/n3 ) );
  XOR \ADD_/FAINST[6].FA_/U2  ( .A(b[6]), .B(\ADD_/c[6] ), .Z(
        \ADD_/FAINST[6].FA_/n2 ) );
  XOR \ADD_/FAINST[6].FA_/U1  ( .A(a[6]), .B(\ADD_/c[6] ), .Z(
        \ADD_/FAINST[6].FA_/n1 ) );
  XOR \ADD_/FAINST[5].FA_/U5  ( .A(\ADD_/FAINST[5].FA_/n3 ), .B(\ADD_/c[5] ), 
        .Z(\ADD_/c[6] ) );
  XOR \ADD_/FAINST[5].FA_/U4  ( .A(\ADD_/FAINST[5].FA_/n1 ), .B(b[5]), .Z(c[5]) );
  AND \ADD_/FAINST[5].FA_/U3  ( .A(\ADD_/FAINST[5].FA_/n1 ), .B(
        \ADD_/FAINST[5].FA_/n2 ), .Z(\ADD_/FAINST[5].FA_/n3 ) );
  XOR \ADD_/FAINST[5].FA_/U2  ( .A(b[5]), .B(\ADD_/c[5] ), .Z(
        \ADD_/FAINST[5].FA_/n2 ) );
  XOR \ADD_/FAINST[5].FA_/U1  ( .A(a[5]), .B(\ADD_/c[5] ), .Z(
        \ADD_/FAINST[5].FA_/n1 ) );
  XOR \ADD_/FAINST[4].FA_/U5  ( .A(\ADD_/FAINST[4].FA_/n3 ), .B(\ADD_/c[4] ), 
        .Z(\ADD_/c[5] ) );
  XOR \ADD_/FAINST[4].FA_/U4  ( .A(\ADD_/FAINST[4].FA_/n1 ), .B(b[4]), .Z(c[4]) );
  AND \ADD_/FAINST[4].FA_/U3  ( .A(\ADD_/FAINST[4].FA_/n1 ), .B(
        \ADD_/FAINST[4].FA_/n2 ), .Z(\ADD_/FAINST[4].FA_/n3 ) );
  XOR \ADD_/FAINST[4].FA_/U2  ( .A(b[4]), .B(\ADD_/c[4] ), .Z(
        \ADD_/FAINST[4].FA_/n2 ) );
  XOR \ADD_/FAINST[4].FA_/U1  ( .A(a[4]), .B(\ADD_/c[4] ), .Z(
        \ADD_/FAINST[4].FA_/n1 ) );
  XOR \ADD_/FAINST[3].FA_/U5  ( .A(\ADD_/FAINST[3].FA_/n3 ), .B(\ADD_/c[3] ), 
        .Z(\ADD_/c[4] ) );
  XOR \ADD_/FAINST[3].FA_/U4  ( .A(\ADD_/FAINST[3].FA_/n1 ), .B(b[3]), .Z(c[3]) );
  AND \ADD_/FAINST[3].FA_/U3  ( .A(\ADD_/FAINST[3].FA_/n1 ), .B(
        \ADD_/FAINST[3].FA_/n2 ), .Z(\ADD_/FAINST[3].FA_/n3 ) );
  XOR \ADD_/FAINST[3].FA_/U2  ( .A(b[3]), .B(\ADD_/c[3] ), .Z(
        \ADD_/FAINST[3].FA_/n2 ) );
  XOR \ADD_/FAINST[3].FA_/U1  ( .A(a[3]), .B(\ADD_/c[3] ), .Z(
        \ADD_/FAINST[3].FA_/n1 ) );
  XOR \ADD_/FAINST[2].FA_/U5  ( .A(\ADD_/FAINST[2].FA_/n3 ), .B(\ADD_/c[2] ), 
        .Z(\ADD_/c[3] ) );
  XOR \ADD_/FAINST[2].FA_/U4  ( .A(\ADD_/FAINST[2].FA_/n1 ), .B(b[2]), .Z(c[2]) );
  AND \ADD_/FAINST[2].FA_/U3  ( .A(\ADD_/FAINST[2].FA_/n1 ), .B(
        \ADD_/FAINST[2].FA_/n2 ), .Z(\ADD_/FAINST[2].FA_/n3 ) );
  XOR \ADD_/FAINST[2].FA_/U2  ( .A(b[2]), .B(\ADD_/c[2] ), .Z(
        \ADD_/FAINST[2].FA_/n2 ) );
  XOR \ADD_/FAINST[2].FA_/U1  ( .A(a[2]), .B(\ADD_/c[2] ), .Z(
        \ADD_/FAINST[2].FA_/n1 ) );
  XOR \ADD_/FAINST[1].FA_/U5  ( .A(\ADD_/FAINST[1].FA_/n3 ), .B(\ADD_/c[1] ), 
        .Z(\ADD_/c[2] ) );
  XOR \ADD_/FAINST[1].FA_/U4  ( .A(\ADD_/FAINST[1].FA_/n1 ), .B(b[1]), .Z(c[1]) );
  AND \ADD_/FAINST[1].FA_/U3  ( .A(\ADD_/FAINST[1].FA_/n1 ), .B(
        \ADD_/FAINST[1].FA_/n2 ), .Z(\ADD_/FAINST[1].FA_/n3 ) );
  XOR \ADD_/FAINST[1].FA_/U2  ( .A(b[1]), .B(\ADD_/c[1] ), .Z(
        \ADD_/FAINST[1].FA_/n2 ) );
  XOR \ADD_/FAINST[1].FA_/U1  ( .A(a[1]), .B(\ADD_/c[1] ), .Z(
        \ADD_/FAINST[1].FA_/n1 ) );
endmodule

