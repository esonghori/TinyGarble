
module sum_N16384_CC128 ( clk, rst, a, b, c );
  input [127:0] a;
  input [127:0] b;
  output [127:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        carry_on) );
  XOR U4 ( .A(n2), .B(n3), .Z(carry_on_d) );
  ANDN U5 ( .B(n4), .A(n5), .Z(n2) );
  XOR U6 ( .A(b[127]), .B(n3), .Z(n4) );
  XNOR U7 ( .A(b[9]), .B(n6), .Z(c[9]) );
  XNOR U8 ( .A(b[99]), .B(n7), .Z(c[99]) );
  XNOR U9 ( .A(b[98]), .B(n8), .Z(c[98]) );
  XNOR U10 ( .A(b[97]), .B(n9), .Z(c[97]) );
  XNOR U11 ( .A(b[96]), .B(n10), .Z(c[96]) );
  XNOR U12 ( .A(b[95]), .B(n11), .Z(c[95]) );
  XNOR U13 ( .A(b[94]), .B(n12), .Z(c[94]) );
  XNOR U14 ( .A(b[93]), .B(n13), .Z(c[93]) );
  XNOR U15 ( .A(b[92]), .B(n14), .Z(c[92]) );
  XNOR U16 ( .A(b[91]), .B(n15), .Z(c[91]) );
  XNOR U17 ( .A(b[90]), .B(n16), .Z(c[90]) );
  XNOR U18 ( .A(b[8]), .B(n17), .Z(c[8]) );
  XNOR U19 ( .A(b[89]), .B(n18), .Z(c[89]) );
  XNOR U20 ( .A(b[88]), .B(n19), .Z(c[88]) );
  XNOR U21 ( .A(b[87]), .B(n20), .Z(c[87]) );
  XNOR U22 ( .A(b[86]), .B(n21), .Z(c[86]) );
  XNOR U23 ( .A(b[85]), .B(n22), .Z(c[85]) );
  XNOR U24 ( .A(b[84]), .B(n23), .Z(c[84]) );
  XNOR U25 ( .A(b[83]), .B(n24), .Z(c[83]) );
  XNOR U26 ( .A(b[82]), .B(n25), .Z(c[82]) );
  XNOR U27 ( .A(b[81]), .B(n26), .Z(c[81]) );
  XNOR U28 ( .A(b[80]), .B(n27), .Z(c[80]) );
  XNOR U29 ( .A(b[7]), .B(n28), .Z(c[7]) );
  XNOR U30 ( .A(b[79]), .B(n29), .Z(c[79]) );
  XNOR U31 ( .A(b[78]), .B(n30), .Z(c[78]) );
  XNOR U32 ( .A(b[77]), .B(n31), .Z(c[77]) );
  XNOR U33 ( .A(b[76]), .B(n32), .Z(c[76]) );
  XNOR U34 ( .A(b[75]), .B(n33), .Z(c[75]) );
  XNOR U35 ( .A(b[74]), .B(n34), .Z(c[74]) );
  XNOR U36 ( .A(b[73]), .B(n35), .Z(c[73]) );
  XNOR U37 ( .A(b[72]), .B(n36), .Z(c[72]) );
  XNOR U38 ( .A(b[71]), .B(n37), .Z(c[71]) );
  XNOR U39 ( .A(b[70]), .B(n38), .Z(c[70]) );
  XNOR U40 ( .A(b[6]), .B(n39), .Z(c[6]) );
  XNOR U41 ( .A(b[69]), .B(n40), .Z(c[69]) );
  XNOR U42 ( .A(b[68]), .B(n41), .Z(c[68]) );
  XNOR U43 ( .A(b[67]), .B(n42), .Z(c[67]) );
  XNOR U44 ( .A(b[66]), .B(n43), .Z(c[66]) );
  XNOR U45 ( .A(b[65]), .B(n44), .Z(c[65]) );
  XNOR U46 ( .A(b[64]), .B(n45), .Z(c[64]) );
  XNOR U47 ( .A(b[63]), .B(n46), .Z(c[63]) );
  XNOR U48 ( .A(b[62]), .B(n47), .Z(c[62]) );
  XNOR U49 ( .A(b[61]), .B(n48), .Z(c[61]) );
  XNOR U50 ( .A(b[60]), .B(n49), .Z(c[60]) );
  XNOR U51 ( .A(b[5]), .B(n50), .Z(c[5]) );
  XNOR U52 ( .A(b[59]), .B(n51), .Z(c[59]) );
  XNOR U53 ( .A(b[58]), .B(n52), .Z(c[58]) );
  XNOR U54 ( .A(b[57]), .B(n53), .Z(c[57]) );
  XNOR U55 ( .A(b[56]), .B(n54), .Z(c[56]) );
  XNOR U56 ( .A(b[55]), .B(n55), .Z(c[55]) );
  XNOR U57 ( .A(b[54]), .B(n56), .Z(c[54]) );
  XNOR U58 ( .A(b[53]), .B(n57), .Z(c[53]) );
  XNOR U59 ( .A(b[52]), .B(n58), .Z(c[52]) );
  XNOR U60 ( .A(b[51]), .B(n59), .Z(c[51]) );
  XNOR U61 ( .A(b[50]), .B(n60), .Z(c[50]) );
  XNOR U62 ( .A(b[4]), .B(n61), .Z(c[4]) );
  XNOR U63 ( .A(b[49]), .B(n62), .Z(c[49]) );
  XNOR U64 ( .A(b[48]), .B(n63), .Z(c[48]) );
  XNOR U65 ( .A(b[47]), .B(n64), .Z(c[47]) );
  XNOR U66 ( .A(b[46]), .B(n65), .Z(c[46]) );
  XNOR U67 ( .A(b[45]), .B(n66), .Z(c[45]) );
  XNOR U68 ( .A(b[44]), .B(n67), .Z(c[44]) );
  XNOR U69 ( .A(b[43]), .B(n68), .Z(c[43]) );
  XNOR U70 ( .A(b[42]), .B(n69), .Z(c[42]) );
  XNOR U71 ( .A(b[41]), .B(n70), .Z(c[41]) );
  XNOR U72 ( .A(b[40]), .B(n71), .Z(c[40]) );
  XNOR U73 ( .A(b[3]), .B(n72), .Z(c[3]) );
  XNOR U74 ( .A(b[39]), .B(n73), .Z(c[39]) );
  XNOR U75 ( .A(b[38]), .B(n74), .Z(c[38]) );
  XNOR U76 ( .A(b[37]), .B(n75), .Z(c[37]) );
  XNOR U77 ( .A(b[36]), .B(n76), .Z(c[36]) );
  XNOR U78 ( .A(b[35]), .B(n77), .Z(c[35]) );
  XNOR U79 ( .A(b[34]), .B(n78), .Z(c[34]) );
  XNOR U80 ( .A(b[33]), .B(n79), .Z(c[33]) );
  XNOR U81 ( .A(b[32]), .B(n80), .Z(c[32]) );
  XNOR U82 ( .A(b[31]), .B(n81), .Z(c[31]) );
  XNOR U83 ( .A(b[30]), .B(n82), .Z(c[30]) );
  XNOR U84 ( .A(b[2]), .B(n83), .Z(c[2]) );
  XNOR U85 ( .A(b[29]), .B(n84), .Z(c[29]) );
  XNOR U86 ( .A(b[28]), .B(n85), .Z(c[28]) );
  XNOR U87 ( .A(b[27]), .B(n86), .Z(c[27]) );
  XNOR U88 ( .A(b[26]), .B(n87), .Z(c[26]) );
  XNOR U89 ( .A(b[25]), .B(n88), .Z(c[25]) );
  XNOR U90 ( .A(b[24]), .B(n89), .Z(c[24]) );
  XNOR U91 ( .A(b[23]), .B(n90), .Z(c[23]) );
  XNOR U92 ( .A(b[22]), .B(n91), .Z(c[22]) );
  XNOR U93 ( .A(b[21]), .B(n92), .Z(c[21]) );
  XNOR U94 ( .A(b[20]), .B(n93), .Z(c[20]) );
  XNOR U95 ( .A(b[1]), .B(n94), .Z(c[1]) );
  XNOR U96 ( .A(b[19]), .B(n95), .Z(c[19]) );
  XNOR U97 ( .A(b[18]), .B(n96), .Z(c[18]) );
  XNOR U98 ( .A(b[17]), .B(n97), .Z(c[17]) );
  XNOR U99 ( .A(b[16]), .B(n98), .Z(c[16]) );
  XNOR U100 ( .A(b[15]), .B(n99), .Z(c[15]) );
  XNOR U101 ( .A(b[14]), .B(n100), .Z(c[14]) );
  XNOR U102 ( .A(b[13]), .B(n101), .Z(c[13]) );
  XNOR U103 ( .A(b[12]), .B(n102), .Z(c[12]) );
  XNOR U104 ( .A(b[127]), .B(n5), .Z(c[127]) );
  XNOR U105 ( .A(a[127]), .B(n3), .Z(n5) );
  XNOR U106 ( .A(n103), .B(n104), .Z(n3) );
  ANDN U107 ( .B(n105), .A(n106), .Z(n103) );
  XNOR U108 ( .A(b[126]), .B(n104), .Z(n105) );
  XNOR U109 ( .A(b[126]), .B(n106), .Z(c[126]) );
  XNOR U110 ( .A(a[126]), .B(n107), .Z(n106) );
  IV U111 ( .A(n104), .Z(n107) );
  XOR U112 ( .A(n108), .B(n109), .Z(n104) );
  ANDN U113 ( .B(n110), .A(n111), .Z(n108) );
  XNOR U114 ( .A(b[125]), .B(n109), .Z(n110) );
  XNOR U115 ( .A(b[125]), .B(n111), .Z(c[125]) );
  XNOR U116 ( .A(a[125]), .B(n112), .Z(n111) );
  IV U117 ( .A(n109), .Z(n112) );
  XOR U118 ( .A(n113), .B(n114), .Z(n109) );
  ANDN U119 ( .B(n115), .A(n116), .Z(n113) );
  XNOR U120 ( .A(b[124]), .B(n114), .Z(n115) );
  XNOR U121 ( .A(b[124]), .B(n116), .Z(c[124]) );
  XNOR U122 ( .A(a[124]), .B(n117), .Z(n116) );
  IV U123 ( .A(n114), .Z(n117) );
  XOR U124 ( .A(n118), .B(n119), .Z(n114) );
  ANDN U125 ( .B(n120), .A(n121), .Z(n118) );
  XNOR U126 ( .A(b[123]), .B(n119), .Z(n120) );
  XNOR U127 ( .A(b[123]), .B(n121), .Z(c[123]) );
  XNOR U128 ( .A(a[123]), .B(n122), .Z(n121) );
  IV U129 ( .A(n119), .Z(n122) );
  XOR U130 ( .A(n123), .B(n124), .Z(n119) );
  ANDN U131 ( .B(n125), .A(n126), .Z(n123) );
  XNOR U132 ( .A(b[122]), .B(n124), .Z(n125) );
  XNOR U133 ( .A(b[122]), .B(n126), .Z(c[122]) );
  XNOR U134 ( .A(a[122]), .B(n127), .Z(n126) );
  IV U135 ( .A(n124), .Z(n127) );
  XOR U136 ( .A(n128), .B(n129), .Z(n124) );
  ANDN U137 ( .B(n130), .A(n131), .Z(n128) );
  XNOR U138 ( .A(b[121]), .B(n129), .Z(n130) );
  XNOR U139 ( .A(b[121]), .B(n131), .Z(c[121]) );
  XNOR U140 ( .A(a[121]), .B(n132), .Z(n131) );
  IV U141 ( .A(n129), .Z(n132) );
  XOR U142 ( .A(n133), .B(n134), .Z(n129) );
  ANDN U143 ( .B(n135), .A(n136), .Z(n133) );
  XNOR U144 ( .A(b[120]), .B(n134), .Z(n135) );
  XNOR U145 ( .A(b[120]), .B(n136), .Z(c[120]) );
  XNOR U146 ( .A(a[120]), .B(n137), .Z(n136) );
  IV U147 ( .A(n134), .Z(n137) );
  XOR U148 ( .A(n138), .B(n139), .Z(n134) );
  ANDN U149 ( .B(n140), .A(n141), .Z(n138) );
  XNOR U150 ( .A(b[119]), .B(n139), .Z(n140) );
  XNOR U151 ( .A(b[11]), .B(n142), .Z(c[11]) );
  XNOR U152 ( .A(b[119]), .B(n141), .Z(c[119]) );
  XNOR U153 ( .A(a[119]), .B(n143), .Z(n141) );
  IV U154 ( .A(n139), .Z(n143) );
  XOR U155 ( .A(n144), .B(n145), .Z(n139) );
  ANDN U156 ( .B(n146), .A(n147), .Z(n144) );
  XNOR U157 ( .A(b[118]), .B(n145), .Z(n146) );
  XNOR U158 ( .A(b[118]), .B(n147), .Z(c[118]) );
  XNOR U159 ( .A(a[118]), .B(n148), .Z(n147) );
  IV U160 ( .A(n145), .Z(n148) );
  XOR U161 ( .A(n149), .B(n150), .Z(n145) );
  ANDN U162 ( .B(n151), .A(n152), .Z(n149) );
  XNOR U163 ( .A(b[117]), .B(n150), .Z(n151) );
  XNOR U164 ( .A(b[117]), .B(n152), .Z(c[117]) );
  XNOR U165 ( .A(a[117]), .B(n153), .Z(n152) );
  IV U166 ( .A(n150), .Z(n153) );
  XOR U167 ( .A(n154), .B(n155), .Z(n150) );
  ANDN U168 ( .B(n156), .A(n157), .Z(n154) );
  XNOR U169 ( .A(b[116]), .B(n155), .Z(n156) );
  XNOR U170 ( .A(b[116]), .B(n157), .Z(c[116]) );
  XNOR U171 ( .A(a[116]), .B(n158), .Z(n157) );
  IV U172 ( .A(n155), .Z(n158) );
  XOR U173 ( .A(n159), .B(n160), .Z(n155) );
  ANDN U174 ( .B(n161), .A(n162), .Z(n159) );
  XNOR U175 ( .A(b[115]), .B(n160), .Z(n161) );
  XNOR U176 ( .A(b[115]), .B(n162), .Z(c[115]) );
  XNOR U177 ( .A(a[115]), .B(n163), .Z(n162) );
  IV U178 ( .A(n160), .Z(n163) );
  XOR U179 ( .A(n164), .B(n165), .Z(n160) );
  ANDN U180 ( .B(n166), .A(n167), .Z(n164) );
  XNOR U181 ( .A(b[114]), .B(n165), .Z(n166) );
  XNOR U182 ( .A(b[114]), .B(n167), .Z(c[114]) );
  XNOR U183 ( .A(a[114]), .B(n168), .Z(n167) );
  IV U184 ( .A(n165), .Z(n168) );
  XOR U185 ( .A(n169), .B(n170), .Z(n165) );
  ANDN U186 ( .B(n171), .A(n172), .Z(n169) );
  XNOR U187 ( .A(b[113]), .B(n170), .Z(n171) );
  XNOR U188 ( .A(b[113]), .B(n172), .Z(c[113]) );
  XNOR U189 ( .A(a[113]), .B(n173), .Z(n172) );
  IV U190 ( .A(n170), .Z(n173) );
  XOR U191 ( .A(n174), .B(n175), .Z(n170) );
  ANDN U192 ( .B(n176), .A(n177), .Z(n174) );
  XNOR U193 ( .A(b[112]), .B(n175), .Z(n176) );
  XNOR U194 ( .A(b[112]), .B(n177), .Z(c[112]) );
  XNOR U195 ( .A(a[112]), .B(n178), .Z(n177) );
  IV U196 ( .A(n175), .Z(n178) );
  XOR U197 ( .A(n179), .B(n180), .Z(n175) );
  ANDN U198 ( .B(n181), .A(n182), .Z(n179) );
  XNOR U199 ( .A(b[111]), .B(n180), .Z(n181) );
  XNOR U200 ( .A(b[111]), .B(n182), .Z(c[111]) );
  XNOR U201 ( .A(a[111]), .B(n183), .Z(n182) );
  IV U202 ( .A(n180), .Z(n183) );
  XOR U203 ( .A(n184), .B(n185), .Z(n180) );
  ANDN U204 ( .B(n186), .A(n187), .Z(n184) );
  XNOR U205 ( .A(b[110]), .B(n185), .Z(n186) );
  XNOR U206 ( .A(b[110]), .B(n187), .Z(c[110]) );
  XNOR U207 ( .A(a[110]), .B(n188), .Z(n187) );
  IV U208 ( .A(n185), .Z(n188) );
  XOR U209 ( .A(n189), .B(n190), .Z(n185) );
  ANDN U210 ( .B(n191), .A(n192), .Z(n189) );
  XNOR U211 ( .A(b[109]), .B(n190), .Z(n191) );
  XNOR U212 ( .A(b[10]), .B(n193), .Z(c[10]) );
  XNOR U213 ( .A(b[109]), .B(n192), .Z(c[109]) );
  XNOR U214 ( .A(a[109]), .B(n194), .Z(n192) );
  IV U215 ( .A(n190), .Z(n194) );
  XOR U216 ( .A(n195), .B(n196), .Z(n190) );
  ANDN U217 ( .B(n197), .A(n198), .Z(n195) );
  XNOR U218 ( .A(b[108]), .B(n196), .Z(n197) );
  XNOR U219 ( .A(b[108]), .B(n198), .Z(c[108]) );
  XNOR U220 ( .A(a[108]), .B(n199), .Z(n198) );
  IV U221 ( .A(n196), .Z(n199) );
  XOR U222 ( .A(n200), .B(n201), .Z(n196) );
  ANDN U223 ( .B(n202), .A(n203), .Z(n200) );
  XNOR U224 ( .A(b[107]), .B(n201), .Z(n202) );
  XNOR U225 ( .A(b[107]), .B(n203), .Z(c[107]) );
  XNOR U226 ( .A(a[107]), .B(n204), .Z(n203) );
  IV U227 ( .A(n201), .Z(n204) );
  XOR U228 ( .A(n205), .B(n206), .Z(n201) );
  ANDN U229 ( .B(n207), .A(n208), .Z(n205) );
  XNOR U230 ( .A(b[106]), .B(n206), .Z(n207) );
  XNOR U231 ( .A(b[106]), .B(n208), .Z(c[106]) );
  XNOR U232 ( .A(a[106]), .B(n209), .Z(n208) );
  IV U233 ( .A(n206), .Z(n209) );
  XOR U234 ( .A(n210), .B(n211), .Z(n206) );
  ANDN U235 ( .B(n212), .A(n213), .Z(n210) );
  XNOR U236 ( .A(b[105]), .B(n211), .Z(n212) );
  XNOR U237 ( .A(b[105]), .B(n213), .Z(c[105]) );
  XNOR U238 ( .A(a[105]), .B(n214), .Z(n213) );
  IV U239 ( .A(n211), .Z(n214) );
  XOR U240 ( .A(n215), .B(n216), .Z(n211) );
  ANDN U241 ( .B(n217), .A(n218), .Z(n215) );
  XNOR U242 ( .A(b[104]), .B(n216), .Z(n217) );
  XNOR U243 ( .A(b[104]), .B(n218), .Z(c[104]) );
  XNOR U244 ( .A(a[104]), .B(n219), .Z(n218) );
  IV U245 ( .A(n216), .Z(n219) );
  XOR U246 ( .A(n220), .B(n221), .Z(n216) );
  ANDN U247 ( .B(n222), .A(n223), .Z(n220) );
  XNOR U248 ( .A(b[103]), .B(n221), .Z(n222) );
  XNOR U249 ( .A(b[103]), .B(n223), .Z(c[103]) );
  XNOR U250 ( .A(a[103]), .B(n224), .Z(n223) );
  IV U251 ( .A(n221), .Z(n224) );
  XOR U252 ( .A(n225), .B(n226), .Z(n221) );
  ANDN U253 ( .B(n227), .A(n228), .Z(n225) );
  XNOR U254 ( .A(b[102]), .B(n226), .Z(n227) );
  XNOR U255 ( .A(b[102]), .B(n228), .Z(c[102]) );
  XNOR U256 ( .A(a[102]), .B(n229), .Z(n228) );
  IV U257 ( .A(n226), .Z(n229) );
  XOR U258 ( .A(n230), .B(n231), .Z(n226) );
  ANDN U259 ( .B(n232), .A(n233), .Z(n230) );
  XNOR U260 ( .A(b[101]), .B(n231), .Z(n232) );
  XNOR U261 ( .A(b[101]), .B(n233), .Z(c[101]) );
  XNOR U262 ( .A(a[101]), .B(n234), .Z(n233) );
  IV U263 ( .A(n231), .Z(n234) );
  XOR U264 ( .A(n235), .B(n236), .Z(n231) );
  ANDN U265 ( .B(n237), .A(n238), .Z(n235) );
  XNOR U266 ( .A(b[100]), .B(n236), .Z(n237) );
  XNOR U267 ( .A(b[100]), .B(n238), .Z(c[100]) );
  XNOR U268 ( .A(a[100]), .B(n239), .Z(n238) );
  IV U269 ( .A(n236), .Z(n239) );
  XOR U270 ( .A(n240), .B(n241), .Z(n236) );
  ANDN U271 ( .B(n242), .A(n7), .Z(n240) );
  XNOR U272 ( .A(a[99]), .B(n243), .Z(n7) );
  IV U273 ( .A(n241), .Z(n243) );
  XNOR U274 ( .A(b[99]), .B(n241), .Z(n242) );
  XOR U275 ( .A(n244), .B(n245), .Z(n241) );
  ANDN U276 ( .B(n246), .A(n8), .Z(n244) );
  XNOR U277 ( .A(a[98]), .B(n247), .Z(n8) );
  IV U278 ( .A(n245), .Z(n247) );
  XNOR U279 ( .A(b[98]), .B(n245), .Z(n246) );
  XOR U280 ( .A(n248), .B(n249), .Z(n245) );
  ANDN U281 ( .B(n250), .A(n9), .Z(n248) );
  XNOR U282 ( .A(a[97]), .B(n251), .Z(n9) );
  IV U283 ( .A(n249), .Z(n251) );
  XNOR U284 ( .A(b[97]), .B(n249), .Z(n250) );
  XOR U285 ( .A(n252), .B(n253), .Z(n249) );
  ANDN U286 ( .B(n254), .A(n10), .Z(n252) );
  XNOR U287 ( .A(a[96]), .B(n255), .Z(n10) );
  IV U288 ( .A(n253), .Z(n255) );
  XNOR U289 ( .A(b[96]), .B(n253), .Z(n254) );
  XOR U290 ( .A(n256), .B(n257), .Z(n253) );
  ANDN U291 ( .B(n258), .A(n11), .Z(n256) );
  XNOR U292 ( .A(a[95]), .B(n259), .Z(n11) );
  IV U293 ( .A(n257), .Z(n259) );
  XNOR U294 ( .A(b[95]), .B(n257), .Z(n258) );
  XOR U295 ( .A(n260), .B(n261), .Z(n257) );
  ANDN U296 ( .B(n262), .A(n12), .Z(n260) );
  XNOR U297 ( .A(a[94]), .B(n263), .Z(n12) );
  IV U298 ( .A(n261), .Z(n263) );
  XNOR U299 ( .A(b[94]), .B(n261), .Z(n262) );
  XOR U300 ( .A(n264), .B(n265), .Z(n261) );
  ANDN U301 ( .B(n266), .A(n13), .Z(n264) );
  XNOR U302 ( .A(a[93]), .B(n267), .Z(n13) );
  IV U303 ( .A(n265), .Z(n267) );
  XNOR U304 ( .A(b[93]), .B(n265), .Z(n266) );
  XOR U305 ( .A(n268), .B(n269), .Z(n265) );
  ANDN U306 ( .B(n270), .A(n14), .Z(n268) );
  XNOR U307 ( .A(a[92]), .B(n271), .Z(n14) );
  IV U308 ( .A(n269), .Z(n271) );
  XNOR U309 ( .A(b[92]), .B(n269), .Z(n270) );
  XOR U310 ( .A(n272), .B(n273), .Z(n269) );
  ANDN U311 ( .B(n274), .A(n15), .Z(n272) );
  XNOR U312 ( .A(a[91]), .B(n275), .Z(n15) );
  IV U313 ( .A(n273), .Z(n275) );
  XNOR U314 ( .A(b[91]), .B(n273), .Z(n274) );
  XOR U315 ( .A(n276), .B(n277), .Z(n273) );
  ANDN U316 ( .B(n278), .A(n16), .Z(n276) );
  XNOR U317 ( .A(a[90]), .B(n279), .Z(n16) );
  IV U318 ( .A(n277), .Z(n279) );
  XNOR U319 ( .A(b[90]), .B(n277), .Z(n278) );
  XOR U320 ( .A(n280), .B(n281), .Z(n277) );
  ANDN U321 ( .B(n282), .A(n18), .Z(n280) );
  XNOR U322 ( .A(a[89]), .B(n283), .Z(n18) );
  IV U323 ( .A(n281), .Z(n283) );
  XNOR U324 ( .A(b[89]), .B(n281), .Z(n282) );
  XOR U325 ( .A(n284), .B(n285), .Z(n281) );
  ANDN U326 ( .B(n286), .A(n19), .Z(n284) );
  XNOR U327 ( .A(a[88]), .B(n287), .Z(n19) );
  IV U328 ( .A(n285), .Z(n287) );
  XNOR U329 ( .A(b[88]), .B(n285), .Z(n286) );
  XOR U330 ( .A(n288), .B(n289), .Z(n285) );
  ANDN U331 ( .B(n290), .A(n20), .Z(n288) );
  XNOR U332 ( .A(a[87]), .B(n291), .Z(n20) );
  IV U333 ( .A(n289), .Z(n291) );
  XNOR U334 ( .A(b[87]), .B(n289), .Z(n290) );
  XOR U335 ( .A(n292), .B(n293), .Z(n289) );
  ANDN U336 ( .B(n294), .A(n21), .Z(n292) );
  XNOR U337 ( .A(a[86]), .B(n295), .Z(n21) );
  IV U338 ( .A(n293), .Z(n295) );
  XNOR U339 ( .A(b[86]), .B(n293), .Z(n294) );
  XOR U340 ( .A(n296), .B(n297), .Z(n293) );
  ANDN U341 ( .B(n298), .A(n22), .Z(n296) );
  XNOR U342 ( .A(a[85]), .B(n299), .Z(n22) );
  IV U343 ( .A(n297), .Z(n299) );
  XNOR U344 ( .A(b[85]), .B(n297), .Z(n298) );
  XOR U345 ( .A(n300), .B(n301), .Z(n297) );
  ANDN U346 ( .B(n302), .A(n23), .Z(n300) );
  XNOR U347 ( .A(a[84]), .B(n303), .Z(n23) );
  IV U348 ( .A(n301), .Z(n303) );
  XNOR U349 ( .A(b[84]), .B(n301), .Z(n302) );
  XOR U350 ( .A(n304), .B(n305), .Z(n301) );
  ANDN U351 ( .B(n306), .A(n24), .Z(n304) );
  XNOR U352 ( .A(a[83]), .B(n307), .Z(n24) );
  IV U353 ( .A(n305), .Z(n307) );
  XNOR U354 ( .A(b[83]), .B(n305), .Z(n306) );
  XOR U355 ( .A(n308), .B(n309), .Z(n305) );
  ANDN U356 ( .B(n310), .A(n25), .Z(n308) );
  XNOR U357 ( .A(a[82]), .B(n311), .Z(n25) );
  IV U358 ( .A(n309), .Z(n311) );
  XNOR U359 ( .A(b[82]), .B(n309), .Z(n310) );
  XOR U360 ( .A(n312), .B(n313), .Z(n309) );
  ANDN U361 ( .B(n314), .A(n26), .Z(n312) );
  XNOR U362 ( .A(a[81]), .B(n315), .Z(n26) );
  IV U363 ( .A(n313), .Z(n315) );
  XNOR U364 ( .A(b[81]), .B(n313), .Z(n314) );
  XOR U365 ( .A(n316), .B(n317), .Z(n313) );
  ANDN U366 ( .B(n318), .A(n27), .Z(n316) );
  XNOR U367 ( .A(a[80]), .B(n319), .Z(n27) );
  IV U368 ( .A(n317), .Z(n319) );
  XNOR U369 ( .A(b[80]), .B(n317), .Z(n318) );
  XOR U370 ( .A(n320), .B(n321), .Z(n317) );
  ANDN U371 ( .B(n322), .A(n29), .Z(n320) );
  XNOR U372 ( .A(a[79]), .B(n323), .Z(n29) );
  IV U373 ( .A(n321), .Z(n323) );
  XNOR U374 ( .A(b[79]), .B(n321), .Z(n322) );
  XOR U375 ( .A(n324), .B(n325), .Z(n321) );
  ANDN U376 ( .B(n326), .A(n30), .Z(n324) );
  XNOR U377 ( .A(a[78]), .B(n327), .Z(n30) );
  IV U378 ( .A(n325), .Z(n327) );
  XNOR U379 ( .A(b[78]), .B(n325), .Z(n326) );
  XOR U380 ( .A(n328), .B(n329), .Z(n325) );
  ANDN U381 ( .B(n330), .A(n31), .Z(n328) );
  XNOR U382 ( .A(a[77]), .B(n331), .Z(n31) );
  IV U383 ( .A(n329), .Z(n331) );
  XNOR U384 ( .A(b[77]), .B(n329), .Z(n330) );
  XOR U385 ( .A(n332), .B(n333), .Z(n329) );
  ANDN U386 ( .B(n334), .A(n32), .Z(n332) );
  XNOR U387 ( .A(a[76]), .B(n335), .Z(n32) );
  IV U388 ( .A(n333), .Z(n335) );
  XNOR U389 ( .A(b[76]), .B(n333), .Z(n334) );
  XOR U390 ( .A(n336), .B(n337), .Z(n333) );
  ANDN U391 ( .B(n338), .A(n33), .Z(n336) );
  XNOR U392 ( .A(a[75]), .B(n339), .Z(n33) );
  IV U393 ( .A(n337), .Z(n339) );
  XNOR U394 ( .A(b[75]), .B(n337), .Z(n338) );
  XOR U395 ( .A(n340), .B(n341), .Z(n337) );
  ANDN U396 ( .B(n342), .A(n34), .Z(n340) );
  XNOR U397 ( .A(a[74]), .B(n343), .Z(n34) );
  IV U398 ( .A(n341), .Z(n343) );
  XNOR U399 ( .A(b[74]), .B(n341), .Z(n342) );
  XOR U400 ( .A(n344), .B(n345), .Z(n341) );
  ANDN U401 ( .B(n346), .A(n35), .Z(n344) );
  XNOR U402 ( .A(a[73]), .B(n347), .Z(n35) );
  IV U403 ( .A(n345), .Z(n347) );
  XNOR U404 ( .A(b[73]), .B(n345), .Z(n346) );
  XOR U405 ( .A(n348), .B(n349), .Z(n345) );
  ANDN U406 ( .B(n350), .A(n36), .Z(n348) );
  XNOR U407 ( .A(a[72]), .B(n351), .Z(n36) );
  IV U408 ( .A(n349), .Z(n351) );
  XNOR U409 ( .A(b[72]), .B(n349), .Z(n350) );
  XOR U410 ( .A(n352), .B(n353), .Z(n349) );
  ANDN U411 ( .B(n354), .A(n37), .Z(n352) );
  XNOR U412 ( .A(a[71]), .B(n355), .Z(n37) );
  IV U413 ( .A(n353), .Z(n355) );
  XNOR U414 ( .A(b[71]), .B(n353), .Z(n354) );
  XOR U415 ( .A(n356), .B(n357), .Z(n353) );
  ANDN U416 ( .B(n358), .A(n38), .Z(n356) );
  XNOR U417 ( .A(a[70]), .B(n359), .Z(n38) );
  IV U418 ( .A(n357), .Z(n359) );
  XNOR U419 ( .A(b[70]), .B(n357), .Z(n358) );
  XOR U420 ( .A(n360), .B(n361), .Z(n357) );
  ANDN U421 ( .B(n362), .A(n40), .Z(n360) );
  XNOR U422 ( .A(a[69]), .B(n363), .Z(n40) );
  IV U423 ( .A(n361), .Z(n363) );
  XNOR U424 ( .A(b[69]), .B(n361), .Z(n362) );
  XOR U425 ( .A(n364), .B(n365), .Z(n361) );
  ANDN U426 ( .B(n366), .A(n41), .Z(n364) );
  XNOR U427 ( .A(a[68]), .B(n367), .Z(n41) );
  IV U428 ( .A(n365), .Z(n367) );
  XNOR U429 ( .A(b[68]), .B(n365), .Z(n366) );
  XOR U430 ( .A(n368), .B(n369), .Z(n365) );
  ANDN U431 ( .B(n370), .A(n42), .Z(n368) );
  XNOR U432 ( .A(a[67]), .B(n371), .Z(n42) );
  IV U433 ( .A(n369), .Z(n371) );
  XNOR U434 ( .A(b[67]), .B(n369), .Z(n370) );
  XOR U435 ( .A(n372), .B(n373), .Z(n369) );
  ANDN U436 ( .B(n374), .A(n43), .Z(n372) );
  XNOR U437 ( .A(a[66]), .B(n375), .Z(n43) );
  IV U438 ( .A(n373), .Z(n375) );
  XNOR U439 ( .A(b[66]), .B(n373), .Z(n374) );
  XOR U440 ( .A(n376), .B(n377), .Z(n373) );
  ANDN U441 ( .B(n378), .A(n44), .Z(n376) );
  XNOR U442 ( .A(a[65]), .B(n379), .Z(n44) );
  IV U443 ( .A(n377), .Z(n379) );
  XNOR U444 ( .A(b[65]), .B(n377), .Z(n378) );
  XOR U445 ( .A(n380), .B(n381), .Z(n377) );
  ANDN U446 ( .B(n382), .A(n45), .Z(n380) );
  XNOR U447 ( .A(a[64]), .B(n383), .Z(n45) );
  IV U448 ( .A(n381), .Z(n383) );
  XNOR U449 ( .A(b[64]), .B(n381), .Z(n382) );
  XOR U450 ( .A(n384), .B(n385), .Z(n381) );
  ANDN U451 ( .B(n386), .A(n46), .Z(n384) );
  XNOR U452 ( .A(a[63]), .B(n387), .Z(n46) );
  IV U453 ( .A(n385), .Z(n387) );
  XNOR U454 ( .A(b[63]), .B(n385), .Z(n386) );
  XOR U455 ( .A(n388), .B(n389), .Z(n385) );
  ANDN U456 ( .B(n390), .A(n47), .Z(n388) );
  XNOR U457 ( .A(a[62]), .B(n391), .Z(n47) );
  IV U458 ( .A(n389), .Z(n391) );
  XNOR U459 ( .A(b[62]), .B(n389), .Z(n390) );
  XOR U460 ( .A(n392), .B(n393), .Z(n389) );
  ANDN U461 ( .B(n394), .A(n48), .Z(n392) );
  XNOR U462 ( .A(a[61]), .B(n395), .Z(n48) );
  IV U463 ( .A(n393), .Z(n395) );
  XNOR U464 ( .A(b[61]), .B(n393), .Z(n394) );
  XOR U465 ( .A(n396), .B(n397), .Z(n393) );
  ANDN U466 ( .B(n398), .A(n49), .Z(n396) );
  XNOR U467 ( .A(a[60]), .B(n399), .Z(n49) );
  IV U468 ( .A(n397), .Z(n399) );
  XNOR U469 ( .A(b[60]), .B(n397), .Z(n398) );
  XOR U470 ( .A(n400), .B(n401), .Z(n397) );
  ANDN U471 ( .B(n402), .A(n51), .Z(n400) );
  XNOR U472 ( .A(a[59]), .B(n403), .Z(n51) );
  IV U473 ( .A(n401), .Z(n403) );
  XNOR U474 ( .A(b[59]), .B(n401), .Z(n402) );
  XOR U475 ( .A(n404), .B(n405), .Z(n401) );
  ANDN U476 ( .B(n406), .A(n52), .Z(n404) );
  XNOR U477 ( .A(a[58]), .B(n407), .Z(n52) );
  IV U478 ( .A(n405), .Z(n407) );
  XNOR U479 ( .A(b[58]), .B(n405), .Z(n406) );
  XOR U480 ( .A(n408), .B(n409), .Z(n405) );
  ANDN U481 ( .B(n410), .A(n53), .Z(n408) );
  XNOR U482 ( .A(a[57]), .B(n411), .Z(n53) );
  IV U483 ( .A(n409), .Z(n411) );
  XNOR U484 ( .A(b[57]), .B(n409), .Z(n410) );
  XOR U485 ( .A(n412), .B(n413), .Z(n409) );
  ANDN U486 ( .B(n414), .A(n54), .Z(n412) );
  XNOR U487 ( .A(a[56]), .B(n415), .Z(n54) );
  IV U488 ( .A(n413), .Z(n415) );
  XNOR U489 ( .A(b[56]), .B(n413), .Z(n414) );
  XOR U490 ( .A(n416), .B(n417), .Z(n413) );
  ANDN U491 ( .B(n418), .A(n55), .Z(n416) );
  XNOR U492 ( .A(a[55]), .B(n419), .Z(n55) );
  IV U493 ( .A(n417), .Z(n419) );
  XNOR U494 ( .A(b[55]), .B(n417), .Z(n418) );
  XOR U495 ( .A(n420), .B(n421), .Z(n417) );
  ANDN U496 ( .B(n422), .A(n56), .Z(n420) );
  XNOR U497 ( .A(a[54]), .B(n423), .Z(n56) );
  IV U498 ( .A(n421), .Z(n423) );
  XNOR U499 ( .A(b[54]), .B(n421), .Z(n422) );
  XOR U500 ( .A(n424), .B(n425), .Z(n421) );
  ANDN U501 ( .B(n426), .A(n57), .Z(n424) );
  XNOR U502 ( .A(a[53]), .B(n427), .Z(n57) );
  IV U503 ( .A(n425), .Z(n427) );
  XNOR U504 ( .A(b[53]), .B(n425), .Z(n426) );
  XOR U505 ( .A(n428), .B(n429), .Z(n425) );
  ANDN U506 ( .B(n430), .A(n58), .Z(n428) );
  XNOR U507 ( .A(a[52]), .B(n431), .Z(n58) );
  IV U508 ( .A(n429), .Z(n431) );
  XNOR U509 ( .A(b[52]), .B(n429), .Z(n430) );
  XOR U510 ( .A(n432), .B(n433), .Z(n429) );
  ANDN U511 ( .B(n434), .A(n59), .Z(n432) );
  XNOR U512 ( .A(a[51]), .B(n435), .Z(n59) );
  IV U513 ( .A(n433), .Z(n435) );
  XNOR U514 ( .A(b[51]), .B(n433), .Z(n434) );
  XOR U515 ( .A(n436), .B(n437), .Z(n433) );
  ANDN U516 ( .B(n438), .A(n60), .Z(n436) );
  XNOR U517 ( .A(a[50]), .B(n439), .Z(n60) );
  IV U518 ( .A(n437), .Z(n439) );
  XNOR U519 ( .A(b[50]), .B(n437), .Z(n438) );
  XOR U520 ( .A(n440), .B(n441), .Z(n437) );
  ANDN U521 ( .B(n442), .A(n62), .Z(n440) );
  XNOR U522 ( .A(a[49]), .B(n443), .Z(n62) );
  IV U523 ( .A(n441), .Z(n443) );
  XNOR U524 ( .A(b[49]), .B(n441), .Z(n442) );
  XOR U525 ( .A(n444), .B(n445), .Z(n441) );
  ANDN U526 ( .B(n446), .A(n63), .Z(n444) );
  XNOR U527 ( .A(a[48]), .B(n447), .Z(n63) );
  IV U528 ( .A(n445), .Z(n447) );
  XNOR U529 ( .A(b[48]), .B(n445), .Z(n446) );
  XOR U530 ( .A(n448), .B(n449), .Z(n445) );
  ANDN U531 ( .B(n450), .A(n64), .Z(n448) );
  XNOR U532 ( .A(a[47]), .B(n451), .Z(n64) );
  IV U533 ( .A(n449), .Z(n451) );
  XNOR U534 ( .A(b[47]), .B(n449), .Z(n450) );
  XOR U535 ( .A(n452), .B(n453), .Z(n449) );
  ANDN U536 ( .B(n454), .A(n65), .Z(n452) );
  XNOR U537 ( .A(a[46]), .B(n455), .Z(n65) );
  IV U538 ( .A(n453), .Z(n455) );
  XNOR U539 ( .A(b[46]), .B(n453), .Z(n454) );
  XOR U540 ( .A(n456), .B(n457), .Z(n453) );
  ANDN U541 ( .B(n458), .A(n66), .Z(n456) );
  XNOR U542 ( .A(a[45]), .B(n459), .Z(n66) );
  IV U543 ( .A(n457), .Z(n459) );
  XNOR U544 ( .A(b[45]), .B(n457), .Z(n458) );
  XOR U545 ( .A(n460), .B(n461), .Z(n457) );
  ANDN U546 ( .B(n462), .A(n67), .Z(n460) );
  XNOR U547 ( .A(a[44]), .B(n463), .Z(n67) );
  IV U548 ( .A(n461), .Z(n463) );
  XNOR U549 ( .A(b[44]), .B(n461), .Z(n462) );
  XOR U550 ( .A(n464), .B(n465), .Z(n461) );
  ANDN U551 ( .B(n466), .A(n68), .Z(n464) );
  XNOR U552 ( .A(a[43]), .B(n467), .Z(n68) );
  IV U553 ( .A(n465), .Z(n467) );
  XNOR U554 ( .A(b[43]), .B(n465), .Z(n466) );
  XOR U555 ( .A(n468), .B(n469), .Z(n465) );
  ANDN U556 ( .B(n470), .A(n69), .Z(n468) );
  XNOR U557 ( .A(a[42]), .B(n471), .Z(n69) );
  IV U558 ( .A(n469), .Z(n471) );
  XNOR U559 ( .A(b[42]), .B(n469), .Z(n470) );
  XOR U560 ( .A(n472), .B(n473), .Z(n469) );
  ANDN U561 ( .B(n474), .A(n70), .Z(n472) );
  XNOR U562 ( .A(a[41]), .B(n475), .Z(n70) );
  IV U563 ( .A(n473), .Z(n475) );
  XNOR U564 ( .A(b[41]), .B(n473), .Z(n474) );
  XOR U565 ( .A(n476), .B(n477), .Z(n473) );
  ANDN U566 ( .B(n478), .A(n71), .Z(n476) );
  XNOR U567 ( .A(a[40]), .B(n479), .Z(n71) );
  IV U568 ( .A(n477), .Z(n479) );
  XNOR U569 ( .A(b[40]), .B(n477), .Z(n478) );
  XOR U570 ( .A(n480), .B(n481), .Z(n477) );
  ANDN U571 ( .B(n482), .A(n73), .Z(n480) );
  XNOR U572 ( .A(a[39]), .B(n483), .Z(n73) );
  IV U573 ( .A(n481), .Z(n483) );
  XNOR U574 ( .A(b[39]), .B(n481), .Z(n482) );
  XOR U575 ( .A(n484), .B(n485), .Z(n481) );
  ANDN U576 ( .B(n486), .A(n74), .Z(n484) );
  XNOR U577 ( .A(a[38]), .B(n487), .Z(n74) );
  IV U578 ( .A(n485), .Z(n487) );
  XNOR U579 ( .A(b[38]), .B(n485), .Z(n486) );
  XOR U580 ( .A(n488), .B(n489), .Z(n485) );
  ANDN U581 ( .B(n490), .A(n75), .Z(n488) );
  XNOR U582 ( .A(a[37]), .B(n491), .Z(n75) );
  IV U583 ( .A(n489), .Z(n491) );
  XNOR U584 ( .A(b[37]), .B(n489), .Z(n490) );
  XOR U585 ( .A(n492), .B(n493), .Z(n489) );
  ANDN U586 ( .B(n494), .A(n76), .Z(n492) );
  XNOR U587 ( .A(a[36]), .B(n495), .Z(n76) );
  IV U588 ( .A(n493), .Z(n495) );
  XNOR U589 ( .A(b[36]), .B(n493), .Z(n494) );
  XOR U590 ( .A(n496), .B(n497), .Z(n493) );
  ANDN U591 ( .B(n498), .A(n77), .Z(n496) );
  XNOR U592 ( .A(a[35]), .B(n499), .Z(n77) );
  IV U593 ( .A(n497), .Z(n499) );
  XNOR U594 ( .A(b[35]), .B(n497), .Z(n498) );
  XOR U595 ( .A(n500), .B(n501), .Z(n497) );
  ANDN U596 ( .B(n502), .A(n78), .Z(n500) );
  XNOR U597 ( .A(a[34]), .B(n503), .Z(n78) );
  IV U598 ( .A(n501), .Z(n503) );
  XNOR U599 ( .A(b[34]), .B(n501), .Z(n502) );
  XOR U600 ( .A(n504), .B(n505), .Z(n501) );
  ANDN U601 ( .B(n506), .A(n79), .Z(n504) );
  XNOR U602 ( .A(a[33]), .B(n507), .Z(n79) );
  IV U603 ( .A(n505), .Z(n507) );
  XNOR U604 ( .A(b[33]), .B(n505), .Z(n506) );
  XOR U605 ( .A(n508), .B(n509), .Z(n505) );
  ANDN U606 ( .B(n510), .A(n80), .Z(n508) );
  XNOR U607 ( .A(a[32]), .B(n511), .Z(n80) );
  IV U608 ( .A(n509), .Z(n511) );
  XNOR U609 ( .A(b[32]), .B(n509), .Z(n510) );
  XOR U610 ( .A(n512), .B(n513), .Z(n509) );
  ANDN U611 ( .B(n514), .A(n81), .Z(n512) );
  XNOR U612 ( .A(a[31]), .B(n515), .Z(n81) );
  IV U613 ( .A(n513), .Z(n515) );
  XNOR U614 ( .A(b[31]), .B(n513), .Z(n514) );
  XOR U615 ( .A(n516), .B(n517), .Z(n513) );
  ANDN U616 ( .B(n518), .A(n82), .Z(n516) );
  XNOR U617 ( .A(a[30]), .B(n519), .Z(n82) );
  IV U618 ( .A(n517), .Z(n519) );
  XNOR U619 ( .A(b[30]), .B(n517), .Z(n518) );
  XOR U620 ( .A(n520), .B(n521), .Z(n517) );
  ANDN U621 ( .B(n522), .A(n84), .Z(n520) );
  XNOR U622 ( .A(a[29]), .B(n523), .Z(n84) );
  IV U623 ( .A(n521), .Z(n523) );
  XNOR U624 ( .A(b[29]), .B(n521), .Z(n522) );
  XOR U625 ( .A(n524), .B(n525), .Z(n521) );
  ANDN U626 ( .B(n526), .A(n85), .Z(n524) );
  XNOR U627 ( .A(a[28]), .B(n527), .Z(n85) );
  IV U628 ( .A(n525), .Z(n527) );
  XNOR U629 ( .A(b[28]), .B(n525), .Z(n526) );
  XOR U630 ( .A(n528), .B(n529), .Z(n525) );
  ANDN U631 ( .B(n530), .A(n86), .Z(n528) );
  XNOR U632 ( .A(a[27]), .B(n531), .Z(n86) );
  IV U633 ( .A(n529), .Z(n531) );
  XNOR U634 ( .A(b[27]), .B(n529), .Z(n530) );
  XOR U635 ( .A(n532), .B(n533), .Z(n529) );
  ANDN U636 ( .B(n534), .A(n87), .Z(n532) );
  XNOR U637 ( .A(a[26]), .B(n535), .Z(n87) );
  IV U638 ( .A(n533), .Z(n535) );
  XNOR U639 ( .A(b[26]), .B(n533), .Z(n534) );
  XOR U640 ( .A(n536), .B(n537), .Z(n533) );
  ANDN U641 ( .B(n538), .A(n88), .Z(n536) );
  XNOR U642 ( .A(a[25]), .B(n539), .Z(n88) );
  IV U643 ( .A(n537), .Z(n539) );
  XNOR U644 ( .A(b[25]), .B(n537), .Z(n538) );
  XOR U645 ( .A(n540), .B(n541), .Z(n537) );
  ANDN U646 ( .B(n542), .A(n89), .Z(n540) );
  XNOR U647 ( .A(a[24]), .B(n543), .Z(n89) );
  IV U648 ( .A(n541), .Z(n543) );
  XNOR U649 ( .A(b[24]), .B(n541), .Z(n542) );
  XOR U650 ( .A(n544), .B(n545), .Z(n541) );
  ANDN U651 ( .B(n546), .A(n90), .Z(n544) );
  XNOR U652 ( .A(a[23]), .B(n547), .Z(n90) );
  IV U653 ( .A(n545), .Z(n547) );
  XNOR U654 ( .A(b[23]), .B(n545), .Z(n546) );
  XOR U655 ( .A(n548), .B(n549), .Z(n545) );
  ANDN U656 ( .B(n550), .A(n91), .Z(n548) );
  XNOR U657 ( .A(a[22]), .B(n551), .Z(n91) );
  IV U658 ( .A(n549), .Z(n551) );
  XNOR U659 ( .A(b[22]), .B(n549), .Z(n550) );
  XOR U660 ( .A(n552), .B(n553), .Z(n549) );
  ANDN U661 ( .B(n554), .A(n92), .Z(n552) );
  XNOR U662 ( .A(a[21]), .B(n555), .Z(n92) );
  IV U663 ( .A(n553), .Z(n555) );
  XNOR U664 ( .A(b[21]), .B(n553), .Z(n554) );
  XOR U665 ( .A(n556), .B(n557), .Z(n553) );
  ANDN U666 ( .B(n558), .A(n93), .Z(n556) );
  XNOR U667 ( .A(a[20]), .B(n559), .Z(n93) );
  IV U668 ( .A(n557), .Z(n559) );
  XNOR U669 ( .A(b[20]), .B(n557), .Z(n558) );
  XOR U670 ( .A(n560), .B(n561), .Z(n557) );
  ANDN U671 ( .B(n562), .A(n95), .Z(n560) );
  XNOR U672 ( .A(a[19]), .B(n563), .Z(n95) );
  IV U673 ( .A(n561), .Z(n563) );
  XNOR U674 ( .A(b[19]), .B(n561), .Z(n562) );
  XOR U675 ( .A(n564), .B(n565), .Z(n561) );
  ANDN U676 ( .B(n566), .A(n96), .Z(n564) );
  XNOR U677 ( .A(a[18]), .B(n567), .Z(n96) );
  IV U678 ( .A(n565), .Z(n567) );
  XNOR U679 ( .A(b[18]), .B(n565), .Z(n566) );
  XOR U680 ( .A(n568), .B(n569), .Z(n565) );
  ANDN U681 ( .B(n570), .A(n97), .Z(n568) );
  XNOR U682 ( .A(a[17]), .B(n571), .Z(n97) );
  IV U683 ( .A(n569), .Z(n571) );
  XNOR U684 ( .A(b[17]), .B(n569), .Z(n570) );
  XOR U685 ( .A(n572), .B(n573), .Z(n569) );
  ANDN U686 ( .B(n574), .A(n98), .Z(n572) );
  XNOR U687 ( .A(a[16]), .B(n575), .Z(n98) );
  IV U688 ( .A(n573), .Z(n575) );
  XNOR U689 ( .A(b[16]), .B(n573), .Z(n574) );
  XOR U690 ( .A(n576), .B(n577), .Z(n573) );
  ANDN U691 ( .B(n578), .A(n99), .Z(n576) );
  XNOR U692 ( .A(a[15]), .B(n579), .Z(n99) );
  IV U693 ( .A(n577), .Z(n579) );
  XNOR U694 ( .A(b[15]), .B(n577), .Z(n578) );
  XOR U695 ( .A(n580), .B(n581), .Z(n577) );
  ANDN U696 ( .B(n582), .A(n100), .Z(n580) );
  XNOR U697 ( .A(a[14]), .B(n583), .Z(n100) );
  IV U698 ( .A(n581), .Z(n583) );
  XNOR U699 ( .A(b[14]), .B(n581), .Z(n582) );
  XOR U700 ( .A(n584), .B(n585), .Z(n581) );
  ANDN U701 ( .B(n586), .A(n101), .Z(n584) );
  XNOR U702 ( .A(a[13]), .B(n587), .Z(n101) );
  IV U703 ( .A(n585), .Z(n587) );
  XNOR U704 ( .A(b[13]), .B(n585), .Z(n586) );
  XOR U705 ( .A(n588), .B(n589), .Z(n585) );
  ANDN U706 ( .B(n590), .A(n102), .Z(n588) );
  XNOR U707 ( .A(a[12]), .B(n591), .Z(n102) );
  IV U708 ( .A(n589), .Z(n591) );
  XNOR U709 ( .A(b[12]), .B(n589), .Z(n590) );
  XOR U710 ( .A(n592), .B(n593), .Z(n589) );
  ANDN U711 ( .B(n594), .A(n142), .Z(n592) );
  XNOR U712 ( .A(a[11]), .B(n595), .Z(n142) );
  IV U713 ( .A(n593), .Z(n595) );
  XNOR U714 ( .A(b[11]), .B(n593), .Z(n594) );
  XOR U715 ( .A(n596), .B(n597), .Z(n593) );
  ANDN U716 ( .B(n598), .A(n193), .Z(n596) );
  XNOR U717 ( .A(a[10]), .B(n599), .Z(n193) );
  IV U718 ( .A(n597), .Z(n599) );
  XNOR U719 ( .A(b[10]), .B(n597), .Z(n598) );
  XOR U720 ( .A(n600), .B(n601), .Z(n597) );
  ANDN U721 ( .B(n602), .A(n6), .Z(n600) );
  XNOR U722 ( .A(a[9]), .B(n603), .Z(n6) );
  IV U723 ( .A(n601), .Z(n603) );
  XNOR U724 ( .A(b[9]), .B(n601), .Z(n602) );
  XOR U725 ( .A(n604), .B(n605), .Z(n601) );
  ANDN U726 ( .B(n606), .A(n17), .Z(n604) );
  XNOR U727 ( .A(a[8]), .B(n607), .Z(n17) );
  IV U728 ( .A(n605), .Z(n607) );
  XNOR U729 ( .A(b[8]), .B(n605), .Z(n606) );
  XOR U730 ( .A(n608), .B(n609), .Z(n605) );
  ANDN U731 ( .B(n610), .A(n28), .Z(n608) );
  XNOR U732 ( .A(a[7]), .B(n611), .Z(n28) );
  IV U733 ( .A(n609), .Z(n611) );
  XNOR U734 ( .A(b[7]), .B(n609), .Z(n610) );
  XOR U735 ( .A(n612), .B(n613), .Z(n609) );
  ANDN U736 ( .B(n614), .A(n39), .Z(n612) );
  XNOR U737 ( .A(a[6]), .B(n615), .Z(n39) );
  IV U738 ( .A(n613), .Z(n615) );
  XNOR U739 ( .A(b[6]), .B(n613), .Z(n614) );
  XOR U740 ( .A(n616), .B(n617), .Z(n613) );
  ANDN U741 ( .B(n618), .A(n50), .Z(n616) );
  XNOR U742 ( .A(a[5]), .B(n619), .Z(n50) );
  IV U743 ( .A(n617), .Z(n619) );
  XNOR U744 ( .A(b[5]), .B(n617), .Z(n618) );
  XOR U745 ( .A(n620), .B(n621), .Z(n617) );
  ANDN U746 ( .B(n622), .A(n61), .Z(n620) );
  XNOR U747 ( .A(a[4]), .B(n623), .Z(n61) );
  IV U748 ( .A(n621), .Z(n623) );
  XNOR U749 ( .A(b[4]), .B(n621), .Z(n622) );
  XOR U750 ( .A(n624), .B(n625), .Z(n621) );
  ANDN U751 ( .B(n626), .A(n72), .Z(n624) );
  XNOR U752 ( .A(a[3]), .B(n627), .Z(n72) );
  IV U753 ( .A(n625), .Z(n627) );
  XNOR U754 ( .A(b[3]), .B(n625), .Z(n626) );
  XOR U755 ( .A(n628), .B(n629), .Z(n625) );
  ANDN U756 ( .B(n630), .A(n83), .Z(n628) );
  XNOR U757 ( .A(a[2]), .B(n631), .Z(n83) );
  IV U758 ( .A(n629), .Z(n631) );
  XNOR U759 ( .A(b[2]), .B(n629), .Z(n630) );
  XOR U760 ( .A(n632), .B(n633), .Z(n629) );
  ANDN U761 ( .B(n634), .A(n94), .Z(n632) );
  XNOR U762 ( .A(a[1]), .B(n635), .Z(n94) );
  IV U763 ( .A(n633), .Z(n635) );
  XNOR U764 ( .A(b[1]), .B(n633), .Z(n634) );
  XOR U765 ( .A(carry_on), .B(n636), .Z(n633) );
  NANDN U766 ( .A(n637), .B(n638), .Z(n636) );
  XOR U767 ( .A(carry_on), .B(b[0]), .Z(n638) );
  XNOR U768 ( .A(b[0]), .B(n637), .Z(c[0]) );
  XNOR U769 ( .A(a[0]), .B(carry_on), .Z(n637) );
endmodule

