
module compare_N16384_CC512 ( clk, rst, x, y, g, e );
  input [31:0] x;
  input [31:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  NANDN U10 ( .A(n143), .B(n142), .Z(n8) );
  AND U11 ( .A(n144), .B(n8), .Z(n9) );
  ANDN U12 ( .B(n145), .A(n9), .Z(n10) );
  NANDN U13 ( .A(y[7]), .B(x[7]), .Z(n11) );
  AND U14 ( .A(n10), .B(n11), .Z(n12) );
  NANDN U15 ( .A(y[9]), .B(x[9]), .Z(n13) );
  NANDN U16 ( .A(n12), .B(n146), .Z(n14) );
  NAND U17 ( .A(n13), .B(n14), .Z(n15) );
  NANDN U18 ( .A(n15), .B(n147), .Z(n16) );
  AND U19 ( .A(n148), .B(n16), .Z(n17) );
  ANDN U20 ( .B(n149), .A(n17), .Z(n18) );
  NANDN U21 ( .A(y[11]), .B(x[11]), .Z(n19) );
  AND U22 ( .A(n18), .B(n19), .Z(n20) );
  NANDN U23 ( .A(n20), .B(n150), .Z(n21) );
  NANDN U24 ( .A(y[13]), .B(x[13]), .Z(n22) );
  AND U25 ( .A(n21), .B(n22), .Z(n23) );
  NAND U26 ( .A(n151), .B(n23), .Z(n24) );
  NAND U27 ( .A(n152), .B(n24), .Z(n153) );
  NOR U28 ( .A(n156), .B(n154), .Z(n25) );
  NAND U29 ( .A(n153), .B(n25), .Z(n26) );
  NAND U30 ( .A(n157), .B(n26), .Z(n27) );
  AND U31 ( .A(n27), .B(n136), .Z(n28) );
  NANDN U32 ( .A(y[17]), .B(x[17]), .Z(n29) );
  AND U33 ( .A(n28), .B(n29), .Z(n30) );
  NANDN U34 ( .A(n30), .B(n158), .Z(n31) );
  AND U35 ( .A(n159), .B(n31), .Z(n32) );
  NANDN U36 ( .A(y[19]), .B(x[19]), .Z(n33) );
  NAND U37 ( .A(n32), .B(n33), .Z(n34) );
  AND U38 ( .A(n160), .B(n34), .Z(n35) );
  ANDN U39 ( .B(n161), .A(n35), .Z(n36) );
  NANDN U40 ( .A(y[21]), .B(x[21]), .Z(n37) );
  NAND U41 ( .A(n36), .B(n37), .Z(n38) );
  AND U42 ( .A(n162), .B(n38), .Z(n39) );
  ANDN U43 ( .B(n135), .A(n39), .Z(n40) );
  NANDN U44 ( .A(y[23]), .B(x[23]), .Z(n41) );
  NAND U45 ( .A(n40), .B(n41), .Z(n163) );
  XNOR U46 ( .A(x[1]), .B(n137), .Z(n42) );
  NANDN U47 ( .A(y[1]), .B(n42), .Z(n43) );
  AND U48 ( .A(n43), .B(n138), .Z(n44) );
  NANDN U49 ( .A(n137), .B(x[1]), .Z(n45) );
  AND U50 ( .A(n44), .B(n45), .Z(n46) );
  NANDN U51 ( .A(n46), .B(n139), .Z(n47) );
  NANDN U52 ( .A(y[3]), .B(x[3]), .Z(n48) );
  AND U53 ( .A(n47), .B(n48), .Z(n49) );
  ANDN U54 ( .B(x[5]), .A(y[5]), .Z(n50) );
  NAND U55 ( .A(n140), .B(n49), .Z(n51) );
  NAND U56 ( .A(n141), .B(n51), .Z(n52) );
  NANDN U57 ( .A(n50), .B(n52), .Z(n143) );
  AND U58 ( .A(e), .B(n170), .Z(n53) );
  NAND U59 ( .A(n164), .B(n163), .Z(n54) );
  AND U60 ( .A(n134), .B(n54), .Z(n55) );
  NANDN U61 ( .A(y[25]), .B(x[25]), .Z(n56) );
  NAND U62 ( .A(n55), .B(n56), .Z(n57) );
  NAND U63 ( .A(n165), .B(n57), .Z(n58) );
  AND U64 ( .A(n58), .B(n166), .Z(n59) );
  NANDN U65 ( .A(y[27]), .B(x[27]), .Z(n60) );
  AND U66 ( .A(n59), .B(n60), .Z(n61) );
  NANDN U67 ( .A(n61), .B(n167), .Z(n62) );
  AND U68 ( .A(n168), .B(n62), .Z(n63) );
  NANDN U69 ( .A(y[29]), .B(x[29]), .Z(n64) );
  AND U70 ( .A(n63), .B(n64), .Z(n65) );
  NANDN U71 ( .A(y[31]), .B(x[31]), .Z(n66) );
  NANDN U72 ( .A(n65), .B(n169), .Z(n67) );
  NAND U73 ( .A(n66), .B(n67), .Z(n68) );
  NAND U74 ( .A(n68), .B(n53), .Z(n69) );
  NANDN U75 ( .A(n53), .B(g), .Z(n70) );
  NAND U76 ( .A(n69), .B(n70), .Z(n4) );
  IV U77 ( .A(ebreg), .Z(e) );
  XNOR U78 ( .A(x[23]), .B(y[23]), .Z(n72) );
  NANDN U79 ( .A(x[22]), .B(y[22]), .Z(n71) );
  AND U80 ( .A(n72), .B(n71), .Z(n162) );
  XNOR U81 ( .A(x[17]), .B(y[17]), .Z(n74) );
  NANDN U82 ( .A(x[16]), .B(y[16]), .Z(n73) );
  AND U83 ( .A(n74), .B(n73), .Z(n157) );
  AND U84 ( .A(n162), .B(n157), .Z(n80) );
  XNOR U85 ( .A(x[21]), .B(y[21]), .Z(n76) );
  NANDN U86 ( .A(x[20]), .B(y[20]), .Z(n75) );
  AND U87 ( .A(n76), .B(n75), .Z(n160) );
  XNOR U88 ( .A(x[19]), .B(y[19]), .Z(n78) );
  NANDN U89 ( .A(x[18]), .B(y[18]), .Z(n77) );
  AND U90 ( .A(n78), .B(n77), .Z(n158) );
  AND U91 ( .A(n160), .B(n158), .Z(n79) );
  AND U92 ( .A(n80), .B(n79), .Z(n133) );
  XNOR U93 ( .A(y[11]), .B(x[11]), .Z(n82) );
  NANDN U94 ( .A(x[10]), .B(y[10]), .Z(n81) );
  AND U95 ( .A(n82), .B(n81), .Z(n148) );
  XNOR U96 ( .A(y[5]), .B(x[5]), .Z(n84) );
  NANDN U97 ( .A(x[4]), .B(y[4]), .Z(n83) );
  AND U98 ( .A(n84), .B(n83), .Z(n141) );
  AND U99 ( .A(n148), .B(n141), .Z(n90) );
  XNOR U100 ( .A(y[9]), .B(x[9]), .Z(n86) );
  NANDN U101 ( .A(x[8]), .B(y[8]), .Z(n85) );
  AND U102 ( .A(n86), .B(n85), .Z(n146) );
  XNOR U103 ( .A(y[7]), .B(x[7]), .Z(n88) );
  NANDN U104 ( .A(x[6]), .B(y[6]), .Z(n87) );
  AND U105 ( .A(n88), .B(n87), .Z(n144) );
  AND U106 ( .A(n146), .B(n144), .Z(n89) );
  AND U107 ( .A(n90), .B(n89), .Z(n102) );
  XNOR U108 ( .A(x[31]), .B(y[31]), .Z(n92) );
  NANDN U109 ( .A(x[30]), .B(y[30]), .Z(n91) );
  AND U110 ( .A(n92), .B(n91), .Z(n169) );
  XNOR U111 ( .A(x[25]), .B(y[25]), .Z(n94) );
  NANDN U112 ( .A(x[24]), .B(y[24]), .Z(n93) );
  AND U113 ( .A(n94), .B(n93), .Z(n164) );
  AND U114 ( .A(n169), .B(n164), .Z(n100) );
  XNOR U115 ( .A(x[29]), .B(y[29]), .Z(n96) );
  NANDN U116 ( .A(x[28]), .B(y[28]), .Z(n95) );
  AND U117 ( .A(n96), .B(n95), .Z(n167) );
  XNOR U118 ( .A(x[27]), .B(y[27]), .Z(n98) );
  NANDN U119 ( .A(x[26]), .B(y[26]), .Z(n97) );
  AND U120 ( .A(n98), .B(n97), .Z(n165) );
  AND U121 ( .A(n167), .B(n165), .Z(n99) );
  AND U122 ( .A(n100), .B(n99), .Z(n101) );
  AND U123 ( .A(n102), .B(n101), .Z(n131) );
  XNOR U124 ( .A(y[1]), .B(x[1]), .Z(n104) );
  NANDN U125 ( .A(x[0]), .B(y[0]), .Z(n103) );
  AND U126 ( .A(n104), .B(n103), .Z(n107) );
  XNOR U127 ( .A(y[13]), .B(x[13]), .Z(n106) );
  NANDN U128 ( .A(x[12]), .B(y[12]), .Z(n105) );
  AND U129 ( .A(n106), .B(n105), .Z(n150) );
  AND U130 ( .A(n107), .B(n150), .Z(n113) );
  XNOR U131 ( .A(y[3]), .B(x[3]), .Z(n109) );
  NANDN U132 ( .A(x[2]), .B(y[2]), .Z(n108) );
  AND U133 ( .A(n109), .B(n108), .Z(n139) );
  XNOR U134 ( .A(y[15]), .B(x[15]), .Z(n111) );
  NANDN U135 ( .A(x[14]), .B(y[14]), .Z(n110) );
  AND U136 ( .A(n111), .B(n110), .Z(n152) );
  AND U137 ( .A(n139), .B(n152), .Z(n112) );
  AND U138 ( .A(n113), .B(n112), .Z(n129) );
  NANDN U139 ( .A(y[30]), .B(x[30]), .Z(n168) );
  NANDN U140 ( .A(y[24]), .B(x[24]), .Z(n135) );
  AND U141 ( .A(n168), .B(n135), .Z(n115) );
  NANDN U142 ( .A(y[28]), .B(x[28]), .Z(n166) );
  NANDN U143 ( .A(y[26]), .B(x[26]), .Z(n134) );
  AND U144 ( .A(n166), .B(n134), .Z(n114) );
  AND U145 ( .A(n115), .B(n114), .Z(n119) );
  NANDN U146 ( .A(y[6]), .B(x[6]), .Z(n142) );
  NANDN U147 ( .A(y[4]), .B(x[4]), .Z(n140) );
  AND U148 ( .A(n142), .B(n140), .Z(n117) );
  NANDN U149 ( .A(y[2]), .B(x[2]), .Z(n138) );
  NANDN U150 ( .A(y[0]), .B(x[0]), .Z(n137) );
  AND U151 ( .A(n138), .B(n137), .Z(n116) );
  AND U152 ( .A(n117), .B(n116), .Z(n118) );
  AND U153 ( .A(n119), .B(n118), .Z(n127) );
  NANDN U154 ( .A(y[22]), .B(x[22]), .Z(n161) );
  NANDN U155 ( .A(y[16]), .B(x[16]), .Z(n155) );
  AND U156 ( .A(n161), .B(n155), .Z(n121) );
  NANDN U157 ( .A(y[20]), .B(x[20]), .Z(n159) );
  NANDN U158 ( .A(y[18]), .B(x[18]), .Z(n136) );
  AND U159 ( .A(n159), .B(n136), .Z(n120) );
  AND U160 ( .A(n121), .B(n120), .Z(n125) );
  NANDN U161 ( .A(y[14]), .B(x[14]), .Z(n151) );
  NANDN U162 ( .A(y[8]), .B(x[8]), .Z(n145) );
  AND U163 ( .A(n151), .B(n145), .Z(n123) );
  NANDN U164 ( .A(y[12]), .B(x[12]), .Z(n149) );
  NANDN U165 ( .A(y[10]), .B(x[10]), .Z(n147) );
  AND U166 ( .A(n149), .B(n147), .Z(n122) );
  AND U167 ( .A(n123), .B(n122), .Z(n124) );
  AND U168 ( .A(n125), .B(n124), .Z(n126) );
  AND U169 ( .A(n127), .B(n126), .Z(n128) );
  AND U170 ( .A(n129), .B(n128), .Z(n130) );
  AND U171 ( .A(n131), .B(n130), .Z(n132) );
  NAND U172 ( .A(n133), .B(n132), .Z(n170) );
  NANDN U173 ( .A(n170), .B(e), .Z(n5) );
  ANDN U174 ( .B(x[15]), .A(y[15]), .Z(n154) );
  IV U175 ( .A(n155), .Z(n156) );
endmodule

