
module sum_N262144_CC64 ( clk, rst, a, b, c );
  input [4095:0] a;
  input [4095:0] b;
  output [4095:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        carry_on) );
  XOR U4 ( .A(a[3]), .B(n16374), .Z(n1056) );
  XOR U5 ( .A(a[6]), .B(n16365), .Z(n339) );
  XOR U6 ( .A(a[9]), .B(n16356), .Z(n6) );
  XOR U7 ( .A(a[12]), .B(n16347), .Z(n12156) );
  XOR U8 ( .A(a[15]), .B(n16338), .Z(n10923) );
  XOR U9 ( .A(a[18]), .B(n16329), .Z(n9690) );
  XOR U10 ( .A(a[21]), .B(n16320), .Z(n8456) );
  XOR U11 ( .A(a[24]), .B(n16311), .Z(n7223) );
  XOR U12 ( .A(a[27]), .B(n16302), .Z(n5990) );
  XOR U13 ( .A(a[30]), .B(n16293), .Z(n4756) );
  XOR U14 ( .A(a[33]), .B(n16284), .Z(n3523) );
  XOR U15 ( .A(a[36]), .B(n16275), .Z(n2290) );
  XOR U16 ( .A(a[39]), .B(n16266), .Z(n1057) );
  XOR U17 ( .A(a[42]), .B(n16257), .Z(n639) );
  XOR U18 ( .A(a[45]), .B(n16248), .Z(n606) );
  XOR U19 ( .A(a[48]), .B(n16239), .Z(n573) );
  XOR U20 ( .A(a[51]), .B(n16230), .Z(n539) );
  XOR U21 ( .A(a[54]), .B(n16221), .Z(n506) );
  XOR U22 ( .A(a[57]), .B(n16212), .Z(n473) );
  XOR U23 ( .A(a[60]), .B(n16203), .Z(n439) );
  XOR U24 ( .A(a[63]), .B(n16194), .Z(n406) );
  XOR U25 ( .A(a[66]), .B(n16185), .Z(n373) );
  XOR U26 ( .A(a[69]), .B(n16176), .Z(n340) );
  XOR U27 ( .A(a[72]), .B(n16167), .Z(n306) );
  XOR U28 ( .A(a[75]), .B(n16158), .Z(n273) );
  XOR U29 ( .A(a[78]), .B(n16149), .Z(n240) );
  XOR U30 ( .A(a[81]), .B(n16140), .Z(n206) );
  XOR U31 ( .A(a[84]), .B(n16131), .Z(n173) );
  XOR U32 ( .A(a[87]), .B(n16122), .Z(n140) );
  XOR U33 ( .A(a[90]), .B(n16113), .Z(n106) );
  XOR U34 ( .A(a[93]), .B(n16104), .Z(n73) );
  XOR U35 ( .A(a[96]), .B(n16095), .Z(n40) );
  XOR U36 ( .A(a[99]), .B(n16086), .Z(n7) );
  XOR U37 ( .A(a[102]), .B(n16077), .Z(n13266) );
  XOR U38 ( .A(a[105]), .B(n16068), .Z(n13143) );
  XOR U39 ( .A(a[108]), .B(n16059), .Z(n13020) );
  XOR U40 ( .A(a[111]), .B(n16050), .Z(n12896) );
  XOR U41 ( .A(a[114]), .B(n16041), .Z(n12773) );
  XOR U42 ( .A(a[117]), .B(n16032), .Z(n12650) );
  XOR U43 ( .A(a[120]), .B(n16023), .Z(n12526) );
  XOR U44 ( .A(a[123]), .B(n16014), .Z(n12403) );
  XOR U45 ( .A(a[126]), .B(n16005), .Z(n12280) );
  XOR U46 ( .A(a[129]), .B(n15996), .Z(n12157) );
  XOR U47 ( .A(a[132]), .B(n15987), .Z(n12033) );
  XOR U48 ( .A(a[135]), .B(n15978), .Z(n11910) );
  XOR U49 ( .A(a[138]), .B(n15969), .Z(n11787) );
  XOR U50 ( .A(a[141]), .B(n15960), .Z(n11663) );
  XOR U51 ( .A(a[144]), .B(n15951), .Z(n11540) );
  XOR U52 ( .A(a[147]), .B(n15942), .Z(n11417) );
  XOR U53 ( .A(a[150]), .B(n15933), .Z(n11293) );
  XOR U54 ( .A(a[153]), .B(n15924), .Z(n11170) );
  XOR U55 ( .A(a[156]), .B(n15915), .Z(n11047) );
  XOR U56 ( .A(a[159]), .B(n15906), .Z(n10924) );
  XOR U57 ( .A(a[162]), .B(n15897), .Z(n10800) );
  XOR U58 ( .A(a[165]), .B(n15888), .Z(n10677) );
  XOR U59 ( .A(a[168]), .B(n15879), .Z(n10554) );
  XOR U60 ( .A(a[171]), .B(n15870), .Z(n10430) );
  XOR U61 ( .A(a[174]), .B(n15861), .Z(n10307) );
  XOR U62 ( .A(a[177]), .B(n15852), .Z(n10184) );
  XOR U63 ( .A(a[180]), .B(n15843), .Z(n10060) );
  XOR U64 ( .A(a[183]), .B(n15834), .Z(n9937) );
  XOR U65 ( .A(a[186]), .B(n15825), .Z(n9814) );
  XOR U66 ( .A(a[189]), .B(n15816), .Z(n9691) );
  XOR U67 ( .A(a[192]), .B(n15807), .Z(n9567) );
  XOR U68 ( .A(a[195]), .B(n15798), .Z(n9444) );
  XOR U69 ( .A(a[198]), .B(n15789), .Z(n9321) );
  XOR U70 ( .A(a[201]), .B(n15780), .Z(n9196) );
  XOR U71 ( .A(a[204]), .B(n15771), .Z(n9073) );
  XOR U72 ( .A(a[207]), .B(n15762), .Z(n8950) );
  XOR U73 ( .A(a[210]), .B(n15753), .Z(n8826) );
  XOR U74 ( .A(a[213]), .B(n15744), .Z(n8703) );
  XOR U75 ( .A(a[216]), .B(n15735), .Z(n8580) );
  XOR U76 ( .A(a[219]), .B(n15726), .Z(n8457) );
  XOR U77 ( .A(a[222]), .B(n15717), .Z(n8333) );
  XOR U78 ( .A(a[225]), .B(n15708), .Z(n8210) );
  XOR U79 ( .A(a[228]), .B(n15699), .Z(n8087) );
  XOR U80 ( .A(a[231]), .B(n15690), .Z(n7963) );
  XOR U81 ( .A(a[234]), .B(n15681), .Z(n7840) );
  XOR U82 ( .A(a[237]), .B(n15672), .Z(n7717) );
  XOR U83 ( .A(a[240]), .B(n15663), .Z(n7593) );
  XOR U84 ( .A(a[243]), .B(n15654), .Z(n7470) );
  XOR U85 ( .A(a[246]), .B(n15645), .Z(n7347) );
  XOR U86 ( .A(a[249]), .B(n15636), .Z(n7224) );
  XOR U87 ( .A(a[252]), .B(n15627), .Z(n7100) );
  XOR U88 ( .A(a[255]), .B(n15618), .Z(n6977) );
  XOR U89 ( .A(a[258]), .B(n15609), .Z(n6854) );
  XOR U90 ( .A(a[261]), .B(n15600), .Z(n6730) );
  XOR U91 ( .A(a[264]), .B(n15591), .Z(n6607) );
  XOR U92 ( .A(a[267]), .B(n15582), .Z(n6484) );
  XOR U93 ( .A(a[270]), .B(n15573), .Z(n6360) );
  XOR U94 ( .A(a[273]), .B(n15564), .Z(n6237) );
  XOR U95 ( .A(a[276]), .B(n15555), .Z(n6114) );
  XOR U96 ( .A(a[279]), .B(n15546), .Z(n5991) );
  XOR U97 ( .A(a[282]), .B(n15537), .Z(n5867) );
  XOR U98 ( .A(a[285]), .B(n15528), .Z(n5744) );
  XOR U99 ( .A(a[288]), .B(n15519), .Z(n5621) );
  XOR U100 ( .A(a[291]), .B(n15510), .Z(n5497) );
  XOR U101 ( .A(a[294]), .B(n15501), .Z(n5374) );
  XOR U102 ( .A(a[297]), .B(n15492), .Z(n5251) );
  XOR U103 ( .A(a[300]), .B(n15483), .Z(n5126) );
  XOR U104 ( .A(a[303]), .B(n15474), .Z(n5003) );
  XOR U105 ( .A(a[306]), .B(n15465), .Z(n4880) );
  XOR U106 ( .A(a[309]), .B(n15456), .Z(n4757) );
  XOR U107 ( .A(a[312]), .B(n15447), .Z(n4633) );
  XOR U108 ( .A(a[315]), .B(n15438), .Z(n4510) );
  XOR U109 ( .A(a[318]), .B(n15429), .Z(n4387) );
  XOR U110 ( .A(a[321]), .B(n15420), .Z(n4263) );
  XOR U111 ( .A(a[324]), .B(n15411), .Z(n4140) );
  XOR U112 ( .A(a[327]), .B(n15402), .Z(n4017) );
  XOR U113 ( .A(a[330]), .B(n15393), .Z(n3893) );
  XOR U114 ( .A(a[333]), .B(n15384), .Z(n3770) );
  XOR U115 ( .A(a[336]), .B(n15375), .Z(n3647) );
  XOR U116 ( .A(a[339]), .B(n15366), .Z(n3524) );
  XOR U117 ( .A(a[342]), .B(n15357), .Z(n3400) );
  XOR U118 ( .A(a[345]), .B(n15348), .Z(n3277) );
  XOR U119 ( .A(a[348]), .B(n15339), .Z(n3154) );
  XOR U120 ( .A(a[351]), .B(n15330), .Z(n3030) );
  XOR U121 ( .A(a[354]), .B(n15321), .Z(n2907) );
  XOR U122 ( .A(a[357]), .B(n15312), .Z(n2784) );
  XOR U123 ( .A(a[360]), .B(n15303), .Z(n2660) );
  XOR U124 ( .A(a[363]), .B(n15294), .Z(n2537) );
  XOR U125 ( .A(a[366]), .B(n15285), .Z(n2414) );
  XOR U126 ( .A(a[369]), .B(n15276), .Z(n2291) );
  XOR U127 ( .A(a[372]), .B(n15267), .Z(n2167) );
  XOR U128 ( .A(a[375]), .B(n15258), .Z(n2044) );
  XOR U129 ( .A(a[378]), .B(n15249), .Z(n1921) );
  XOR U130 ( .A(a[381]), .B(n15240), .Z(n1797) );
  XOR U131 ( .A(a[384]), .B(n15231), .Z(n1674) );
  XOR U132 ( .A(a[387]), .B(n15222), .Z(n1551) );
  XOR U133 ( .A(a[390]), .B(n15213), .Z(n1427) );
  XOR U134 ( .A(a[393]), .B(n15204), .Z(n1304) );
  XOR U135 ( .A(a[396]), .B(n15195), .Z(n1181) );
  XOR U136 ( .A(a[399]), .B(n15186), .Z(n1058) );
  XOR U137 ( .A(a[402]), .B(n15177), .Z(n933) );
  XOR U138 ( .A(a[405]), .B(n15168), .Z(n810) );
  XOR U139 ( .A(a[408]), .B(n15159), .Z(n687) );
  XOR U140 ( .A(a[411]), .B(n15150), .Z(n659) );
  XOR U141 ( .A(a[414]), .B(n15141), .Z(n656) );
  XOR U142 ( .A(a[417]), .B(n15132), .Z(n653) );
  XOR U143 ( .A(a[420]), .B(n15123), .Z(n649) );
  XOR U144 ( .A(a[423]), .B(n15114), .Z(n646) );
  XOR U145 ( .A(a[426]), .B(n15105), .Z(n643) );
  XOR U146 ( .A(a[429]), .B(n15096), .Z(n640) );
  XOR U147 ( .A(a[432]), .B(n15087), .Z(n636) );
  XOR U148 ( .A(a[435]), .B(n15078), .Z(n633) );
  XOR U149 ( .A(a[438]), .B(n15069), .Z(n630) );
  XOR U150 ( .A(a[441]), .B(n15060), .Z(n626) );
  XOR U151 ( .A(a[444]), .B(n15051), .Z(n623) );
  XOR U152 ( .A(a[447]), .B(n15042), .Z(n620) );
  XOR U153 ( .A(a[450]), .B(n15033), .Z(n616) );
  XOR U154 ( .A(a[453]), .B(n15024), .Z(n613) );
  XOR U155 ( .A(a[456]), .B(n15015), .Z(n610) );
  XOR U156 ( .A(a[459]), .B(n15006), .Z(n607) );
  XOR U157 ( .A(a[462]), .B(n14997), .Z(n603) );
  XOR U158 ( .A(a[465]), .B(n14988), .Z(n600) );
  XOR U159 ( .A(a[468]), .B(n14979), .Z(n597) );
  XOR U160 ( .A(a[471]), .B(n14970), .Z(n593) );
  XOR U161 ( .A(a[474]), .B(n14961), .Z(n590) );
  XOR U162 ( .A(a[477]), .B(n14952), .Z(n587) );
  XOR U163 ( .A(a[480]), .B(n14943), .Z(n583) );
  XOR U164 ( .A(a[483]), .B(n14934), .Z(n580) );
  XOR U165 ( .A(a[486]), .B(n14925), .Z(n577) );
  XOR U166 ( .A(a[489]), .B(n14916), .Z(n574) );
  XOR U167 ( .A(a[492]), .B(n14907), .Z(n570) );
  XOR U168 ( .A(a[495]), .B(n14898), .Z(n567) );
  XOR U169 ( .A(a[498]), .B(n14889), .Z(n564) );
  XOR U170 ( .A(a[501]), .B(n14880), .Z(n559) );
  XOR U171 ( .A(a[504]), .B(n14871), .Z(n556) );
  XOR U172 ( .A(a[507]), .B(n14862), .Z(n553) );
  XOR U173 ( .A(a[510]), .B(n14853), .Z(n549) );
  XOR U174 ( .A(a[513]), .B(n14844), .Z(n546) );
  XOR U175 ( .A(a[516]), .B(n14835), .Z(n543) );
  XOR U176 ( .A(a[519]), .B(n14826), .Z(n540) );
  XOR U177 ( .A(a[522]), .B(n14817), .Z(n536) );
  XOR U178 ( .A(a[525]), .B(n14808), .Z(n533) );
  XOR U179 ( .A(a[528]), .B(n14799), .Z(n530) );
  XOR U180 ( .A(a[531]), .B(n14790), .Z(n526) );
  XOR U181 ( .A(a[534]), .B(n14781), .Z(n523) );
  XOR U182 ( .A(a[537]), .B(n14772), .Z(n520) );
  XOR U183 ( .A(a[540]), .B(n14763), .Z(n516) );
  XOR U184 ( .A(a[543]), .B(n14754), .Z(n513) );
  XOR U185 ( .A(a[546]), .B(n14745), .Z(n510) );
  XOR U186 ( .A(a[549]), .B(n14736), .Z(n507) );
  XOR U187 ( .A(a[552]), .B(n14727), .Z(n503) );
  XOR U188 ( .A(a[555]), .B(n14718), .Z(n500) );
  XOR U189 ( .A(a[558]), .B(n14709), .Z(n497) );
  XOR U190 ( .A(a[561]), .B(n14700), .Z(n493) );
  XOR U191 ( .A(a[564]), .B(n14691), .Z(n490) );
  XOR U192 ( .A(a[567]), .B(n14682), .Z(n487) );
  XOR U193 ( .A(a[570]), .B(n14673), .Z(n483) );
  XOR U194 ( .A(a[573]), .B(n14664), .Z(n480) );
  XOR U195 ( .A(a[576]), .B(n14655), .Z(n477) );
  XOR U196 ( .A(a[579]), .B(n14646), .Z(n474) );
  XOR U197 ( .A(a[582]), .B(n14637), .Z(n470) );
  XOR U198 ( .A(a[585]), .B(n14628), .Z(n467) );
  XOR U199 ( .A(a[588]), .B(n14619), .Z(n464) );
  XOR U200 ( .A(a[591]), .B(n14610), .Z(n460) );
  XOR U201 ( .A(a[594]), .B(n14601), .Z(n457) );
  XOR U202 ( .A(a[597]), .B(n14592), .Z(n454) );
  XOR U203 ( .A(a[600]), .B(n14583), .Z(n449) );
  XOR U204 ( .A(a[603]), .B(n14574), .Z(n446) );
  XOR U205 ( .A(a[606]), .B(n14565), .Z(n443) );
  XOR U206 ( .A(a[609]), .B(n14556), .Z(n440) );
  XOR U207 ( .A(a[612]), .B(n14547), .Z(n436) );
  XOR U208 ( .A(a[615]), .B(n14538), .Z(n433) );
  XOR U209 ( .A(a[618]), .B(n14529), .Z(n430) );
  XOR U210 ( .A(a[621]), .B(n14520), .Z(n426) );
  XOR U211 ( .A(a[624]), .B(n14511), .Z(n423) );
  XOR U212 ( .A(a[627]), .B(n14502), .Z(n420) );
  XOR U213 ( .A(a[630]), .B(n14493), .Z(n416) );
  XOR U214 ( .A(a[633]), .B(n14484), .Z(n413) );
  XOR U215 ( .A(a[636]), .B(n14475), .Z(n410) );
  XOR U216 ( .A(a[639]), .B(n14466), .Z(n407) );
  XOR U217 ( .A(a[642]), .B(n14457), .Z(n403) );
  XOR U218 ( .A(a[645]), .B(n14448), .Z(n400) );
  XOR U219 ( .A(a[648]), .B(n14439), .Z(n397) );
  XOR U220 ( .A(a[651]), .B(n14430), .Z(n393) );
  XOR U221 ( .A(a[654]), .B(n14421), .Z(n390) );
  XOR U222 ( .A(a[657]), .B(n14412), .Z(n387) );
  XOR U223 ( .A(a[660]), .B(n14403), .Z(n383) );
  XOR U224 ( .A(a[663]), .B(n14394), .Z(n380) );
  XOR U225 ( .A(a[666]), .B(n14385), .Z(n377) );
  XOR U226 ( .A(a[669]), .B(n14376), .Z(n374) );
  XOR U227 ( .A(a[672]), .B(n14367), .Z(n370) );
  XOR U228 ( .A(a[675]), .B(n14358), .Z(n367) );
  XOR U229 ( .A(a[678]), .B(n14349), .Z(n364) );
  XOR U230 ( .A(a[681]), .B(n14340), .Z(n360) );
  XOR U231 ( .A(a[684]), .B(n14331), .Z(n357) );
  XOR U232 ( .A(a[687]), .B(n14322), .Z(n354) );
  XOR U233 ( .A(a[690]), .B(n14313), .Z(n350) );
  XOR U234 ( .A(a[693]), .B(n14304), .Z(n347) );
  XOR U235 ( .A(a[696]), .B(n14295), .Z(n344) );
  XOR U236 ( .A(a[699]), .B(n14286), .Z(n341) );
  XOR U237 ( .A(a[702]), .B(n14277), .Z(n336) );
  XOR U238 ( .A(a[705]), .B(n14268), .Z(n333) );
  XOR U239 ( .A(a[708]), .B(n14259), .Z(n330) );
  XOR U240 ( .A(a[711]), .B(n14250), .Z(n326) );
  XOR U241 ( .A(a[714]), .B(n14241), .Z(n323) );
  XOR U242 ( .A(a[717]), .B(n14232), .Z(n320) );
  XOR U243 ( .A(a[720]), .B(n14223), .Z(n316) );
  XOR U244 ( .A(a[723]), .B(n14214), .Z(n313) );
  XOR U245 ( .A(a[726]), .B(n14205), .Z(n310) );
  XOR U246 ( .A(a[729]), .B(n14196), .Z(n307) );
  XOR U247 ( .A(a[732]), .B(n14187), .Z(n303) );
  XOR U248 ( .A(a[735]), .B(n14178), .Z(n300) );
  XOR U249 ( .A(a[738]), .B(n14169), .Z(n297) );
  XOR U250 ( .A(a[741]), .B(n14160), .Z(n293) );
  XOR U251 ( .A(a[744]), .B(n14151), .Z(n290) );
  XOR U252 ( .A(a[747]), .B(n14142), .Z(n287) );
  XOR U253 ( .A(a[750]), .B(n14133), .Z(n283) );
  XOR U254 ( .A(a[753]), .B(n14124), .Z(n280) );
  XOR U255 ( .A(a[756]), .B(n14115), .Z(n277) );
  XOR U256 ( .A(a[759]), .B(n14106), .Z(n274) );
  XOR U257 ( .A(a[762]), .B(n14097), .Z(n270) );
  XOR U258 ( .A(a[765]), .B(n14088), .Z(n267) );
  XOR U259 ( .A(a[768]), .B(n14079), .Z(n264) );
  XOR U260 ( .A(a[771]), .B(n14070), .Z(n260) );
  XOR U261 ( .A(a[774]), .B(n14061), .Z(n257) );
  XOR U262 ( .A(a[777]), .B(n14052), .Z(n254) );
  XOR U263 ( .A(a[780]), .B(n14043), .Z(n250) );
  XOR U264 ( .A(a[783]), .B(n14034), .Z(n247) );
  XOR U265 ( .A(a[786]), .B(n14025), .Z(n244) );
  XOR U266 ( .A(a[789]), .B(n14016), .Z(n241) );
  XOR U267 ( .A(a[792]), .B(n14007), .Z(n237) );
  XOR U268 ( .A(a[795]), .B(n13998), .Z(n234) );
  XOR U269 ( .A(a[798]), .B(n13989), .Z(n231) );
  XOR U270 ( .A(a[801]), .B(n13980), .Z(n226) );
  XOR U271 ( .A(a[804]), .B(n13971), .Z(n223) );
  XOR U272 ( .A(a[807]), .B(n13962), .Z(n220) );
  XOR U273 ( .A(a[810]), .B(n13953), .Z(n216) );
  XOR U274 ( .A(a[813]), .B(n13944), .Z(n213) );
  XOR U275 ( .A(a[816]), .B(n13935), .Z(n210) );
  XOR U276 ( .A(a[819]), .B(n13926), .Z(n207) );
  XOR U277 ( .A(a[822]), .B(n13917), .Z(n203) );
  XOR U278 ( .A(a[825]), .B(n13908), .Z(n200) );
  XOR U279 ( .A(a[828]), .B(n13899), .Z(n197) );
  XOR U280 ( .A(a[831]), .B(n13890), .Z(n193) );
  XOR U281 ( .A(a[834]), .B(n13881), .Z(n190) );
  XOR U282 ( .A(a[837]), .B(n13872), .Z(n187) );
  XOR U283 ( .A(a[840]), .B(n13863), .Z(n183) );
  XOR U284 ( .A(a[843]), .B(n13854), .Z(n180) );
  XOR U285 ( .A(a[846]), .B(n13845), .Z(n177) );
  XOR U286 ( .A(a[849]), .B(n13836), .Z(n174) );
  XOR U287 ( .A(a[852]), .B(n13827), .Z(n170) );
  XOR U288 ( .A(a[855]), .B(n13818), .Z(n167) );
  XOR U289 ( .A(a[858]), .B(n13809), .Z(n164) );
  XOR U290 ( .A(a[861]), .B(n13800), .Z(n160) );
  XOR U291 ( .A(a[864]), .B(n13791), .Z(n157) );
  XOR U292 ( .A(a[867]), .B(n13782), .Z(n154) );
  XOR U293 ( .A(a[870]), .B(n13773), .Z(n150) );
  XOR U294 ( .A(a[873]), .B(n13764), .Z(n147) );
  XOR U295 ( .A(a[876]), .B(n13755), .Z(n144) );
  XOR U296 ( .A(a[879]), .B(n13746), .Z(n141) );
  XOR U297 ( .A(a[882]), .B(n13737), .Z(n137) );
  XOR U298 ( .A(a[885]), .B(n13728), .Z(n134) );
  XOR U299 ( .A(a[888]), .B(n13719), .Z(n131) );
  XOR U300 ( .A(a[891]), .B(n13710), .Z(n127) );
  XOR U301 ( .A(a[894]), .B(n13701), .Z(n124) );
  XOR U302 ( .A(a[897]), .B(n13692), .Z(n121) );
  XOR U303 ( .A(a[900]), .B(n13683), .Z(n116) );
  XOR U304 ( .A(a[903]), .B(n13674), .Z(n113) );
  XOR U305 ( .A(a[906]), .B(n13665), .Z(n110) );
  XOR U306 ( .A(a[909]), .B(n13656), .Z(n107) );
  XOR U307 ( .A(a[912]), .B(n13647), .Z(n103) );
  XOR U308 ( .A(a[915]), .B(n13638), .Z(n100) );
  XOR U309 ( .A(a[918]), .B(n13629), .Z(n97) );
  XOR U310 ( .A(a[921]), .B(n13620), .Z(n93) );
  XOR U311 ( .A(a[924]), .B(n13611), .Z(n90) );
  XOR U312 ( .A(a[927]), .B(n13602), .Z(n87) );
  XOR U313 ( .A(a[930]), .B(n13593), .Z(n83) );
  XOR U314 ( .A(a[933]), .B(n13584), .Z(n80) );
  XOR U315 ( .A(a[936]), .B(n13575), .Z(n77) );
  XOR U316 ( .A(a[939]), .B(n13566), .Z(n74) );
  XOR U317 ( .A(a[942]), .B(n13557), .Z(n70) );
  XOR U318 ( .A(a[945]), .B(n13548), .Z(n67) );
  XOR U319 ( .A(a[948]), .B(n13539), .Z(n64) );
  XOR U320 ( .A(a[951]), .B(n13530), .Z(n60) );
  XOR U321 ( .A(a[954]), .B(n13521), .Z(n57) );
  XOR U322 ( .A(a[957]), .B(n13512), .Z(n54) );
  XOR U323 ( .A(a[960]), .B(n13503), .Z(n50) );
  XOR U324 ( .A(a[963]), .B(n13494), .Z(n47) );
  XOR U325 ( .A(a[966]), .B(n13485), .Z(n44) );
  XOR U326 ( .A(a[969]), .B(n13476), .Z(n41) );
  XOR U327 ( .A(a[972]), .B(n13467), .Z(n37) );
  XOR U328 ( .A(a[975]), .B(n13458), .Z(n34) );
  XOR U329 ( .A(a[978]), .B(n13449), .Z(n31) );
  XOR U330 ( .A(a[981]), .B(n13440), .Z(n27) );
  XOR U331 ( .A(a[984]), .B(n13431), .Z(n24) );
  XOR U332 ( .A(a[987]), .B(n13422), .Z(n21) );
  XOR U333 ( .A(a[990]), .B(n13413), .Z(n17) );
  XOR U334 ( .A(a[993]), .B(n13404), .Z(n14) );
  XOR U335 ( .A(a[996]), .B(n13395), .Z(n11) );
  XOR U336 ( .A(a[999]), .B(n13386), .Z(n8) );
  XOR U337 ( .A(a[1002]), .B(n13374), .Z(n13376) );
  XOR U338 ( .A(a[1005]), .B(n13362), .Z(n13364) );
  XOR U339 ( .A(a[1008]), .B(n13350), .Z(n13352) );
  XOR U340 ( .A(a[1011]), .B(n13337), .Z(n13339) );
  XOR U341 ( .A(a[1014]), .B(n13325), .Z(n13327) );
  XOR U342 ( .A(a[1017]), .B(n13313), .Z(n13315) );
  XOR U343 ( .A(a[1020]), .B(n13300), .Z(n13302) );
  XOR U344 ( .A(a[1023]), .B(n13288), .Z(n13290) );
  XOR U345 ( .A(a[1026]), .B(n13276), .Z(n13278) );
  XOR U346 ( .A(a[1029]), .B(n13263), .Z(n13265) );
  XOR U347 ( .A(a[1032]), .B(n13251), .Z(n13253) );
  XOR U348 ( .A(a[1035]), .B(n13239), .Z(n13241) );
  XOR U349 ( .A(a[1038]), .B(n13227), .Z(n13229) );
  XOR U350 ( .A(a[1041]), .B(n13214), .Z(n13216) );
  XOR U351 ( .A(a[1044]), .B(n13202), .Z(n13204) );
  XOR U352 ( .A(a[1047]), .B(n13190), .Z(n13192) );
  XOR U353 ( .A(a[1050]), .B(n13177), .Z(n13179) );
  XOR U354 ( .A(a[1053]), .B(n13165), .Z(n13167) );
  XOR U355 ( .A(a[1056]), .B(n13153), .Z(n13155) );
  XOR U356 ( .A(a[1059]), .B(n13140), .Z(n13142) );
  XOR U357 ( .A(a[1062]), .B(n13128), .Z(n13130) );
  XOR U358 ( .A(a[1065]), .B(n13116), .Z(n13118) );
  XOR U359 ( .A(a[1068]), .B(n13104), .Z(n13106) );
  XOR U360 ( .A(a[1071]), .B(n13091), .Z(n13093) );
  XOR U361 ( .A(a[1074]), .B(n13079), .Z(n13081) );
  XOR U362 ( .A(a[1077]), .B(n13067), .Z(n13069) );
  XOR U363 ( .A(a[1080]), .B(n13054), .Z(n13056) );
  XOR U364 ( .A(a[1083]), .B(n13042), .Z(n13044) );
  XOR U365 ( .A(a[1086]), .B(n13030), .Z(n13032) );
  XOR U366 ( .A(a[1089]), .B(n13017), .Z(n13019) );
  XOR U367 ( .A(a[1092]), .B(n13005), .Z(n13007) );
  XOR U368 ( .A(a[1095]), .B(n12993), .Z(n12995) );
  XOR U369 ( .A(a[1098]), .B(n12981), .Z(n12983) );
  XOR U370 ( .A(a[1101]), .B(n12967), .Z(n12969) );
  XOR U371 ( .A(a[1104]), .B(n12955), .Z(n12957) );
  XOR U372 ( .A(a[1107]), .B(n12943), .Z(n12945) );
  XOR U373 ( .A(a[1110]), .B(n12930), .Z(n12932) );
  XOR U374 ( .A(a[1113]), .B(n12918), .Z(n12920) );
  XOR U375 ( .A(a[1116]), .B(n12906), .Z(n12908) );
  XOR U376 ( .A(a[1119]), .B(n12893), .Z(n12895) );
  XOR U377 ( .A(a[1122]), .B(n12881), .Z(n12883) );
  XOR U378 ( .A(a[1125]), .B(n12869), .Z(n12871) );
  XOR U379 ( .A(a[1128]), .B(n12857), .Z(n12859) );
  XOR U380 ( .A(a[1131]), .B(n12844), .Z(n12846) );
  XOR U381 ( .A(a[1134]), .B(n12832), .Z(n12834) );
  XOR U382 ( .A(a[1137]), .B(n12820), .Z(n12822) );
  XOR U383 ( .A(a[1140]), .B(n12807), .Z(n12809) );
  XOR U384 ( .A(a[1143]), .B(n12795), .Z(n12797) );
  XOR U385 ( .A(a[1146]), .B(n12783), .Z(n12785) );
  XOR U386 ( .A(a[1149]), .B(n12770), .Z(n12772) );
  XOR U387 ( .A(a[1152]), .B(n12758), .Z(n12760) );
  XOR U388 ( .A(a[1155]), .B(n12746), .Z(n12748) );
  XOR U389 ( .A(a[1158]), .B(n12734), .Z(n12736) );
  XOR U390 ( .A(a[1161]), .B(n12721), .Z(n12723) );
  XOR U391 ( .A(a[1164]), .B(n12709), .Z(n12711) );
  XOR U392 ( .A(a[1167]), .B(n12697), .Z(n12699) );
  XOR U393 ( .A(a[1170]), .B(n12684), .Z(n12686) );
  XOR U394 ( .A(a[1173]), .B(n12672), .Z(n12674) );
  XOR U395 ( .A(a[1176]), .B(n12660), .Z(n12662) );
  XOR U396 ( .A(a[1179]), .B(n12647), .Z(n12649) );
  XOR U397 ( .A(a[1182]), .B(n12635), .Z(n12637) );
  XOR U398 ( .A(a[1185]), .B(n12623), .Z(n12625) );
  XOR U399 ( .A(a[1188]), .B(n12611), .Z(n12613) );
  XOR U400 ( .A(a[1191]), .B(n12598), .Z(n12600) );
  XOR U401 ( .A(a[1194]), .B(n12586), .Z(n12588) );
  XOR U402 ( .A(a[1197]), .B(n12574), .Z(n12576) );
  XOR U403 ( .A(a[1200]), .B(n12560), .Z(n12562) );
  XOR U404 ( .A(a[1203]), .B(n12548), .Z(n12550) );
  XOR U405 ( .A(a[1206]), .B(n12536), .Z(n12538) );
  XOR U406 ( .A(a[1209]), .B(n12523), .Z(n12525) );
  XOR U407 ( .A(a[1212]), .B(n12511), .Z(n12513) );
  XOR U408 ( .A(a[1215]), .B(n12499), .Z(n12501) );
  XOR U409 ( .A(a[1218]), .B(n12487), .Z(n12489) );
  XOR U410 ( .A(a[1221]), .B(n12474), .Z(n12476) );
  XOR U411 ( .A(a[1224]), .B(n12462), .Z(n12464) );
  XOR U412 ( .A(a[1227]), .B(n12450), .Z(n12452) );
  XOR U413 ( .A(a[1230]), .B(n12437), .Z(n12439) );
  XOR U414 ( .A(a[1233]), .B(n12425), .Z(n12427) );
  XOR U415 ( .A(a[1236]), .B(n12413), .Z(n12415) );
  XOR U416 ( .A(a[1239]), .B(n12400), .Z(n12402) );
  XOR U417 ( .A(a[1242]), .B(n12388), .Z(n12390) );
  XOR U418 ( .A(a[1245]), .B(n12376), .Z(n12378) );
  XOR U419 ( .A(a[1248]), .B(n12364), .Z(n12366) );
  XOR U420 ( .A(a[1251]), .B(n12351), .Z(n12353) );
  XOR U421 ( .A(a[1254]), .B(n12339), .Z(n12341) );
  XOR U422 ( .A(a[1257]), .B(n12327), .Z(n12329) );
  XOR U423 ( .A(a[1260]), .B(n12314), .Z(n12316) );
  XOR U424 ( .A(a[1263]), .B(n12302), .Z(n12304) );
  XOR U425 ( .A(a[1266]), .B(n12290), .Z(n12292) );
  XOR U426 ( .A(a[1269]), .B(n12277), .Z(n12279) );
  XOR U427 ( .A(a[1272]), .B(n12265), .Z(n12267) );
  XOR U428 ( .A(a[1275]), .B(n12253), .Z(n12255) );
  XOR U429 ( .A(a[1278]), .B(n12241), .Z(n12243) );
  XOR U430 ( .A(a[1281]), .B(n12228), .Z(n12230) );
  XOR U431 ( .A(a[1284]), .B(n12216), .Z(n12218) );
  XOR U432 ( .A(a[1287]), .B(n12204), .Z(n12206) );
  XOR U433 ( .A(a[1290]), .B(n12191), .Z(n12193) );
  XOR U434 ( .A(a[1293]), .B(n12179), .Z(n12181) );
  XOR U435 ( .A(a[1296]), .B(n12167), .Z(n12169) );
  XOR U436 ( .A(a[1299]), .B(n12153), .Z(n12155) );
  XOR U437 ( .A(a[1302]), .B(n12141), .Z(n12143) );
  XOR U438 ( .A(a[1305]), .B(n12129), .Z(n12131) );
  XOR U439 ( .A(a[1308]), .B(n12117), .Z(n12119) );
  XOR U440 ( .A(a[1311]), .B(n12104), .Z(n12106) );
  XOR U441 ( .A(a[1314]), .B(n12092), .Z(n12094) );
  XOR U442 ( .A(a[1317]), .B(n12080), .Z(n12082) );
  XOR U443 ( .A(a[1320]), .B(n12067), .Z(n12069) );
  XOR U444 ( .A(a[1323]), .B(n12055), .Z(n12057) );
  XOR U445 ( .A(a[1326]), .B(n12043), .Z(n12045) );
  XOR U446 ( .A(a[1329]), .B(n12030), .Z(n12032) );
  XOR U447 ( .A(a[1332]), .B(n12018), .Z(n12020) );
  XOR U448 ( .A(a[1335]), .B(n12006), .Z(n12008) );
  XOR U449 ( .A(a[1338]), .B(n11994), .Z(n11996) );
  XOR U450 ( .A(a[1341]), .B(n11981), .Z(n11983) );
  XOR U451 ( .A(a[1344]), .B(n11969), .Z(n11971) );
  XOR U452 ( .A(a[1347]), .B(n11957), .Z(n11959) );
  XOR U453 ( .A(a[1350]), .B(n11944), .Z(n11946) );
  XOR U454 ( .A(a[1353]), .B(n11932), .Z(n11934) );
  XOR U455 ( .A(a[1356]), .B(n11920), .Z(n11922) );
  XOR U456 ( .A(a[1359]), .B(n11907), .Z(n11909) );
  XOR U457 ( .A(a[1362]), .B(n11895), .Z(n11897) );
  XOR U458 ( .A(a[1365]), .B(n11883), .Z(n11885) );
  XOR U459 ( .A(a[1368]), .B(n11871), .Z(n11873) );
  XOR U460 ( .A(a[1371]), .B(n11858), .Z(n11860) );
  XOR U461 ( .A(a[1374]), .B(n11846), .Z(n11848) );
  XOR U462 ( .A(a[1377]), .B(n11834), .Z(n11836) );
  XOR U463 ( .A(a[1380]), .B(n11821), .Z(n11823) );
  XOR U464 ( .A(a[1383]), .B(n11809), .Z(n11811) );
  XOR U465 ( .A(a[1386]), .B(n11797), .Z(n11799) );
  XOR U466 ( .A(a[1389]), .B(n11784), .Z(n11786) );
  XOR U467 ( .A(a[1392]), .B(n11772), .Z(n11774) );
  XOR U468 ( .A(a[1395]), .B(n11760), .Z(n11762) );
  XOR U469 ( .A(a[1398]), .B(n11748), .Z(n11750) );
  XOR U470 ( .A(a[1401]), .B(n11734), .Z(n11736) );
  XOR U471 ( .A(a[1404]), .B(n11722), .Z(n11724) );
  XOR U472 ( .A(a[1407]), .B(n11710), .Z(n11712) );
  XOR U473 ( .A(a[1410]), .B(n11697), .Z(n11699) );
  XOR U474 ( .A(a[1413]), .B(n11685), .Z(n11687) );
  XOR U475 ( .A(a[1416]), .B(n11673), .Z(n11675) );
  XOR U476 ( .A(a[1419]), .B(n11660), .Z(n11662) );
  XOR U477 ( .A(a[1422]), .B(n11648), .Z(n11650) );
  XOR U478 ( .A(a[1425]), .B(n11636), .Z(n11638) );
  XOR U479 ( .A(a[1428]), .B(n11624), .Z(n11626) );
  XOR U480 ( .A(a[1431]), .B(n11611), .Z(n11613) );
  XOR U481 ( .A(a[1434]), .B(n11599), .Z(n11601) );
  XOR U482 ( .A(a[1437]), .B(n11587), .Z(n11589) );
  XOR U483 ( .A(a[1440]), .B(n11574), .Z(n11576) );
  XOR U484 ( .A(a[1443]), .B(n11562), .Z(n11564) );
  XOR U485 ( .A(a[1446]), .B(n11550), .Z(n11552) );
  XOR U486 ( .A(a[1449]), .B(n11537), .Z(n11539) );
  XOR U487 ( .A(a[1452]), .B(n11525), .Z(n11527) );
  XOR U488 ( .A(a[1455]), .B(n11513), .Z(n11515) );
  XOR U489 ( .A(a[1458]), .B(n11501), .Z(n11503) );
  XOR U490 ( .A(a[1461]), .B(n11488), .Z(n11490) );
  XOR U491 ( .A(a[1464]), .B(n11476), .Z(n11478) );
  XOR U492 ( .A(a[1467]), .B(n11464), .Z(n11466) );
  XOR U493 ( .A(a[1470]), .B(n11451), .Z(n11453) );
  XOR U494 ( .A(a[1473]), .B(n11439), .Z(n11441) );
  XOR U495 ( .A(a[1476]), .B(n11427), .Z(n11429) );
  XOR U496 ( .A(a[1479]), .B(n11414), .Z(n11416) );
  XOR U497 ( .A(a[1482]), .B(n11402), .Z(n11404) );
  XOR U498 ( .A(a[1485]), .B(n11390), .Z(n11392) );
  XOR U499 ( .A(a[1488]), .B(n11378), .Z(n11380) );
  XOR U500 ( .A(a[1491]), .B(n11365), .Z(n11367) );
  XOR U501 ( .A(a[1494]), .B(n11353), .Z(n11355) );
  XOR U502 ( .A(a[1497]), .B(n11341), .Z(n11343) );
  XOR U503 ( .A(a[1500]), .B(n11327), .Z(n11329) );
  XOR U504 ( .A(a[1503]), .B(n11315), .Z(n11317) );
  XOR U505 ( .A(a[1506]), .B(n11303), .Z(n11305) );
  XOR U506 ( .A(a[1509]), .B(n11290), .Z(n11292) );
  XOR U507 ( .A(a[1512]), .B(n11278), .Z(n11280) );
  XOR U508 ( .A(a[1515]), .B(n11266), .Z(n11268) );
  XOR U509 ( .A(a[1518]), .B(n11254), .Z(n11256) );
  XOR U510 ( .A(a[1521]), .B(n11241), .Z(n11243) );
  XOR U511 ( .A(a[1524]), .B(n11229), .Z(n11231) );
  XOR U512 ( .A(a[1527]), .B(n11217), .Z(n11219) );
  XOR U513 ( .A(a[1530]), .B(n11204), .Z(n11206) );
  XOR U514 ( .A(a[1533]), .B(n11192), .Z(n11194) );
  XOR U515 ( .A(a[1536]), .B(n11180), .Z(n11182) );
  XOR U516 ( .A(a[1539]), .B(n11167), .Z(n11169) );
  XOR U517 ( .A(a[1542]), .B(n11155), .Z(n11157) );
  XOR U518 ( .A(a[1545]), .B(n11143), .Z(n11145) );
  XOR U519 ( .A(a[1548]), .B(n11131), .Z(n11133) );
  XOR U520 ( .A(a[1551]), .B(n11118), .Z(n11120) );
  XOR U521 ( .A(a[1554]), .B(n11106), .Z(n11108) );
  XOR U522 ( .A(a[1557]), .B(n11094), .Z(n11096) );
  XOR U523 ( .A(a[1560]), .B(n11081), .Z(n11083) );
  XOR U524 ( .A(a[1563]), .B(n11069), .Z(n11071) );
  XOR U525 ( .A(a[1566]), .B(n11057), .Z(n11059) );
  XOR U526 ( .A(a[1569]), .B(n11044), .Z(n11046) );
  XOR U527 ( .A(a[1572]), .B(n11032), .Z(n11034) );
  XOR U528 ( .A(a[1575]), .B(n11020), .Z(n11022) );
  XOR U529 ( .A(a[1578]), .B(n11008), .Z(n11010) );
  XOR U530 ( .A(a[1581]), .B(n10995), .Z(n10997) );
  XOR U531 ( .A(a[1584]), .B(n10983), .Z(n10985) );
  XOR U532 ( .A(a[1587]), .B(n10971), .Z(n10973) );
  XOR U533 ( .A(a[1590]), .B(n10958), .Z(n10960) );
  XOR U534 ( .A(a[1593]), .B(n10946), .Z(n10948) );
  XOR U535 ( .A(a[1596]), .B(n10934), .Z(n10936) );
  XOR U536 ( .A(a[1599]), .B(n10920), .Z(n10922) );
  XOR U537 ( .A(a[1602]), .B(n10908), .Z(n10910) );
  XOR U538 ( .A(a[1605]), .B(n10896), .Z(n10898) );
  XOR U539 ( .A(a[1608]), .B(n10884), .Z(n10886) );
  XOR U540 ( .A(a[1611]), .B(n10871), .Z(n10873) );
  XOR U541 ( .A(a[1614]), .B(n10859), .Z(n10861) );
  XOR U542 ( .A(a[1617]), .B(n10847), .Z(n10849) );
  XOR U543 ( .A(a[1620]), .B(n10834), .Z(n10836) );
  XOR U544 ( .A(a[1623]), .B(n10822), .Z(n10824) );
  XOR U545 ( .A(a[1626]), .B(n10810), .Z(n10812) );
  XOR U546 ( .A(a[1629]), .B(n10797), .Z(n10799) );
  XOR U547 ( .A(a[1632]), .B(n10785), .Z(n10787) );
  XOR U548 ( .A(a[1635]), .B(n10773), .Z(n10775) );
  XOR U549 ( .A(a[1638]), .B(n10761), .Z(n10763) );
  XOR U550 ( .A(a[1641]), .B(n10748), .Z(n10750) );
  XOR U551 ( .A(a[1644]), .B(n10736), .Z(n10738) );
  XOR U552 ( .A(a[1647]), .B(n10724), .Z(n10726) );
  XOR U553 ( .A(a[1650]), .B(n10711), .Z(n10713) );
  XOR U554 ( .A(a[1653]), .B(n10699), .Z(n10701) );
  XOR U555 ( .A(a[1656]), .B(n10687), .Z(n10689) );
  XOR U556 ( .A(a[1659]), .B(n10674), .Z(n10676) );
  XOR U557 ( .A(a[1662]), .B(n10662), .Z(n10664) );
  XOR U558 ( .A(a[1665]), .B(n10650), .Z(n10652) );
  XOR U559 ( .A(a[1668]), .B(n10638), .Z(n10640) );
  XOR U560 ( .A(a[1671]), .B(n10625), .Z(n10627) );
  XOR U561 ( .A(a[1674]), .B(n10613), .Z(n10615) );
  XOR U562 ( .A(a[1677]), .B(n10601), .Z(n10603) );
  XOR U563 ( .A(a[1680]), .B(n10588), .Z(n10590) );
  XOR U564 ( .A(a[1683]), .B(n10576), .Z(n10578) );
  XOR U565 ( .A(a[1686]), .B(n10564), .Z(n10566) );
  XOR U566 ( .A(a[1689]), .B(n10551), .Z(n10553) );
  XOR U567 ( .A(a[1692]), .B(n10539), .Z(n10541) );
  XOR U568 ( .A(a[1695]), .B(n10527), .Z(n10529) );
  XOR U569 ( .A(a[1698]), .B(n10515), .Z(n10517) );
  XOR U570 ( .A(a[1701]), .B(n10501), .Z(n10503) );
  XOR U571 ( .A(a[1704]), .B(n10489), .Z(n10491) );
  XOR U572 ( .A(a[1707]), .B(n10477), .Z(n10479) );
  XOR U573 ( .A(a[1710]), .B(n10464), .Z(n10466) );
  XOR U574 ( .A(a[1713]), .B(n10452), .Z(n10454) );
  XOR U575 ( .A(a[1716]), .B(n10440), .Z(n10442) );
  XOR U576 ( .A(a[1719]), .B(n10427), .Z(n10429) );
  XOR U577 ( .A(a[1722]), .B(n10415), .Z(n10417) );
  XOR U578 ( .A(a[1725]), .B(n10403), .Z(n10405) );
  XOR U579 ( .A(a[1728]), .B(n10391), .Z(n10393) );
  XOR U580 ( .A(a[1731]), .B(n10378), .Z(n10380) );
  XOR U581 ( .A(a[1734]), .B(n10366), .Z(n10368) );
  XOR U582 ( .A(a[1737]), .B(n10354), .Z(n10356) );
  XOR U583 ( .A(a[1740]), .B(n10341), .Z(n10343) );
  XOR U584 ( .A(a[1743]), .B(n10329), .Z(n10331) );
  XOR U585 ( .A(a[1746]), .B(n10317), .Z(n10319) );
  XOR U586 ( .A(a[1749]), .B(n10304), .Z(n10306) );
  XOR U587 ( .A(a[1752]), .B(n10292), .Z(n10294) );
  XOR U588 ( .A(a[1755]), .B(n10280), .Z(n10282) );
  XOR U589 ( .A(a[1758]), .B(n10268), .Z(n10270) );
  XOR U590 ( .A(a[1761]), .B(n10255), .Z(n10257) );
  XOR U591 ( .A(a[1764]), .B(n10243), .Z(n10245) );
  XOR U592 ( .A(a[1767]), .B(n10231), .Z(n10233) );
  XOR U593 ( .A(a[1770]), .B(n10218), .Z(n10220) );
  XOR U594 ( .A(a[1773]), .B(n10206), .Z(n10208) );
  XOR U595 ( .A(a[1776]), .B(n10194), .Z(n10196) );
  XOR U596 ( .A(a[1779]), .B(n10181), .Z(n10183) );
  XOR U597 ( .A(a[1782]), .B(n10169), .Z(n10171) );
  XOR U598 ( .A(a[1785]), .B(n10157), .Z(n10159) );
  XOR U599 ( .A(a[1788]), .B(n10145), .Z(n10147) );
  XOR U600 ( .A(a[1791]), .B(n10132), .Z(n10134) );
  XOR U601 ( .A(a[1794]), .B(n10120), .Z(n10122) );
  XOR U602 ( .A(a[1797]), .B(n10108), .Z(n10110) );
  XOR U603 ( .A(a[1800]), .B(n10094), .Z(n10096) );
  XOR U604 ( .A(a[1803]), .B(n10082), .Z(n10084) );
  XOR U605 ( .A(a[1806]), .B(n10070), .Z(n10072) );
  XOR U606 ( .A(a[1809]), .B(n10057), .Z(n10059) );
  XOR U607 ( .A(a[1812]), .B(n10045), .Z(n10047) );
  XOR U608 ( .A(a[1815]), .B(n10033), .Z(n10035) );
  XOR U609 ( .A(a[1818]), .B(n10021), .Z(n10023) );
  XOR U610 ( .A(a[1821]), .B(n10008), .Z(n10010) );
  XOR U611 ( .A(a[1824]), .B(n9996), .Z(n9998) );
  XOR U612 ( .A(a[1827]), .B(n9984), .Z(n9986) );
  XOR U613 ( .A(a[1830]), .B(n9971), .Z(n9973) );
  XOR U614 ( .A(a[1833]), .B(n9959), .Z(n9961) );
  XOR U615 ( .A(a[1836]), .B(n9947), .Z(n9949) );
  XOR U616 ( .A(a[1839]), .B(n9934), .Z(n9936) );
  XOR U617 ( .A(a[1842]), .B(n9922), .Z(n9924) );
  XOR U618 ( .A(a[1845]), .B(n9910), .Z(n9912) );
  XOR U619 ( .A(a[1848]), .B(n9898), .Z(n9900) );
  XOR U620 ( .A(a[1851]), .B(n9885), .Z(n9887) );
  XOR U621 ( .A(a[1854]), .B(n9873), .Z(n9875) );
  XOR U622 ( .A(a[1857]), .B(n9861), .Z(n9863) );
  XOR U623 ( .A(a[1860]), .B(n9848), .Z(n9850) );
  XOR U624 ( .A(a[1863]), .B(n9836), .Z(n9838) );
  XOR U625 ( .A(a[1866]), .B(n9824), .Z(n9826) );
  XOR U626 ( .A(a[1869]), .B(n9811), .Z(n9813) );
  XOR U627 ( .A(a[1872]), .B(n9799), .Z(n9801) );
  XOR U628 ( .A(a[1875]), .B(n9787), .Z(n9789) );
  XOR U629 ( .A(a[1878]), .B(n9775), .Z(n9777) );
  XOR U630 ( .A(a[1881]), .B(n9762), .Z(n9764) );
  XOR U631 ( .A(a[1884]), .B(n9750), .Z(n9752) );
  XOR U632 ( .A(a[1887]), .B(n9738), .Z(n9740) );
  XOR U633 ( .A(a[1890]), .B(n9725), .Z(n9727) );
  XOR U634 ( .A(a[1893]), .B(n9713), .Z(n9715) );
  XOR U635 ( .A(a[1896]), .B(n9701), .Z(n9703) );
  XOR U636 ( .A(a[1899]), .B(n9687), .Z(n9689) );
  XOR U637 ( .A(a[1902]), .B(n9675), .Z(n9677) );
  XOR U638 ( .A(a[1905]), .B(n9663), .Z(n9665) );
  XOR U639 ( .A(a[1908]), .B(n9651), .Z(n9653) );
  XOR U640 ( .A(a[1911]), .B(n9638), .Z(n9640) );
  XOR U641 ( .A(a[1914]), .B(n9626), .Z(n9628) );
  XOR U642 ( .A(a[1917]), .B(n9614), .Z(n9616) );
  XOR U643 ( .A(a[1920]), .B(n9601), .Z(n9603) );
  XOR U644 ( .A(a[1923]), .B(n9589), .Z(n9591) );
  XOR U645 ( .A(a[1926]), .B(n9577), .Z(n9579) );
  XOR U646 ( .A(a[1929]), .B(n9564), .Z(n9566) );
  XOR U647 ( .A(a[1932]), .B(n9552), .Z(n9554) );
  XOR U648 ( .A(a[1935]), .B(n9540), .Z(n9542) );
  XOR U649 ( .A(a[1938]), .B(n9528), .Z(n9530) );
  XOR U650 ( .A(a[1941]), .B(n9515), .Z(n9517) );
  XOR U651 ( .A(a[1944]), .B(n9503), .Z(n9505) );
  XOR U652 ( .A(a[1947]), .B(n9491), .Z(n9493) );
  XOR U653 ( .A(a[1950]), .B(n9478), .Z(n9480) );
  XOR U654 ( .A(a[1953]), .B(n9466), .Z(n9468) );
  XOR U655 ( .A(a[1956]), .B(n9454), .Z(n9456) );
  XOR U656 ( .A(a[1959]), .B(n9441), .Z(n9443) );
  XOR U657 ( .A(a[1962]), .B(n9429), .Z(n9431) );
  XOR U658 ( .A(a[1965]), .B(n9417), .Z(n9419) );
  XOR U659 ( .A(a[1968]), .B(n9405), .Z(n9407) );
  XOR U660 ( .A(a[1971]), .B(n9392), .Z(n9394) );
  XOR U661 ( .A(a[1974]), .B(n9380), .Z(n9382) );
  XOR U662 ( .A(a[1977]), .B(n9368), .Z(n9370) );
  XOR U663 ( .A(a[1980]), .B(n9355), .Z(n9357) );
  XOR U664 ( .A(a[1983]), .B(n9343), .Z(n9345) );
  XOR U665 ( .A(a[1986]), .B(n9331), .Z(n9333) );
  XOR U666 ( .A(a[1989]), .B(n9318), .Z(n9320) );
  XOR U667 ( .A(a[1992]), .B(n9306), .Z(n9308) );
  XOR U668 ( .A(a[1995]), .B(n9294), .Z(n9296) );
  XOR U669 ( .A(a[1998]), .B(n9282), .Z(n9284) );
  XOR U670 ( .A(a[2001]), .B(n9267), .Z(n9269) );
  XOR U671 ( .A(a[2004]), .B(n9255), .Z(n9257) );
  XOR U672 ( .A(a[2007]), .B(n9243), .Z(n9245) );
  XOR U673 ( .A(a[2010]), .B(n9230), .Z(n9232) );
  XOR U674 ( .A(a[2013]), .B(n9218), .Z(n9220) );
  XOR U675 ( .A(a[2016]), .B(n9206), .Z(n9208) );
  XOR U676 ( .A(a[2019]), .B(n9193), .Z(n9195) );
  XOR U677 ( .A(a[2022]), .B(n9181), .Z(n9183) );
  XOR U678 ( .A(a[2025]), .B(n9169), .Z(n9171) );
  XOR U679 ( .A(a[2028]), .B(n9157), .Z(n9159) );
  XOR U680 ( .A(a[2031]), .B(n9144), .Z(n9146) );
  XOR U681 ( .A(a[2034]), .B(n9132), .Z(n9134) );
  XOR U682 ( .A(a[2037]), .B(n9120), .Z(n9122) );
  XOR U683 ( .A(a[2040]), .B(n9107), .Z(n9109) );
  XOR U684 ( .A(a[2043]), .B(n9095), .Z(n9097) );
  XOR U685 ( .A(a[2046]), .B(n9083), .Z(n9085) );
  XOR U686 ( .A(a[2049]), .B(n9070), .Z(n9072) );
  XOR U687 ( .A(a[2052]), .B(n9058), .Z(n9060) );
  XOR U688 ( .A(a[2055]), .B(n9046), .Z(n9048) );
  XOR U689 ( .A(a[2058]), .B(n9034), .Z(n9036) );
  XOR U690 ( .A(a[2061]), .B(n9021), .Z(n9023) );
  XOR U691 ( .A(a[2064]), .B(n9009), .Z(n9011) );
  XOR U692 ( .A(a[2067]), .B(n8997), .Z(n8999) );
  XOR U693 ( .A(a[2070]), .B(n8984), .Z(n8986) );
  XOR U694 ( .A(a[2073]), .B(n8972), .Z(n8974) );
  XOR U695 ( .A(a[2076]), .B(n8960), .Z(n8962) );
  XOR U696 ( .A(a[2079]), .B(n8947), .Z(n8949) );
  XOR U697 ( .A(a[2082]), .B(n8935), .Z(n8937) );
  XOR U698 ( .A(a[2085]), .B(n8923), .Z(n8925) );
  XOR U699 ( .A(a[2088]), .B(n8911), .Z(n8913) );
  XOR U700 ( .A(a[2091]), .B(n8898), .Z(n8900) );
  XOR U701 ( .A(a[2094]), .B(n8886), .Z(n8888) );
  XOR U702 ( .A(a[2097]), .B(n8874), .Z(n8876) );
  XOR U703 ( .A(a[2100]), .B(n8860), .Z(n8862) );
  XOR U704 ( .A(a[2103]), .B(n8848), .Z(n8850) );
  XOR U705 ( .A(a[2106]), .B(n8836), .Z(n8838) );
  XOR U706 ( .A(a[2109]), .B(n8823), .Z(n8825) );
  XOR U707 ( .A(a[2112]), .B(n8811), .Z(n8813) );
  XOR U708 ( .A(a[2115]), .B(n8799), .Z(n8801) );
  XOR U709 ( .A(a[2118]), .B(n8787), .Z(n8789) );
  XOR U710 ( .A(a[2121]), .B(n8774), .Z(n8776) );
  XOR U711 ( .A(a[2124]), .B(n8762), .Z(n8764) );
  XOR U712 ( .A(a[2127]), .B(n8750), .Z(n8752) );
  XOR U713 ( .A(a[2130]), .B(n8737), .Z(n8739) );
  XOR U714 ( .A(a[2133]), .B(n8725), .Z(n8727) );
  XOR U715 ( .A(a[2136]), .B(n8713), .Z(n8715) );
  XOR U716 ( .A(a[2139]), .B(n8700), .Z(n8702) );
  XOR U717 ( .A(a[2142]), .B(n8688), .Z(n8690) );
  XOR U718 ( .A(a[2145]), .B(n8676), .Z(n8678) );
  XOR U719 ( .A(a[2148]), .B(n8664), .Z(n8666) );
  XOR U720 ( .A(a[2151]), .B(n8651), .Z(n8653) );
  XOR U721 ( .A(a[2154]), .B(n8639), .Z(n8641) );
  XOR U722 ( .A(a[2157]), .B(n8627), .Z(n8629) );
  XOR U723 ( .A(a[2160]), .B(n8614), .Z(n8616) );
  XOR U724 ( .A(a[2163]), .B(n8602), .Z(n8604) );
  XOR U725 ( .A(a[2166]), .B(n8590), .Z(n8592) );
  XOR U726 ( .A(a[2169]), .B(n8577), .Z(n8579) );
  XOR U727 ( .A(a[2172]), .B(n8565), .Z(n8567) );
  XOR U728 ( .A(a[2175]), .B(n8553), .Z(n8555) );
  XOR U729 ( .A(a[2178]), .B(n8541), .Z(n8543) );
  XOR U730 ( .A(a[2181]), .B(n8528), .Z(n8530) );
  XOR U731 ( .A(a[2184]), .B(n8516), .Z(n8518) );
  XOR U732 ( .A(a[2187]), .B(n8504), .Z(n8506) );
  XOR U733 ( .A(a[2190]), .B(n8491), .Z(n8493) );
  XOR U734 ( .A(a[2193]), .B(n8479), .Z(n8481) );
  XOR U735 ( .A(a[2196]), .B(n8467), .Z(n8469) );
  XOR U736 ( .A(a[2199]), .B(n8453), .Z(n8455) );
  XOR U737 ( .A(a[2202]), .B(n8441), .Z(n8443) );
  XOR U738 ( .A(a[2205]), .B(n8429), .Z(n8431) );
  XOR U739 ( .A(a[2208]), .B(n8417), .Z(n8419) );
  XOR U740 ( .A(a[2211]), .B(n8404), .Z(n8406) );
  XOR U741 ( .A(a[2214]), .B(n8392), .Z(n8394) );
  XOR U742 ( .A(a[2217]), .B(n8380), .Z(n8382) );
  XOR U743 ( .A(a[2220]), .B(n8367), .Z(n8369) );
  XOR U744 ( .A(a[2223]), .B(n8355), .Z(n8357) );
  XOR U745 ( .A(a[2226]), .B(n8343), .Z(n8345) );
  XOR U746 ( .A(a[2229]), .B(n8330), .Z(n8332) );
  XOR U747 ( .A(a[2232]), .B(n8318), .Z(n8320) );
  XOR U748 ( .A(a[2235]), .B(n8306), .Z(n8308) );
  XOR U749 ( .A(a[2238]), .B(n8294), .Z(n8296) );
  XOR U750 ( .A(a[2241]), .B(n8281), .Z(n8283) );
  XOR U751 ( .A(a[2244]), .B(n8269), .Z(n8271) );
  XOR U752 ( .A(a[2247]), .B(n8257), .Z(n8259) );
  XOR U753 ( .A(a[2250]), .B(n8244), .Z(n8246) );
  XOR U754 ( .A(a[2253]), .B(n8232), .Z(n8234) );
  XOR U755 ( .A(a[2256]), .B(n8220), .Z(n8222) );
  XOR U756 ( .A(a[2259]), .B(n8207), .Z(n8209) );
  XOR U757 ( .A(a[2262]), .B(n8195), .Z(n8197) );
  XOR U758 ( .A(a[2265]), .B(n8183), .Z(n8185) );
  XOR U759 ( .A(a[2268]), .B(n8171), .Z(n8173) );
  XOR U760 ( .A(a[2271]), .B(n8158), .Z(n8160) );
  XOR U761 ( .A(a[2274]), .B(n8146), .Z(n8148) );
  XOR U762 ( .A(a[2277]), .B(n8134), .Z(n8136) );
  XOR U763 ( .A(a[2280]), .B(n8121), .Z(n8123) );
  XOR U764 ( .A(a[2283]), .B(n8109), .Z(n8111) );
  XOR U765 ( .A(a[2286]), .B(n8097), .Z(n8099) );
  XOR U766 ( .A(a[2289]), .B(n8084), .Z(n8086) );
  XOR U767 ( .A(a[2292]), .B(n8072), .Z(n8074) );
  XOR U768 ( .A(a[2295]), .B(n8060), .Z(n8062) );
  XOR U769 ( .A(a[2298]), .B(n8048), .Z(n8050) );
  XOR U770 ( .A(a[2301]), .B(n8034), .Z(n8036) );
  XOR U771 ( .A(a[2304]), .B(n8022), .Z(n8024) );
  XOR U772 ( .A(a[2307]), .B(n8010), .Z(n8012) );
  XOR U773 ( .A(a[2310]), .B(n7997), .Z(n7999) );
  XOR U774 ( .A(a[2313]), .B(n7985), .Z(n7987) );
  XOR U775 ( .A(a[2316]), .B(n7973), .Z(n7975) );
  XOR U776 ( .A(a[2319]), .B(n7960), .Z(n7962) );
  XOR U777 ( .A(a[2322]), .B(n7948), .Z(n7950) );
  XOR U778 ( .A(a[2325]), .B(n7936), .Z(n7938) );
  XOR U779 ( .A(a[2328]), .B(n7924), .Z(n7926) );
  XOR U780 ( .A(a[2331]), .B(n7911), .Z(n7913) );
  XOR U781 ( .A(a[2334]), .B(n7899), .Z(n7901) );
  XOR U782 ( .A(a[2337]), .B(n7887), .Z(n7889) );
  XOR U783 ( .A(a[2340]), .B(n7874), .Z(n7876) );
  XOR U784 ( .A(a[2343]), .B(n7862), .Z(n7864) );
  XOR U785 ( .A(a[2346]), .B(n7850), .Z(n7852) );
  XOR U786 ( .A(a[2349]), .B(n7837), .Z(n7839) );
  XOR U787 ( .A(a[2352]), .B(n7825), .Z(n7827) );
  XOR U788 ( .A(a[2355]), .B(n7813), .Z(n7815) );
  XOR U789 ( .A(a[2358]), .B(n7801), .Z(n7803) );
  XOR U790 ( .A(a[2361]), .B(n7788), .Z(n7790) );
  XOR U791 ( .A(a[2364]), .B(n7776), .Z(n7778) );
  XOR U792 ( .A(a[2367]), .B(n7764), .Z(n7766) );
  XOR U793 ( .A(a[2370]), .B(n7751), .Z(n7753) );
  XOR U794 ( .A(a[2373]), .B(n7739), .Z(n7741) );
  XOR U795 ( .A(a[2376]), .B(n7727), .Z(n7729) );
  XOR U796 ( .A(a[2379]), .B(n7714), .Z(n7716) );
  XOR U797 ( .A(a[2382]), .B(n7702), .Z(n7704) );
  XOR U798 ( .A(a[2385]), .B(n7690), .Z(n7692) );
  XOR U799 ( .A(a[2388]), .B(n7678), .Z(n7680) );
  XOR U800 ( .A(a[2391]), .B(n7665), .Z(n7667) );
  XOR U801 ( .A(a[2394]), .B(n7653), .Z(n7655) );
  XOR U802 ( .A(a[2397]), .B(n7641), .Z(n7643) );
  XOR U803 ( .A(a[2400]), .B(n7627), .Z(n7629) );
  XOR U804 ( .A(a[2403]), .B(n7615), .Z(n7617) );
  XOR U805 ( .A(a[2406]), .B(n7603), .Z(n7605) );
  XOR U806 ( .A(a[2409]), .B(n7590), .Z(n7592) );
  XOR U807 ( .A(a[2412]), .B(n7578), .Z(n7580) );
  XOR U808 ( .A(a[2415]), .B(n7566), .Z(n7568) );
  XOR U809 ( .A(a[2418]), .B(n7554), .Z(n7556) );
  XOR U810 ( .A(a[2421]), .B(n7541), .Z(n7543) );
  XOR U811 ( .A(a[2424]), .B(n7529), .Z(n7531) );
  XOR U812 ( .A(a[2427]), .B(n7517), .Z(n7519) );
  XOR U813 ( .A(a[2430]), .B(n7504), .Z(n7506) );
  XOR U814 ( .A(a[2433]), .B(n7492), .Z(n7494) );
  XOR U815 ( .A(a[2436]), .B(n7480), .Z(n7482) );
  XOR U816 ( .A(a[2439]), .B(n7467), .Z(n7469) );
  XOR U817 ( .A(a[2442]), .B(n7455), .Z(n7457) );
  XOR U818 ( .A(a[2445]), .B(n7443), .Z(n7445) );
  XOR U819 ( .A(a[2448]), .B(n7431), .Z(n7433) );
  XOR U820 ( .A(a[2451]), .B(n7418), .Z(n7420) );
  XOR U821 ( .A(a[2454]), .B(n7406), .Z(n7408) );
  XOR U822 ( .A(a[2457]), .B(n7394), .Z(n7396) );
  XOR U823 ( .A(a[2460]), .B(n7381), .Z(n7383) );
  XOR U824 ( .A(a[2463]), .B(n7369), .Z(n7371) );
  XOR U825 ( .A(a[2466]), .B(n7357), .Z(n7359) );
  XOR U826 ( .A(a[2469]), .B(n7344), .Z(n7346) );
  XOR U827 ( .A(a[2472]), .B(n7332), .Z(n7334) );
  XOR U828 ( .A(a[2475]), .B(n7320), .Z(n7322) );
  XOR U829 ( .A(a[2478]), .B(n7308), .Z(n7310) );
  XOR U830 ( .A(a[2481]), .B(n7295), .Z(n7297) );
  XOR U831 ( .A(a[2484]), .B(n7283), .Z(n7285) );
  XOR U832 ( .A(a[2487]), .B(n7271), .Z(n7273) );
  XOR U833 ( .A(a[2490]), .B(n7258), .Z(n7260) );
  XOR U834 ( .A(a[2493]), .B(n7246), .Z(n7248) );
  XOR U835 ( .A(a[2496]), .B(n7234), .Z(n7236) );
  XOR U836 ( .A(a[2499]), .B(n7220), .Z(n7222) );
  XOR U837 ( .A(a[2502]), .B(n7208), .Z(n7210) );
  XOR U838 ( .A(a[2505]), .B(n7196), .Z(n7198) );
  XOR U839 ( .A(a[2508]), .B(n7184), .Z(n7186) );
  XOR U840 ( .A(a[2511]), .B(n7171), .Z(n7173) );
  XOR U841 ( .A(a[2514]), .B(n7159), .Z(n7161) );
  XOR U842 ( .A(a[2517]), .B(n7147), .Z(n7149) );
  XOR U843 ( .A(a[2520]), .B(n7134), .Z(n7136) );
  XOR U844 ( .A(a[2523]), .B(n7122), .Z(n7124) );
  XOR U845 ( .A(a[2526]), .B(n7110), .Z(n7112) );
  XOR U846 ( .A(a[2529]), .B(n7097), .Z(n7099) );
  XOR U847 ( .A(a[2532]), .B(n7085), .Z(n7087) );
  XOR U848 ( .A(a[2535]), .B(n7073), .Z(n7075) );
  XOR U849 ( .A(a[2538]), .B(n7061), .Z(n7063) );
  XOR U850 ( .A(a[2541]), .B(n7048), .Z(n7050) );
  XOR U851 ( .A(a[2544]), .B(n7036), .Z(n7038) );
  XOR U852 ( .A(a[2547]), .B(n7024), .Z(n7026) );
  XOR U853 ( .A(a[2550]), .B(n7011), .Z(n7013) );
  XOR U854 ( .A(a[2553]), .B(n6999), .Z(n7001) );
  XOR U855 ( .A(a[2556]), .B(n6987), .Z(n6989) );
  XOR U856 ( .A(a[2559]), .B(n6974), .Z(n6976) );
  XOR U857 ( .A(a[2562]), .B(n6962), .Z(n6964) );
  XOR U858 ( .A(a[2565]), .B(n6950), .Z(n6952) );
  XOR U859 ( .A(a[2568]), .B(n6938), .Z(n6940) );
  XOR U860 ( .A(a[2571]), .B(n6925), .Z(n6927) );
  XOR U861 ( .A(a[2574]), .B(n6913), .Z(n6915) );
  XOR U862 ( .A(a[2577]), .B(n6901), .Z(n6903) );
  XOR U863 ( .A(a[2580]), .B(n6888), .Z(n6890) );
  XOR U864 ( .A(a[2583]), .B(n6876), .Z(n6878) );
  XOR U865 ( .A(a[2586]), .B(n6864), .Z(n6866) );
  XOR U866 ( .A(a[2589]), .B(n6851), .Z(n6853) );
  XOR U867 ( .A(a[2592]), .B(n6839), .Z(n6841) );
  XOR U868 ( .A(a[2595]), .B(n6827), .Z(n6829) );
  XOR U869 ( .A(a[2598]), .B(n6815), .Z(n6817) );
  XOR U870 ( .A(a[2601]), .B(n6801), .Z(n6803) );
  XOR U871 ( .A(a[2604]), .B(n6789), .Z(n6791) );
  XOR U872 ( .A(a[2607]), .B(n6777), .Z(n6779) );
  XOR U873 ( .A(a[2610]), .B(n6764), .Z(n6766) );
  XOR U874 ( .A(a[2613]), .B(n6752), .Z(n6754) );
  XOR U875 ( .A(a[2616]), .B(n6740), .Z(n6742) );
  XOR U876 ( .A(a[2619]), .B(n6727), .Z(n6729) );
  XOR U877 ( .A(a[2622]), .B(n6715), .Z(n6717) );
  XOR U878 ( .A(a[2625]), .B(n6703), .Z(n6705) );
  XOR U879 ( .A(a[2628]), .B(n6691), .Z(n6693) );
  XOR U880 ( .A(a[2631]), .B(n6678), .Z(n6680) );
  XOR U881 ( .A(a[2634]), .B(n6666), .Z(n6668) );
  XOR U882 ( .A(a[2637]), .B(n6654), .Z(n6656) );
  XOR U883 ( .A(a[2640]), .B(n6641), .Z(n6643) );
  XOR U884 ( .A(a[2643]), .B(n6629), .Z(n6631) );
  XOR U885 ( .A(a[2646]), .B(n6617), .Z(n6619) );
  XOR U886 ( .A(a[2649]), .B(n6604), .Z(n6606) );
  XOR U887 ( .A(a[2652]), .B(n6592), .Z(n6594) );
  XOR U888 ( .A(a[2655]), .B(n6580), .Z(n6582) );
  XOR U889 ( .A(a[2658]), .B(n6568), .Z(n6570) );
  XOR U890 ( .A(a[2661]), .B(n6555), .Z(n6557) );
  XOR U891 ( .A(a[2664]), .B(n6543), .Z(n6545) );
  XOR U892 ( .A(a[2667]), .B(n6531), .Z(n6533) );
  XOR U893 ( .A(a[2670]), .B(n6518), .Z(n6520) );
  XOR U894 ( .A(a[2673]), .B(n6506), .Z(n6508) );
  XOR U895 ( .A(a[2676]), .B(n6494), .Z(n6496) );
  XOR U896 ( .A(a[2679]), .B(n6481), .Z(n6483) );
  XOR U897 ( .A(a[2682]), .B(n6469), .Z(n6471) );
  XOR U898 ( .A(a[2685]), .B(n6457), .Z(n6459) );
  XOR U899 ( .A(a[2688]), .B(n6445), .Z(n6447) );
  XOR U900 ( .A(a[2691]), .B(n6432), .Z(n6434) );
  XOR U901 ( .A(a[2694]), .B(n6420), .Z(n6422) );
  XOR U902 ( .A(a[2697]), .B(n6408), .Z(n6410) );
  XOR U903 ( .A(a[2700]), .B(n6394), .Z(n6396) );
  XOR U904 ( .A(a[2703]), .B(n6382), .Z(n6384) );
  XOR U905 ( .A(a[2706]), .B(n6370), .Z(n6372) );
  XOR U906 ( .A(a[2709]), .B(n6357), .Z(n6359) );
  XOR U907 ( .A(a[2712]), .B(n6345), .Z(n6347) );
  XOR U908 ( .A(a[2715]), .B(n6333), .Z(n6335) );
  XOR U909 ( .A(a[2718]), .B(n6321), .Z(n6323) );
  XOR U910 ( .A(a[2721]), .B(n6308), .Z(n6310) );
  XOR U911 ( .A(a[2724]), .B(n6296), .Z(n6298) );
  XOR U912 ( .A(a[2727]), .B(n6284), .Z(n6286) );
  XOR U913 ( .A(a[2730]), .B(n6271), .Z(n6273) );
  XOR U914 ( .A(a[2733]), .B(n6259), .Z(n6261) );
  XOR U915 ( .A(a[2736]), .B(n6247), .Z(n6249) );
  XOR U916 ( .A(a[2739]), .B(n6234), .Z(n6236) );
  XOR U917 ( .A(a[2742]), .B(n6222), .Z(n6224) );
  XOR U918 ( .A(a[2745]), .B(n6210), .Z(n6212) );
  XOR U919 ( .A(a[2748]), .B(n6198), .Z(n6200) );
  XOR U920 ( .A(a[2751]), .B(n6185), .Z(n6187) );
  XOR U921 ( .A(a[2754]), .B(n6173), .Z(n6175) );
  XOR U922 ( .A(a[2757]), .B(n6161), .Z(n6163) );
  XOR U923 ( .A(a[2760]), .B(n6148), .Z(n6150) );
  XOR U924 ( .A(a[2763]), .B(n6136), .Z(n6138) );
  XOR U925 ( .A(a[2766]), .B(n6124), .Z(n6126) );
  XOR U926 ( .A(a[2769]), .B(n6111), .Z(n6113) );
  XOR U927 ( .A(a[2772]), .B(n6099), .Z(n6101) );
  XOR U928 ( .A(a[2775]), .B(n6087), .Z(n6089) );
  XOR U929 ( .A(a[2778]), .B(n6075), .Z(n6077) );
  XOR U930 ( .A(a[2781]), .B(n6062), .Z(n6064) );
  XOR U931 ( .A(a[2784]), .B(n6050), .Z(n6052) );
  XOR U932 ( .A(a[2787]), .B(n6038), .Z(n6040) );
  XOR U933 ( .A(a[2790]), .B(n6025), .Z(n6027) );
  XOR U934 ( .A(a[2793]), .B(n6013), .Z(n6015) );
  XOR U935 ( .A(a[2796]), .B(n6001), .Z(n6003) );
  XOR U936 ( .A(a[2799]), .B(n5987), .Z(n5989) );
  XOR U937 ( .A(a[2802]), .B(n5975), .Z(n5977) );
  XOR U938 ( .A(a[2805]), .B(n5963), .Z(n5965) );
  XOR U939 ( .A(a[2808]), .B(n5951), .Z(n5953) );
  XOR U940 ( .A(a[2811]), .B(n5938), .Z(n5940) );
  XOR U941 ( .A(a[2814]), .B(n5926), .Z(n5928) );
  XOR U942 ( .A(a[2817]), .B(n5914), .Z(n5916) );
  XOR U943 ( .A(a[2820]), .B(n5901), .Z(n5903) );
  XOR U944 ( .A(a[2823]), .B(n5889), .Z(n5891) );
  XOR U945 ( .A(a[2826]), .B(n5877), .Z(n5879) );
  XOR U946 ( .A(a[2829]), .B(n5864), .Z(n5866) );
  XOR U947 ( .A(a[2832]), .B(n5852), .Z(n5854) );
  XOR U948 ( .A(a[2835]), .B(n5840), .Z(n5842) );
  XOR U949 ( .A(a[2838]), .B(n5828), .Z(n5830) );
  XOR U950 ( .A(a[2841]), .B(n5815), .Z(n5817) );
  XOR U951 ( .A(a[2844]), .B(n5803), .Z(n5805) );
  XOR U952 ( .A(a[2847]), .B(n5791), .Z(n5793) );
  XOR U953 ( .A(a[2850]), .B(n5778), .Z(n5780) );
  XOR U954 ( .A(a[2853]), .B(n5766), .Z(n5768) );
  XOR U955 ( .A(a[2856]), .B(n5754), .Z(n5756) );
  XOR U956 ( .A(a[2859]), .B(n5741), .Z(n5743) );
  XOR U957 ( .A(a[2862]), .B(n5729), .Z(n5731) );
  XOR U958 ( .A(a[2865]), .B(n5717), .Z(n5719) );
  XOR U959 ( .A(a[2868]), .B(n5705), .Z(n5707) );
  XOR U960 ( .A(a[2871]), .B(n5692), .Z(n5694) );
  XOR U961 ( .A(a[2874]), .B(n5680), .Z(n5682) );
  XOR U962 ( .A(a[2877]), .B(n5668), .Z(n5670) );
  XOR U963 ( .A(a[2880]), .B(n5655), .Z(n5657) );
  XOR U964 ( .A(a[2883]), .B(n5643), .Z(n5645) );
  XOR U965 ( .A(a[2886]), .B(n5631), .Z(n5633) );
  XOR U966 ( .A(a[2889]), .B(n5618), .Z(n5620) );
  XOR U967 ( .A(a[2892]), .B(n5606), .Z(n5608) );
  XOR U968 ( .A(a[2895]), .B(n5594), .Z(n5596) );
  XOR U969 ( .A(a[2898]), .B(n5582), .Z(n5584) );
  XOR U970 ( .A(a[2901]), .B(n5568), .Z(n5570) );
  XOR U971 ( .A(a[2904]), .B(n5556), .Z(n5558) );
  XOR U972 ( .A(a[2907]), .B(n5544), .Z(n5546) );
  XOR U973 ( .A(a[2910]), .B(n5531), .Z(n5533) );
  XOR U974 ( .A(a[2913]), .B(n5519), .Z(n5521) );
  XOR U975 ( .A(a[2916]), .B(n5507), .Z(n5509) );
  XOR U976 ( .A(a[2919]), .B(n5494), .Z(n5496) );
  XOR U977 ( .A(a[2922]), .B(n5482), .Z(n5484) );
  XOR U978 ( .A(a[2925]), .B(n5470), .Z(n5472) );
  XOR U979 ( .A(a[2928]), .B(n5458), .Z(n5460) );
  XOR U980 ( .A(a[2931]), .B(n5445), .Z(n5447) );
  XOR U981 ( .A(a[2934]), .B(n5433), .Z(n5435) );
  XOR U982 ( .A(a[2937]), .B(n5421), .Z(n5423) );
  XOR U983 ( .A(a[2940]), .B(n5408), .Z(n5410) );
  XOR U984 ( .A(a[2943]), .B(n5396), .Z(n5398) );
  XOR U985 ( .A(a[2946]), .B(n5384), .Z(n5386) );
  XOR U986 ( .A(a[2949]), .B(n5371), .Z(n5373) );
  XOR U987 ( .A(a[2952]), .B(n5359), .Z(n5361) );
  XOR U988 ( .A(a[2955]), .B(n5347), .Z(n5349) );
  XOR U989 ( .A(a[2958]), .B(n5335), .Z(n5337) );
  XOR U990 ( .A(a[2961]), .B(n5322), .Z(n5324) );
  XOR U991 ( .A(a[2964]), .B(n5310), .Z(n5312) );
  XOR U992 ( .A(a[2967]), .B(n5298), .Z(n5300) );
  XOR U993 ( .A(a[2970]), .B(n5285), .Z(n5287) );
  XOR U994 ( .A(a[2973]), .B(n5273), .Z(n5275) );
  XOR U995 ( .A(a[2976]), .B(n5261), .Z(n5263) );
  XOR U996 ( .A(a[2979]), .B(n5248), .Z(n5250) );
  XOR U997 ( .A(a[2982]), .B(n5236), .Z(n5238) );
  XOR U998 ( .A(a[2985]), .B(n5224), .Z(n5226) );
  XOR U999 ( .A(a[2988]), .B(n5212), .Z(n5214) );
  XOR U1000 ( .A(a[2991]), .B(n5199), .Z(n5201) );
  XOR U1001 ( .A(a[2994]), .B(n5187), .Z(n5189) );
  XOR U1002 ( .A(a[2997]), .B(n5175), .Z(n5177) );
  XOR U1003 ( .A(a[3000]), .B(n5160), .Z(n5162) );
  XOR U1004 ( .A(a[3003]), .B(n5148), .Z(n5150) );
  XOR U1005 ( .A(a[3006]), .B(n5136), .Z(n5138) );
  XOR U1006 ( .A(a[3009]), .B(n5123), .Z(n5125) );
  XOR U1007 ( .A(a[3012]), .B(n5111), .Z(n5113) );
  XOR U1008 ( .A(a[3015]), .B(n5099), .Z(n5101) );
  XOR U1009 ( .A(a[3018]), .B(n5087), .Z(n5089) );
  XOR U1010 ( .A(a[3021]), .B(n5074), .Z(n5076) );
  XOR U1011 ( .A(a[3024]), .B(n5062), .Z(n5064) );
  XOR U1012 ( .A(a[3027]), .B(n5050), .Z(n5052) );
  XOR U1013 ( .A(a[3030]), .B(n5037), .Z(n5039) );
  XOR U1014 ( .A(a[3033]), .B(n5025), .Z(n5027) );
  XOR U1015 ( .A(a[3036]), .B(n5013), .Z(n5015) );
  XOR U1016 ( .A(a[3039]), .B(n5000), .Z(n5002) );
  XOR U1017 ( .A(a[3042]), .B(n4988), .Z(n4990) );
  XOR U1018 ( .A(a[3045]), .B(n4976), .Z(n4978) );
  XOR U1019 ( .A(a[3048]), .B(n4964), .Z(n4966) );
  XOR U1020 ( .A(a[3051]), .B(n4951), .Z(n4953) );
  XOR U1021 ( .A(a[3054]), .B(n4939), .Z(n4941) );
  XOR U1022 ( .A(a[3057]), .B(n4927), .Z(n4929) );
  XOR U1023 ( .A(a[3060]), .B(n4914), .Z(n4916) );
  XOR U1024 ( .A(a[3063]), .B(n4902), .Z(n4904) );
  XOR U1025 ( .A(a[3066]), .B(n4890), .Z(n4892) );
  XOR U1026 ( .A(a[3069]), .B(n4877), .Z(n4879) );
  XOR U1027 ( .A(a[3072]), .B(n4865), .Z(n4867) );
  XOR U1028 ( .A(a[3075]), .B(n4853), .Z(n4855) );
  XOR U1029 ( .A(a[3078]), .B(n4841), .Z(n4843) );
  XOR U1030 ( .A(a[3081]), .B(n4828), .Z(n4830) );
  XOR U1031 ( .A(a[3084]), .B(n4816), .Z(n4818) );
  XOR U1032 ( .A(a[3087]), .B(n4804), .Z(n4806) );
  XOR U1033 ( .A(a[3090]), .B(n4791), .Z(n4793) );
  XOR U1034 ( .A(a[3093]), .B(n4779), .Z(n4781) );
  XOR U1035 ( .A(a[3096]), .B(n4767), .Z(n4769) );
  XOR U1036 ( .A(a[3099]), .B(n4753), .Z(n4755) );
  XOR U1037 ( .A(a[3102]), .B(n4741), .Z(n4743) );
  XOR U1038 ( .A(a[3105]), .B(n4729), .Z(n4731) );
  XOR U1039 ( .A(a[3108]), .B(n4717), .Z(n4719) );
  XOR U1040 ( .A(a[3111]), .B(n4704), .Z(n4706) );
  XOR U1041 ( .A(a[3114]), .B(n4692), .Z(n4694) );
  XOR U1042 ( .A(a[3117]), .B(n4680), .Z(n4682) );
  XOR U1043 ( .A(a[3120]), .B(n4667), .Z(n4669) );
  XOR U1044 ( .A(a[3123]), .B(n4655), .Z(n4657) );
  XOR U1045 ( .A(a[3126]), .B(n4643), .Z(n4645) );
  XOR U1046 ( .A(a[3129]), .B(n4630), .Z(n4632) );
  XOR U1047 ( .A(a[3132]), .B(n4618), .Z(n4620) );
  XOR U1048 ( .A(a[3135]), .B(n4606), .Z(n4608) );
  XOR U1049 ( .A(a[3138]), .B(n4594), .Z(n4596) );
  XOR U1050 ( .A(a[3141]), .B(n4581), .Z(n4583) );
  XOR U1051 ( .A(a[3144]), .B(n4569), .Z(n4571) );
  XOR U1052 ( .A(a[3147]), .B(n4557), .Z(n4559) );
  XOR U1053 ( .A(a[3150]), .B(n4544), .Z(n4546) );
  XOR U1054 ( .A(a[3153]), .B(n4532), .Z(n4534) );
  XOR U1055 ( .A(a[3156]), .B(n4520), .Z(n4522) );
  XOR U1056 ( .A(a[3159]), .B(n4507), .Z(n4509) );
  XOR U1057 ( .A(a[3162]), .B(n4495), .Z(n4497) );
  XOR U1058 ( .A(a[3165]), .B(n4483), .Z(n4485) );
  XOR U1059 ( .A(a[3168]), .B(n4471), .Z(n4473) );
  XOR U1060 ( .A(a[3171]), .B(n4458), .Z(n4460) );
  XOR U1061 ( .A(a[3174]), .B(n4446), .Z(n4448) );
  XOR U1062 ( .A(a[3177]), .B(n4434), .Z(n4436) );
  XOR U1063 ( .A(a[3180]), .B(n4421), .Z(n4423) );
  XOR U1064 ( .A(a[3183]), .B(n4409), .Z(n4411) );
  XOR U1065 ( .A(a[3186]), .B(n4397), .Z(n4399) );
  XOR U1066 ( .A(a[3189]), .B(n4384), .Z(n4386) );
  XOR U1067 ( .A(a[3192]), .B(n4372), .Z(n4374) );
  XOR U1068 ( .A(a[3195]), .B(n4360), .Z(n4362) );
  XOR U1069 ( .A(a[3198]), .B(n4348), .Z(n4350) );
  XOR U1070 ( .A(a[3201]), .B(n4334), .Z(n4336) );
  XOR U1071 ( .A(a[3204]), .B(n4322), .Z(n4324) );
  XOR U1072 ( .A(a[3207]), .B(n4310), .Z(n4312) );
  XOR U1073 ( .A(a[3210]), .B(n4297), .Z(n4299) );
  XOR U1074 ( .A(a[3213]), .B(n4285), .Z(n4287) );
  XOR U1075 ( .A(a[3216]), .B(n4273), .Z(n4275) );
  XOR U1076 ( .A(a[3219]), .B(n4260), .Z(n4262) );
  XOR U1077 ( .A(a[3222]), .B(n4248), .Z(n4250) );
  XOR U1078 ( .A(a[3225]), .B(n4236), .Z(n4238) );
  XOR U1079 ( .A(a[3228]), .B(n4224), .Z(n4226) );
  XOR U1080 ( .A(a[3231]), .B(n4211), .Z(n4213) );
  XOR U1081 ( .A(a[3234]), .B(n4199), .Z(n4201) );
  XOR U1082 ( .A(a[3237]), .B(n4187), .Z(n4189) );
  XOR U1083 ( .A(a[3240]), .B(n4174), .Z(n4176) );
  XOR U1084 ( .A(a[3243]), .B(n4162), .Z(n4164) );
  XOR U1085 ( .A(a[3246]), .B(n4150), .Z(n4152) );
  XOR U1086 ( .A(a[3249]), .B(n4137), .Z(n4139) );
  XOR U1087 ( .A(a[3252]), .B(n4125), .Z(n4127) );
  XOR U1088 ( .A(a[3255]), .B(n4113), .Z(n4115) );
  XOR U1089 ( .A(a[3258]), .B(n4101), .Z(n4103) );
  XOR U1090 ( .A(a[3261]), .B(n4088), .Z(n4090) );
  XOR U1091 ( .A(a[3264]), .B(n4076), .Z(n4078) );
  XOR U1092 ( .A(a[3267]), .B(n4064), .Z(n4066) );
  XOR U1093 ( .A(a[3270]), .B(n4051), .Z(n4053) );
  XOR U1094 ( .A(a[3273]), .B(n4039), .Z(n4041) );
  XOR U1095 ( .A(a[3276]), .B(n4027), .Z(n4029) );
  XOR U1096 ( .A(a[3279]), .B(n4014), .Z(n4016) );
  XOR U1097 ( .A(a[3282]), .B(n4002), .Z(n4004) );
  XOR U1098 ( .A(a[3285]), .B(n3990), .Z(n3992) );
  XOR U1099 ( .A(a[3288]), .B(n3978), .Z(n3980) );
  XOR U1100 ( .A(a[3291]), .B(n3965), .Z(n3967) );
  XOR U1101 ( .A(a[3294]), .B(n3953), .Z(n3955) );
  XOR U1102 ( .A(a[3297]), .B(n3941), .Z(n3943) );
  XOR U1103 ( .A(a[3300]), .B(n3927), .Z(n3929) );
  XOR U1104 ( .A(a[3303]), .B(n3915), .Z(n3917) );
  XOR U1105 ( .A(a[3306]), .B(n3903), .Z(n3905) );
  XOR U1106 ( .A(a[3309]), .B(n3890), .Z(n3892) );
  XOR U1107 ( .A(a[3312]), .B(n3878), .Z(n3880) );
  XOR U1108 ( .A(a[3315]), .B(n3866), .Z(n3868) );
  XOR U1109 ( .A(a[3318]), .B(n3854), .Z(n3856) );
  XOR U1110 ( .A(a[3321]), .B(n3841), .Z(n3843) );
  XOR U1111 ( .A(a[3324]), .B(n3829), .Z(n3831) );
  XOR U1112 ( .A(a[3327]), .B(n3817), .Z(n3819) );
  XOR U1113 ( .A(a[3330]), .B(n3804), .Z(n3806) );
  XOR U1114 ( .A(a[3333]), .B(n3792), .Z(n3794) );
  XOR U1115 ( .A(a[3336]), .B(n3780), .Z(n3782) );
  XOR U1116 ( .A(a[3339]), .B(n3767), .Z(n3769) );
  XOR U1117 ( .A(a[3342]), .B(n3755), .Z(n3757) );
  XOR U1118 ( .A(a[3345]), .B(n3743), .Z(n3745) );
  XOR U1119 ( .A(a[3348]), .B(n3731), .Z(n3733) );
  XOR U1120 ( .A(a[3351]), .B(n3718), .Z(n3720) );
  XOR U1121 ( .A(a[3354]), .B(n3706), .Z(n3708) );
  XOR U1122 ( .A(a[3357]), .B(n3694), .Z(n3696) );
  XOR U1123 ( .A(a[3360]), .B(n3681), .Z(n3683) );
  XOR U1124 ( .A(a[3363]), .B(n3669), .Z(n3671) );
  XOR U1125 ( .A(a[3366]), .B(n3657), .Z(n3659) );
  XOR U1126 ( .A(a[3369]), .B(n3644), .Z(n3646) );
  XOR U1127 ( .A(a[3372]), .B(n3632), .Z(n3634) );
  XOR U1128 ( .A(a[3375]), .B(n3620), .Z(n3622) );
  XOR U1129 ( .A(a[3378]), .B(n3608), .Z(n3610) );
  XOR U1130 ( .A(a[3381]), .B(n3595), .Z(n3597) );
  XOR U1131 ( .A(a[3384]), .B(n3583), .Z(n3585) );
  XOR U1132 ( .A(a[3387]), .B(n3571), .Z(n3573) );
  XOR U1133 ( .A(a[3390]), .B(n3558), .Z(n3560) );
  XOR U1134 ( .A(a[3393]), .B(n3546), .Z(n3548) );
  XOR U1135 ( .A(a[3396]), .B(n3534), .Z(n3536) );
  XOR U1136 ( .A(a[3399]), .B(n3520), .Z(n3522) );
  XOR U1137 ( .A(a[3402]), .B(n3508), .Z(n3510) );
  XOR U1138 ( .A(a[3405]), .B(n3496), .Z(n3498) );
  XOR U1139 ( .A(a[3408]), .B(n3484), .Z(n3486) );
  XOR U1140 ( .A(a[3411]), .B(n3471), .Z(n3473) );
  XOR U1141 ( .A(a[3414]), .B(n3459), .Z(n3461) );
  XOR U1142 ( .A(a[3417]), .B(n3447), .Z(n3449) );
  XOR U1143 ( .A(a[3420]), .B(n3434), .Z(n3436) );
  XOR U1144 ( .A(a[3423]), .B(n3422), .Z(n3424) );
  XOR U1145 ( .A(a[3426]), .B(n3410), .Z(n3412) );
  XOR U1146 ( .A(a[3429]), .B(n3397), .Z(n3399) );
  XOR U1147 ( .A(a[3432]), .B(n3385), .Z(n3387) );
  XOR U1148 ( .A(a[3435]), .B(n3373), .Z(n3375) );
  XOR U1149 ( .A(a[3438]), .B(n3361), .Z(n3363) );
  XOR U1150 ( .A(a[3441]), .B(n3348), .Z(n3350) );
  XOR U1151 ( .A(a[3444]), .B(n3336), .Z(n3338) );
  XOR U1152 ( .A(a[3447]), .B(n3324), .Z(n3326) );
  XOR U1153 ( .A(a[3450]), .B(n3311), .Z(n3313) );
  XOR U1154 ( .A(a[3453]), .B(n3299), .Z(n3301) );
  XOR U1155 ( .A(a[3456]), .B(n3287), .Z(n3289) );
  XOR U1156 ( .A(a[3459]), .B(n3274), .Z(n3276) );
  XOR U1157 ( .A(a[3462]), .B(n3262), .Z(n3264) );
  XOR U1158 ( .A(a[3465]), .B(n3250), .Z(n3252) );
  XOR U1159 ( .A(a[3468]), .B(n3238), .Z(n3240) );
  XOR U1160 ( .A(a[3471]), .B(n3225), .Z(n3227) );
  XOR U1161 ( .A(a[3474]), .B(n3213), .Z(n3215) );
  XOR U1162 ( .A(a[3477]), .B(n3201), .Z(n3203) );
  XOR U1163 ( .A(a[3480]), .B(n3188), .Z(n3190) );
  XOR U1164 ( .A(a[3483]), .B(n3176), .Z(n3178) );
  XOR U1165 ( .A(a[3486]), .B(n3164), .Z(n3166) );
  XOR U1166 ( .A(a[3489]), .B(n3151), .Z(n3153) );
  XOR U1167 ( .A(a[3492]), .B(n3139), .Z(n3141) );
  XOR U1168 ( .A(a[3495]), .B(n3127), .Z(n3129) );
  XOR U1169 ( .A(a[3498]), .B(n3115), .Z(n3117) );
  XOR U1170 ( .A(a[3501]), .B(n3101), .Z(n3103) );
  XOR U1171 ( .A(a[3504]), .B(n3089), .Z(n3091) );
  XOR U1172 ( .A(a[3507]), .B(n3077), .Z(n3079) );
  XOR U1173 ( .A(a[3510]), .B(n3064), .Z(n3066) );
  XOR U1174 ( .A(a[3513]), .B(n3052), .Z(n3054) );
  XOR U1175 ( .A(a[3516]), .B(n3040), .Z(n3042) );
  XOR U1176 ( .A(a[3519]), .B(n3027), .Z(n3029) );
  XOR U1177 ( .A(a[3522]), .B(n3015), .Z(n3017) );
  XOR U1178 ( .A(a[3525]), .B(n3003), .Z(n3005) );
  XOR U1179 ( .A(a[3528]), .B(n2991), .Z(n2993) );
  XOR U1180 ( .A(a[3531]), .B(n2978), .Z(n2980) );
  XOR U1181 ( .A(a[3534]), .B(n2966), .Z(n2968) );
  XOR U1182 ( .A(a[3537]), .B(n2954), .Z(n2956) );
  XOR U1183 ( .A(a[3540]), .B(n2941), .Z(n2943) );
  XOR U1184 ( .A(a[3543]), .B(n2929), .Z(n2931) );
  XOR U1185 ( .A(a[3546]), .B(n2917), .Z(n2919) );
  XOR U1186 ( .A(a[3549]), .B(n2904), .Z(n2906) );
  XOR U1187 ( .A(a[3552]), .B(n2892), .Z(n2894) );
  XOR U1188 ( .A(a[3555]), .B(n2880), .Z(n2882) );
  XOR U1189 ( .A(a[3558]), .B(n2868), .Z(n2870) );
  XOR U1190 ( .A(a[3561]), .B(n2855), .Z(n2857) );
  XOR U1191 ( .A(a[3564]), .B(n2843), .Z(n2845) );
  XOR U1192 ( .A(a[3567]), .B(n2831), .Z(n2833) );
  XOR U1193 ( .A(a[3570]), .B(n2818), .Z(n2820) );
  XOR U1194 ( .A(a[3573]), .B(n2806), .Z(n2808) );
  XOR U1195 ( .A(a[3576]), .B(n2794), .Z(n2796) );
  XOR U1196 ( .A(a[3579]), .B(n2781), .Z(n2783) );
  XOR U1197 ( .A(a[3582]), .B(n2769), .Z(n2771) );
  XOR U1198 ( .A(a[3585]), .B(n2757), .Z(n2759) );
  XOR U1199 ( .A(a[3588]), .B(n2745), .Z(n2747) );
  XOR U1200 ( .A(a[3591]), .B(n2732), .Z(n2734) );
  XOR U1201 ( .A(a[3594]), .B(n2720), .Z(n2722) );
  XOR U1202 ( .A(a[3597]), .B(n2708), .Z(n2710) );
  XOR U1203 ( .A(a[3600]), .B(n2694), .Z(n2696) );
  XOR U1204 ( .A(a[3603]), .B(n2682), .Z(n2684) );
  XOR U1205 ( .A(a[3606]), .B(n2670), .Z(n2672) );
  XOR U1206 ( .A(a[3609]), .B(n2657), .Z(n2659) );
  XOR U1207 ( .A(a[3612]), .B(n2645), .Z(n2647) );
  XOR U1208 ( .A(a[3615]), .B(n2633), .Z(n2635) );
  XOR U1209 ( .A(a[3618]), .B(n2621), .Z(n2623) );
  XOR U1210 ( .A(a[3621]), .B(n2608), .Z(n2610) );
  XOR U1211 ( .A(a[3624]), .B(n2596), .Z(n2598) );
  XOR U1212 ( .A(a[3627]), .B(n2584), .Z(n2586) );
  XOR U1213 ( .A(a[3630]), .B(n2571), .Z(n2573) );
  XOR U1214 ( .A(a[3633]), .B(n2559), .Z(n2561) );
  XOR U1215 ( .A(a[3636]), .B(n2547), .Z(n2549) );
  XOR U1216 ( .A(a[3639]), .B(n2534), .Z(n2536) );
  XOR U1217 ( .A(a[3642]), .B(n2522), .Z(n2524) );
  XOR U1218 ( .A(a[3645]), .B(n2510), .Z(n2512) );
  XOR U1219 ( .A(a[3648]), .B(n2498), .Z(n2500) );
  XOR U1220 ( .A(a[3651]), .B(n2485), .Z(n2487) );
  XOR U1221 ( .A(a[3654]), .B(n2473), .Z(n2475) );
  XOR U1222 ( .A(a[3657]), .B(n2461), .Z(n2463) );
  XOR U1223 ( .A(a[3660]), .B(n2448), .Z(n2450) );
  XOR U1224 ( .A(a[3663]), .B(n2436), .Z(n2438) );
  XOR U1225 ( .A(a[3666]), .B(n2424), .Z(n2426) );
  XOR U1226 ( .A(a[3669]), .B(n2411), .Z(n2413) );
  XOR U1227 ( .A(a[3672]), .B(n2399), .Z(n2401) );
  XOR U1228 ( .A(a[3675]), .B(n2387), .Z(n2389) );
  XOR U1229 ( .A(a[3678]), .B(n2375), .Z(n2377) );
  XOR U1230 ( .A(a[3681]), .B(n2362), .Z(n2364) );
  XOR U1231 ( .A(a[3684]), .B(n2350), .Z(n2352) );
  XOR U1232 ( .A(a[3687]), .B(n2338), .Z(n2340) );
  XOR U1233 ( .A(a[3690]), .B(n2325), .Z(n2327) );
  XOR U1234 ( .A(a[3693]), .B(n2313), .Z(n2315) );
  XOR U1235 ( .A(a[3696]), .B(n2301), .Z(n2303) );
  XOR U1236 ( .A(a[3699]), .B(n2287), .Z(n2289) );
  XOR U1237 ( .A(a[3702]), .B(n2275), .Z(n2277) );
  XOR U1238 ( .A(a[3705]), .B(n2263), .Z(n2265) );
  XOR U1239 ( .A(a[3708]), .B(n2251), .Z(n2253) );
  XOR U1240 ( .A(a[3711]), .B(n2238), .Z(n2240) );
  XOR U1241 ( .A(a[3714]), .B(n2226), .Z(n2228) );
  XOR U1242 ( .A(a[3717]), .B(n2214), .Z(n2216) );
  XOR U1243 ( .A(a[3720]), .B(n2201), .Z(n2203) );
  XOR U1244 ( .A(a[3723]), .B(n2189), .Z(n2191) );
  XOR U1245 ( .A(a[3726]), .B(n2177), .Z(n2179) );
  XOR U1246 ( .A(a[3729]), .B(n2164), .Z(n2166) );
  XOR U1247 ( .A(a[3732]), .B(n2152), .Z(n2154) );
  XOR U1248 ( .A(a[3735]), .B(n2140), .Z(n2142) );
  XOR U1249 ( .A(a[3738]), .B(n2128), .Z(n2130) );
  XOR U1250 ( .A(a[3741]), .B(n2115), .Z(n2117) );
  XOR U1251 ( .A(a[3744]), .B(n2103), .Z(n2105) );
  XOR U1252 ( .A(a[3747]), .B(n2091), .Z(n2093) );
  XOR U1253 ( .A(a[3750]), .B(n2078), .Z(n2080) );
  XOR U1254 ( .A(a[3753]), .B(n2066), .Z(n2068) );
  XOR U1255 ( .A(a[3756]), .B(n2054), .Z(n2056) );
  XOR U1256 ( .A(a[3759]), .B(n2041), .Z(n2043) );
  XOR U1257 ( .A(a[3762]), .B(n2029), .Z(n2031) );
  XOR U1258 ( .A(a[3765]), .B(n2017), .Z(n2019) );
  XOR U1259 ( .A(a[3768]), .B(n2005), .Z(n2007) );
  XOR U1260 ( .A(a[3771]), .B(n1992), .Z(n1994) );
  XOR U1261 ( .A(a[3774]), .B(n1980), .Z(n1982) );
  XOR U1262 ( .A(a[3777]), .B(n1968), .Z(n1970) );
  XOR U1263 ( .A(a[3780]), .B(n1955), .Z(n1957) );
  XOR U1264 ( .A(a[3783]), .B(n1943), .Z(n1945) );
  XOR U1265 ( .A(a[3786]), .B(n1931), .Z(n1933) );
  XOR U1266 ( .A(a[3789]), .B(n1918), .Z(n1920) );
  XOR U1267 ( .A(a[3792]), .B(n1906), .Z(n1908) );
  XOR U1268 ( .A(a[3795]), .B(n1894), .Z(n1896) );
  XOR U1269 ( .A(a[3798]), .B(n1882), .Z(n1884) );
  XOR U1270 ( .A(a[3801]), .B(n1868), .Z(n1870) );
  XOR U1271 ( .A(a[3804]), .B(n1856), .Z(n1858) );
  XOR U1272 ( .A(a[3807]), .B(n1844), .Z(n1846) );
  XOR U1273 ( .A(a[3810]), .B(n1831), .Z(n1833) );
  XOR U1274 ( .A(a[3813]), .B(n1819), .Z(n1821) );
  XOR U1275 ( .A(a[3816]), .B(n1807), .Z(n1809) );
  XOR U1276 ( .A(a[3819]), .B(n1794), .Z(n1796) );
  XOR U1277 ( .A(a[3822]), .B(n1782), .Z(n1784) );
  XOR U1278 ( .A(a[3825]), .B(n1770), .Z(n1772) );
  XOR U1279 ( .A(a[3828]), .B(n1758), .Z(n1760) );
  XOR U1280 ( .A(a[3831]), .B(n1745), .Z(n1747) );
  XOR U1281 ( .A(a[3834]), .B(n1733), .Z(n1735) );
  XOR U1282 ( .A(a[3837]), .B(n1721), .Z(n1723) );
  XOR U1283 ( .A(a[3840]), .B(n1708), .Z(n1710) );
  XOR U1284 ( .A(a[3843]), .B(n1696), .Z(n1698) );
  XOR U1285 ( .A(a[3846]), .B(n1684), .Z(n1686) );
  XOR U1286 ( .A(a[3849]), .B(n1671), .Z(n1673) );
  XOR U1287 ( .A(a[3852]), .B(n1659), .Z(n1661) );
  XOR U1288 ( .A(a[3855]), .B(n1647), .Z(n1649) );
  XOR U1289 ( .A(a[3858]), .B(n1635), .Z(n1637) );
  XOR U1290 ( .A(a[3861]), .B(n1622), .Z(n1624) );
  XOR U1291 ( .A(a[3864]), .B(n1610), .Z(n1612) );
  XOR U1292 ( .A(a[3867]), .B(n1598), .Z(n1600) );
  XOR U1293 ( .A(a[3870]), .B(n1585), .Z(n1587) );
  XOR U1294 ( .A(a[3873]), .B(n1573), .Z(n1575) );
  XOR U1295 ( .A(a[3876]), .B(n1561), .Z(n1563) );
  XOR U1296 ( .A(a[3879]), .B(n1548), .Z(n1550) );
  XOR U1297 ( .A(a[3882]), .B(n1536), .Z(n1538) );
  XOR U1298 ( .A(a[3885]), .B(n1524), .Z(n1526) );
  XOR U1299 ( .A(a[3888]), .B(n1512), .Z(n1514) );
  XOR U1300 ( .A(a[3891]), .B(n1499), .Z(n1501) );
  XOR U1301 ( .A(a[3894]), .B(n1487), .Z(n1489) );
  XOR U1302 ( .A(a[3897]), .B(n1475), .Z(n1477) );
  XOR U1303 ( .A(a[3900]), .B(n1461), .Z(n1463) );
  XOR U1304 ( .A(a[3903]), .B(n1449), .Z(n1451) );
  XOR U1305 ( .A(a[3906]), .B(n1437), .Z(n1439) );
  XOR U1306 ( .A(a[3909]), .B(n1424), .Z(n1426) );
  XOR U1307 ( .A(a[3912]), .B(n1412), .Z(n1414) );
  XOR U1308 ( .A(a[3915]), .B(n1400), .Z(n1402) );
  XOR U1309 ( .A(a[3918]), .B(n1388), .Z(n1390) );
  XOR U1310 ( .A(a[3921]), .B(n1375), .Z(n1377) );
  XOR U1311 ( .A(a[3924]), .B(n1363), .Z(n1365) );
  XOR U1312 ( .A(a[3927]), .B(n1351), .Z(n1353) );
  XOR U1313 ( .A(a[3930]), .B(n1338), .Z(n1340) );
  XOR U1314 ( .A(a[3933]), .B(n1326), .Z(n1328) );
  XOR U1315 ( .A(a[3936]), .B(n1314), .Z(n1316) );
  XOR U1316 ( .A(a[3939]), .B(n1301), .Z(n1303) );
  XOR U1317 ( .A(a[3942]), .B(n1289), .Z(n1291) );
  XOR U1318 ( .A(a[3945]), .B(n1277), .Z(n1279) );
  XOR U1319 ( .A(a[3948]), .B(n1265), .Z(n1267) );
  XOR U1320 ( .A(a[3951]), .B(n1252), .Z(n1254) );
  XOR U1321 ( .A(a[3954]), .B(n1240), .Z(n1242) );
  XOR U1322 ( .A(a[3957]), .B(n1228), .Z(n1230) );
  XOR U1323 ( .A(a[3960]), .B(n1215), .Z(n1217) );
  XOR U1324 ( .A(a[3963]), .B(n1203), .Z(n1205) );
  XOR U1325 ( .A(a[3966]), .B(n1191), .Z(n1193) );
  XOR U1326 ( .A(a[3969]), .B(n1178), .Z(n1180) );
  XOR U1327 ( .A(a[3972]), .B(n1166), .Z(n1168) );
  XOR U1328 ( .A(a[3975]), .B(n1154), .Z(n1156) );
  XOR U1329 ( .A(a[3978]), .B(n1142), .Z(n1144) );
  XOR U1330 ( .A(a[3981]), .B(n1129), .Z(n1131) );
  XOR U1331 ( .A(a[3984]), .B(n1117), .Z(n1119) );
  XOR U1332 ( .A(a[3987]), .B(n1105), .Z(n1107) );
  XOR U1333 ( .A(a[3990]), .B(n1092), .Z(n1094) );
  XOR U1334 ( .A(a[3993]), .B(n1080), .Z(n1082) );
  XOR U1335 ( .A(a[3996]), .B(n1068), .Z(n1070) );
  XOR U1336 ( .A(a[3999]), .B(n1053), .Z(n1055) );
  XOR U1337 ( .A(a[4002]), .B(n1041), .Z(n1043) );
  XOR U1338 ( .A(a[4005]), .B(n1029), .Z(n1031) );
  XOR U1339 ( .A(a[4008]), .B(n1017), .Z(n1019) );
  XOR U1340 ( .A(a[4011]), .B(n1004), .Z(n1006) );
  XOR U1341 ( .A(a[4014]), .B(n992), .Z(n994) );
  XOR U1342 ( .A(a[4017]), .B(n980), .Z(n982) );
  XOR U1343 ( .A(a[4020]), .B(n967), .Z(n969) );
  XOR U1344 ( .A(a[4023]), .B(n955), .Z(n957) );
  XOR U1345 ( .A(a[4026]), .B(n943), .Z(n945) );
  XOR U1346 ( .A(a[4029]), .B(n930), .Z(n932) );
  XOR U1347 ( .A(a[4032]), .B(n918), .Z(n920) );
  XOR U1348 ( .A(a[4035]), .B(n906), .Z(n908) );
  XOR U1349 ( .A(a[4038]), .B(n894), .Z(n896) );
  XOR U1350 ( .A(a[4041]), .B(n881), .Z(n883) );
  XOR U1351 ( .A(a[4044]), .B(n869), .Z(n871) );
  XOR U1352 ( .A(a[4047]), .B(n857), .Z(n859) );
  XOR U1353 ( .A(a[4050]), .B(n844), .Z(n846) );
  XOR U1354 ( .A(a[4053]), .B(n832), .Z(n834) );
  XOR U1355 ( .A(a[4056]), .B(n820), .Z(n822) );
  XOR U1356 ( .A(a[4059]), .B(n807), .Z(n809) );
  XOR U1357 ( .A(a[4062]), .B(n795), .Z(n797) );
  XOR U1358 ( .A(a[4065]), .B(n783), .Z(n785) );
  XOR U1359 ( .A(a[4068]), .B(n771), .Z(n773) );
  XOR U1360 ( .A(a[4071]), .B(n758), .Z(n760) );
  XOR U1361 ( .A(a[4074]), .B(n746), .Z(n748) );
  XOR U1362 ( .A(a[4077]), .B(n734), .Z(n736) );
  XOR U1363 ( .A(a[4080]), .B(n721), .Z(n723) );
  XOR U1364 ( .A(a[4083]), .B(n709), .Z(n711) );
  XOR U1365 ( .A(a[4086]), .B(n697), .Z(n699) );
  XOR U1366 ( .A(a[4089]), .B(n684), .Z(n686) );
  XOR U1367 ( .A(a[4092]), .B(n672), .Z(n674) );
  XOR U1368 ( .A(a[1]), .B(n16380), .Z(n9278) );
  XOR U1369 ( .A(a[4]), .B(n16371), .Z(n561) );
  XOR U1370 ( .A(a[7]), .B(n16362), .Z(n228) );
  XOR U1371 ( .A(a[10]), .B(n16353), .Z(n12978) );
  XOR U1372 ( .A(a[13]), .B(n16344), .Z(n11745) );
  XOR U1373 ( .A(a[16]), .B(n16335), .Z(n10512) );
  XOR U1374 ( .A(a[19]), .B(n16326), .Z(n9279) );
  XOR U1375 ( .A(a[22]), .B(n16317), .Z(n8045) );
  XOR U1376 ( .A(a[25]), .B(n16308), .Z(n6812) );
  XOR U1377 ( .A(a[28]), .B(n16299), .Z(n5579) );
  XOR U1378 ( .A(a[31]), .B(n16290), .Z(n4345) );
  XOR U1379 ( .A(a[34]), .B(n16281), .Z(n3112) );
  XOR U1380 ( .A(a[37]), .B(n16272), .Z(n1879) );
  XOR U1381 ( .A(a[40]), .B(n16263), .Z(n661) );
  XOR U1382 ( .A(a[43]), .B(n16254), .Z(n628) );
  XOR U1383 ( .A(a[46]), .B(n16245), .Z(n595) );
  XOR U1384 ( .A(a[49]), .B(n16236), .Z(n562) );
  XOR U1385 ( .A(a[52]), .B(n16227), .Z(n528) );
  XOR U1386 ( .A(a[55]), .B(n16218), .Z(n495) );
  XOR U1387 ( .A(a[58]), .B(n16209), .Z(n462) );
  XOR U1388 ( .A(a[61]), .B(n16200), .Z(n428) );
  XOR U1389 ( .A(a[64]), .B(n16191), .Z(n395) );
  XOR U1390 ( .A(a[67]), .B(n16182), .Z(n362) );
  XOR U1391 ( .A(a[70]), .B(n16173), .Z(n328) );
  XOR U1392 ( .A(a[73]), .B(n16164), .Z(n295) );
  XOR U1393 ( .A(a[76]), .B(n16155), .Z(n262) );
  XOR U1394 ( .A(a[79]), .B(n16146), .Z(n229) );
  XOR U1395 ( .A(a[82]), .B(n16137), .Z(n195) );
  XOR U1396 ( .A(a[85]), .B(n16128), .Z(n162) );
  XOR U1397 ( .A(a[88]), .B(n16119), .Z(n129) );
  XOR U1398 ( .A(a[91]), .B(n16110), .Z(n95) );
  XOR U1399 ( .A(a[94]), .B(n16101), .Z(n62) );
  XOR U1400 ( .A(a[97]), .B(n16092), .Z(n29) );
  XOR U1401 ( .A(a[100]), .B(n16083), .Z(n13348) );
  XOR U1402 ( .A(a[103]), .B(n16074), .Z(n13225) );
  XOR U1403 ( .A(a[106]), .B(n16065), .Z(n13102) );
  XOR U1404 ( .A(a[109]), .B(n16056), .Z(n12979) );
  XOR U1405 ( .A(a[112]), .B(n16047), .Z(n12855) );
  XOR U1406 ( .A(a[115]), .B(n16038), .Z(n12732) );
  XOR U1407 ( .A(a[118]), .B(n16029), .Z(n12609) );
  XOR U1408 ( .A(a[121]), .B(n16020), .Z(n12485) );
  XOR U1409 ( .A(a[124]), .B(n16011), .Z(n12362) );
  XOR U1410 ( .A(a[127]), .B(n16002), .Z(n12239) );
  XOR U1411 ( .A(a[130]), .B(n15993), .Z(n12115) );
  XOR U1412 ( .A(a[133]), .B(n15984), .Z(n11992) );
  XOR U1413 ( .A(a[136]), .B(n15975), .Z(n11869) );
  XOR U1414 ( .A(a[139]), .B(n15966), .Z(n11746) );
  XOR U1415 ( .A(a[142]), .B(n15957), .Z(n11622) );
  XOR U1416 ( .A(a[145]), .B(n15948), .Z(n11499) );
  XOR U1417 ( .A(a[148]), .B(n15939), .Z(n11376) );
  XOR U1418 ( .A(a[151]), .B(n15930), .Z(n11252) );
  XOR U1419 ( .A(a[154]), .B(n15921), .Z(n11129) );
  XOR U1420 ( .A(a[157]), .B(n15912), .Z(n11006) );
  XOR U1421 ( .A(a[160]), .B(n15903), .Z(n10882) );
  XOR U1422 ( .A(a[163]), .B(n15894), .Z(n10759) );
  XOR U1423 ( .A(a[166]), .B(n15885), .Z(n10636) );
  XOR U1424 ( .A(a[169]), .B(n15876), .Z(n10513) );
  XOR U1425 ( .A(a[172]), .B(n15867), .Z(n10389) );
  XOR U1426 ( .A(a[175]), .B(n15858), .Z(n10266) );
  XOR U1427 ( .A(a[178]), .B(n15849), .Z(n10143) );
  XOR U1428 ( .A(a[181]), .B(n15840), .Z(n10019) );
  XOR U1429 ( .A(a[184]), .B(n15831), .Z(n9896) );
  XOR U1430 ( .A(a[187]), .B(n15822), .Z(n9773) );
  XOR U1431 ( .A(a[190]), .B(n15813), .Z(n9649) );
  XOR U1432 ( .A(a[193]), .B(n15804), .Z(n9526) );
  XOR U1433 ( .A(a[196]), .B(n15795), .Z(n9403) );
  XOR U1434 ( .A(a[199]), .B(n15786), .Z(n9280) );
  XOR U1435 ( .A(a[202]), .B(n15777), .Z(n9155) );
  XOR U1436 ( .A(a[205]), .B(n15768), .Z(n9032) );
  XOR U1437 ( .A(a[208]), .B(n15759), .Z(n8909) );
  XOR U1438 ( .A(a[211]), .B(n15750), .Z(n8785) );
  XOR U1439 ( .A(a[214]), .B(n15741), .Z(n8662) );
  XOR U1440 ( .A(a[217]), .B(n15732), .Z(n8539) );
  XOR U1441 ( .A(a[220]), .B(n15723), .Z(n8415) );
  XOR U1442 ( .A(a[223]), .B(n15714), .Z(n8292) );
  XOR U1443 ( .A(a[226]), .B(n15705), .Z(n8169) );
  XOR U1444 ( .A(a[229]), .B(n15696), .Z(n8046) );
  XOR U1445 ( .A(a[232]), .B(n15687), .Z(n7922) );
  XOR U1446 ( .A(a[235]), .B(n15678), .Z(n7799) );
  XOR U1447 ( .A(a[238]), .B(n15669), .Z(n7676) );
  XOR U1448 ( .A(a[241]), .B(n15660), .Z(n7552) );
  XOR U1449 ( .A(a[244]), .B(n15651), .Z(n7429) );
  XOR U1450 ( .A(a[247]), .B(n15642), .Z(n7306) );
  XOR U1451 ( .A(a[250]), .B(n15633), .Z(n7182) );
  XOR U1452 ( .A(a[253]), .B(n15624), .Z(n7059) );
  XOR U1453 ( .A(a[256]), .B(n15615), .Z(n6936) );
  XOR U1454 ( .A(a[259]), .B(n15606), .Z(n6813) );
  XOR U1455 ( .A(a[262]), .B(n15597), .Z(n6689) );
  XOR U1456 ( .A(a[265]), .B(n15588), .Z(n6566) );
  XOR U1457 ( .A(a[268]), .B(n15579), .Z(n6443) );
  XOR U1458 ( .A(a[271]), .B(n15570), .Z(n6319) );
  XOR U1459 ( .A(a[274]), .B(n15561), .Z(n6196) );
  XOR U1460 ( .A(a[277]), .B(n15552), .Z(n6073) );
  XOR U1461 ( .A(a[280]), .B(n15543), .Z(n5949) );
  XOR U1462 ( .A(a[283]), .B(n15534), .Z(n5826) );
  XOR U1463 ( .A(a[286]), .B(n15525), .Z(n5703) );
  XOR U1464 ( .A(a[289]), .B(n15516), .Z(n5580) );
  XOR U1465 ( .A(a[292]), .B(n15507), .Z(n5456) );
  XOR U1466 ( .A(a[295]), .B(n15498), .Z(n5333) );
  XOR U1467 ( .A(a[298]), .B(n15489), .Z(n5210) );
  XOR U1468 ( .A(a[301]), .B(n15480), .Z(n5085) );
  XOR U1469 ( .A(a[304]), .B(n15471), .Z(n4962) );
  XOR U1470 ( .A(a[307]), .B(n15462), .Z(n4839) );
  XOR U1471 ( .A(a[310]), .B(n15453), .Z(n4715) );
  XOR U1472 ( .A(a[313]), .B(n15444), .Z(n4592) );
  XOR U1473 ( .A(a[316]), .B(n15435), .Z(n4469) );
  XOR U1474 ( .A(a[319]), .B(n15426), .Z(n4346) );
  XOR U1475 ( .A(a[322]), .B(n15417), .Z(n4222) );
  XOR U1476 ( .A(a[325]), .B(n15408), .Z(n4099) );
  XOR U1477 ( .A(a[328]), .B(n15399), .Z(n3976) );
  XOR U1478 ( .A(a[331]), .B(n15390), .Z(n3852) );
  XOR U1479 ( .A(a[334]), .B(n15381), .Z(n3729) );
  XOR U1480 ( .A(a[337]), .B(n15372), .Z(n3606) );
  XOR U1481 ( .A(a[340]), .B(n15363), .Z(n3482) );
  XOR U1482 ( .A(a[343]), .B(n15354), .Z(n3359) );
  XOR U1483 ( .A(a[346]), .B(n15345), .Z(n3236) );
  XOR U1484 ( .A(a[349]), .B(n15336), .Z(n3113) );
  XOR U1485 ( .A(a[352]), .B(n15327), .Z(n2989) );
  XOR U1486 ( .A(a[355]), .B(n15318), .Z(n2866) );
  XOR U1487 ( .A(a[358]), .B(n15309), .Z(n2743) );
  XOR U1488 ( .A(a[361]), .B(n15300), .Z(n2619) );
  XOR U1489 ( .A(a[364]), .B(n15291), .Z(n2496) );
  XOR U1490 ( .A(a[367]), .B(n15282), .Z(n2373) );
  XOR U1491 ( .A(a[370]), .B(n15273), .Z(n2249) );
  XOR U1492 ( .A(a[373]), .B(n15264), .Z(n2126) );
  XOR U1493 ( .A(a[376]), .B(n15255), .Z(n2003) );
  XOR U1494 ( .A(a[379]), .B(n15246), .Z(n1880) );
  XOR U1495 ( .A(a[382]), .B(n15237), .Z(n1756) );
  XOR U1496 ( .A(a[385]), .B(n15228), .Z(n1633) );
  XOR U1497 ( .A(a[388]), .B(n15219), .Z(n1510) );
  XOR U1498 ( .A(a[391]), .B(n15210), .Z(n1386) );
  XOR U1499 ( .A(a[394]), .B(n15201), .Z(n1263) );
  XOR U1500 ( .A(a[397]), .B(n15192), .Z(n1140) );
  XOR U1501 ( .A(a[400]), .B(n15183), .Z(n1015) );
  XOR U1502 ( .A(a[403]), .B(n15174), .Z(n892) );
  XOR U1503 ( .A(a[406]), .B(n15165), .Z(n769) );
  XOR U1504 ( .A(a[409]), .B(n15156), .Z(n662) );
  XOR U1505 ( .A(a[412]), .B(n15147), .Z(n658) );
  XOR U1506 ( .A(a[415]), .B(n15138), .Z(n655) );
  XOR U1507 ( .A(a[418]), .B(n15129), .Z(n652) );
  XOR U1508 ( .A(a[421]), .B(n15120), .Z(n648) );
  XOR U1509 ( .A(a[424]), .B(n15111), .Z(n645) );
  XOR U1510 ( .A(a[427]), .B(n15102), .Z(n642) );
  XOR U1511 ( .A(a[430]), .B(n15093), .Z(n638) );
  XOR U1512 ( .A(a[433]), .B(n15084), .Z(n635) );
  XOR U1513 ( .A(a[436]), .B(n15075), .Z(n632) );
  XOR U1514 ( .A(a[439]), .B(n15066), .Z(n629) );
  XOR U1515 ( .A(a[442]), .B(n15057), .Z(n625) );
  XOR U1516 ( .A(a[445]), .B(n15048), .Z(n622) );
  XOR U1517 ( .A(a[448]), .B(n15039), .Z(n619) );
  XOR U1518 ( .A(a[451]), .B(n15030), .Z(n615) );
  XOR U1519 ( .A(a[454]), .B(n15021), .Z(n612) );
  XOR U1520 ( .A(a[457]), .B(n15012), .Z(n609) );
  XOR U1521 ( .A(a[460]), .B(n15003), .Z(n605) );
  XOR U1522 ( .A(a[463]), .B(n14994), .Z(n602) );
  XOR U1523 ( .A(a[466]), .B(n14985), .Z(n599) );
  XOR U1524 ( .A(a[469]), .B(n14976), .Z(n596) );
  XOR U1525 ( .A(a[472]), .B(n14967), .Z(n592) );
  XOR U1526 ( .A(a[475]), .B(n14958), .Z(n589) );
  XOR U1527 ( .A(a[478]), .B(n14949), .Z(n586) );
  XOR U1528 ( .A(a[481]), .B(n14940), .Z(n582) );
  XOR U1529 ( .A(a[484]), .B(n14931), .Z(n579) );
  XOR U1530 ( .A(a[487]), .B(n14922), .Z(n576) );
  XOR U1531 ( .A(a[490]), .B(n14913), .Z(n572) );
  XOR U1532 ( .A(a[493]), .B(n14904), .Z(n569) );
  XOR U1533 ( .A(a[496]), .B(n14895), .Z(n566) );
  XOR U1534 ( .A(a[499]), .B(n14886), .Z(n563) );
  XOR U1535 ( .A(a[502]), .B(n14877), .Z(n558) );
  XOR U1536 ( .A(a[505]), .B(n14868), .Z(n555) );
  XOR U1537 ( .A(a[508]), .B(n14859), .Z(n552) );
  XOR U1538 ( .A(a[511]), .B(n14850), .Z(n548) );
  XOR U1539 ( .A(a[514]), .B(n14841), .Z(n545) );
  XOR U1540 ( .A(a[517]), .B(n14832), .Z(n542) );
  XOR U1541 ( .A(a[520]), .B(n14823), .Z(n538) );
  XOR U1542 ( .A(a[523]), .B(n14814), .Z(n535) );
  XOR U1543 ( .A(a[526]), .B(n14805), .Z(n532) );
  XOR U1544 ( .A(a[529]), .B(n14796), .Z(n529) );
  XOR U1545 ( .A(a[532]), .B(n14787), .Z(n525) );
  XOR U1546 ( .A(a[535]), .B(n14778), .Z(n522) );
  XOR U1547 ( .A(a[538]), .B(n14769), .Z(n519) );
  XOR U1548 ( .A(a[541]), .B(n14760), .Z(n515) );
  XOR U1549 ( .A(a[544]), .B(n14751), .Z(n512) );
  XOR U1550 ( .A(a[547]), .B(n14742), .Z(n509) );
  XOR U1551 ( .A(a[550]), .B(n14733), .Z(n505) );
  XOR U1552 ( .A(a[553]), .B(n14724), .Z(n502) );
  XOR U1553 ( .A(a[556]), .B(n14715), .Z(n499) );
  XOR U1554 ( .A(a[559]), .B(n14706), .Z(n496) );
  XOR U1555 ( .A(a[562]), .B(n14697), .Z(n492) );
  XOR U1556 ( .A(a[565]), .B(n14688), .Z(n489) );
  XOR U1557 ( .A(a[568]), .B(n14679), .Z(n486) );
  XOR U1558 ( .A(a[571]), .B(n14670), .Z(n482) );
  XOR U1559 ( .A(a[574]), .B(n14661), .Z(n479) );
  XOR U1560 ( .A(a[577]), .B(n14652), .Z(n476) );
  XOR U1561 ( .A(a[580]), .B(n14643), .Z(n472) );
  XOR U1562 ( .A(a[583]), .B(n14634), .Z(n469) );
  XOR U1563 ( .A(a[586]), .B(n14625), .Z(n466) );
  XOR U1564 ( .A(a[589]), .B(n14616), .Z(n463) );
  XOR U1565 ( .A(a[592]), .B(n14607), .Z(n459) );
  XOR U1566 ( .A(a[595]), .B(n14598), .Z(n456) );
  XOR U1567 ( .A(a[598]), .B(n14589), .Z(n453) );
  XOR U1568 ( .A(a[601]), .B(n14580), .Z(n448) );
  XOR U1569 ( .A(a[604]), .B(n14571), .Z(n445) );
  XOR U1570 ( .A(a[607]), .B(n14562), .Z(n442) );
  XOR U1571 ( .A(a[610]), .B(n14553), .Z(n438) );
  XOR U1572 ( .A(a[613]), .B(n14544), .Z(n435) );
  XOR U1573 ( .A(a[616]), .B(n14535), .Z(n432) );
  XOR U1574 ( .A(a[619]), .B(n14526), .Z(n429) );
  XOR U1575 ( .A(a[622]), .B(n14517), .Z(n425) );
  XOR U1576 ( .A(a[625]), .B(n14508), .Z(n422) );
  XOR U1577 ( .A(a[628]), .B(n14499), .Z(n419) );
  XOR U1578 ( .A(a[631]), .B(n14490), .Z(n415) );
  XOR U1579 ( .A(a[634]), .B(n14481), .Z(n412) );
  XOR U1580 ( .A(a[637]), .B(n14472), .Z(n409) );
  XOR U1581 ( .A(a[640]), .B(n14463), .Z(n405) );
  XOR U1582 ( .A(a[643]), .B(n14454), .Z(n402) );
  XOR U1583 ( .A(a[646]), .B(n14445), .Z(n399) );
  XOR U1584 ( .A(a[649]), .B(n14436), .Z(n396) );
  XOR U1585 ( .A(a[652]), .B(n14427), .Z(n392) );
  XOR U1586 ( .A(a[655]), .B(n14418), .Z(n389) );
  XOR U1587 ( .A(a[658]), .B(n14409), .Z(n386) );
  XOR U1588 ( .A(a[661]), .B(n14400), .Z(n382) );
  XOR U1589 ( .A(a[664]), .B(n14391), .Z(n379) );
  XOR U1590 ( .A(a[667]), .B(n14382), .Z(n376) );
  XOR U1591 ( .A(a[670]), .B(n14373), .Z(n372) );
  XOR U1592 ( .A(a[673]), .B(n14364), .Z(n369) );
  XOR U1593 ( .A(a[676]), .B(n14355), .Z(n366) );
  XOR U1594 ( .A(a[679]), .B(n14346), .Z(n363) );
  XOR U1595 ( .A(a[682]), .B(n14337), .Z(n359) );
  XOR U1596 ( .A(a[685]), .B(n14328), .Z(n356) );
  XOR U1597 ( .A(a[688]), .B(n14319), .Z(n353) );
  XOR U1598 ( .A(a[691]), .B(n14310), .Z(n349) );
  XOR U1599 ( .A(a[694]), .B(n14301), .Z(n346) );
  XOR U1600 ( .A(a[697]), .B(n14292), .Z(n343) );
  XOR U1601 ( .A(a[700]), .B(n14283), .Z(n338) );
  XOR U1602 ( .A(a[703]), .B(n14274), .Z(n335) );
  XOR U1603 ( .A(a[706]), .B(n14265), .Z(n332) );
  XOR U1604 ( .A(a[709]), .B(n14256), .Z(n329) );
  XOR U1605 ( .A(a[712]), .B(n14247), .Z(n325) );
  XOR U1606 ( .A(a[715]), .B(n14238), .Z(n322) );
  XOR U1607 ( .A(a[718]), .B(n14229), .Z(n319) );
  XOR U1608 ( .A(a[721]), .B(n14220), .Z(n315) );
  XOR U1609 ( .A(a[724]), .B(n14211), .Z(n312) );
  XOR U1610 ( .A(a[727]), .B(n14202), .Z(n309) );
  XOR U1611 ( .A(a[730]), .B(n14193), .Z(n305) );
  XOR U1612 ( .A(a[733]), .B(n14184), .Z(n302) );
  XOR U1613 ( .A(a[736]), .B(n14175), .Z(n299) );
  XOR U1614 ( .A(a[739]), .B(n14166), .Z(n296) );
  XOR U1615 ( .A(a[742]), .B(n14157), .Z(n292) );
  XOR U1616 ( .A(a[745]), .B(n14148), .Z(n289) );
  XOR U1617 ( .A(a[748]), .B(n14139), .Z(n286) );
  XOR U1618 ( .A(a[751]), .B(n14130), .Z(n282) );
  XOR U1619 ( .A(a[754]), .B(n14121), .Z(n279) );
  XOR U1620 ( .A(a[757]), .B(n14112), .Z(n276) );
  XOR U1621 ( .A(a[760]), .B(n14103), .Z(n272) );
  XOR U1622 ( .A(a[763]), .B(n14094), .Z(n269) );
  XOR U1623 ( .A(a[766]), .B(n14085), .Z(n266) );
  XOR U1624 ( .A(a[769]), .B(n14076), .Z(n263) );
  XOR U1625 ( .A(a[772]), .B(n14067), .Z(n259) );
  XOR U1626 ( .A(a[775]), .B(n14058), .Z(n256) );
  XOR U1627 ( .A(a[778]), .B(n14049), .Z(n253) );
  XOR U1628 ( .A(a[781]), .B(n14040), .Z(n249) );
  XOR U1629 ( .A(a[784]), .B(n14031), .Z(n246) );
  XOR U1630 ( .A(a[787]), .B(n14022), .Z(n243) );
  XOR U1631 ( .A(a[790]), .B(n14013), .Z(n239) );
  XOR U1632 ( .A(a[793]), .B(n14004), .Z(n236) );
  XOR U1633 ( .A(a[796]), .B(n13995), .Z(n233) );
  XOR U1634 ( .A(a[799]), .B(n13986), .Z(n230) );
  XOR U1635 ( .A(a[802]), .B(n13977), .Z(n225) );
  XOR U1636 ( .A(a[805]), .B(n13968), .Z(n222) );
  XOR U1637 ( .A(a[808]), .B(n13959), .Z(n219) );
  XOR U1638 ( .A(a[811]), .B(n13950), .Z(n215) );
  XOR U1639 ( .A(a[814]), .B(n13941), .Z(n212) );
  XOR U1640 ( .A(a[817]), .B(n13932), .Z(n209) );
  XOR U1641 ( .A(a[820]), .B(n13923), .Z(n205) );
  XOR U1642 ( .A(a[823]), .B(n13914), .Z(n202) );
  XOR U1643 ( .A(a[826]), .B(n13905), .Z(n199) );
  XOR U1644 ( .A(a[829]), .B(n13896), .Z(n196) );
  XOR U1645 ( .A(a[832]), .B(n13887), .Z(n192) );
  XOR U1646 ( .A(a[835]), .B(n13878), .Z(n189) );
  XOR U1647 ( .A(a[838]), .B(n13869), .Z(n186) );
  XOR U1648 ( .A(a[841]), .B(n13860), .Z(n182) );
  XOR U1649 ( .A(a[844]), .B(n13851), .Z(n179) );
  XOR U1650 ( .A(a[847]), .B(n13842), .Z(n176) );
  XOR U1651 ( .A(a[850]), .B(n13833), .Z(n172) );
  XOR U1652 ( .A(a[853]), .B(n13824), .Z(n169) );
  XOR U1653 ( .A(a[856]), .B(n13815), .Z(n166) );
  XOR U1654 ( .A(a[859]), .B(n13806), .Z(n163) );
  XOR U1655 ( .A(a[862]), .B(n13797), .Z(n159) );
  XOR U1656 ( .A(a[865]), .B(n13788), .Z(n156) );
  XOR U1657 ( .A(a[868]), .B(n13779), .Z(n153) );
  XOR U1658 ( .A(a[871]), .B(n13770), .Z(n149) );
  XOR U1659 ( .A(a[874]), .B(n13761), .Z(n146) );
  XOR U1660 ( .A(a[877]), .B(n13752), .Z(n143) );
  XOR U1661 ( .A(a[880]), .B(n13743), .Z(n139) );
  XOR U1662 ( .A(a[883]), .B(n13734), .Z(n136) );
  XOR U1663 ( .A(a[886]), .B(n13725), .Z(n133) );
  XOR U1664 ( .A(a[889]), .B(n13716), .Z(n130) );
  XOR U1665 ( .A(a[892]), .B(n13707), .Z(n126) );
  XOR U1666 ( .A(a[895]), .B(n13698), .Z(n123) );
  XOR U1667 ( .A(a[898]), .B(n13689), .Z(n120) );
  XOR U1668 ( .A(a[901]), .B(n13680), .Z(n115) );
  XOR U1669 ( .A(a[904]), .B(n13671), .Z(n112) );
  XOR U1670 ( .A(a[907]), .B(n13662), .Z(n109) );
  XOR U1671 ( .A(a[910]), .B(n13653), .Z(n105) );
  XOR U1672 ( .A(a[913]), .B(n13644), .Z(n102) );
  XOR U1673 ( .A(a[916]), .B(n13635), .Z(n99) );
  XOR U1674 ( .A(a[919]), .B(n13626), .Z(n96) );
  XOR U1675 ( .A(a[922]), .B(n13617), .Z(n92) );
  XOR U1676 ( .A(a[925]), .B(n13608), .Z(n89) );
  XOR U1677 ( .A(a[928]), .B(n13599), .Z(n86) );
  XOR U1678 ( .A(a[931]), .B(n13590), .Z(n82) );
  XOR U1679 ( .A(a[934]), .B(n13581), .Z(n79) );
  XOR U1680 ( .A(a[937]), .B(n13572), .Z(n76) );
  XOR U1681 ( .A(a[940]), .B(n13563), .Z(n72) );
  XOR U1682 ( .A(a[943]), .B(n13554), .Z(n69) );
  XOR U1683 ( .A(a[946]), .B(n13545), .Z(n66) );
  XOR U1684 ( .A(a[949]), .B(n13536), .Z(n63) );
  XOR U1685 ( .A(a[952]), .B(n13527), .Z(n59) );
  XOR U1686 ( .A(a[955]), .B(n13518), .Z(n56) );
  XOR U1687 ( .A(a[958]), .B(n13509), .Z(n53) );
  XOR U1688 ( .A(a[961]), .B(n13500), .Z(n49) );
  XOR U1689 ( .A(a[964]), .B(n13491), .Z(n46) );
  XOR U1690 ( .A(a[967]), .B(n13482), .Z(n43) );
  XOR U1691 ( .A(a[970]), .B(n13473), .Z(n39) );
  XOR U1692 ( .A(a[973]), .B(n13464), .Z(n36) );
  XOR U1693 ( .A(a[976]), .B(n13455), .Z(n33) );
  XOR U1694 ( .A(a[979]), .B(n13446), .Z(n30) );
  XOR U1695 ( .A(a[982]), .B(n13437), .Z(n26) );
  XOR U1696 ( .A(a[985]), .B(n13428), .Z(n23) );
  XOR U1697 ( .A(a[988]), .B(n13419), .Z(n20) );
  XOR U1698 ( .A(a[991]), .B(n13410), .Z(n16) );
  XOR U1699 ( .A(a[994]), .B(n13401), .Z(n13) );
  XOR U1700 ( .A(a[997]), .B(n13392), .Z(n10) );
  XOR U1701 ( .A(a[1000]), .B(n13382), .Z(n13384) );
  XOR U1702 ( .A(a[1003]), .B(n13370), .Z(n13372) );
  XOR U1703 ( .A(a[1006]), .B(n13358), .Z(n13360) );
  XOR U1704 ( .A(a[1009]), .B(n13345), .Z(n13347) );
  XOR U1705 ( .A(a[1012]), .B(n13333), .Z(n13335) );
  XOR U1706 ( .A(a[1015]), .B(n13321), .Z(n13323) );
  XOR U1707 ( .A(a[1018]), .B(n13309), .Z(n13311) );
  XOR U1708 ( .A(a[1021]), .B(n13296), .Z(n13298) );
  XOR U1709 ( .A(a[1024]), .B(n13284), .Z(n13286) );
  XOR U1710 ( .A(a[1027]), .B(n13272), .Z(n13274) );
  XOR U1711 ( .A(a[1030]), .B(n13259), .Z(n13261) );
  XOR U1712 ( .A(a[1033]), .B(n13247), .Z(n13249) );
  XOR U1713 ( .A(a[1036]), .B(n13235), .Z(n13237) );
  XOR U1714 ( .A(a[1039]), .B(n13222), .Z(n13224) );
  XOR U1715 ( .A(a[1042]), .B(n13210), .Z(n13212) );
  XOR U1716 ( .A(a[1045]), .B(n13198), .Z(n13200) );
  XOR U1717 ( .A(a[1048]), .B(n13186), .Z(n13188) );
  XOR U1718 ( .A(a[1051]), .B(n13173), .Z(n13175) );
  XOR U1719 ( .A(a[1054]), .B(n13161), .Z(n13163) );
  XOR U1720 ( .A(a[1057]), .B(n13149), .Z(n13151) );
  XOR U1721 ( .A(a[1060]), .B(n13136), .Z(n13138) );
  XOR U1722 ( .A(a[1063]), .B(n13124), .Z(n13126) );
  XOR U1723 ( .A(a[1066]), .B(n13112), .Z(n13114) );
  XOR U1724 ( .A(a[1069]), .B(n13099), .Z(n13101) );
  XOR U1725 ( .A(a[1072]), .B(n13087), .Z(n13089) );
  XOR U1726 ( .A(a[1075]), .B(n13075), .Z(n13077) );
  XOR U1727 ( .A(a[1078]), .B(n13063), .Z(n13065) );
  XOR U1728 ( .A(a[1081]), .B(n13050), .Z(n13052) );
  XOR U1729 ( .A(a[1084]), .B(n13038), .Z(n13040) );
  XOR U1730 ( .A(a[1087]), .B(n13026), .Z(n13028) );
  XOR U1731 ( .A(a[1090]), .B(n13013), .Z(n13015) );
  XOR U1732 ( .A(a[1093]), .B(n13001), .Z(n13003) );
  XOR U1733 ( .A(a[1096]), .B(n12989), .Z(n12991) );
  XOR U1734 ( .A(a[1099]), .B(n12975), .Z(n12977) );
  XOR U1735 ( .A(a[1102]), .B(n12963), .Z(n12965) );
  XOR U1736 ( .A(a[1105]), .B(n12951), .Z(n12953) );
  XOR U1737 ( .A(a[1108]), .B(n12939), .Z(n12941) );
  XOR U1738 ( .A(a[1111]), .B(n12926), .Z(n12928) );
  XOR U1739 ( .A(a[1114]), .B(n12914), .Z(n12916) );
  XOR U1740 ( .A(a[1117]), .B(n12902), .Z(n12904) );
  XOR U1741 ( .A(a[1120]), .B(n12889), .Z(n12891) );
  XOR U1742 ( .A(a[1123]), .B(n12877), .Z(n12879) );
  XOR U1743 ( .A(a[1126]), .B(n12865), .Z(n12867) );
  XOR U1744 ( .A(a[1129]), .B(n12852), .Z(n12854) );
  XOR U1745 ( .A(a[1132]), .B(n12840), .Z(n12842) );
  XOR U1746 ( .A(a[1135]), .B(n12828), .Z(n12830) );
  XOR U1747 ( .A(a[1138]), .B(n12816), .Z(n12818) );
  XOR U1748 ( .A(a[1141]), .B(n12803), .Z(n12805) );
  XOR U1749 ( .A(a[1144]), .B(n12791), .Z(n12793) );
  XOR U1750 ( .A(a[1147]), .B(n12779), .Z(n12781) );
  XOR U1751 ( .A(a[1150]), .B(n12766), .Z(n12768) );
  XOR U1752 ( .A(a[1153]), .B(n12754), .Z(n12756) );
  XOR U1753 ( .A(a[1156]), .B(n12742), .Z(n12744) );
  XOR U1754 ( .A(a[1159]), .B(n12729), .Z(n12731) );
  XOR U1755 ( .A(a[1162]), .B(n12717), .Z(n12719) );
  XOR U1756 ( .A(a[1165]), .B(n12705), .Z(n12707) );
  XOR U1757 ( .A(a[1168]), .B(n12693), .Z(n12695) );
  XOR U1758 ( .A(a[1171]), .B(n12680), .Z(n12682) );
  XOR U1759 ( .A(a[1174]), .B(n12668), .Z(n12670) );
  XOR U1760 ( .A(a[1177]), .B(n12656), .Z(n12658) );
  XOR U1761 ( .A(a[1180]), .B(n12643), .Z(n12645) );
  XOR U1762 ( .A(a[1183]), .B(n12631), .Z(n12633) );
  XOR U1763 ( .A(a[1186]), .B(n12619), .Z(n12621) );
  XOR U1764 ( .A(a[1189]), .B(n12606), .Z(n12608) );
  XOR U1765 ( .A(a[1192]), .B(n12594), .Z(n12596) );
  XOR U1766 ( .A(a[1195]), .B(n12582), .Z(n12584) );
  XOR U1767 ( .A(a[1198]), .B(n12570), .Z(n12572) );
  XOR U1768 ( .A(a[1201]), .B(n12556), .Z(n12558) );
  XOR U1769 ( .A(a[1204]), .B(n12544), .Z(n12546) );
  XOR U1770 ( .A(a[1207]), .B(n12532), .Z(n12534) );
  XOR U1771 ( .A(a[1210]), .B(n12519), .Z(n12521) );
  XOR U1772 ( .A(a[1213]), .B(n12507), .Z(n12509) );
  XOR U1773 ( .A(a[1216]), .B(n12495), .Z(n12497) );
  XOR U1774 ( .A(a[1219]), .B(n12482), .Z(n12484) );
  XOR U1775 ( .A(a[1222]), .B(n12470), .Z(n12472) );
  XOR U1776 ( .A(a[1225]), .B(n12458), .Z(n12460) );
  XOR U1777 ( .A(a[1228]), .B(n12446), .Z(n12448) );
  XOR U1778 ( .A(a[1231]), .B(n12433), .Z(n12435) );
  XOR U1779 ( .A(a[1234]), .B(n12421), .Z(n12423) );
  XOR U1780 ( .A(a[1237]), .B(n12409), .Z(n12411) );
  XOR U1781 ( .A(a[1240]), .B(n12396), .Z(n12398) );
  XOR U1782 ( .A(a[1243]), .B(n12384), .Z(n12386) );
  XOR U1783 ( .A(a[1246]), .B(n12372), .Z(n12374) );
  XOR U1784 ( .A(a[1249]), .B(n12359), .Z(n12361) );
  XOR U1785 ( .A(a[1252]), .B(n12347), .Z(n12349) );
  XOR U1786 ( .A(a[1255]), .B(n12335), .Z(n12337) );
  XOR U1787 ( .A(a[1258]), .B(n12323), .Z(n12325) );
  XOR U1788 ( .A(a[1261]), .B(n12310), .Z(n12312) );
  XOR U1789 ( .A(a[1264]), .B(n12298), .Z(n12300) );
  XOR U1790 ( .A(a[1267]), .B(n12286), .Z(n12288) );
  XOR U1791 ( .A(a[1270]), .B(n12273), .Z(n12275) );
  XOR U1792 ( .A(a[1273]), .B(n12261), .Z(n12263) );
  XOR U1793 ( .A(a[1276]), .B(n12249), .Z(n12251) );
  XOR U1794 ( .A(a[1279]), .B(n12236), .Z(n12238) );
  XOR U1795 ( .A(a[1282]), .B(n12224), .Z(n12226) );
  XOR U1796 ( .A(a[1285]), .B(n12212), .Z(n12214) );
  XOR U1797 ( .A(a[1288]), .B(n12200), .Z(n12202) );
  XOR U1798 ( .A(a[1291]), .B(n12187), .Z(n12189) );
  XOR U1799 ( .A(a[1294]), .B(n12175), .Z(n12177) );
  XOR U1800 ( .A(a[1297]), .B(n12163), .Z(n12165) );
  XOR U1801 ( .A(a[1300]), .B(n12149), .Z(n12151) );
  XOR U1802 ( .A(a[1303]), .B(n12137), .Z(n12139) );
  XOR U1803 ( .A(a[1306]), .B(n12125), .Z(n12127) );
  XOR U1804 ( .A(a[1309]), .B(n12112), .Z(n12114) );
  XOR U1805 ( .A(a[1312]), .B(n12100), .Z(n12102) );
  XOR U1806 ( .A(a[1315]), .B(n12088), .Z(n12090) );
  XOR U1807 ( .A(a[1318]), .B(n12076), .Z(n12078) );
  XOR U1808 ( .A(a[1321]), .B(n12063), .Z(n12065) );
  XOR U1809 ( .A(a[1324]), .B(n12051), .Z(n12053) );
  XOR U1810 ( .A(a[1327]), .B(n12039), .Z(n12041) );
  XOR U1811 ( .A(a[1330]), .B(n12026), .Z(n12028) );
  XOR U1812 ( .A(a[1333]), .B(n12014), .Z(n12016) );
  XOR U1813 ( .A(a[1336]), .B(n12002), .Z(n12004) );
  XOR U1814 ( .A(a[1339]), .B(n11989), .Z(n11991) );
  XOR U1815 ( .A(a[1342]), .B(n11977), .Z(n11979) );
  XOR U1816 ( .A(a[1345]), .B(n11965), .Z(n11967) );
  XOR U1817 ( .A(a[1348]), .B(n11953), .Z(n11955) );
  XOR U1818 ( .A(a[1351]), .B(n11940), .Z(n11942) );
  XOR U1819 ( .A(a[1354]), .B(n11928), .Z(n11930) );
  XOR U1820 ( .A(a[1357]), .B(n11916), .Z(n11918) );
  XOR U1821 ( .A(a[1360]), .B(n11903), .Z(n11905) );
  XOR U1822 ( .A(a[1363]), .B(n11891), .Z(n11893) );
  XOR U1823 ( .A(a[1366]), .B(n11879), .Z(n11881) );
  XOR U1824 ( .A(a[1369]), .B(n11866), .Z(n11868) );
  XOR U1825 ( .A(a[1372]), .B(n11854), .Z(n11856) );
  XOR U1826 ( .A(a[1375]), .B(n11842), .Z(n11844) );
  XOR U1827 ( .A(a[1378]), .B(n11830), .Z(n11832) );
  XOR U1828 ( .A(a[1381]), .B(n11817), .Z(n11819) );
  XOR U1829 ( .A(a[1384]), .B(n11805), .Z(n11807) );
  XOR U1830 ( .A(a[1387]), .B(n11793), .Z(n11795) );
  XOR U1831 ( .A(a[1390]), .B(n11780), .Z(n11782) );
  XOR U1832 ( .A(a[1393]), .B(n11768), .Z(n11770) );
  XOR U1833 ( .A(a[1396]), .B(n11756), .Z(n11758) );
  XOR U1834 ( .A(a[1399]), .B(n11742), .Z(n11744) );
  XOR U1835 ( .A(a[1402]), .B(n11730), .Z(n11732) );
  XOR U1836 ( .A(a[1405]), .B(n11718), .Z(n11720) );
  XOR U1837 ( .A(a[1408]), .B(n11706), .Z(n11708) );
  XOR U1838 ( .A(a[1411]), .B(n11693), .Z(n11695) );
  XOR U1839 ( .A(a[1414]), .B(n11681), .Z(n11683) );
  XOR U1840 ( .A(a[1417]), .B(n11669), .Z(n11671) );
  XOR U1841 ( .A(a[1420]), .B(n11656), .Z(n11658) );
  XOR U1842 ( .A(a[1423]), .B(n11644), .Z(n11646) );
  XOR U1843 ( .A(a[1426]), .B(n11632), .Z(n11634) );
  XOR U1844 ( .A(a[1429]), .B(n11619), .Z(n11621) );
  XOR U1845 ( .A(a[1432]), .B(n11607), .Z(n11609) );
  XOR U1846 ( .A(a[1435]), .B(n11595), .Z(n11597) );
  XOR U1847 ( .A(a[1438]), .B(n11583), .Z(n11585) );
  XOR U1848 ( .A(a[1441]), .B(n11570), .Z(n11572) );
  XOR U1849 ( .A(a[1444]), .B(n11558), .Z(n11560) );
  XOR U1850 ( .A(a[1447]), .B(n11546), .Z(n11548) );
  XOR U1851 ( .A(a[1450]), .B(n11533), .Z(n11535) );
  XOR U1852 ( .A(a[1453]), .B(n11521), .Z(n11523) );
  XOR U1853 ( .A(a[1456]), .B(n11509), .Z(n11511) );
  XOR U1854 ( .A(a[1459]), .B(n11496), .Z(n11498) );
  XOR U1855 ( .A(a[1462]), .B(n11484), .Z(n11486) );
  XOR U1856 ( .A(a[1465]), .B(n11472), .Z(n11474) );
  XOR U1857 ( .A(a[1468]), .B(n11460), .Z(n11462) );
  XOR U1858 ( .A(a[1471]), .B(n11447), .Z(n11449) );
  XOR U1859 ( .A(a[1474]), .B(n11435), .Z(n11437) );
  XOR U1860 ( .A(a[1477]), .B(n11423), .Z(n11425) );
  XOR U1861 ( .A(a[1480]), .B(n11410), .Z(n11412) );
  XOR U1862 ( .A(a[1483]), .B(n11398), .Z(n11400) );
  XOR U1863 ( .A(a[1486]), .B(n11386), .Z(n11388) );
  XOR U1864 ( .A(a[1489]), .B(n11373), .Z(n11375) );
  XOR U1865 ( .A(a[1492]), .B(n11361), .Z(n11363) );
  XOR U1866 ( .A(a[1495]), .B(n11349), .Z(n11351) );
  XOR U1867 ( .A(a[1498]), .B(n11337), .Z(n11339) );
  XOR U1868 ( .A(a[1501]), .B(n11323), .Z(n11325) );
  XOR U1869 ( .A(a[1504]), .B(n11311), .Z(n11313) );
  XOR U1870 ( .A(a[1507]), .B(n11299), .Z(n11301) );
  XOR U1871 ( .A(a[1510]), .B(n11286), .Z(n11288) );
  XOR U1872 ( .A(a[1513]), .B(n11274), .Z(n11276) );
  XOR U1873 ( .A(a[1516]), .B(n11262), .Z(n11264) );
  XOR U1874 ( .A(a[1519]), .B(n11249), .Z(n11251) );
  XOR U1875 ( .A(a[1522]), .B(n11237), .Z(n11239) );
  XOR U1876 ( .A(a[1525]), .B(n11225), .Z(n11227) );
  XOR U1877 ( .A(a[1528]), .B(n11213), .Z(n11215) );
  XOR U1878 ( .A(a[1531]), .B(n11200), .Z(n11202) );
  XOR U1879 ( .A(a[1534]), .B(n11188), .Z(n11190) );
  XOR U1880 ( .A(a[1537]), .B(n11176), .Z(n11178) );
  XOR U1881 ( .A(a[1540]), .B(n11163), .Z(n11165) );
  XOR U1882 ( .A(a[1543]), .B(n11151), .Z(n11153) );
  XOR U1883 ( .A(a[1546]), .B(n11139), .Z(n11141) );
  XOR U1884 ( .A(a[1549]), .B(n11126), .Z(n11128) );
  XOR U1885 ( .A(a[1552]), .B(n11114), .Z(n11116) );
  XOR U1886 ( .A(a[1555]), .B(n11102), .Z(n11104) );
  XOR U1887 ( .A(a[1558]), .B(n11090), .Z(n11092) );
  XOR U1888 ( .A(a[1561]), .B(n11077), .Z(n11079) );
  XOR U1889 ( .A(a[1564]), .B(n11065), .Z(n11067) );
  XOR U1890 ( .A(a[1567]), .B(n11053), .Z(n11055) );
  XOR U1891 ( .A(a[1570]), .B(n11040), .Z(n11042) );
  XOR U1892 ( .A(a[1573]), .B(n11028), .Z(n11030) );
  XOR U1893 ( .A(a[1576]), .B(n11016), .Z(n11018) );
  XOR U1894 ( .A(a[1579]), .B(n11003), .Z(n11005) );
  XOR U1895 ( .A(a[1582]), .B(n10991), .Z(n10993) );
  XOR U1896 ( .A(a[1585]), .B(n10979), .Z(n10981) );
  XOR U1897 ( .A(a[1588]), .B(n10967), .Z(n10969) );
  XOR U1898 ( .A(a[1591]), .B(n10954), .Z(n10956) );
  XOR U1899 ( .A(a[1594]), .B(n10942), .Z(n10944) );
  XOR U1900 ( .A(a[1597]), .B(n10930), .Z(n10932) );
  XOR U1901 ( .A(a[1600]), .B(n10916), .Z(n10918) );
  XOR U1902 ( .A(a[1603]), .B(n10904), .Z(n10906) );
  XOR U1903 ( .A(a[1606]), .B(n10892), .Z(n10894) );
  XOR U1904 ( .A(a[1609]), .B(n10879), .Z(n10881) );
  XOR U1905 ( .A(a[1612]), .B(n10867), .Z(n10869) );
  XOR U1906 ( .A(a[1615]), .B(n10855), .Z(n10857) );
  XOR U1907 ( .A(a[1618]), .B(n10843), .Z(n10845) );
  XOR U1908 ( .A(a[1621]), .B(n10830), .Z(n10832) );
  XOR U1909 ( .A(a[1624]), .B(n10818), .Z(n10820) );
  XOR U1910 ( .A(a[1627]), .B(n10806), .Z(n10808) );
  XOR U1911 ( .A(a[1630]), .B(n10793), .Z(n10795) );
  XOR U1912 ( .A(a[1633]), .B(n10781), .Z(n10783) );
  XOR U1913 ( .A(a[1636]), .B(n10769), .Z(n10771) );
  XOR U1914 ( .A(a[1639]), .B(n10756), .Z(n10758) );
  XOR U1915 ( .A(a[1642]), .B(n10744), .Z(n10746) );
  XOR U1916 ( .A(a[1645]), .B(n10732), .Z(n10734) );
  XOR U1917 ( .A(a[1648]), .B(n10720), .Z(n10722) );
  XOR U1918 ( .A(a[1651]), .B(n10707), .Z(n10709) );
  XOR U1919 ( .A(a[1654]), .B(n10695), .Z(n10697) );
  XOR U1920 ( .A(a[1657]), .B(n10683), .Z(n10685) );
  XOR U1921 ( .A(a[1660]), .B(n10670), .Z(n10672) );
  XOR U1922 ( .A(a[1663]), .B(n10658), .Z(n10660) );
  XOR U1923 ( .A(a[1666]), .B(n10646), .Z(n10648) );
  XOR U1924 ( .A(a[1669]), .B(n10633), .Z(n10635) );
  XOR U1925 ( .A(a[1672]), .B(n10621), .Z(n10623) );
  XOR U1926 ( .A(a[1675]), .B(n10609), .Z(n10611) );
  XOR U1927 ( .A(a[1678]), .B(n10597), .Z(n10599) );
  XOR U1928 ( .A(a[1681]), .B(n10584), .Z(n10586) );
  XOR U1929 ( .A(a[1684]), .B(n10572), .Z(n10574) );
  XOR U1930 ( .A(a[1687]), .B(n10560), .Z(n10562) );
  XOR U1931 ( .A(a[1690]), .B(n10547), .Z(n10549) );
  XOR U1932 ( .A(a[1693]), .B(n10535), .Z(n10537) );
  XOR U1933 ( .A(a[1696]), .B(n10523), .Z(n10525) );
  XOR U1934 ( .A(a[1699]), .B(n10509), .Z(n10511) );
  XOR U1935 ( .A(a[1702]), .B(n10497), .Z(n10499) );
  XOR U1936 ( .A(a[1705]), .B(n10485), .Z(n10487) );
  XOR U1937 ( .A(a[1708]), .B(n10473), .Z(n10475) );
  XOR U1938 ( .A(a[1711]), .B(n10460), .Z(n10462) );
  XOR U1939 ( .A(a[1714]), .B(n10448), .Z(n10450) );
  XOR U1940 ( .A(a[1717]), .B(n10436), .Z(n10438) );
  XOR U1941 ( .A(a[1720]), .B(n10423), .Z(n10425) );
  XOR U1942 ( .A(a[1723]), .B(n10411), .Z(n10413) );
  XOR U1943 ( .A(a[1726]), .B(n10399), .Z(n10401) );
  XOR U1944 ( .A(a[1729]), .B(n10386), .Z(n10388) );
  XOR U1945 ( .A(a[1732]), .B(n10374), .Z(n10376) );
  XOR U1946 ( .A(a[1735]), .B(n10362), .Z(n10364) );
  XOR U1947 ( .A(a[1738]), .B(n10350), .Z(n10352) );
  XOR U1948 ( .A(a[1741]), .B(n10337), .Z(n10339) );
  XOR U1949 ( .A(a[1744]), .B(n10325), .Z(n10327) );
  XOR U1950 ( .A(a[1747]), .B(n10313), .Z(n10315) );
  XOR U1951 ( .A(a[1750]), .B(n10300), .Z(n10302) );
  XOR U1952 ( .A(a[1753]), .B(n10288), .Z(n10290) );
  XOR U1953 ( .A(a[1756]), .B(n10276), .Z(n10278) );
  XOR U1954 ( .A(a[1759]), .B(n10263), .Z(n10265) );
  XOR U1955 ( .A(a[1762]), .B(n10251), .Z(n10253) );
  XOR U1956 ( .A(a[1765]), .B(n10239), .Z(n10241) );
  XOR U1957 ( .A(a[1768]), .B(n10227), .Z(n10229) );
  XOR U1958 ( .A(a[1771]), .B(n10214), .Z(n10216) );
  XOR U1959 ( .A(a[1774]), .B(n10202), .Z(n10204) );
  XOR U1960 ( .A(a[1777]), .B(n10190), .Z(n10192) );
  XOR U1961 ( .A(a[1780]), .B(n10177), .Z(n10179) );
  XOR U1962 ( .A(a[1783]), .B(n10165), .Z(n10167) );
  XOR U1963 ( .A(a[1786]), .B(n10153), .Z(n10155) );
  XOR U1964 ( .A(a[1789]), .B(n10140), .Z(n10142) );
  XOR U1965 ( .A(a[1792]), .B(n10128), .Z(n10130) );
  XOR U1966 ( .A(a[1795]), .B(n10116), .Z(n10118) );
  XOR U1967 ( .A(a[1798]), .B(n10104), .Z(n10106) );
  XOR U1968 ( .A(a[1801]), .B(n10090), .Z(n10092) );
  XOR U1969 ( .A(a[1804]), .B(n10078), .Z(n10080) );
  XOR U1970 ( .A(a[1807]), .B(n10066), .Z(n10068) );
  XOR U1971 ( .A(a[1810]), .B(n10053), .Z(n10055) );
  XOR U1972 ( .A(a[1813]), .B(n10041), .Z(n10043) );
  XOR U1973 ( .A(a[1816]), .B(n10029), .Z(n10031) );
  XOR U1974 ( .A(a[1819]), .B(n10016), .Z(n10018) );
  XOR U1975 ( .A(a[1822]), .B(n10004), .Z(n10006) );
  XOR U1976 ( .A(a[1825]), .B(n9992), .Z(n9994) );
  XOR U1977 ( .A(a[1828]), .B(n9980), .Z(n9982) );
  XOR U1978 ( .A(a[1831]), .B(n9967), .Z(n9969) );
  XOR U1979 ( .A(a[1834]), .B(n9955), .Z(n9957) );
  XOR U1980 ( .A(a[1837]), .B(n9943), .Z(n9945) );
  XOR U1981 ( .A(a[1840]), .B(n9930), .Z(n9932) );
  XOR U1982 ( .A(a[1843]), .B(n9918), .Z(n9920) );
  XOR U1983 ( .A(a[1846]), .B(n9906), .Z(n9908) );
  XOR U1984 ( .A(a[1849]), .B(n9893), .Z(n9895) );
  XOR U1985 ( .A(a[1852]), .B(n9881), .Z(n9883) );
  XOR U1986 ( .A(a[1855]), .B(n9869), .Z(n9871) );
  XOR U1987 ( .A(a[1858]), .B(n9857), .Z(n9859) );
  XOR U1988 ( .A(a[1861]), .B(n9844), .Z(n9846) );
  XOR U1989 ( .A(a[1864]), .B(n9832), .Z(n9834) );
  XOR U1990 ( .A(a[1867]), .B(n9820), .Z(n9822) );
  XOR U1991 ( .A(a[1870]), .B(n9807), .Z(n9809) );
  XOR U1992 ( .A(a[1873]), .B(n9795), .Z(n9797) );
  XOR U1993 ( .A(a[1876]), .B(n9783), .Z(n9785) );
  XOR U1994 ( .A(a[1879]), .B(n9770), .Z(n9772) );
  XOR U1995 ( .A(a[1882]), .B(n9758), .Z(n9760) );
  XOR U1996 ( .A(a[1885]), .B(n9746), .Z(n9748) );
  XOR U1997 ( .A(a[1888]), .B(n9734), .Z(n9736) );
  XOR U1998 ( .A(a[1891]), .B(n9721), .Z(n9723) );
  XOR U1999 ( .A(a[1894]), .B(n9709), .Z(n9711) );
  XOR U2000 ( .A(a[1897]), .B(n9697), .Z(n9699) );
  XOR U2001 ( .A(a[1900]), .B(n9683), .Z(n9685) );
  XOR U2002 ( .A(a[1903]), .B(n9671), .Z(n9673) );
  XOR U2003 ( .A(a[1906]), .B(n9659), .Z(n9661) );
  XOR U2004 ( .A(a[1909]), .B(n9646), .Z(n9648) );
  XOR U2005 ( .A(a[1912]), .B(n9634), .Z(n9636) );
  XOR U2006 ( .A(a[1915]), .B(n9622), .Z(n9624) );
  XOR U2007 ( .A(a[1918]), .B(n9610), .Z(n9612) );
  XOR U2008 ( .A(a[1921]), .B(n9597), .Z(n9599) );
  XOR U2009 ( .A(a[1924]), .B(n9585), .Z(n9587) );
  XOR U2010 ( .A(a[1927]), .B(n9573), .Z(n9575) );
  XOR U2011 ( .A(a[1930]), .B(n9560), .Z(n9562) );
  XOR U2012 ( .A(a[1933]), .B(n9548), .Z(n9550) );
  XOR U2013 ( .A(a[1936]), .B(n9536), .Z(n9538) );
  XOR U2014 ( .A(a[1939]), .B(n9523), .Z(n9525) );
  XOR U2015 ( .A(a[1942]), .B(n9511), .Z(n9513) );
  XOR U2016 ( .A(a[1945]), .B(n9499), .Z(n9501) );
  XOR U2017 ( .A(a[1948]), .B(n9487), .Z(n9489) );
  XOR U2018 ( .A(a[1951]), .B(n9474), .Z(n9476) );
  XOR U2019 ( .A(a[1954]), .B(n9462), .Z(n9464) );
  XOR U2020 ( .A(a[1957]), .B(n9450), .Z(n9452) );
  XOR U2021 ( .A(a[1960]), .B(n9437), .Z(n9439) );
  XOR U2022 ( .A(a[1963]), .B(n9425), .Z(n9427) );
  XOR U2023 ( .A(a[1966]), .B(n9413), .Z(n9415) );
  XOR U2024 ( .A(a[1969]), .B(n9400), .Z(n9402) );
  XOR U2025 ( .A(a[1972]), .B(n9388), .Z(n9390) );
  XOR U2026 ( .A(a[1975]), .B(n9376), .Z(n9378) );
  XOR U2027 ( .A(a[1978]), .B(n9364), .Z(n9366) );
  XOR U2028 ( .A(a[1981]), .B(n9351), .Z(n9353) );
  XOR U2029 ( .A(a[1984]), .B(n9339), .Z(n9341) );
  XOR U2030 ( .A(a[1987]), .B(n9327), .Z(n9329) );
  XOR U2031 ( .A(a[1990]), .B(n9314), .Z(n9316) );
  XOR U2032 ( .A(a[1993]), .B(n9302), .Z(n9304) );
  XOR U2033 ( .A(a[1996]), .B(n9290), .Z(n9292) );
  XOR U2034 ( .A(a[1999]), .B(n9275), .Z(n9277) );
  XOR U2035 ( .A(a[2002]), .B(n9263), .Z(n9265) );
  XOR U2036 ( .A(a[2005]), .B(n9251), .Z(n9253) );
  XOR U2037 ( .A(a[2008]), .B(n9239), .Z(n9241) );
  XOR U2038 ( .A(a[2011]), .B(n9226), .Z(n9228) );
  XOR U2039 ( .A(a[2014]), .B(n9214), .Z(n9216) );
  XOR U2040 ( .A(a[2017]), .B(n9202), .Z(n9204) );
  XOR U2041 ( .A(a[2020]), .B(n9189), .Z(n9191) );
  XOR U2042 ( .A(a[2023]), .B(n9177), .Z(n9179) );
  XOR U2043 ( .A(a[2026]), .B(n9165), .Z(n9167) );
  XOR U2044 ( .A(a[2029]), .B(n9152), .Z(n9154) );
  XOR U2045 ( .A(a[2032]), .B(n9140), .Z(n9142) );
  XOR U2046 ( .A(a[2035]), .B(n9128), .Z(n9130) );
  XOR U2047 ( .A(a[2038]), .B(n9116), .Z(n9118) );
  XOR U2048 ( .A(a[2041]), .B(n9103), .Z(n9105) );
  XOR U2049 ( .A(a[2044]), .B(n9091), .Z(n9093) );
  XOR U2050 ( .A(a[2047]), .B(n9079), .Z(n9081) );
  XOR U2051 ( .A(a[2050]), .B(n9066), .Z(n9068) );
  XOR U2052 ( .A(a[2053]), .B(n9054), .Z(n9056) );
  XOR U2053 ( .A(a[2056]), .B(n9042), .Z(n9044) );
  XOR U2054 ( .A(a[2059]), .B(n9029), .Z(n9031) );
  XOR U2055 ( .A(a[2062]), .B(n9017), .Z(n9019) );
  XOR U2056 ( .A(a[2065]), .B(n9005), .Z(n9007) );
  XOR U2057 ( .A(a[2068]), .B(n8993), .Z(n8995) );
  XOR U2058 ( .A(a[2071]), .B(n8980), .Z(n8982) );
  XOR U2059 ( .A(a[2074]), .B(n8968), .Z(n8970) );
  XOR U2060 ( .A(a[2077]), .B(n8956), .Z(n8958) );
  XOR U2061 ( .A(a[2080]), .B(n8943), .Z(n8945) );
  XOR U2062 ( .A(a[2083]), .B(n8931), .Z(n8933) );
  XOR U2063 ( .A(a[2086]), .B(n8919), .Z(n8921) );
  XOR U2064 ( .A(a[2089]), .B(n8906), .Z(n8908) );
  XOR U2065 ( .A(a[2092]), .B(n8894), .Z(n8896) );
  XOR U2066 ( .A(a[2095]), .B(n8882), .Z(n8884) );
  XOR U2067 ( .A(a[2098]), .B(n8870), .Z(n8872) );
  XOR U2068 ( .A(a[2101]), .B(n8856), .Z(n8858) );
  XOR U2069 ( .A(a[2104]), .B(n8844), .Z(n8846) );
  XOR U2070 ( .A(a[2107]), .B(n8832), .Z(n8834) );
  XOR U2071 ( .A(a[2110]), .B(n8819), .Z(n8821) );
  XOR U2072 ( .A(a[2113]), .B(n8807), .Z(n8809) );
  XOR U2073 ( .A(a[2116]), .B(n8795), .Z(n8797) );
  XOR U2074 ( .A(a[2119]), .B(n8782), .Z(n8784) );
  XOR U2075 ( .A(a[2122]), .B(n8770), .Z(n8772) );
  XOR U2076 ( .A(a[2125]), .B(n8758), .Z(n8760) );
  XOR U2077 ( .A(a[2128]), .B(n8746), .Z(n8748) );
  XOR U2078 ( .A(a[2131]), .B(n8733), .Z(n8735) );
  XOR U2079 ( .A(a[2134]), .B(n8721), .Z(n8723) );
  XOR U2080 ( .A(a[2137]), .B(n8709), .Z(n8711) );
  XOR U2081 ( .A(a[2140]), .B(n8696), .Z(n8698) );
  XOR U2082 ( .A(a[2143]), .B(n8684), .Z(n8686) );
  XOR U2083 ( .A(a[2146]), .B(n8672), .Z(n8674) );
  XOR U2084 ( .A(a[2149]), .B(n8659), .Z(n8661) );
  XOR U2085 ( .A(a[2152]), .B(n8647), .Z(n8649) );
  XOR U2086 ( .A(a[2155]), .B(n8635), .Z(n8637) );
  XOR U2087 ( .A(a[2158]), .B(n8623), .Z(n8625) );
  XOR U2088 ( .A(a[2161]), .B(n8610), .Z(n8612) );
  XOR U2089 ( .A(a[2164]), .B(n8598), .Z(n8600) );
  XOR U2090 ( .A(a[2167]), .B(n8586), .Z(n8588) );
  XOR U2091 ( .A(a[2170]), .B(n8573), .Z(n8575) );
  XOR U2092 ( .A(a[2173]), .B(n8561), .Z(n8563) );
  XOR U2093 ( .A(a[2176]), .B(n8549), .Z(n8551) );
  XOR U2094 ( .A(a[2179]), .B(n8536), .Z(n8538) );
  XOR U2095 ( .A(a[2182]), .B(n8524), .Z(n8526) );
  XOR U2096 ( .A(a[2185]), .B(n8512), .Z(n8514) );
  XOR U2097 ( .A(a[2188]), .B(n8500), .Z(n8502) );
  XOR U2098 ( .A(a[2191]), .B(n8487), .Z(n8489) );
  XOR U2099 ( .A(a[2194]), .B(n8475), .Z(n8477) );
  XOR U2100 ( .A(a[2197]), .B(n8463), .Z(n8465) );
  XOR U2101 ( .A(a[2200]), .B(n8449), .Z(n8451) );
  XOR U2102 ( .A(a[2203]), .B(n8437), .Z(n8439) );
  XOR U2103 ( .A(a[2206]), .B(n8425), .Z(n8427) );
  XOR U2104 ( .A(a[2209]), .B(n8412), .Z(n8414) );
  XOR U2105 ( .A(a[2212]), .B(n8400), .Z(n8402) );
  XOR U2106 ( .A(a[2215]), .B(n8388), .Z(n8390) );
  XOR U2107 ( .A(a[2218]), .B(n8376), .Z(n8378) );
  XOR U2108 ( .A(a[2221]), .B(n8363), .Z(n8365) );
  XOR U2109 ( .A(a[2224]), .B(n8351), .Z(n8353) );
  XOR U2110 ( .A(a[2227]), .B(n8339), .Z(n8341) );
  XOR U2111 ( .A(a[2230]), .B(n8326), .Z(n8328) );
  XOR U2112 ( .A(a[2233]), .B(n8314), .Z(n8316) );
  XOR U2113 ( .A(a[2236]), .B(n8302), .Z(n8304) );
  XOR U2114 ( .A(a[2239]), .B(n8289), .Z(n8291) );
  XOR U2115 ( .A(a[2242]), .B(n8277), .Z(n8279) );
  XOR U2116 ( .A(a[2245]), .B(n8265), .Z(n8267) );
  XOR U2117 ( .A(a[2248]), .B(n8253), .Z(n8255) );
  XOR U2118 ( .A(a[2251]), .B(n8240), .Z(n8242) );
  XOR U2119 ( .A(a[2254]), .B(n8228), .Z(n8230) );
  XOR U2120 ( .A(a[2257]), .B(n8216), .Z(n8218) );
  XOR U2121 ( .A(a[2260]), .B(n8203), .Z(n8205) );
  XOR U2122 ( .A(a[2263]), .B(n8191), .Z(n8193) );
  XOR U2123 ( .A(a[2266]), .B(n8179), .Z(n8181) );
  XOR U2124 ( .A(a[2269]), .B(n8166), .Z(n8168) );
  XOR U2125 ( .A(a[2272]), .B(n8154), .Z(n8156) );
  XOR U2126 ( .A(a[2275]), .B(n8142), .Z(n8144) );
  XOR U2127 ( .A(a[2278]), .B(n8130), .Z(n8132) );
  XOR U2128 ( .A(a[2281]), .B(n8117), .Z(n8119) );
  XOR U2129 ( .A(a[2284]), .B(n8105), .Z(n8107) );
  XOR U2130 ( .A(a[2287]), .B(n8093), .Z(n8095) );
  XOR U2131 ( .A(a[2290]), .B(n8080), .Z(n8082) );
  XOR U2132 ( .A(a[2293]), .B(n8068), .Z(n8070) );
  XOR U2133 ( .A(a[2296]), .B(n8056), .Z(n8058) );
  XOR U2134 ( .A(a[2299]), .B(n8042), .Z(n8044) );
  XOR U2135 ( .A(a[2302]), .B(n8030), .Z(n8032) );
  XOR U2136 ( .A(a[2305]), .B(n8018), .Z(n8020) );
  XOR U2137 ( .A(a[2308]), .B(n8006), .Z(n8008) );
  XOR U2138 ( .A(a[2311]), .B(n7993), .Z(n7995) );
  XOR U2139 ( .A(a[2314]), .B(n7981), .Z(n7983) );
  XOR U2140 ( .A(a[2317]), .B(n7969), .Z(n7971) );
  XOR U2141 ( .A(a[2320]), .B(n7956), .Z(n7958) );
  XOR U2142 ( .A(a[2323]), .B(n7944), .Z(n7946) );
  XOR U2143 ( .A(a[2326]), .B(n7932), .Z(n7934) );
  XOR U2144 ( .A(a[2329]), .B(n7919), .Z(n7921) );
  XOR U2145 ( .A(a[2332]), .B(n7907), .Z(n7909) );
  XOR U2146 ( .A(a[2335]), .B(n7895), .Z(n7897) );
  XOR U2147 ( .A(a[2338]), .B(n7883), .Z(n7885) );
  XOR U2148 ( .A(a[2341]), .B(n7870), .Z(n7872) );
  XOR U2149 ( .A(a[2344]), .B(n7858), .Z(n7860) );
  XOR U2150 ( .A(a[2347]), .B(n7846), .Z(n7848) );
  XOR U2151 ( .A(a[2350]), .B(n7833), .Z(n7835) );
  XOR U2152 ( .A(a[2353]), .B(n7821), .Z(n7823) );
  XOR U2153 ( .A(a[2356]), .B(n7809), .Z(n7811) );
  XOR U2154 ( .A(a[2359]), .B(n7796), .Z(n7798) );
  XOR U2155 ( .A(a[2362]), .B(n7784), .Z(n7786) );
  XOR U2156 ( .A(a[2365]), .B(n7772), .Z(n7774) );
  XOR U2157 ( .A(a[2368]), .B(n7760), .Z(n7762) );
  XOR U2158 ( .A(a[2371]), .B(n7747), .Z(n7749) );
  XOR U2159 ( .A(a[2374]), .B(n7735), .Z(n7737) );
  XOR U2160 ( .A(a[2377]), .B(n7723), .Z(n7725) );
  XOR U2161 ( .A(a[2380]), .B(n7710), .Z(n7712) );
  XOR U2162 ( .A(a[2383]), .B(n7698), .Z(n7700) );
  XOR U2163 ( .A(a[2386]), .B(n7686), .Z(n7688) );
  XOR U2164 ( .A(a[2389]), .B(n7673), .Z(n7675) );
  XOR U2165 ( .A(a[2392]), .B(n7661), .Z(n7663) );
  XOR U2166 ( .A(a[2395]), .B(n7649), .Z(n7651) );
  XOR U2167 ( .A(a[2398]), .B(n7637), .Z(n7639) );
  XOR U2168 ( .A(a[2401]), .B(n7623), .Z(n7625) );
  XOR U2169 ( .A(a[2404]), .B(n7611), .Z(n7613) );
  XOR U2170 ( .A(a[2407]), .B(n7599), .Z(n7601) );
  XOR U2171 ( .A(a[2410]), .B(n7586), .Z(n7588) );
  XOR U2172 ( .A(a[2413]), .B(n7574), .Z(n7576) );
  XOR U2173 ( .A(a[2416]), .B(n7562), .Z(n7564) );
  XOR U2174 ( .A(a[2419]), .B(n7549), .Z(n7551) );
  XOR U2175 ( .A(a[2422]), .B(n7537), .Z(n7539) );
  XOR U2176 ( .A(a[2425]), .B(n7525), .Z(n7527) );
  XOR U2177 ( .A(a[2428]), .B(n7513), .Z(n7515) );
  XOR U2178 ( .A(a[2431]), .B(n7500), .Z(n7502) );
  XOR U2179 ( .A(a[2434]), .B(n7488), .Z(n7490) );
  XOR U2180 ( .A(a[2437]), .B(n7476), .Z(n7478) );
  XOR U2181 ( .A(a[2440]), .B(n7463), .Z(n7465) );
  XOR U2182 ( .A(a[2443]), .B(n7451), .Z(n7453) );
  XOR U2183 ( .A(a[2446]), .B(n7439), .Z(n7441) );
  XOR U2184 ( .A(a[2449]), .B(n7426), .Z(n7428) );
  XOR U2185 ( .A(a[2452]), .B(n7414), .Z(n7416) );
  XOR U2186 ( .A(a[2455]), .B(n7402), .Z(n7404) );
  XOR U2187 ( .A(a[2458]), .B(n7390), .Z(n7392) );
  XOR U2188 ( .A(a[2461]), .B(n7377), .Z(n7379) );
  XOR U2189 ( .A(a[2464]), .B(n7365), .Z(n7367) );
  XOR U2190 ( .A(a[2467]), .B(n7353), .Z(n7355) );
  XOR U2191 ( .A(a[2470]), .B(n7340), .Z(n7342) );
  XOR U2192 ( .A(a[2473]), .B(n7328), .Z(n7330) );
  XOR U2193 ( .A(a[2476]), .B(n7316), .Z(n7318) );
  XOR U2194 ( .A(a[2479]), .B(n7303), .Z(n7305) );
  XOR U2195 ( .A(a[2482]), .B(n7291), .Z(n7293) );
  XOR U2196 ( .A(a[2485]), .B(n7279), .Z(n7281) );
  XOR U2197 ( .A(a[2488]), .B(n7267), .Z(n7269) );
  XOR U2198 ( .A(a[2491]), .B(n7254), .Z(n7256) );
  XOR U2199 ( .A(a[2494]), .B(n7242), .Z(n7244) );
  XOR U2200 ( .A(a[2497]), .B(n7230), .Z(n7232) );
  XOR U2201 ( .A(a[2500]), .B(n7216), .Z(n7218) );
  XOR U2202 ( .A(a[2503]), .B(n7204), .Z(n7206) );
  XOR U2203 ( .A(a[2506]), .B(n7192), .Z(n7194) );
  XOR U2204 ( .A(a[2509]), .B(n7179), .Z(n7181) );
  XOR U2205 ( .A(a[2512]), .B(n7167), .Z(n7169) );
  XOR U2206 ( .A(a[2515]), .B(n7155), .Z(n7157) );
  XOR U2207 ( .A(a[2518]), .B(n7143), .Z(n7145) );
  XOR U2208 ( .A(a[2521]), .B(n7130), .Z(n7132) );
  XOR U2209 ( .A(a[2524]), .B(n7118), .Z(n7120) );
  XOR U2210 ( .A(a[2527]), .B(n7106), .Z(n7108) );
  XOR U2211 ( .A(a[2530]), .B(n7093), .Z(n7095) );
  XOR U2212 ( .A(a[2533]), .B(n7081), .Z(n7083) );
  XOR U2213 ( .A(a[2536]), .B(n7069), .Z(n7071) );
  XOR U2214 ( .A(a[2539]), .B(n7056), .Z(n7058) );
  XOR U2215 ( .A(a[2542]), .B(n7044), .Z(n7046) );
  XOR U2216 ( .A(a[2545]), .B(n7032), .Z(n7034) );
  XOR U2217 ( .A(a[2548]), .B(n7020), .Z(n7022) );
  XOR U2218 ( .A(a[2551]), .B(n7007), .Z(n7009) );
  XOR U2219 ( .A(a[2554]), .B(n6995), .Z(n6997) );
  XOR U2220 ( .A(a[2557]), .B(n6983), .Z(n6985) );
  XOR U2221 ( .A(a[2560]), .B(n6970), .Z(n6972) );
  XOR U2222 ( .A(a[2563]), .B(n6958), .Z(n6960) );
  XOR U2223 ( .A(a[2566]), .B(n6946), .Z(n6948) );
  XOR U2224 ( .A(a[2569]), .B(n6933), .Z(n6935) );
  XOR U2225 ( .A(a[2572]), .B(n6921), .Z(n6923) );
  XOR U2226 ( .A(a[2575]), .B(n6909), .Z(n6911) );
  XOR U2227 ( .A(a[2578]), .B(n6897), .Z(n6899) );
  XOR U2228 ( .A(a[2581]), .B(n6884), .Z(n6886) );
  XOR U2229 ( .A(a[2584]), .B(n6872), .Z(n6874) );
  XOR U2230 ( .A(a[2587]), .B(n6860), .Z(n6862) );
  XOR U2231 ( .A(a[2590]), .B(n6847), .Z(n6849) );
  XOR U2232 ( .A(a[2593]), .B(n6835), .Z(n6837) );
  XOR U2233 ( .A(a[2596]), .B(n6823), .Z(n6825) );
  XOR U2234 ( .A(a[2599]), .B(n6809), .Z(n6811) );
  XOR U2235 ( .A(a[2602]), .B(n6797), .Z(n6799) );
  XOR U2236 ( .A(a[2605]), .B(n6785), .Z(n6787) );
  XOR U2237 ( .A(a[2608]), .B(n6773), .Z(n6775) );
  XOR U2238 ( .A(a[2611]), .B(n6760), .Z(n6762) );
  XOR U2239 ( .A(a[2614]), .B(n6748), .Z(n6750) );
  XOR U2240 ( .A(a[2617]), .B(n6736), .Z(n6738) );
  XOR U2241 ( .A(a[2620]), .B(n6723), .Z(n6725) );
  XOR U2242 ( .A(a[2623]), .B(n6711), .Z(n6713) );
  XOR U2243 ( .A(a[2626]), .B(n6699), .Z(n6701) );
  XOR U2244 ( .A(a[2629]), .B(n6686), .Z(n6688) );
  XOR U2245 ( .A(a[2632]), .B(n6674), .Z(n6676) );
  XOR U2246 ( .A(a[2635]), .B(n6662), .Z(n6664) );
  XOR U2247 ( .A(a[2638]), .B(n6650), .Z(n6652) );
  XOR U2248 ( .A(a[2641]), .B(n6637), .Z(n6639) );
  XOR U2249 ( .A(a[2644]), .B(n6625), .Z(n6627) );
  XOR U2250 ( .A(a[2647]), .B(n6613), .Z(n6615) );
  XOR U2251 ( .A(a[2650]), .B(n6600), .Z(n6602) );
  XOR U2252 ( .A(a[2653]), .B(n6588), .Z(n6590) );
  XOR U2253 ( .A(a[2656]), .B(n6576), .Z(n6578) );
  XOR U2254 ( .A(a[2659]), .B(n6563), .Z(n6565) );
  XOR U2255 ( .A(a[2662]), .B(n6551), .Z(n6553) );
  XOR U2256 ( .A(a[2665]), .B(n6539), .Z(n6541) );
  XOR U2257 ( .A(a[2668]), .B(n6527), .Z(n6529) );
  XOR U2258 ( .A(a[2671]), .B(n6514), .Z(n6516) );
  XOR U2259 ( .A(a[2674]), .B(n6502), .Z(n6504) );
  XOR U2260 ( .A(a[2677]), .B(n6490), .Z(n6492) );
  XOR U2261 ( .A(a[2680]), .B(n6477), .Z(n6479) );
  XOR U2262 ( .A(a[2683]), .B(n6465), .Z(n6467) );
  XOR U2263 ( .A(a[2686]), .B(n6453), .Z(n6455) );
  XOR U2264 ( .A(a[2689]), .B(n6440), .Z(n6442) );
  XOR U2265 ( .A(a[2692]), .B(n6428), .Z(n6430) );
  XOR U2266 ( .A(a[2695]), .B(n6416), .Z(n6418) );
  XOR U2267 ( .A(a[2698]), .B(n6404), .Z(n6406) );
  XOR U2268 ( .A(a[2701]), .B(n6390), .Z(n6392) );
  XOR U2269 ( .A(a[2704]), .B(n6378), .Z(n6380) );
  XOR U2270 ( .A(a[2707]), .B(n6366), .Z(n6368) );
  XOR U2271 ( .A(a[2710]), .B(n6353), .Z(n6355) );
  XOR U2272 ( .A(a[2713]), .B(n6341), .Z(n6343) );
  XOR U2273 ( .A(a[2716]), .B(n6329), .Z(n6331) );
  XOR U2274 ( .A(a[2719]), .B(n6316), .Z(n6318) );
  XOR U2275 ( .A(a[2722]), .B(n6304), .Z(n6306) );
  XOR U2276 ( .A(a[2725]), .B(n6292), .Z(n6294) );
  XOR U2277 ( .A(a[2728]), .B(n6280), .Z(n6282) );
  XOR U2278 ( .A(a[2731]), .B(n6267), .Z(n6269) );
  XOR U2279 ( .A(a[2734]), .B(n6255), .Z(n6257) );
  XOR U2280 ( .A(a[2737]), .B(n6243), .Z(n6245) );
  XOR U2281 ( .A(a[2740]), .B(n6230), .Z(n6232) );
  XOR U2282 ( .A(a[2743]), .B(n6218), .Z(n6220) );
  XOR U2283 ( .A(a[2746]), .B(n6206), .Z(n6208) );
  XOR U2284 ( .A(a[2749]), .B(n6193), .Z(n6195) );
  XOR U2285 ( .A(a[2752]), .B(n6181), .Z(n6183) );
  XOR U2286 ( .A(a[2755]), .B(n6169), .Z(n6171) );
  XOR U2287 ( .A(a[2758]), .B(n6157), .Z(n6159) );
  XOR U2288 ( .A(a[2761]), .B(n6144), .Z(n6146) );
  XOR U2289 ( .A(a[2764]), .B(n6132), .Z(n6134) );
  XOR U2290 ( .A(a[2767]), .B(n6120), .Z(n6122) );
  XOR U2291 ( .A(a[2770]), .B(n6107), .Z(n6109) );
  XOR U2292 ( .A(a[2773]), .B(n6095), .Z(n6097) );
  XOR U2293 ( .A(a[2776]), .B(n6083), .Z(n6085) );
  XOR U2294 ( .A(a[2779]), .B(n6070), .Z(n6072) );
  XOR U2295 ( .A(a[2782]), .B(n6058), .Z(n6060) );
  XOR U2296 ( .A(a[2785]), .B(n6046), .Z(n6048) );
  XOR U2297 ( .A(a[2788]), .B(n6034), .Z(n6036) );
  XOR U2298 ( .A(a[2791]), .B(n6021), .Z(n6023) );
  XOR U2299 ( .A(a[2794]), .B(n6009), .Z(n6011) );
  XOR U2300 ( .A(a[2797]), .B(n5997), .Z(n5999) );
  XOR U2301 ( .A(a[2800]), .B(n5983), .Z(n5985) );
  XOR U2302 ( .A(a[2803]), .B(n5971), .Z(n5973) );
  XOR U2303 ( .A(a[2806]), .B(n5959), .Z(n5961) );
  XOR U2304 ( .A(a[2809]), .B(n5946), .Z(n5948) );
  XOR U2305 ( .A(a[2812]), .B(n5934), .Z(n5936) );
  XOR U2306 ( .A(a[2815]), .B(n5922), .Z(n5924) );
  XOR U2307 ( .A(a[2818]), .B(n5910), .Z(n5912) );
  XOR U2308 ( .A(a[2821]), .B(n5897), .Z(n5899) );
  XOR U2309 ( .A(a[2824]), .B(n5885), .Z(n5887) );
  XOR U2310 ( .A(a[2827]), .B(n5873), .Z(n5875) );
  XOR U2311 ( .A(a[2830]), .B(n5860), .Z(n5862) );
  XOR U2312 ( .A(a[2833]), .B(n5848), .Z(n5850) );
  XOR U2313 ( .A(a[2836]), .B(n5836), .Z(n5838) );
  XOR U2314 ( .A(a[2839]), .B(n5823), .Z(n5825) );
  XOR U2315 ( .A(a[2842]), .B(n5811), .Z(n5813) );
  XOR U2316 ( .A(a[2845]), .B(n5799), .Z(n5801) );
  XOR U2317 ( .A(a[2848]), .B(n5787), .Z(n5789) );
  XOR U2318 ( .A(a[2851]), .B(n5774), .Z(n5776) );
  XOR U2319 ( .A(a[2854]), .B(n5762), .Z(n5764) );
  XOR U2320 ( .A(a[2857]), .B(n5750), .Z(n5752) );
  XOR U2321 ( .A(a[2860]), .B(n5737), .Z(n5739) );
  XOR U2322 ( .A(a[2863]), .B(n5725), .Z(n5727) );
  XOR U2323 ( .A(a[2866]), .B(n5713), .Z(n5715) );
  XOR U2324 ( .A(a[2869]), .B(n5700), .Z(n5702) );
  XOR U2325 ( .A(a[2872]), .B(n5688), .Z(n5690) );
  XOR U2326 ( .A(a[2875]), .B(n5676), .Z(n5678) );
  XOR U2327 ( .A(a[2878]), .B(n5664), .Z(n5666) );
  XOR U2328 ( .A(a[2881]), .B(n5651), .Z(n5653) );
  XOR U2329 ( .A(a[2884]), .B(n5639), .Z(n5641) );
  XOR U2330 ( .A(a[2887]), .B(n5627), .Z(n5629) );
  XOR U2331 ( .A(a[2890]), .B(n5614), .Z(n5616) );
  XOR U2332 ( .A(a[2893]), .B(n5602), .Z(n5604) );
  XOR U2333 ( .A(a[2896]), .B(n5590), .Z(n5592) );
  XOR U2334 ( .A(a[2899]), .B(n5576), .Z(n5578) );
  XOR U2335 ( .A(a[2902]), .B(n5564), .Z(n5566) );
  XOR U2336 ( .A(a[2905]), .B(n5552), .Z(n5554) );
  XOR U2337 ( .A(a[2908]), .B(n5540), .Z(n5542) );
  XOR U2338 ( .A(a[2911]), .B(n5527), .Z(n5529) );
  XOR U2339 ( .A(a[2914]), .B(n5515), .Z(n5517) );
  XOR U2340 ( .A(a[2917]), .B(n5503), .Z(n5505) );
  XOR U2341 ( .A(a[2920]), .B(n5490), .Z(n5492) );
  XOR U2342 ( .A(a[2923]), .B(n5478), .Z(n5480) );
  XOR U2343 ( .A(a[2926]), .B(n5466), .Z(n5468) );
  XOR U2344 ( .A(a[2929]), .B(n5453), .Z(n5455) );
  XOR U2345 ( .A(a[2932]), .B(n5441), .Z(n5443) );
  XOR U2346 ( .A(a[2935]), .B(n5429), .Z(n5431) );
  XOR U2347 ( .A(a[2938]), .B(n5417), .Z(n5419) );
  XOR U2348 ( .A(a[2941]), .B(n5404), .Z(n5406) );
  XOR U2349 ( .A(a[2944]), .B(n5392), .Z(n5394) );
  XOR U2350 ( .A(a[2947]), .B(n5380), .Z(n5382) );
  XOR U2351 ( .A(a[2950]), .B(n5367), .Z(n5369) );
  XOR U2352 ( .A(a[2953]), .B(n5355), .Z(n5357) );
  XOR U2353 ( .A(a[2956]), .B(n5343), .Z(n5345) );
  XOR U2354 ( .A(a[2959]), .B(n5330), .Z(n5332) );
  XOR U2355 ( .A(a[2962]), .B(n5318), .Z(n5320) );
  XOR U2356 ( .A(a[2965]), .B(n5306), .Z(n5308) );
  XOR U2357 ( .A(a[2968]), .B(n5294), .Z(n5296) );
  XOR U2358 ( .A(a[2971]), .B(n5281), .Z(n5283) );
  XOR U2359 ( .A(a[2974]), .B(n5269), .Z(n5271) );
  XOR U2360 ( .A(a[2977]), .B(n5257), .Z(n5259) );
  XOR U2361 ( .A(a[2980]), .B(n5244), .Z(n5246) );
  XOR U2362 ( .A(a[2983]), .B(n5232), .Z(n5234) );
  XOR U2363 ( .A(a[2986]), .B(n5220), .Z(n5222) );
  XOR U2364 ( .A(a[2989]), .B(n5207), .Z(n5209) );
  XOR U2365 ( .A(a[2992]), .B(n5195), .Z(n5197) );
  XOR U2366 ( .A(a[2995]), .B(n5183), .Z(n5185) );
  XOR U2367 ( .A(a[2998]), .B(n5171), .Z(n5173) );
  XOR U2368 ( .A(a[3001]), .B(n5156), .Z(n5158) );
  XOR U2369 ( .A(a[3004]), .B(n5144), .Z(n5146) );
  XOR U2370 ( .A(a[3007]), .B(n5132), .Z(n5134) );
  XOR U2371 ( .A(a[3010]), .B(n5119), .Z(n5121) );
  XOR U2372 ( .A(a[3013]), .B(n5107), .Z(n5109) );
  XOR U2373 ( .A(a[3016]), .B(n5095), .Z(n5097) );
  XOR U2374 ( .A(a[3019]), .B(n5082), .Z(n5084) );
  XOR U2375 ( .A(a[3022]), .B(n5070), .Z(n5072) );
  XOR U2376 ( .A(a[3025]), .B(n5058), .Z(n5060) );
  XOR U2377 ( .A(a[3028]), .B(n5046), .Z(n5048) );
  XOR U2378 ( .A(a[3031]), .B(n5033), .Z(n5035) );
  XOR U2379 ( .A(a[3034]), .B(n5021), .Z(n5023) );
  XOR U2380 ( .A(a[3037]), .B(n5009), .Z(n5011) );
  XOR U2381 ( .A(a[3040]), .B(n4996), .Z(n4998) );
  XOR U2382 ( .A(a[3043]), .B(n4984), .Z(n4986) );
  XOR U2383 ( .A(a[3046]), .B(n4972), .Z(n4974) );
  XOR U2384 ( .A(a[3049]), .B(n4959), .Z(n4961) );
  XOR U2385 ( .A(a[3052]), .B(n4947), .Z(n4949) );
  XOR U2386 ( .A(a[3055]), .B(n4935), .Z(n4937) );
  XOR U2387 ( .A(a[3058]), .B(n4923), .Z(n4925) );
  XOR U2388 ( .A(a[3061]), .B(n4910), .Z(n4912) );
  XOR U2389 ( .A(a[3064]), .B(n4898), .Z(n4900) );
  XOR U2390 ( .A(a[3067]), .B(n4886), .Z(n4888) );
  XOR U2391 ( .A(a[3070]), .B(n4873), .Z(n4875) );
  XOR U2392 ( .A(a[3073]), .B(n4861), .Z(n4863) );
  XOR U2393 ( .A(a[3076]), .B(n4849), .Z(n4851) );
  XOR U2394 ( .A(a[3079]), .B(n4836), .Z(n4838) );
  XOR U2395 ( .A(a[3082]), .B(n4824), .Z(n4826) );
  XOR U2396 ( .A(a[3085]), .B(n4812), .Z(n4814) );
  XOR U2397 ( .A(a[3088]), .B(n4800), .Z(n4802) );
  XOR U2398 ( .A(a[3091]), .B(n4787), .Z(n4789) );
  XOR U2399 ( .A(a[3094]), .B(n4775), .Z(n4777) );
  XOR U2400 ( .A(a[3097]), .B(n4763), .Z(n4765) );
  XOR U2401 ( .A(a[3100]), .B(n4749), .Z(n4751) );
  XOR U2402 ( .A(a[3103]), .B(n4737), .Z(n4739) );
  XOR U2403 ( .A(a[3106]), .B(n4725), .Z(n4727) );
  XOR U2404 ( .A(a[3109]), .B(n4712), .Z(n4714) );
  XOR U2405 ( .A(a[3112]), .B(n4700), .Z(n4702) );
  XOR U2406 ( .A(a[3115]), .B(n4688), .Z(n4690) );
  XOR U2407 ( .A(a[3118]), .B(n4676), .Z(n4678) );
  XOR U2408 ( .A(a[3121]), .B(n4663), .Z(n4665) );
  XOR U2409 ( .A(a[3124]), .B(n4651), .Z(n4653) );
  XOR U2410 ( .A(a[3127]), .B(n4639), .Z(n4641) );
  XOR U2411 ( .A(a[3130]), .B(n4626), .Z(n4628) );
  XOR U2412 ( .A(a[3133]), .B(n4614), .Z(n4616) );
  XOR U2413 ( .A(a[3136]), .B(n4602), .Z(n4604) );
  XOR U2414 ( .A(a[3139]), .B(n4589), .Z(n4591) );
  XOR U2415 ( .A(a[3142]), .B(n4577), .Z(n4579) );
  XOR U2416 ( .A(a[3145]), .B(n4565), .Z(n4567) );
  XOR U2417 ( .A(a[3148]), .B(n4553), .Z(n4555) );
  XOR U2418 ( .A(a[3151]), .B(n4540), .Z(n4542) );
  XOR U2419 ( .A(a[3154]), .B(n4528), .Z(n4530) );
  XOR U2420 ( .A(a[3157]), .B(n4516), .Z(n4518) );
  XOR U2421 ( .A(a[3160]), .B(n4503), .Z(n4505) );
  XOR U2422 ( .A(a[3163]), .B(n4491), .Z(n4493) );
  XOR U2423 ( .A(a[3166]), .B(n4479), .Z(n4481) );
  XOR U2424 ( .A(a[3169]), .B(n4466), .Z(n4468) );
  XOR U2425 ( .A(a[3172]), .B(n4454), .Z(n4456) );
  XOR U2426 ( .A(a[3175]), .B(n4442), .Z(n4444) );
  XOR U2427 ( .A(a[3178]), .B(n4430), .Z(n4432) );
  XOR U2428 ( .A(a[3181]), .B(n4417), .Z(n4419) );
  XOR U2429 ( .A(a[3184]), .B(n4405), .Z(n4407) );
  XOR U2430 ( .A(a[3187]), .B(n4393), .Z(n4395) );
  XOR U2431 ( .A(a[3190]), .B(n4380), .Z(n4382) );
  XOR U2432 ( .A(a[3193]), .B(n4368), .Z(n4370) );
  XOR U2433 ( .A(a[3196]), .B(n4356), .Z(n4358) );
  XOR U2434 ( .A(a[3199]), .B(n4342), .Z(n4344) );
  XOR U2435 ( .A(a[3202]), .B(n4330), .Z(n4332) );
  XOR U2436 ( .A(a[3205]), .B(n4318), .Z(n4320) );
  XOR U2437 ( .A(a[3208]), .B(n4306), .Z(n4308) );
  XOR U2438 ( .A(a[3211]), .B(n4293), .Z(n4295) );
  XOR U2439 ( .A(a[3214]), .B(n4281), .Z(n4283) );
  XOR U2440 ( .A(a[3217]), .B(n4269), .Z(n4271) );
  XOR U2441 ( .A(a[3220]), .B(n4256), .Z(n4258) );
  XOR U2442 ( .A(a[3223]), .B(n4244), .Z(n4246) );
  XOR U2443 ( .A(a[3226]), .B(n4232), .Z(n4234) );
  XOR U2444 ( .A(a[3229]), .B(n4219), .Z(n4221) );
  XOR U2445 ( .A(a[3232]), .B(n4207), .Z(n4209) );
  XOR U2446 ( .A(a[3235]), .B(n4195), .Z(n4197) );
  XOR U2447 ( .A(a[3238]), .B(n4183), .Z(n4185) );
  XOR U2448 ( .A(a[3241]), .B(n4170), .Z(n4172) );
  XOR U2449 ( .A(a[3244]), .B(n4158), .Z(n4160) );
  XOR U2450 ( .A(a[3247]), .B(n4146), .Z(n4148) );
  XOR U2451 ( .A(a[3250]), .B(n4133), .Z(n4135) );
  XOR U2452 ( .A(a[3253]), .B(n4121), .Z(n4123) );
  XOR U2453 ( .A(a[3256]), .B(n4109), .Z(n4111) );
  XOR U2454 ( .A(a[3259]), .B(n4096), .Z(n4098) );
  XOR U2455 ( .A(a[3262]), .B(n4084), .Z(n4086) );
  XOR U2456 ( .A(a[3265]), .B(n4072), .Z(n4074) );
  XOR U2457 ( .A(a[3268]), .B(n4060), .Z(n4062) );
  XOR U2458 ( .A(a[3271]), .B(n4047), .Z(n4049) );
  XOR U2459 ( .A(a[3274]), .B(n4035), .Z(n4037) );
  XOR U2460 ( .A(a[3277]), .B(n4023), .Z(n4025) );
  XOR U2461 ( .A(a[3280]), .B(n4010), .Z(n4012) );
  XOR U2462 ( .A(a[3283]), .B(n3998), .Z(n4000) );
  XOR U2463 ( .A(a[3286]), .B(n3986), .Z(n3988) );
  XOR U2464 ( .A(a[3289]), .B(n3973), .Z(n3975) );
  XOR U2465 ( .A(a[3292]), .B(n3961), .Z(n3963) );
  XOR U2466 ( .A(a[3295]), .B(n3949), .Z(n3951) );
  XOR U2467 ( .A(a[3298]), .B(n3937), .Z(n3939) );
  XOR U2468 ( .A(a[3301]), .B(n3923), .Z(n3925) );
  XOR U2469 ( .A(a[3304]), .B(n3911), .Z(n3913) );
  XOR U2470 ( .A(a[3307]), .B(n3899), .Z(n3901) );
  XOR U2471 ( .A(a[3310]), .B(n3886), .Z(n3888) );
  XOR U2472 ( .A(a[3313]), .B(n3874), .Z(n3876) );
  XOR U2473 ( .A(a[3316]), .B(n3862), .Z(n3864) );
  XOR U2474 ( .A(a[3319]), .B(n3849), .Z(n3851) );
  XOR U2475 ( .A(a[3322]), .B(n3837), .Z(n3839) );
  XOR U2476 ( .A(a[3325]), .B(n3825), .Z(n3827) );
  XOR U2477 ( .A(a[3328]), .B(n3813), .Z(n3815) );
  XOR U2478 ( .A(a[3331]), .B(n3800), .Z(n3802) );
  XOR U2479 ( .A(a[3334]), .B(n3788), .Z(n3790) );
  XOR U2480 ( .A(a[3337]), .B(n3776), .Z(n3778) );
  XOR U2481 ( .A(a[3340]), .B(n3763), .Z(n3765) );
  XOR U2482 ( .A(a[3343]), .B(n3751), .Z(n3753) );
  XOR U2483 ( .A(a[3346]), .B(n3739), .Z(n3741) );
  XOR U2484 ( .A(a[3349]), .B(n3726), .Z(n3728) );
  XOR U2485 ( .A(a[3352]), .B(n3714), .Z(n3716) );
  XOR U2486 ( .A(a[3355]), .B(n3702), .Z(n3704) );
  XOR U2487 ( .A(a[3358]), .B(n3690), .Z(n3692) );
  XOR U2488 ( .A(a[3361]), .B(n3677), .Z(n3679) );
  XOR U2489 ( .A(a[3364]), .B(n3665), .Z(n3667) );
  XOR U2490 ( .A(a[3367]), .B(n3653), .Z(n3655) );
  XOR U2491 ( .A(a[3370]), .B(n3640), .Z(n3642) );
  XOR U2492 ( .A(a[3373]), .B(n3628), .Z(n3630) );
  XOR U2493 ( .A(a[3376]), .B(n3616), .Z(n3618) );
  XOR U2494 ( .A(a[3379]), .B(n3603), .Z(n3605) );
  XOR U2495 ( .A(a[3382]), .B(n3591), .Z(n3593) );
  XOR U2496 ( .A(a[3385]), .B(n3579), .Z(n3581) );
  XOR U2497 ( .A(a[3388]), .B(n3567), .Z(n3569) );
  XOR U2498 ( .A(a[3391]), .B(n3554), .Z(n3556) );
  XOR U2499 ( .A(a[3394]), .B(n3542), .Z(n3544) );
  XOR U2500 ( .A(a[3397]), .B(n3530), .Z(n3532) );
  XOR U2501 ( .A(a[3400]), .B(n3516), .Z(n3518) );
  XOR U2502 ( .A(a[3403]), .B(n3504), .Z(n3506) );
  XOR U2503 ( .A(a[3406]), .B(n3492), .Z(n3494) );
  XOR U2504 ( .A(a[3409]), .B(n3479), .Z(n3481) );
  XOR U2505 ( .A(a[3412]), .B(n3467), .Z(n3469) );
  XOR U2506 ( .A(a[3415]), .B(n3455), .Z(n3457) );
  XOR U2507 ( .A(a[3418]), .B(n3443), .Z(n3445) );
  XOR U2508 ( .A(a[3421]), .B(n3430), .Z(n3432) );
  XOR U2509 ( .A(a[3424]), .B(n3418), .Z(n3420) );
  XOR U2510 ( .A(a[3427]), .B(n3406), .Z(n3408) );
  XOR U2511 ( .A(a[3430]), .B(n3393), .Z(n3395) );
  XOR U2512 ( .A(a[3433]), .B(n3381), .Z(n3383) );
  XOR U2513 ( .A(a[3436]), .B(n3369), .Z(n3371) );
  XOR U2514 ( .A(a[3439]), .B(n3356), .Z(n3358) );
  XOR U2515 ( .A(a[3442]), .B(n3344), .Z(n3346) );
  XOR U2516 ( .A(a[3445]), .B(n3332), .Z(n3334) );
  XOR U2517 ( .A(a[3448]), .B(n3320), .Z(n3322) );
  XOR U2518 ( .A(a[3451]), .B(n3307), .Z(n3309) );
  XOR U2519 ( .A(a[3454]), .B(n3295), .Z(n3297) );
  XOR U2520 ( .A(a[3457]), .B(n3283), .Z(n3285) );
  XOR U2521 ( .A(a[3460]), .B(n3270), .Z(n3272) );
  XOR U2522 ( .A(a[3463]), .B(n3258), .Z(n3260) );
  XOR U2523 ( .A(a[3466]), .B(n3246), .Z(n3248) );
  XOR U2524 ( .A(a[3469]), .B(n3233), .Z(n3235) );
  XOR U2525 ( .A(a[3472]), .B(n3221), .Z(n3223) );
  XOR U2526 ( .A(a[3475]), .B(n3209), .Z(n3211) );
  XOR U2527 ( .A(a[3478]), .B(n3197), .Z(n3199) );
  XOR U2528 ( .A(a[3481]), .B(n3184), .Z(n3186) );
  XOR U2529 ( .A(a[3484]), .B(n3172), .Z(n3174) );
  XOR U2530 ( .A(a[3487]), .B(n3160), .Z(n3162) );
  XOR U2531 ( .A(a[3490]), .B(n3147), .Z(n3149) );
  XOR U2532 ( .A(a[3493]), .B(n3135), .Z(n3137) );
  XOR U2533 ( .A(a[3496]), .B(n3123), .Z(n3125) );
  XOR U2534 ( .A(a[3499]), .B(n3109), .Z(n3111) );
  XOR U2535 ( .A(a[3502]), .B(n3097), .Z(n3099) );
  XOR U2536 ( .A(a[3505]), .B(n3085), .Z(n3087) );
  XOR U2537 ( .A(a[3508]), .B(n3073), .Z(n3075) );
  XOR U2538 ( .A(a[3511]), .B(n3060), .Z(n3062) );
  XOR U2539 ( .A(a[3514]), .B(n3048), .Z(n3050) );
  XOR U2540 ( .A(a[3517]), .B(n3036), .Z(n3038) );
  XOR U2541 ( .A(a[3520]), .B(n3023), .Z(n3025) );
  XOR U2542 ( .A(a[3523]), .B(n3011), .Z(n3013) );
  XOR U2543 ( .A(a[3526]), .B(n2999), .Z(n3001) );
  XOR U2544 ( .A(a[3529]), .B(n2986), .Z(n2988) );
  XOR U2545 ( .A(a[3532]), .B(n2974), .Z(n2976) );
  XOR U2546 ( .A(a[3535]), .B(n2962), .Z(n2964) );
  XOR U2547 ( .A(a[3538]), .B(n2950), .Z(n2952) );
  XOR U2548 ( .A(a[3541]), .B(n2937), .Z(n2939) );
  XOR U2549 ( .A(a[3544]), .B(n2925), .Z(n2927) );
  XOR U2550 ( .A(a[3547]), .B(n2913), .Z(n2915) );
  XOR U2551 ( .A(a[3550]), .B(n2900), .Z(n2902) );
  XOR U2552 ( .A(a[3553]), .B(n2888), .Z(n2890) );
  XOR U2553 ( .A(a[3556]), .B(n2876), .Z(n2878) );
  XOR U2554 ( .A(a[3559]), .B(n2863), .Z(n2865) );
  XOR U2555 ( .A(a[3562]), .B(n2851), .Z(n2853) );
  XOR U2556 ( .A(a[3565]), .B(n2839), .Z(n2841) );
  XOR U2557 ( .A(a[3568]), .B(n2827), .Z(n2829) );
  XOR U2558 ( .A(a[3571]), .B(n2814), .Z(n2816) );
  XOR U2559 ( .A(a[3574]), .B(n2802), .Z(n2804) );
  XOR U2560 ( .A(a[3577]), .B(n2790), .Z(n2792) );
  XOR U2561 ( .A(a[3580]), .B(n2777), .Z(n2779) );
  XOR U2562 ( .A(a[3583]), .B(n2765), .Z(n2767) );
  XOR U2563 ( .A(a[3586]), .B(n2753), .Z(n2755) );
  XOR U2564 ( .A(a[3589]), .B(n2740), .Z(n2742) );
  XOR U2565 ( .A(a[3592]), .B(n2728), .Z(n2730) );
  XOR U2566 ( .A(a[3595]), .B(n2716), .Z(n2718) );
  XOR U2567 ( .A(a[3598]), .B(n2704), .Z(n2706) );
  XOR U2568 ( .A(a[3601]), .B(n2690), .Z(n2692) );
  XOR U2569 ( .A(a[3604]), .B(n2678), .Z(n2680) );
  XOR U2570 ( .A(a[3607]), .B(n2666), .Z(n2668) );
  XOR U2571 ( .A(a[3610]), .B(n2653), .Z(n2655) );
  XOR U2572 ( .A(a[3613]), .B(n2641), .Z(n2643) );
  XOR U2573 ( .A(a[3616]), .B(n2629), .Z(n2631) );
  XOR U2574 ( .A(a[3619]), .B(n2616), .Z(n2618) );
  XOR U2575 ( .A(a[3622]), .B(n2604), .Z(n2606) );
  XOR U2576 ( .A(a[3625]), .B(n2592), .Z(n2594) );
  XOR U2577 ( .A(a[3628]), .B(n2580), .Z(n2582) );
  XOR U2578 ( .A(a[3631]), .B(n2567), .Z(n2569) );
  XOR U2579 ( .A(a[3634]), .B(n2555), .Z(n2557) );
  XOR U2580 ( .A(a[3637]), .B(n2543), .Z(n2545) );
  XOR U2581 ( .A(a[3640]), .B(n2530), .Z(n2532) );
  XOR U2582 ( .A(a[3643]), .B(n2518), .Z(n2520) );
  XOR U2583 ( .A(a[3646]), .B(n2506), .Z(n2508) );
  XOR U2584 ( .A(a[3649]), .B(n2493), .Z(n2495) );
  XOR U2585 ( .A(a[3652]), .B(n2481), .Z(n2483) );
  XOR U2586 ( .A(a[3655]), .B(n2469), .Z(n2471) );
  XOR U2587 ( .A(a[3658]), .B(n2457), .Z(n2459) );
  XOR U2588 ( .A(a[3661]), .B(n2444), .Z(n2446) );
  XOR U2589 ( .A(a[3664]), .B(n2432), .Z(n2434) );
  XOR U2590 ( .A(a[3667]), .B(n2420), .Z(n2422) );
  XOR U2591 ( .A(a[3670]), .B(n2407), .Z(n2409) );
  XOR U2592 ( .A(a[3673]), .B(n2395), .Z(n2397) );
  XOR U2593 ( .A(a[3676]), .B(n2383), .Z(n2385) );
  XOR U2594 ( .A(a[3679]), .B(n2370), .Z(n2372) );
  XOR U2595 ( .A(a[3682]), .B(n2358), .Z(n2360) );
  XOR U2596 ( .A(a[3685]), .B(n2346), .Z(n2348) );
  XOR U2597 ( .A(a[3688]), .B(n2334), .Z(n2336) );
  XOR U2598 ( .A(a[3691]), .B(n2321), .Z(n2323) );
  XOR U2599 ( .A(a[3694]), .B(n2309), .Z(n2311) );
  XOR U2600 ( .A(a[3697]), .B(n2297), .Z(n2299) );
  XOR U2601 ( .A(a[3700]), .B(n2283), .Z(n2285) );
  XOR U2602 ( .A(a[3703]), .B(n2271), .Z(n2273) );
  XOR U2603 ( .A(a[3706]), .B(n2259), .Z(n2261) );
  XOR U2604 ( .A(a[3709]), .B(n2246), .Z(n2248) );
  XOR U2605 ( .A(a[3712]), .B(n2234), .Z(n2236) );
  XOR U2606 ( .A(a[3715]), .B(n2222), .Z(n2224) );
  XOR U2607 ( .A(a[3718]), .B(n2210), .Z(n2212) );
  XOR U2608 ( .A(a[3721]), .B(n2197), .Z(n2199) );
  XOR U2609 ( .A(a[3724]), .B(n2185), .Z(n2187) );
  XOR U2610 ( .A(a[3727]), .B(n2173), .Z(n2175) );
  XOR U2611 ( .A(a[3730]), .B(n2160), .Z(n2162) );
  XOR U2612 ( .A(a[3733]), .B(n2148), .Z(n2150) );
  XOR U2613 ( .A(a[3736]), .B(n2136), .Z(n2138) );
  XOR U2614 ( .A(a[3739]), .B(n2123), .Z(n2125) );
  XOR U2615 ( .A(a[3742]), .B(n2111), .Z(n2113) );
  XOR U2616 ( .A(a[3745]), .B(n2099), .Z(n2101) );
  XOR U2617 ( .A(a[3748]), .B(n2087), .Z(n2089) );
  XOR U2618 ( .A(a[3751]), .B(n2074), .Z(n2076) );
  XOR U2619 ( .A(a[3754]), .B(n2062), .Z(n2064) );
  XOR U2620 ( .A(a[3757]), .B(n2050), .Z(n2052) );
  XOR U2621 ( .A(a[3760]), .B(n2037), .Z(n2039) );
  XOR U2622 ( .A(a[3763]), .B(n2025), .Z(n2027) );
  XOR U2623 ( .A(a[3766]), .B(n2013), .Z(n2015) );
  XOR U2624 ( .A(a[3769]), .B(n2000), .Z(n2002) );
  XOR U2625 ( .A(a[3772]), .B(n1988), .Z(n1990) );
  XOR U2626 ( .A(a[3775]), .B(n1976), .Z(n1978) );
  XOR U2627 ( .A(a[3778]), .B(n1964), .Z(n1966) );
  XOR U2628 ( .A(a[3781]), .B(n1951), .Z(n1953) );
  XOR U2629 ( .A(a[3784]), .B(n1939), .Z(n1941) );
  XOR U2630 ( .A(a[3787]), .B(n1927), .Z(n1929) );
  XOR U2631 ( .A(a[3790]), .B(n1914), .Z(n1916) );
  XOR U2632 ( .A(a[3793]), .B(n1902), .Z(n1904) );
  XOR U2633 ( .A(a[3796]), .B(n1890), .Z(n1892) );
  XOR U2634 ( .A(a[3799]), .B(n1876), .Z(n1878) );
  XOR U2635 ( .A(a[3802]), .B(n1864), .Z(n1866) );
  XOR U2636 ( .A(a[3805]), .B(n1852), .Z(n1854) );
  XOR U2637 ( .A(a[3808]), .B(n1840), .Z(n1842) );
  XOR U2638 ( .A(a[3811]), .B(n1827), .Z(n1829) );
  XOR U2639 ( .A(a[3814]), .B(n1815), .Z(n1817) );
  XOR U2640 ( .A(a[3817]), .B(n1803), .Z(n1805) );
  XOR U2641 ( .A(a[3820]), .B(n1790), .Z(n1792) );
  XOR U2642 ( .A(a[3823]), .B(n1778), .Z(n1780) );
  XOR U2643 ( .A(a[3826]), .B(n1766), .Z(n1768) );
  XOR U2644 ( .A(a[3829]), .B(n1753), .Z(n1755) );
  XOR U2645 ( .A(a[3832]), .B(n1741), .Z(n1743) );
  XOR U2646 ( .A(a[3835]), .B(n1729), .Z(n1731) );
  XOR U2647 ( .A(a[3838]), .B(n1717), .Z(n1719) );
  XOR U2648 ( .A(a[3841]), .B(n1704), .Z(n1706) );
  XOR U2649 ( .A(a[3844]), .B(n1692), .Z(n1694) );
  XOR U2650 ( .A(a[3847]), .B(n1680), .Z(n1682) );
  XOR U2651 ( .A(a[3850]), .B(n1667), .Z(n1669) );
  XOR U2652 ( .A(a[3853]), .B(n1655), .Z(n1657) );
  XOR U2653 ( .A(a[3856]), .B(n1643), .Z(n1645) );
  XOR U2654 ( .A(a[3859]), .B(n1630), .Z(n1632) );
  XOR U2655 ( .A(a[3862]), .B(n1618), .Z(n1620) );
  XOR U2656 ( .A(a[3865]), .B(n1606), .Z(n1608) );
  XOR U2657 ( .A(a[3868]), .B(n1594), .Z(n1596) );
  XOR U2658 ( .A(a[3871]), .B(n1581), .Z(n1583) );
  XOR U2659 ( .A(a[3874]), .B(n1569), .Z(n1571) );
  XOR U2660 ( .A(a[3877]), .B(n1557), .Z(n1559) );
  XOR U2661 ( .A(a[3880]), .B(n1544), .Z(n1546) );
  XOR U2662 ( .A(a[3883]), .B(n1532), .Z(n1534) );
  XOR U2663 ( .A(a[3886]), .B(n1520), .Z(n1522) );
  XOR U2664 ( .A(a[3889]), .B(n1507), .Z(n1509) );
  XOR U2665 ( .A(a[3892]), .B(n1495), .Z(n1497) );
  XOR U2666 ( .A(a[3895]), .B(n1483), .Z(n1485) );
  XOR U2667 ( .A(a[3898]), .B(n1471), .Z(n1473) );
  XOR U2668 ( .A(a[3901]), .B(n1457), .Z(n1459) );
  XOR U2669 ( .A(a[3904]), .B(n1445), .Z(n1447) );
  XOR U2670 ( .A(a[3907]), .B(n1433), .Z(n1435) );
  XOR U2671 ( .A(a[3910]), .B(n1420), .Z(n1422) );
  XOR U2672 ( .A(a[3913]), .B(n1408), .Z(n1410) );
  XOR U2673 ( .A(a[3916]), .B(n1396), .Z(n1398) );
  XOR U2674 ( .A(a[3919]), .B(n1383), .Z(n1385) );
  XOR U2675 ( .A(a[3922]), .B(n1371), .Z(n1373) );
  XOR U2676 ( .A(a[3925]), .B(n1359), .Z(n1361) );
  XOR U2677 ( .A(a[3928]), .B(n1347), .Z(n1349) );
  XOR U2678 ( .A(a[3931]), .B(n1334), .Z(n1336) );
  XOR U2679 ( .A(a[3934]), .B(n1322), .Z(n1324) );
  XOR U2680 ( .A(a[3937]), .B(n1310), .Z(n1312) );
  XOR U2681 ( .A(a[3940]), .B(n1297), .Z(n1299) );
  XOR U2682 ( .A(a[3943]), .B(n1285), .Z(n1287) );
  XOR U2683 ( .A(a[3946]), .B(n1273), .Z(n1275) );
  XOR U2684 ( .A(a[3949]), .B(n1260), .Z(n1262) );
  XOR U2685 ( .A(a[3952]), .B(n1248), .Z(n1250) );
  XOR U2686 ( .A(a[3955]), .B(n1236), .Z(n1238) );
  XOR U2687 ( .A(a[3958]), .B(n1224), .Z(n1226) );
  XOR U2688 ( .A(a[3961]), .B(n1211), .Z(n1213) );
  XOR U2689 ( .A(a[3964]), .B(n1199), .Z(n1201) );
  XOR U2690 ( .A(a[3967]), .B(n1187), .Z(n1189) );
  XOR U2691 ( .A(a[3970]), .B(n1174), .Z(n1176) );
  XOR U2692 ( .A(a[3973]), .B(n1162), .Z(n1164) );
  XOR U2693 ( .A(a[3976]), .B(n1150), .Z(n1152) );
  XOR U2694 ( .A(a[3979]), .B(n1137), .Z(n1139) );
  XOR U2695 ( .A(a[3982]), .B(n1125), .Z(n1127) );
  XOR U2696 ( .A(a[3985]), .B(n1113), .Z(n1115) );
  XOR U2697 ( .A(a[3988]), .B(n1101), .Z(n1103) );
  XOR U2698 ( .A(a[3991]), .B(n1088), .Z(n1090) );
  XOR U2699 ( .A(a[3994]), .B(n1076), .Z(n1078) );
  XOR U2700 ( .A(a[3997]), .B(n1064), .Z(n1066) );
  XOR U2701 ( .A(a[4000]), .B(n1049), .Z(n1051) );
  XOR U2702 ( .A(a[4003]), .B(n1037), .Z(n1039) );
  XOR U2703 ( .A(a[4006]), .B(n1025), .Z(n1027) );
  XOR U2704 ( .A(a[4009]), .B(n1012), .Z(n1014) );
  XOR U2705 ( .A(a[4012]), .B(n1000), .Z(n1002) );
  XOR U2706 ( .A(a[4015]), .B(n988), .Z(n990) );
  XOR U2707 ( .A(a[4018]), .B(n976), .Z(n978) );
  XOR U2708 ( .A(a[4021]), .B(n963), .Z(n965) );
  XOR U2709 ( .A(a[4024]), .B(n951), .Z(n953) );
  XOR U2710 ( .A(a[4027]), .B(n939), .Z(n941) );
  XOR U2711 ( .A(a[4030]), .B(n926), .Z(n928) );
  XOR U2712 ( .A(a[4033]), .B(n914), .Z(n916) );
  XOR U2713 ( .A(a[4036]), .B(n902), .Z(n904) );
  XOR U2714 ( .A(a[4039]), .B(n889), .Z(n891) );
  XOR U2715 ( .A(a[4042]), .B(n877), .Z(n879) );
  XOR U2716 ( .A(a[4045]), .B(n865), .Z(n867) );
  XOR U2717 ( .A(a[4048]), .B(n853), .Z(n855) );
  XOR U2718 ( .A(a[4051]), .B(n840), .Z(n842) );
  XOR U2719 ( .A(a[4054]), .B(n828), .Z(n830) );
  XOR U2720 ( .A(a[4057]), .B(n816), .Z(n818) );
  XOR U2721 ( .A(a[4060]), .B(n803), .Z(n805) );
  XOR U2722 ( .A(a[4063]), .B(n791), .Z(n793) );
  XOR U2723 ( .A(a[4066]), .B(n779), .Z(n781) );
  XOR U2724 ( .A(a[4069]), .B(n766), .Z(n768) );
  XOR U2725 ( .A(a[4072]), .B(n754), .Z(n756) );
  XOR U2726 ( .A(a[4075]), .B(n742), .Z(n744) );
  XOR U2727 ( .A(a[4078]), .B(n730), .Z(n732) );
  XOR U2728 ( .A(a[4081]), .B(n717), .Z(n719) );
  XOR U2729 ( .A(a[4084]), .B(n705), .Z(n707) );
  XOR U2730 ( .A(a[4087]), .B(n693), .Z(n695) );
  XOR U2731 ( .A(a[4090]), .B(n680), .Z(n682) );
  XOR U2732 ( .A(a[4093]), .B(n668), .Z(n670) );
  XOR U2733 ( .A(a[2]), .B(n16377), .Z(n5167) );
  XOR U2734 ( .A(a[5]), .B(n16368), .Z(n450) );
  XOR U2735 ( .A(a[8]), .B(n16359), .Z(n117) );
  XOR U2736 ( .A(a[11]), .B(n16350), .Z(n12567) );
  XOR U2737 ( .A(a[14]), .B(n16341), .Z(n11334) );
  XOR U2738 ( .A(a[17]), .B(n16332), .Z(n10101) );
  XOR U2739 ( .A(a[20]), .B(n16323), .Z(n8867) );
  XOR U2740 ( .A(a[23]), .B(n16314), .Z(n7634) );
  XOR U2741 ( .A(a[26]), .B(n16305), .Z(n6401) );
  XOR U2742 ( .A(a[29]), .B(n16296), .Z(n5168) );
  XOR U2743 ( .A(a[32]), .B(n16287), .Z(n3934) );
  XOR U2744 ( .A(a[35]), .B(n16278), .Z(n2701) );
  XOR U2745 ( .A(a[38]), .B(n16269), .Z(n1468) );
  XOR U2746 ( .A(a[41]), .B(n16260), .Z(n650) );
  XOR U2747 ( .A(a[44]), .B(n16251), .Z(n617) );
  XOR U2748 ( .A(a[47]), .B(n16242), .Z(n584) );
  XOR U2749 ( .A(a[50]), .B(n16233), .Z(n550) );
  XOR U2750 ( .A(a[53]), .B(n16224), .Z(n517) );
  XOR U2751 ( .A(a[56]), .B(n16215), .Z(n484) );
  XOR U2752 ( .A(a[59]), .B(n16206), .Z(n451) );
  XOR U2753 ( .A(a[62]), .B(n16197), .Z(n417) );
  XOR U2754 ( .A(a[65]), .B(n16188), .Z(n384) );
  XOR U2755 ( .A(a[68]), .B(n16179), .Z(n351) );
  XOR U2756 ( .A(a[71]), .B(n16170), .Z(n317) );
  XOR U2757 ( .A(a[74]), .B(n16161), .Z(n284) );
  XOR U2758 ( .A(a[77]), .B(n16152), .Z(n251) );
  XOR U2759 ( .A(a[80]), .B(n16143), .Z(n217) );
  XOR U2760 ( .A(a[83]), .B(n16134), .Z(n184) );
  XOR U2761 ( .A(a[86]), .B(n16125), .Z(n151) );
  XOR U2762 ( .A(a[89]), .B(n16116), .Z(n118) );
  XOR U2763 ( .A(a[92]), .B(n16107), .Z(n84) );
  XOR U2764 ( .A(a[95]), .B(n16098), .Z(n51) );
  XOR U2765 ( .A(a[98]), .B(n16089), .Z(n18) );
  XOR U2766 ( .A(a[101]), .B(n16080), .Z(n13307) );
  XOR U2767 ( .A(a[104]), .B(n16071), .Z(n13184) );
  XOR U2768 ( .A(a[107]), .B(n16062), .Z(n13061) );
  XOR U2769 ( .A(a[110]), .B(n16053), .Z(n12937) );
  XOR U2770 ( .A(a[113]), .B(n16044), .Z(n12814) );
  XOR U2771 ( .A(a[116]), .B(n16035), .Z(n12691) );
  XOR U2772 ( .A(a[119]), .B(n16026), .Z(n12568) );
  XOR U2773 ( .A(a[122]), .B(n16017), .Z(n12444) );
  XOR U2774 ( .A(a[125]), .B(n16008), .Z(n12321) );
  XOR U2775 ( .A(a[128]), .B(n15999), .Z(n12198) );
  XOR U2776 ( .A(a[131]), .B(n15990), .Z(n12074) );
  XOR U2777 ( .A(a[134]), .B(n15981), .Z(n11951) );
  XOR U2778 ( .A(a[137]), .B(n15972), .Z(n11828) );
  XOR U2779 ( .A(a[140]), .B(n15963), .Z(n11704) );
  XOR U2780 ( .A(a[143]), .B(n15954), .Z(n11581) );
  XOR U2781 ( .A(a[146]), .B(n15945), .Z(n11458) );
  XOR U2782 ( .A(a[149]), .B(n15936), .Z(n11335) );
  XOR U2783 ( .A(a[152]), .B(n15927), .Z(n11211) );
  XOR U2784 ( .A(a[155]), .B(n15918), .Z(n11088) );
  XOR U2785 ( .A(a[158]), .B(n15909), .Z(n10965) );
  XOR U2786 ( .A(a[161]), .B(n15900), .Z(n10841) );
  XOR U2787 ( .A(a[164]), .B(n15891), .Z(n10718) );
  XOR U2788 ( .A(a[167]), .B(n15882), .Z(n10595) );
  XOR U2789 ( .A(a[170]), .B(n15873), .Z(n10471) );
  XOR U2790 ( .A(a[173]), .B(n15864), .Z(n10348) );
  XOR U2791 ( .A(a[176]), .B(n15855), .Z(n10225) );
  XOR U2792 ( .A(a[179]), .B(n15846), .Z(n10102) );
  XOR U2793 ( .A(a[182]), .B(n15837), .Z(n9978) );
  XOR U2794 ( .A(a[185]), .B(n15828), .Z(n9855) );
  XOR U2795 ( .A(a[188]), .B(n15819), .Z(n9732) );
  XOR U2796 ( .A(a[191]), .B(n15810), .Z(n9608) );
  XOR U2797 ( .A(a[194]), .B(n15801), .Z(n9485) );
  XOR U2798 ( .A(a[197]), .B(n15792), .Z(n9362) );
  XOR U2799 ( .A(a[200]), .B(n15783), .Z(n9237) );
  XOR U2800 ( .A(a[203]), .B(n15774), .Z(n9114) );
  XOR U2801 ( .A(a[206]), .B(n15765), .Z(n8991) );
  XOR U2802 ( .A(a[209]), .B(n15756), .Z(n8868) );
  XOR U2803 ( .A(a[212]), .B(n15747), .Z(n8744) );
  XOR U2804 ( .A(a[215]), .B(n15738), .Z(n8621) );
  XOR U2805 ( .A(a[218]), .B(n15729), .Z(n8498) );
  XOR U2806 ( .A(a[221]), .B(n15720), .Z(n8374) );
  XOR U2807 ( .A(a[224]), .B(n15711), .Z(n8251) );
  XOR U2808 ( .A(a[227]), .B(n15702), .Z(n8128) );
  XOR U2809 ( .A(a[230]), .B(n15693), .Z(n8004) );
  XOR U2810 ( .A(a[233]), .B(n15684), .Z(n7881) );
  XOR U2811 ( .A(a[236]), .B(n15675), .Z(n7758) );
  XOR U2812 ( .A(a[239]), .B(n15666), .Z(n7635) );
  XOR U2813 ( .A(a[242]), .B(n15657), .Z(n7511) );
  XOR U2814 ( .A(a[245]), .B(n15648), .Z(n7388) );
  XOR U2815 ( .A(a[248]), .B(n15639), .Z(n7265) );
  XOR U2816 ( .A(a[251]), .B(n15630), .Z(n7141) );
  XOR U2817 ( .A(a[254]), .B(n15621), .Z(n7018) );
  XOR U2818 ( .A(a[257]), .B(n15612), .Z(n6895) );
  XOR U2819 ( .A(a[260]), .B(n15603), .Z(n6771) );
  XOR U2820 ( .A(a[263]), .B(n15594), .Z(n6648) );
  XOR U2821 ( .A(a[266]), .B(n15585), .Z(n6525) );
  XOR U2822 ( .A(a[269]), .B(n15576), .Z(n6402) );
  XOR U2823 ( .A(a[272]), .B(n15567), .Z(n6278) );
  XOR U2824 ( .A(a[275]), .B(n15558), .Z(n6155) );
  XOR U2825 ( .A(a[278]), .B(n15549), .Z(n6032) );
  XOR U2826 ( .A(a[281]), .B(n15540), .Z(n5908) );
  XOR U2827 ( .A(a[284]), .B(n15531), .Z(n5785) );
  XOR U2828 ( .A(a[287]), .B(n15522), .Z(n5662) );
  XOR U2829 ( .A(a[290]), .B(n15513), .Z(n5538) );
  XOR U2830 ( .A(a[293]), .B(n15504), .Z(n5415) );
  XOR U2831 ( .A(a[296]), .B(n15495), .Z(n5292) );
  XOR U2832 ( .A(a[299]), .B(n15486), .Z(n5169) );
  XOR U2833 ( .A(a[302]), .B(n15477), .Z(n5044) );
  XOR U2834 ( .A(a[305]), .B(n15468), .Z(n4921) );
  XOR U2835 ( .A(a[308]), .B(n15459), .Z(n4798) );
  XOR U2836 ( .A(a[311]), .B(n15450), .Z(n4674) );
  XOR U2837 ( .A(a[314]), .B(n15441), .Z(n4551) );
  XOR U2838 ( .A(a[317]), .B(n15432), .Z(n4428) );
  XOR U2839 ( .A(a[320]), .B(n15423), .Z(n4304) );
  XOR U2840 ( .A(a[323]), .B(n15414), .Z(n4181) );
  XOR U2841 ( .A(a[326]), .B(n15405), .Z(n4058) );
  XOR U2842 ( .A(a[329]), .B(n15396), .Z(n3935) );
  XOR U2843 ( .A(a[332]), .B(n15387), .Z(n3811) );
  XOR U2844 ( .A(a[335]), .B(n15378), .Z(n3688) );
  XOR U2845 ( .A(a[338]), .B(n15369), .Z(n3565) );
  XOR U2846 ( .A(a[341]), .B(n15360), .Z(n3441) );
  XOR U2847 ( .A(a[344]), .B(n15351), .Z(n3318) );
  XOR U2848 ( .A(a[347]), .B(n15342), .Z(n3195) );
  XOR U2849 ( .A(a[350]), .B(n15333), .Z(n3071) );
  XOR U2850 ( .A(a[353]), .B(n15324), .Z(n2948) );
  XOR U2851 ( .A(a[356]), .B(n15315), .Z(n2825) );
  XOR U2852 ( .A(a[359]), .B(n15306), .Z(n2702) );
  XOR U2853 ( .A(a[362]), .B(n15297), .Z(n2578) );
  XOR U2854 ( .A(a[365]), .B(n15288), .Z(n2455) );
  XOR U2855 ( .A(a[368]), .B(n15279), .Z(n2332) );
  XOR U2856 ( .A(a[371]), .B(n15270), .Z(n2208) );
  XOR U2857 ( .A(a[374]), .B(n15261), .Z(n2085) );
  XOR U2858 ( .A(a[377]), .B(n15252), .Z(n1962) );
  XOR U2859 ( .A(a[380]), .B(n15243), .Z(n1838) );
  XOR U2860 ( .A(a[383]), .B(n15234), .Z(n1715) );
  XOR U2861 ( .A(a[386]), .B(n15225), .Z(n1592) );
  XOR U2862 ( .A(a[389]), .B(n15216), .Z(n1469) );
  XOR U2863 ( .A(a[392]), .B(n15207), .Z(n1345) );
  XOR U2864 ( .A(a[395]), .B(n15198), .Z(n1222) );
  XOR U2865 ( .A(a[398]), .B(n15189), .Z(n1099) );
  XOR U2866 ( .A(a[401]), .B(n15180), .Z(n974) );
  XOR U2867 ( .A(a[404]), .B(n15171), .Z(n851) );
  XOR U2868 ( .A(a[407]), .B(n15162), .Z(n728) );
  XOR U2869 ( .A(a[410]), .B(n15153), .Z(n660) );
  XOR U2870 ( .A(a[413]), .B(n15144), .Z(n657) );
  XOR U2871 ( .A(a[416]), .B(n15135), .Z(n654) );
  XOR U2872 ( .A(a[419]), .B(n15126), .Z(n651) );
  XOR U2873 ( .A(a[422]), .B(n15117), .Z(n647) );
  XOR U2874 ( .A(a[425]), .B(n15108), .Z(n644) );
  XOR U2875 ( .A(a[428]), .B(n15099), .Z(n641) );
  XOR U2876 ( .A(a[431]), .B(n15090), .Z(n637) );
  XOR U2877 ( .A(a[434]), .B(n15081), .Z(n634) );
  XOR U2878 ( .A(a[437]), .B(n15072), .Z(n631) );
  XOR U2879 ( .A(a[440]), .B(n15063), .Z(n627) );
  XOR U2880 ( .A(a[443]), .B(n15054), .Z(n624) );
  XOR U2881 ( .A(a[446]), .B(n15045), .Z(n621) );
  XOR U2882 ( .A(a[449]), .B(n15036), .Z(n618) );
  XOR U2883 ( .A(a[452]), .B(n15027), .Z(n614) );
  XOR U2884 ( .A(a[455]), .B(n15018), .Z(n611) );
  XOR U2885 ( .A(a[458]), .B(n15009), .Z(n608) );
  XOR U2886 ( .A(a[461]), .B(n15000), .Z(n604) );
  XOR U2887 ( .A(a[464]), .B(n14991), .Z(n601) );
  XOR U2888 ( .A(a[467]), .B(n14982), .Z(n598) );
  XOR U2889 ( .A(a[470]), .B(n14973), .Z(n594) );
  XOR U2890 ( .A(a[473]), .B(n14964), .Z(n591) );
  XOR U2891 ( .A(a[476]), .B(n14955), .Z(n588) );
  XOR U2892 ( .A(a[479]), .B(n14946), .Z(n585) );
  XOR U2893 ( .A(a[482]), .B(n14937), .Z(n581) );
  XOR U2894 ( .A(a[485]), .B(n14928), .Z(n578) );
  XOR U2895 ( .A(a[488]), .B(n14919), .Z(n575) );
  XOR U2896 ( .A(a[491]), .B(n14910), .Z(n571) );
  XOR U2897 ( .A(a[494]), .B(n14901), .Z(n568) );
  XOR U2898 ( .A(a[497]), .B(n14892), .Z(n565) );
  XOR U2899 ( .A(a[500]), .B(n14883), .Z(n560) );
  XOR U2900 ( .A(a[503]), .B(n14874), .Z(n557) );
  XOR U2901 ( .A(a[506]), .B(n14865), .Z(n554) );
  XOR U2902 ( .A(a[509]), .B(n14856), .Z(n551) );
  XOR U2903 ( .A(a[512]), .B(n14847), .Z(n547) );
  XOR U2904 ( .A(a[515]), .B(n14838), .Z(n544) );
  XOR U2905 ( .A(a[518]), .B(n14829), .Z(n541) );
  XOR U2906 ( .A(a[521]), .B(n14820), .Z(n537) );
  XOR U2907 ( .A(a[524]), .B(n14811), .Z(n534) );
  XOR U2908 ( .A(a[527]), .B(n14802), .Z(n531) );
  XOR U2909 ( .A(a[530]), .B(n14793), .Z(n527) );
  XOR U2910 ( .A(a[533]), .B(n14784), .Z(n524) );
  XOR U2911 ( .A(a[536]), .B(n14775), .Z(n521) );
  XOR U2912 ( .A(a[539]), .B(n14766), .Z(n518) );
  XOR U2913 ( .A(a[542]), .B(n14757), .Z(n514) );
  XOR U2914 ( .A(a[545]), .B(n14748), .Z(n511) );
  XOR U2915 ( .A(a[548]), .B(n14739), .Z(n508) );
  XOR U2916 ( .A(a[551]), .B(n14730), .Z(n504) );
  XOR U2917 ( .A(a[554]), .B(n14721), .Z(n501) );
  XOR U2918 ( .A(a[557]), .B(n14712), .Z(n498) );
  XOR U2919 ( .A(a[560]), .B(n14703), .Z(n494) );
  XOR U2920 ( .A(a[563]), .B(n14694), .Z(n491) );
  XOR U2921 ( .A(a[566]), .B(n14685), .Z(n488) );
  XOR U2922 ( .A(a[569]), .B(n14676), .Z(n485) );
  XOR U2923 ( .A(a[572]), .B(n14667), .Z(n481) );
  XOR U2924 ( .A(a[575]), .B(n14658), .Z(n478) );
  XOR U2925 ( .A(a[578]), .B(n14649), .Z(n475) );
  XOR U2926 ( .A(a[581]), .B(n14640), .Z(n471) );
  XOR U2927 ( .A(a[584]), .B(n14631), .Z(n468) );
  XOR U2928 ( .A(a[587]), .B(n14622), .Z(n465) );
  XOR U2929 ( .A(a[590]), .B(n14613), .Z(n461) );
  XOR U2930 ( .A(a[593]), .B(n14604), .Z(n458) );
  XOR U2931 ( .A(a[596]), .B(n14595), .Z(n455) );
  XOR U2932 ( .A(a[599]), .B(n14586), .Z(n452) );
  XOR U2933 ( .A(a[602]), .B(n14577), .Z(n447) );
  XOR U2934 ( .A(a[605]), .B(n14568), .Z(n444) );
  XOR U2935 ( .A(a[608]), .B(n14559), .Z(n441) );
  XOR U2936 ( .A(a[611]), .B(n14550), .Z(n437) );
  XOR U2937 ( .A(a[614]), .B(n14541), .Z(n434) );
  XOR U2938 ( .A(a[617]), .B(n14532), .Z(n431) );
  XOR U2939 ( .A(a[620]), .B(n14523), .Z(n427) );
  XOR U2940 ( .A(a[623]), .B(n14514), .Z(n424) );
  XOR U2941 ( .A(a[626]), .B(n14505), .Z(n421) );
  XOR U2942 ( .A(a[629]), .B(n14496), .Z(n418) );
  XOR U2943 ( .A(a[632]), .B(n14487), .Z(n414) );
  XOR U2944 ( .A(a[635]), .B(n14478), .Z(n411) );
  XOR U2945 ( .A(a[638]), .B(n14469), .Z(n408) );
  XOR U2946 ( .A(a[641]), .B(n14460), .Z(n404) );
  XOR U2947 ( .A(a[644]), .B(n14451), .Z(n401) );
  XOR U2948 ( .A(a[647]), .B(n14442), .Z(n398) );
  XOR U2949 ( .A(a[650]), .B(n14433), .Z(n394) );
  XOR U2950 ( .A(a[653]), .B(n14424), .Z(n391) );
  XOR U2951 ( .A(a[656]), .B(n14415), .Z(n388) );
  XOR U2952 ( .A(a[659]), .B(n14406), .Z(n385) );
  XOR U2953 ( .A(a[662]), .B(n14397), .Z(n381) );
  XOR U2954 ( .A(a[665]), .B(n14388), .Z(n378) );
  XOR U2955 ( .A(a[668]), .B(n14379), .Z(n375) );
  XOR U2956 ( .A(a[671]), .B(n14370), .Z(n371) );
  XOR U2957 ( .A(a[674]), .B(n14361), .Z(n368) );
  XOR U2958 ( .A(a[677]), .B(n14352), .Z(n365) );
  XOR U2959 ( .A(a[680]), .B(n14343), .Z(n361) );
  XOR U2960 ( .A(a[683]), .B(n14334), .Z(n358) );
  XOR U2961 ( .A(a[686]), .B(n14325), .Z(n355) );
  XOR U2962 ( .A(a[689]), .B(n14316), .Z(n352) );
  XOR U2963 ( .A(a[692]), .B(n14307), .Z(n348) );
  XOR U2964 ( .A(a[695]), .B(n14298), .Z(n345) );
  XOR U2965 ( .A(a[698]), .B(n14289), .Z(n342) );
  XOR U2966 ( .A(a[701]), .B(n14280), .Z(n337) );
  XOR U2967 ( .A(a[704]), .B(n14271), .Z(n334) );
  XOR U2968 ( .A(a[707]), .B(n14262), .Z(n331) );
  XOR U2969 ( .A(a[710]), .B(n14253), .Z(n327) );
  XOR U2970 ( .A(a[713]), .B(n14244), .Z(n324) );
  XOR U2971 ( .A(a[716]), .B(n14235), .Z(n321) );
  XOR U2972 ( .A(a[719]), .B(n14226), .Z(n318) );
  XOR U2973 ( .A(a[722]), .B(n14217), .Z(n314) );
  XOR U2974 ( .A(a[725]), .B(n14208), .Z(n311) );
  XOR U2975 ( .A(a[728]), .B(n14199), .Z(n308) );
  XOR U2976 ( .A(a[731]), .B(n14190), .Z(n304) );
  XOR U2977 ( .A(a[734]), .B(n14181), .Z(n301) );
  XOR U2978 ( .A(a[737]), .B(n14172), .Z(n298) );
  XOR U2979 ( .A(a[740]), .B(n14163), .Z(n294) );
  XOR U2980 ( .A(a[743]), .B(n14154), .Z(n291) );
  XOR U2981 ( .A(a[746]), .B(n14145), .Z(n288) );
  XOR U2982 ( .A(a[749]), .B(n14136), .Z(n285) );
  XOR U2983 ( .A(a[752]), .B(n14127), .Z(n281) );
  XOR U2984 ( .A(a[755]), .B(n14118), .Z(n278) );
  XOR U2985 ( .A(a[758]), .B(n14109), .Z(n275) );
  XOR U2986 ( .A(a[761]), .B(n14100), .Z(n271) );
  XOR U2987 ( .A(a[764]), .B(n14091), .Z(n268) );
  XOR U2988 ( .A(a[767]), .B(n14082), .Z(n265) );
  XOR U2989 ( .A(a[770]), .B(n14073), .Z(n261) );
  XOR U2990 ( .A(a[773]), .B(n14064), .Z(n258) );
  XOR U2991 ( .A(a[776]), .B(n14055), .Z(n255) );
  XOR U2992 ( .A(a[779]), .B(n14046), .Z(n252) );
  XOR U2993 ( .A(a[782]), .B(n14037), .Z(n248) );
  XOR U2994 ( .A(a[785]), .B(n14028), .Z(n245) );
  XOR U2995 ( .A(a[788]), .B(n14019), .Z(n242) );
  XOR U2996 ( .A(a[791]), .B(n14010), .Z(n238) );
  XOR U2997 ( .A(a[794]), .B(n14001), .Z(n235) );
  XOR U2998 ( .A(a[797]), .B(n13992), .Z(n232) );
  XOR U2999 ( .A(a[800]), .B(n13983), .Z(n227) );
  XOR U3000 ( .A(a[803]), .B(n13974), .Z(n224) );
  XOR U3001 ( .A(a[806]), .B(n13965), .Z(n221) );
  XOR U3002 ( .A(a[809]), .B(n13956), .Z(n218) );
  XOR U3003 ( .A(a[812]), .B(n13947), .Z(n214) );
  XOR U3004 ( .A(a[815]), .B(n13938), .Z(n211) );
  XOR U3005 ( .A(a[818]), .B(n13929), .Z(n208) );
  XOR U3006 ( .A(a[821]), .B(n13920), .Z(n204) );
  XOR U3007 ( .A(a[824]), .B(n13911), .Z(n201) );
  XOR U3008 ( .A(a[827]), .B(n13902), .Z(n198) );
  XOR U3009 ( .A(a[830]), .B(n13893), .Z(n194) );
  XOR U3010 ( .A(a[833]), .B(n13884), .Z(n191) );
  XOR U3011 ( .A(a[836]), .B(n13875), .Z(n188) );
  XOR U3012 ( .A(a[839]), .B(n13866), .Z(n185) );
  XOR U3013 ( .A(a[842]), .B(n13857), .Z(n181) );
  XOR U3014 ( .A(a[845]), .B(n13848), .Z(n178) );
  XOR U3015 ( .A(a[848]), .B(n13839), .Z(n175) );
  XOR U3016 ( .A(a[851]), .B(n13830), .Z(n171) );
  XOR U3017 ( .A(a[854]), .B(n13821), .Z(n168) );
  XOR U3018 ( .A(a[857]), .B(n13812), .Z(n165) );
  XOR U3019 ( .A(a[860]), .B(n13803), .Z(n161) );
  XOR U3020 ( .A(a[863]), .B(n13794), .Z(n158) );
  XOR U3021 ( .A(a[866]), .B(n13785), .Z(n155) );
  XOR U3022 ( .A(a[869]), .B(n13776), .Z(n152) );
  XOR U3023 ( .A(a[872]), .B(n13767), .Z(n148) );
  XOR U3024 ( .A(a[875]), .B(n13758), .Z(n145) );
  XOR U3025 ( .A(a[878]), .B(n13749), .Z(n142) );
  XOR U3026 ( .A(a[881]), .B(n13740), .Z(n138) );
  XOR U3027 ( .A(a[884]), .B(n13731), .Z(n135) );
  XOR U3028 ( .A(a[887]), .B(n13722), .Z(n132) );
  XOR U3029 ( .A(a[890]), .B(n13713), .Z(n128) );
  XOR U3030 ( .A(a[893]), .B(n13704), .Z(n125) );
  XOR U3031 ( .A(a[896]), .B(n13695), .Z(n122) );
  XOR U3032 ( .A(a[899]), .B(n13686), .Z(n119) );
  XOR U3033 ( .A(a[902]), .B(n13677), .Z(n114) );
  XOR U3034 ( .A(a[905]), .B(n13668), .Z(n111) );
  XOR U3035 ( .A(a[908]), .B(n13659), .Z(n108) );
  XOR U3036 ( .A(a[911]), .B(n13650), .Z(n104) );
  XOR U3037 ( .A(a[914]), .B(n13641), .Z(n101) );
  XOR U3038 ( .A(a[917]), .B(n13632), .Z(n98) );
  XOR U3039 ( .A(a[920]), .B(n13623), .Z(n94) );
  XOR U3040 ( .A(a[923]), .B(n13614), .Z(n91) );
  XOR U3041 ( .A(a[926]), .B(n13605), .Z(n88) );
  XOR U3042 ( .A(a[929]), .B(n13596), .Z(n85) );
  XOR U3043 ( .A(a[932]), .B(n13587), .Z(n81) );
  XOR U3044 ( .A(a[935]), .B(n13578), .Z(n78) );
  XOR U3045 ( .A(a[938]), .B(n13569), .Z(n75) );
  XOR U3046 ( .A(a[941]), .B(n13560), .Z(n71) );
  XOR U3047 ( .A(a[944]), .B(n13551), .Z(n68) );
  XOR U3048 ( .A(a[947]), .B(n13542), .Z(n65) );
  XOR U3049 ( .A(a[950]), .B(n13533), .Z(n61) );
  XOR U3050 ( .A(a[953]), .B(n13524), .Z(n58) );
  XOR U3051 ( .A(a[956]), .B(n13515), .Z(n55) );
  XOR U3052 ( .A(a[959]), .B(n13506), .Z(n52) );
  XOR U3053 ( .A(a[962]), .B(n13497), .Z(n48) );
  XOR U3054 ( .A(a[965]), .B(n13488), .Z(n45) );
  XOR U3055 ( .A(a[968]), .B(n13479), .Z(n42) );
  XOR U3056 ( .A(a[971]), .B(n13470), .Z(n38) );
  XOR U3057 ( .A(a[974]), .B(n13461), .Z(n35) );
  XOR U3058 ( .A(a[977]), .B(n13452), .Z(n32) );
  XOR U3059 ( .A(a[980]), .B(n13443), .Z(n28) );
  XOR U3060 ( .A(a[983]), .B(n13434), .Z(n25) );
  XOR U3061 ( .A(a[986]), .B(n13425), .Z(n22) );
  XOR U3062 ( .A(a[989]), .B(n13416), .Z(n19) );
  XOR U3063 ( .A(a[992]), .B(n13407), .Z(n15) );
  XOR U3064 ( .A(a[995]), .B(n13398), .Z(n12) );
  XOR U3065 ( .A(a[998]), .B(n13389), .Z(n9) );
  XOR U3066 ( .A(a[1001]), .B(n13378), .Z(n13380) );
  XOR U3067 ( .A(a[1004]), .B(n13366), .Z(n13368) );
  XOR U3068 ( .A(a[1007]), .B(n13354), .Z(n13356) );
  XOR U3069 ( .A(a[1010]), .B(n13341), .Z(n13343) );
  XOR U3070 ( .A(a[1013]), .B(n13329), .Z(n13331) );
  XOR U3071 ( .A(a[1016]), .B(n13317), .Z(n13319) );
  XOR U3072 ( .A(a[1019]), .B(n13304), .Z(n13306) );
  XOR U3073 ( .A(a[1022]), .B(n13292), .Z(n13294) );
  XOR U3074 ( .A(a[1025]), .B(n13280), .Z(n13282) );
  XOR U3075 ( .A(a[1028]), .B(n13268), .Z(n13270) );
  XOR U3076 ( .A(a[1031]), .B(n13255), .Z(n13257) );
  XOR U3077 ( .A(a[1034]), .B(n13243), .Z(n13245) );
  XOR U3078 ( .A(a[1037]), .B(n13231), .Z(n13233) );
  XOR U3079 ( .A(a[1040]), .B(n13218), .Z(n13220) );
  XOR U3080 ( .A(a[1043]), .B(n13206), .Z(n13208) );
  XOR U3081 ( .A(a[1046]), .B(n13194), .Z(n13196) );
  XOR U3082 ( .A(a[1049]), .B(n13181), .Z(n13183) );
  XOR U3083 ( .A(a[1052]), .B(n13169), .Z(n13171) );
  XOR U3084 ( .A(a[1055]), .B(n13157), .Z(n13159) );
  XOR U3085 ( .A(a[1058]), .B(n13145), .Z(n13147) );
  XOR U3086 ( .A(a[1061]), .B(n13132), .Z(n13134) );
  XOR U3087 ( .A(a[1064]), .B(n13120), .Z(n13122) );
  XOR U3088 ( .A(a[1067]), .B(n13108), .Z(n13110) );
  XOR U3089 ( .A(a[1070]), .B(n13095), .Z(n13097) );
  XOR U3090 ( .A(a[1073]), .B(n13083), .Z(n13085) );
  XOR U3091 ( .A(a[1076]), .B(n13071), .Z(n13073) );
  XOR U3092 ( .A(a[1079]), .B(n13058), .Z(n13060) );
  XOR U3093 ( .A(a[1082]), .B(n13046), .Z(n13048) );
  XOR U3094 ( .A(a[1085]), .B(n13034), .Z(n13036) );
  XOR U3095 ( .A(a[1088]), .B(n13022), .Z(n13024) );
  XOR U3096 ( .A(a[1091]), .B(n13009), .Z(n13011) );
  XOR U3097 ( .A(a[1094]), .B(n12997), .Z(n12999) );
  XOR U3098 ( .A(a[1097]), .B(n12985), .Z(n12987) );
  XOR U3099 ( .A(a[1100]), .B(n12971), .Z(n12973) );
  XOR U3100 ( .A(a[1103]), .B(n12959), .Z(n12961) );
  XOR U3101 ( .A(a[1106]), .B(n12947), .Z(n12949) );
  XOR U3102 ( .A(a[1109]), .B(n12934), .Z(n12936) );
  XOR U3103 ( .A(a[1112]), .B(n12922), .Z(n12924) );
  XOR U3104 ( .A(a[1115]), .B(n12910), .Z(n12912) );
  XOR U3105 ( .A(a[1118]), .B(n12898), .Z(n12900) );
  XOR U3106 ( .A(a[1121]), .B(n12885), .Z(n12887) );
  XOR U3107 ( .A(a[1124]), .B(n12873), .Z(n12875) );
  XOR U3108 ( .A(a[1127]), .B(n12861), .Z(n12863) );
  XOR U3109 ( .A(a[1130]), .B(n12848), .Z(n12850) );
  XOR U3110 ( .A(a[1133]), .B(n12836), .Z(n12838) );
  XOR U3111 ( .A(a[1136]), .B(n12824), .Z(n12826) );
  XOR U3112 ( .A(a[1139]), .B(n12811), .Z(n12813) );
  XOR U3113 ( .A(a[1142]), .B(n12799), .Z(n12801) );
  XOR U3114 ( .A(a[1145]), .B(n12787), .Z(n12789) );
  XOR U3115 ( .A(a[1148]), .B(n12775), .Z(n12777) );
  XOR U3116 ( .A(a[1151]), .B(n12762), .Z(n12764) );
  XOR U3117 ( .A(a[1154]), .B(n12750), .Z(n12752) );
  XOR U3118 ( .A(a[1157]), .B(n12738), .Z(n12740) );
  XOR U3119 ( .A(a[1160]), .B(n12725), .Z(n12727) );
  XOR U3120 ( .A(a[1163]), .B(n12713), .Z(n12715) );
  XOR U3121 ( .A(a[1166]), .B(n12701), .Z(n12703) );
  XOR U3122 ( .A(a[1169]), .B(n12688), .Z(n12690) );
  XOR U3123 ( .A(a[1172]), .B(n12676), .Z(n12678) );
  XOR U3124 ( .A(a[1175]), .B(n12664), .Z(n12666) );
  XOR U3125 ( .A(a[1178]), .B(n12652), .Z(n12654) );
  XOR U3126 ( .A(a[1181]), .B(n12639), .Z(n12641) );
  XOR U3127 ( .A(a[1184]), .B(n12627), .Z(n12629) );
  XOR U3128 ( .A(a[1187]), .B(n12615), .Z(n12617) );
  XOR U3129 ( .A(a[1190]), .B(n12602), .Z(n12604) );
  XOR U3130 ( .A(a[1193]), .B(n12590), .Z(n12592) );
  XOR U3131 ( .A(a[1196]), .B(n12578), .Z(n12580) );
  XOR U3132 ( .A(a[1199]), .B(n12564), .Z(n12566) );
  XOR U3133 ( .A(a[1202]), .B(n12552), .Z(n12554) );
  XOR U3134 ( .A(a[1205]), .B(n12540), .Z(n12542) );
  XOR U3135 ( .A(a[1208]), .B(n12528), .Z(n12530) );
  XOR U3136 ( .A(a[1211]), .B(n12515), .Z(n12517) );
  XOR U3137 ( .A(a[1214]), .B(n12503), .Z(n12505) );
  XOR U3138 ( .A(a[1217]), .B(n12491), .Z(n12493) );
  XOR U3139 ( .A(a[1220]), .B(n12478), .Z(n12480) );
  XOR U3140 ( .A(a[1223]), .B(n12466), .Z(n12468) );
  XOR U3141 ( .A(a[1226]), .B(n12454), .Z(n12456) );
  XOR U3142 ( .A(a[1229]), .B(n12441), .Z(n12443) );
  XOR U3143 ( .A(a[1232]), .B(n12429), .Z(n12431) );
  XOR U3144 ( .A(a[1235]), .B(n12417), .Z(n12419) );
  XOR U3145 ( .A(a[1238]), .B(n12405), .Z(n12407) );
  XOR U3146 ( .A(a[1241]), .B(n12392), .Z(n12394) );
  XOR U3147 ( .A(a[1244]), .B(n12380), .Z(n12382) );
  XOR U3148 ( .A(a[1247]), .B(n12368), .Z(n12370) );
  XOR U3149 ( .A(a[1250]), .B(n12355), .Z(n12357) );
  XOR U3150 ( .A(a[1253]), .B(n12343), .Z(n12345) );
  XOR U3151 ( .A(a[1256]), .B(n12331), .Z(n12333) );
  XOR U3152 ( .A(a[1259]), .B(n12318), .Z(n12320) );
  XOR U3153 ( .A(a[1262]), .B(n12306), .Z(n12308) );
  XOR U3154 ( .A(a[1265]), .B(n12294), .Z(n12296) );
  XOR U3155 ( .A(a[1268]), .B(n12282), .Z(n12284) );
  XOR U3156 ( .A(a[1271]), .B(n12269), .Z(n12271) );
  XOR U3157 ( .A(a[1274]), .B(n12257), .Z(n12259) );
  XOR U3158 ( .A(a[1277]), .B(n12245), .Z(n12247) );
  XOR U3159 ( .A(a[1280]), .B(n12232), .Z(n12234) );
  XOR U3160 ( .A(a[1283]), .B(n12220), .Z(n12222) );
  XOR U3161 ( .A(a[1286]), .B(n12208), .Z(n12210) );
  XOR U3162 ( .A(a[1289]), .B(n12195), .Z(n12197) );
  XOR U3163 ( .A(a[1292]), .B(n12183), .Z(n12185) );
  XOR U3164 ( .A(a[1295]), .B(n12171), .Z(n12173) );
  XOR U3165 ( .A(a[1298]), .B(n12159), .Z(n12161) );
  XOR U3166 ( .A(a[1301]), .B(n12145), .Z(n12147) );
  XOR U3167 ( .A(a[1304]), .B(n12133), .Z(n12135) );
  XOR U3168 ( .A(a[1307]), .B(n12121), .Z(n12123) );
  XOR U3169 ( .A(a[1310]), .B(n12108), .Z(n12110) );
  XOR U3170 ( .A(a[1313]), .B(n12096), .Z(n12098) );
  XOR U3171 ( .A(a[1316]), .B(n12084), .Z(n12086) );
  XOR U3172 ( .A(a[1319]), .B(n12071), .Z(n12073) );
  XOR U3173 ( .A(a[1322]), .B(n12059), .Z(n12061) );
  XOR U3174 ( .A(a[1325]), .B(n12047), .Z(n12049) );
  XOR U3175 ( .A(a[1328]), .B(n12035), .Z(n12037) );
  XOR U3176 ( .A(a[1331]), .B(n12022), .Z(n12024) );
  XOR U3177 ( .A(a[1334]), .B(n12010), .Z(n12012) );
  XOR U3178 ( .A(a[1337]), .B(n11998), .Z(n12000) );
  XOR U3179 ( .A(a[1340]), .B(n11985), .Z(n11987) );
  XOR U3180 ( .A(a[1343]), .B(n11973), .Z(n11975) );
  XOR U3181 ( .A(a[1346]), .B(n11961), .Z(n11963) );
  XOR U3182 ( .A(a[1349]), .B(n11948), .Z(n11950) );
  XOR U3183 ( .A(a[1352]), .B(n11936), .Z(n11938) );
  XOR U3184 ( .A(a[1355]), .B(n11924), .Z(n11926) );
  XOR U3185 ( .A(a[1358]), .B(n11912), .Z(n11914) );
  XOR U3186 ( .A(a[1361]), .B(n11899), .Z(n11901) );
  XOR U3187 ( .A(a[1364]), .B(n11887), .Z(n11889) );
  XOR U3188 ( .A(a[1367]), .B(n11875), .Z(n11877) );
  XOR U3189 ( .A(a[1370]), .B(n11862), .Z(n11864) );
  XOR U3190 ( .A(a[1373]), .B(n11850), .Z(n11852) );
  XOR U3191 ( .A(a[1376]), .B(n11838), .Z(n11840) );
  XOR U3192 ( .A(a[1379]), .B(n11825), .Z(n11827) );
  XOR U3193 ( .A(a[1382]), .B(n11813), .Z(n11815) );
  XOR U3194 ( .A(a[1385]), .B(n11801), .Z(n11803) );
  XOR U3195 ( .A(a[1388]), .B(n11789), .Z(n11791) );
  XOR U3196 ( .A(a[1391]), .B(n11776), .Z(n11778) );
  XOR U3197 ( .A(a[1394]), .B(n11764), .Z(n11766) );
  XOR U3198 ( .A(a[1397]), .B(n11752), .Z(n11754) );
  XOR U3199 ( .A(a[1400]), .B(n11738), .Z(n11740) );
  XOR U3200 ( .A(a[1403]), .B(n11726), .Z(n11728) );
  XOR U3201 ( .A(a[1406]), .B(n11714), .Z(n11716) );
  XOR U3202 ( .A(a[1409]), .B(n11701), .Z(n11703) );
  XOR U3203 ( .A(a[1412]), .B(n11689), .Z(n11691) );
  XOR U3204 ( .A(a[1415]), .B(n11677), .Z(n11679) );
  XOR U3205 ( .A(a[1418]), .B(n11665), .Z(n11667) );
  XOR U3206 ( .A(a[1421]), .B(n11652), .Z(n11654) );
  XOR U3207 ( .A(a[1424]), .B(n11640), .Z(n11642) );
  XOR U3208 ( .A(a[1427]), .B(n11628), .Z(n11630) );
  XOR U3209 ( .A(a[1430]), .B(n11615), .Z(n11617) );
  XOR U3210 ( .A(a[1433]), .B(n11603), .Z(n11605) );
  XOR U3211 ( .A(a[1436]), .B(n11591), .Z(n11593) );
  XOR U3212 ( .A(a[1439]), .B(n11578), .Z(n11580) );
  XOR U3213 ( .A(a[1442]), .B(n11566), .Z(n11568) );
  XOR U3214 ( .A(a[1445]), .B(n11554), .Z(n11556) );
  XOR U3215 ( .A(a[1448]), .B(n11542), .Z(n11544) );
  XOR U3216 ( .A(a[1451]), .B(n11529), .Z(n11531) );
  XOR U3217 ( .A(a[1454]), .B(n11517), .Z(n11519) );
  XOR U3218 ( .A(a[1457]), .B(n11505), .Z(n11507) );
  XOR U3219 ( .A(a[1460]), .B(n11492), .Z(n11494) );
  XOR U3220 ( .A(a[1463]), .B(n11480), .Z(n11482) );
  XOR U3221 ( .A(a[1466]), .B(n11468), .Z(n11470) );
  XOR U3222 ( .A(a[1469]), .B(n11455), .Z(n11457) );
  XOR U3223 ( .A(a[1472]), .B(n11443), .Z(n11445) );
  XOR U3224 ( .A(a[1475]), .B(n11431), .Z(n11433) );
  XOR U3225 ( .A(a[1478]), .B(n11419), .Z(n11421) );
  XOR U3226 ( .A(a[1481]), .B(n11406), .Z(n11408) );
  XOR U3227 ( .A(a[1484]), .B(n11394), .Z(n11396) );
  XOR U3228 ( .A(a[1487]), .B(n11382), .Z(n11384) );
  XOR U3229 ( .A(a[1490]), .B(n11369), .Z(n11371) );
  XOR U3230 ( .A(a[1493]), .B(n11357), .Z(n11359) );
  XOR U3231 ( .A(a[1496]), .B(n11345), .Z(n11347) );
  XOR U3232 ( .A(a[1499]), .B(n11331), .Z(n11333) );
  XOR U3233 ( .A(a[1502]), .B(n11319), .Z(n11321) );
  XOR U3234 ( .A(a[1505]), .B(n11307), .Z(n11309) );
  XOR U3235 ( .A(a[1508]), .B(n11295), .Z(n11297) );
  XOR U3236 ( .A(a[1511]), .B(n11282), .Z(n11284) );
  XOR U3237 ( .A(a[1514]), .B(n11270), .Z(n11272) );
  XOR U3238 ( .A(a[1517]), .B(n11258), .Z(n11260) );
  XOR U3239 ( .A(a[1520]), .B(n11245), .Z(n11247) );
  XOR U3240 ( .A(a[1523]), .B(n11233), .Z(n11235) );
  XOR U3241 ( .A(a[1526]), .B(n11221), .Z(n11223) );
  XOR U3242 ( .A(a[1529]), .B(n11208), .Z(n11210) );
  XOR U3243 ( .A(a[1532]), .B(n11196), .Z(n11198) );
  XOR U3244 ( .A(a[1535]), .B(n11184), .Z(n11186) );
  XOR U3245 ( .A(a[1538]), .B(n11172), .Z(n11174) );
  XOR U3246 ( .A(a[1541]), .B(n11159), .Z(n11161) );
  XOR U3247 ( .A(a[1544]), .B(n11147), .Z(n11149) );
  XOR U3248 ( .A(a[1547]), .B(n11135), .Z(n11137) );
  XOR U3249 ( .A(a[1550]), .B(n11122), .Z(n11124) );
  XOR U3250 ( .A(a[1553]), .B(n11110), .Z(n11112) );
  XOR U3251 ( .A(a[1556]), .B(n11098), .Z(n11100) );
  XOR U3252 ( .A(a[1559]), .B(n11085), .Z(n11087) );
  XOR U3253 ( .A(a[1562]), .B(n11073), .Z(n11075) );
  XOR U3254 ( .A(a[1565]), .B(n11061), .Z(n11063) );
  XOR U3255 ( .A(a[1568]), .B(n11049), .Z(n11051) );
  XOR U3256 ( .A(a[1571]), .B(n11036), .Z(n11038) );
  XOR U3257 ( .A(a[1574]), .B(n11024), .Z(n11026) );
  XOR U3258 ( .A(a[1577]), .B(n11012), .Z(n11014) );
  XOR U3259 ( .A(a[1580]), .B(n10999), .Z(n11001) );
  XOR U3260 ( .A(a[1583]), .B(n10987), .Z(n10989) );
  XOR U3261 ( .A(a[1586]), .B(n10975), .Z(n10977) );
  XOR U3262 ( .A(a[1589]), .B(n10962), .Z(n10964) );
  XOR U3263 ( .A(a[1592]), .B(n10950), .Z(n10952) );
  XOR U3264 ( .A(a[1595]), .B(n10938), .Z(n10940) );
  XOR U3265 ( .A(a[1598]), .B(n10926), .Z(n10928) );
  XOR U3266 ( .A(a[1601]), .B(n10912), .Z(n10914) );
  XOR U3267 ( .A(a[1604]), .B(n10900), .Z(n10902) );
  XOR U3268 ( .A(a[1607]), .B(n10888), .Z(n10890) );
  XOR U3269 ( .A(a[1610]), .B(n10875), .Z(n10877) );
  XOR U3270 ( .A(a[1613]), .B(n10863), .Z(n10865) );
  XOR U3271 ( .A(a[1616]), .B(n10851), .Z(n10853) );
  XOR U3272 ( .A(a[1619]), .B(n10838), .Z(n10840) );
  XOR U3273 ( .A(a[1622]), .B(n10826), .Z(n10828) );
  XOR U3274 ( .A(a[1625]), .B(n10814), .Z(n10816) );
  XOR U3275 ( .A(a[1628]), .B(n10802), .Z(n10804) );
  XOR U3276 ( .A(a[1631]), .B(n10789), .Z(n10791) );
  XOR U3277 ( .A(a[1634]), .B(n10777), .Z(n10779) );
  XOR U3278 ( .A(a[1637]), .B(n10765), .Z(n10767) );
  XOR U3279 ( .A(a[1640]), .B(n10752), .Z(n10754) );
  XOR U3280 ( .A(a[1643]), .B(n10740), .Z(n10742) );
  XOR U3281 ( .A(a[1646]), .B(n10728), .Z(n10730) );
  XOR U3282 ( .A(a[1649]), .B(n10715), .Z(n10717) );
  XOR U3283 ( .A(a[1652]), .B(n10703), .Z(n10705) );
  XOR U3284 ( .A(a[1655]), .B(n10691), .Z(n10693) );
  XOR U3285 ( .A(a[1658]), .B(n10679), .Z(n10681) );
  XOR U3286 ( .A(a[1661]), .B(n10666), .Z(n10668) );
  XOR U3287 ( .A(a[1664]), .B(n10654), .Z(n10656) );
  XOR U3288 ( .A(a[1667]), .B(n10642), .Z(n10644) );
  XOR U3289 ( .A(a[1670]), .B(n10629), .Z(n10631) );
  XOR U3290 ( .A(a[1673]), .B(n10617), .Z(n10619) );
  XOR U3291 ( .A(a[1676]), .B(n10605), .Z(n10607) );
  XOR U3292 ( .A(a[1679]), .B(n10592), .Z(n10594) );
  XOR U3293 ( .A(a[1682]), .B(n10580), .Z(n10582) );
  XOR U3294 ( .A(a[1685]), .B(n10568), .Z(n10570) );
  XOR U3295 ( .A(a[1688]), .B(n10556), .Z(n10558) );
  XOR U3296 ( .A(a[1691]), .B(n10543), .Z(n10545) );
  XOR U3297 ( .A(a[1694]), .B(n10531), .Z(n10533) );
  XOR U3298 ( .A(a[1697]), .B(n10519), .Z(n10521) );
  XOR U3299 ( .A(a[1700]), .B(n10505), .Z(n10507) );
  XOR U3300 ( .A(a[1703]), .B(n10493), .Z(n10495) );
  XOR U3301 ( .A(a[1706]), .B(n10481), .Z(n10483) );
  XOR U3302 ( .A(a[1709]), .B(n10468), .Z(n10470) );
  XOR U3303 ( .A(a[1712]), .B(n10456), .Z(n10458) );
  XOR U3304 ( .A(a[1715]), .B(n10444), .Z(n10446) );
  XOR U3305 ( .A(a[1718]), .B(n10432), .Z(n10434) );
  XOR U3306 ( .A(a[1721]), .B(n10419), .Z(n10421) );
  XOR U3307 ( .A(a[1724]), .B(n10407), .Z(n10409) );
  XOR U3308 ( .A(a[1727]), .B(n10395), .Z(n10397) );
  XOR U3309 ( .A(a[1730]), .B(n10382), .Z(n10384) );
  XOR U3310 ( .A(a[1733]), .B(n10370), .Z(n10372) );
  XOR U3311 ( .A(a[1736]), .B(n10358), .Z(n10360) );
  XOR U3312 ( .A(a[1739]), .B(n10345), .Z(n10347) );
  XOR U3313 ( .A(a[1742]), .B(n10333), .Z(n10335) );
  XOR U3314 ( .A(a[1745]), .B(n10321), .Z(n10323) );
  XOR U3315 ( .A(a[1748]), .B(n10309), .Z(n10311) );
  XOR U3316 ( .A(a[1751]), .B(n10296), .Z(n10298) );
  XOR U3317 ( .A(a[1754]), .B(n10284), .Z(n10286) );
  XOR U3318 ( .A(a[1757]), .B(n10272), .Z(n10274) );
  XOR U3319 ( .A(a[1760]), .B(n10259), .Z(n10261) );
  XOR U3320 ( .A(a[1763]), .B(n10247), .Z(n10249) );
  XOR U3321 ( .A(a[1766]), .B(n10235), .Z(n10237) );
  XOR U3322 ( .A(a[1769]), .B(n10222), .Z(n10224) );
  XOR U3323 ( .A(a[1772]), .B(n10210), .Z(n10212) );
  XOR U3324 ( .A(a[1775]), .B(n10198), .Z(n10200) );
  XOR U3325 ( .A(a[1778]), .B(n10186), .Z(n10188) );
  XOR U3326 ( .A(a[1781]), .B(n10173), .Z(n10175) );
  XOR U3327 ( .A(a[1784]), .B(n10161), .Z(n10163) );
  XOR U3328 ( .A(a[1787]), .B(n10149), .Z(n10151) );
  XOR U3329 ( .A(a[1790]), .B(n10136), .Z(n10138) );
  XOR U3330 ( .A(a[1793]), .B(n10124), .Z(n10126) );
  XOR U3331 ( .A(a[1796]), .B(n10112), .Z(n10114) );
  XOR U3332 ( .A(a[1799]), .B(n10098), .Z(n10100) );
  XOR U3333 ( .A(a[1802]), .B(n10086), .Z(n10088) );
  XOR U3334 ( .A(a[1805]), .B(n10074), .Z(n10076) );
  XOR U3335 ( .A(a[1808]), .B(n10062), .Z(n10064) );
  XOR U3336 ( .A(a[1811]), .B(n10049), .Z(n10051) );
  XOR U3337 ( .A(a[1814]), .B(n10037), .Z(n10039) );
  XOR U3338 ( .A(a[1817]), .B(n10025), .Z(n10027) );
  XOR U3339 ( .A(a[1820]), .B(n10012), .Z(n10014) );
  XOR U3340 ( .A(a[1823]), .B(n10000), .Z(n10002) );
  XOR U3341 ( .A(a[1826]), .B(n9988), .Z(n9990) );
  XOR U3342 ( .A(a[1829]), .B(n9975), .Z(n9977) );
  XOR U3343 ( .A(a[1832]), .B(n9963), .Z(n9965) );
  XOR U3344 ( .A(a[1835]), .B(n9951), .Z(n9953) );
  XOR U3345 ( .A(a[1838]), .B(n9939), .Z(n9941) );
  XOR U3346 ( .A(a[1841]), .B(n9926), .Z(n9928) );
  XOR U3347 ( .A(a[1844]), .B(n9914), .Z(n9916) );
  XOR U3348 ( .A(a[1847]), .B(n9902), .Z(n9904) );
  XOR U3349 ( .A(a[1850]), .B(n9889), .Z(n9891) );
  XOR U3350 ( .A(a[1853]), .B(n9877), .Z(n9879) );
  XOR U3351 ( .A(a[1856]), .B(n9865), .Z(n9867) );
  XOR U3352 ( .A(a[1859]), .B(n9852), .Z(n9854) );
  XOR U3353 ( .A(a[1862]), .B(n9840), .Z(n9842) );
  XOR U3354 ( .A(a[1865]), .B(n9828), .Z(n9830) );
  XOR U3355 ( .A(a[1868]), .B(n9816), .Z(n9818) );
  XOR U3356 ( .A(a[1871]), .B(n9803), .Z(n9805) );
  XOR U3357 ( .A(a[1874]), .B(n9791), .Z(n9793) );
  XOR U3358 ( .A(a[1877]), .B(n9779), .Z(n9781) );
  XOR U3359 ( .A(a[1880]), .B(n9766), .Z(n9768) );
  XOR U3360 ( .A(a[1883]), .B(n9754), .Z(n9756) );
  XOR U3361 ( .A(a[1886]), .B(n9742), .Z(n9744) );
  XOR U3362 ( .A(a[1889]), .B(n9729), .Z(n9731) );
  XOR U3363 ( .A(a[1892]), .B(n9717), .Z(n9719) );
  XOR U3364 ( .A(a[1895]), .B(n9705), .Z(n9707) );
  XOR U3365 ( .A(a[1898]), .B(n9693), .Z(n9695) );
  XOR U3366 ( .A(a[1901]), .B(n9679), .Z(n9681) );
  XOR U3367 ( .A(a[1904]), .B(n9667), .Z(n9669) );
  XOR U3368 ( .A(a[1907]), .B(n9655), .Z(n9657) );
  XOR U3369 ( .A(a[1910]), .B(n9642), .Z(n9644) );
  XOR U3370 ( .A(a[1913]), .B(n9630), .Z(n9632) );
  XOR U3371 ( .A(a[1916]), .B(n9618), .Z(n9620) );
  XOR U3372 ( .A(a[1919]), .B(n9605), .Z(n9607) );
  XOR U3373 ( .A(a[1922]), .B(n9593), .Z(n9595) );
  XOR U3374 ( .A(a[1925]), .B(n9581), .Z(n9583) );
  XOR U3375 ( .A(a[1928]), .B(n9569), .Z(n9571) );
  XOR U3376 ( .A(a[1931]), .B(n9556), .Z(n9558) );
  XOR U3377 ( .A(a[1934]), .B(n9544), .Z(n9546) );
  XOR U3378 ( .A(a[1937]), .B(n9532), .Z(n9534) );
  XOR U3379 ( .A(a[1940]), .B(n9519), .Z(n9521) );
  XOR U3380 ( .A(a[1943]), .B(n9507), .Z(n9509) );
  XOR U3381 ( .A(a[1946]), .B(n9495), .Z(n9497) );
  XOR U3382 ( .A(a[1949]), .B(n9482), .Z(n9484) );
  XOR U3383 ( .A(a[1952]), .B(n9470), .Z(n9472) );
  XOR U3384 ( .A(a[1955]), .B(n9458), .Z(n9460) );
  XOR U3385 ( .A(a[1958]), .B(n9446), .Z(n9448) );
  XOR U3386 ( .A(a[1961]), .B(n9433), .Z(n9435) );
  XOR U3387 ( .A(a[1964]), .B(n9421), .Z(n9423) );
  XOR U3388 ( .A(a[1967]), .B(n9409), .Z(n9411) );
  XOR U3389 ( .A(a[1970]), .B(n9396), .Z(n9398) );
  XOR U3390 ( .A(a[1973]), .B(n9384), .Z(n9386) );
  XOR U3391 ( .A(a[1976]), .B(n9372), .Z(n9374) );
  XOR U3392 ( .A(a[1979]), .B(n9359), .Z(n9361) );
  XOR U3393 ( .A(a[1982]), .B(n9347), .Z(n9349) );
  XOR U3394 ( .A(a[1985]), .B(n9335), .Z(n9337) );
  XOR U3395 ( .A(a[1988]), .B(n9323), .Z(n9325) );
  XOR U3396 ( .A(a[1991]), .B(n9310), .Z(n9312) );
  XOR U3397 ( .A(a[1994]), .B(n9298), .Z(n9300) );
  XOR U3398 ( .A(a[1997]), .B(n9286), .Z(n9288) );
  XOR U3399 ( .A(a[2000]), .B(n9271), .Z(n9273) );
  XOR U3400 ( .A(a[2003]), .B(n9259), .Z(n9261) );
  XOR U3401 ( .A(a[2006]), .B(n9247), .Z(n9249) );
  XOR U3402 ( .A(a[2009]), .B(n9234), .Z(n9236) );
  XOR U3403 ( .A(a[2012]), .B(n9222), .Z(n9224) );
  XOR U3404 ( .A(a[2015]), .B(n9210), .Z(n9212) );
  XOR U3405 ( .A(a[2018]), .B(n9198), .Z(n9200) );
  XOR U3406 ( .A(a[2021]), .B(n9185), .Z(n9187) );
  XOR U3407 ( .A(a[2024]), .B(n9173), .Z(n9175) );
  XOR U3408 ( .A(a[2027]), .B(n9161), .Z(n9163) );
  XOR U3409 ( .A(a[2030]), .B(n9148), .Z(n9150) );
  XOR U3410 ( .A(a[2033]), .B(n9136), .Z(n9138) );
  XOR U3411 ( .A(a[2036]), .B(n9124), .Z(n9126) );
  XOR U3412 ( .A(a[2039]), .B(n9111), .Z(n9113) );
  XOR U3413 ( .A(a[2042]), .B(n9099), .Z(n9101) );
  XOR U3414 ( .A(a[2045]), .B(n9087), .Z(n9089) );
  XOR U3415 ( .A(a[2048]), .B(n9075), .Z(n9077) );
  XOR U3416 ( .A(a[2051]), .B(n9062), .Z(n9064) );
  XOR U3417 ( .A(a[2054]), .B(n9050), .Z(n9052) );
  XOR U3418 ( .A(a[2057]), .B(n9038), .Z(n9040) );
  XOR U3419 ( .A(a[2060]), .B(n9025), .Z(n9027) );
  XOR U3420 ( .A(a[2063]), .B(n9013), .Z(n9015) );
  XOR U3421 ( .A(a[2066]), .B(n9001), .Z(n9003) );
  XOR U3422 ( .A(a[2069]), .B(n8988), .Z(n8990) );
  XOR U3423 ( .A(a[2072]), .B(n8976), .Z(n8978) );
  XOR U3424 ( .A(a[2075]), .B(n8964), .Z(n8966) );
  XOR U3425 ( .A(a[2078]), .B(n8952), .Z(n8954) );
  XOR U3426 ( .A(a[2081]), .B(n8939), .Z(n8941) );
  XOR U3427 ( .A(a[2084]), .B(n8927), .Z(n8929) );
  XOR U3428 ( .A(a[2087]), .B(n8915), .Z(n8917) );
  XOR U3429 ( .A(a[2090]), .B(n8902), .Z(n8904) );
  XOR U3430 ( .A(a[2093]), .B(n8890), .Z(n8892) );
  XOR U3431 ( .A(a[2096]), .B(n8878), .Z(n8880) );
  XOR U3432 ( .A(a[2099]), .B(n8864), .Z(n8866) );
  XOR U3433 ( .A(a[2102]), .B(n8852), .Z(n8854) );
  XOR U3434 ( .A(a[2105]), .B(n8840), .Z(n8842) );
  XOR U3435 ( .A(a[2108]), .B(n8828), .Z(n8830) );
  XOR U3436 ( .A(a[2111]), .B(n8815), .Z(n8817) );
  XOR U3437 ( .A(a[2114]), .B(n8803), .Z(n8805) );
  XOR U3438 ( .A(a[2117]), .B(n8791), .Z(n8793) );
  XOR U3439 ( .A(a[2120]), .B(n8778), .Z(n8780) );
  XOR U3440 ( .A(a[2123]), .B(n8766), .Z(n8768) );
  XOR U3441 ( .A(a[2126]), .B(n8754), .Z(n8756) );
  XOR U3442 ( .A(a[2129]), .B(n8741), .Z(n8743) );
  XOR U3443 ( .A(a[2132]), .B(n8729), .Z(n8731) );
  XOR U3444 ( .A(a[2135]), .B(n8717), .Z(n8719) );
  XOR U3445 ( .A(a[2138]), .B(n8705), .Z(n8707) );
  XOR U3446 ( .A(a[2141]), .B(n8692), .Z(n8694) );
  XOR U3447 ( .A(a[2144]), .B(n8680), .Z(n8682) );
  XOR U3448 ( .A(a[2147]), .B(n8668), .Z(n8670) );
  XOR U3449 ( .A(a[2150]), .B(n8655), .Z(n8657) );
  XOR U3450 ( .A(a[2153]), .B(n8643), .Z(n8645) );
  XOR U3451 ( .A(a[2156]), .B(n8631), .Z(n8633) );
  XOR U3452 ( .A(a[2159]), .B(n8618), .Z(n8620) );
  XOR U3453 ( .A(a[2162]), .B(n8606), .Z(n8608) );
  XOR U3454 ( .A(a[2165]), .B(n8594), .Z(n8596) );
  XOR U3455 ( .A(a[2168]), .B(n8582), .Z(n8584) );
  XOR U3456 ( .A(a[2171]), .B(n8569), .Z(n8571) );
  XOR U3457 ( .A(a[2174]), .B(n8557), .Z(n8559) );
  XOR U3458 ( .A(a[2177]), .B(n8545), .Z(n8547) );
  XOR U3459 ( .A(a[2180]), .B(n8532), .Z(n8534) );
  XOR U3460 ( .A(a[2183]), .B(n8520), .Z(n8522) );
  XOR U3461 ( .A(a[2186]), .B(n8508), .Z(n8510) );
  XOR U3462 ( .A(a[2189]), .B(n8495), .Z(n8497) );
  XOR U3463 ( .A(a[2192]), .B(n8483), .Z(n8485) );
  XOR U3464 ( .A(a[2195]), .B(n8471), .Z(n8473) );
  XOR U3465 ( .A(a[2198]), .B(n8459), .Z(n8461) );
  XOR U3466 ( .A(a[2201]), .B(n8445), .Z(n8447) );
  XOR U3467 ( .A(a[2204]), .B(n8433), .Z(n8435) );
  XOR U3468 ( .A(a[2207]), .B(n8421), .Z(n8423) );
  XOR U3469 ( .A(a[2210]), .B(n8408), .Z(n8410) );
  XOR U3470 ( .A(a[2213]), .B(n8396), .Z(n8398) );
  XOR U3471 ( .A(a[2216]), .B(n8384), .Z(n8386) );
  XOR U3472 ( .A(a[2219]), .B(n8371), .Z(n8373) );
  XOR U3473 ( .A(a[2222]), .B(n8359), .Z(n8361) );
  XOR U3474 ( .A(a[2225]), .B(n8347), .Z(n8349) );
  XOR U3475 ( .A(a[2228]), .B(n8335), .Z(n8337) );
  XOR U3476 ( .A(a[2231]), .B(n8322), .Z(n8324) );
  XOR U3477 ( .A(a[2234]), .B(n8310), .Z(n8312) );
  XOR U3478 ( .A(a[2237]), .B(n8298), .Z(n8300) );
  XOR U3479 ( .A(a[2240]), .B(n8285), .Z(n8287) );
  XOR U3480 ( .A(a[2243]), .B(n8273), .Z(n8275) );
  XOR U3481 ( .A(a[2246]), .B(n8261), .Z(n8263) );
  XOR U3482 ( .A(a[2249]), .B(n8248), .Z(n8250) );
  XOR U3483 ( .A(a[2252]), .B(n8236), .Z(n8238) );
  XOR U3484 ( .A(a[2255]), .B(n8224), .Z(n8226) );
  XOR U3485 ( .A(a[2258]), .B(n8212), .Z(n8214) );
  XOR U3486 ( .A(a[2261]), .B(n8199), .Z(n8201) );
  XOR U3487 ( .A(a[2264]), .B(n8187), .Z(n8189) );
  XOR U3488 ( .A(a[2267]), .B(n8175), .Z(n8177) );
  XOR U3489 ( .A(a[2270]), .B(n8162), .Z(n8164) );
  XOR U3490 ( .A(a[2273]), .B(n8150), .Z(n8152) );
  XOR U3491 ( .A(a[2276]), .B(n8138), .Z(n8140) );
  XOR U3492 ( .A(a[2279]), .B(n8125), .Z(n8127) );
  XOR U3493 ( .A(a[2282]), .B(n8113), .Z(n8115) );
  XOR U3494 ( .A(a[2285]), .B(n8101), .Z(n8103) );
  XOR U3495 ( .A(a[2288]), .B(n8089), .Z(n8091) );
  XOR U3496 ( .A(a[2291]), .B(n8076), .Z(n8078) );
  XOR U3497 ( .A(a[2294]), .B(n8064), .Z(n8066) );
  XOR U3498 ( .A(a[2297]), .B(n8052), .Z(n8054) );
  XOR U3499 ( .A(a[2300]), .B(n8038), .Z(n8040) );
  XOR U3500 ( .A(a[2303]), .B(n8026), .Z(n8028) );
  XOR U3501 ( .A(a[2306]), .B(n8014), .Z(n8016) );
  XOR U3502 ( .A(a[2309]), .B(n8001), .Z(n8003) );
  XOR U3503 ( .A(a[2312]), .B(n7989), .Z(n7991) );
  XOR U3504 ( .A(a[2315]), .B(n7977), .Z(n7979) );
  XOR U3505 ( .A(a[2318]), .B(n7965), .Z(n7967) );
  XOR U3506 ( .A(a[2321]), .B(n7952), .Z(n7954) );
  XOR U3507 ( .A(a[2324]), .B(n7940), .Z(n7942) );
  XOR U3508 ( .A(a[2327]), .B(n7928), .Z(n7930) );
  XOR U3509 ( .A(a[2330]), .B(n7915), .Z(n7917) );
  XOR U3510 ( .A(a[2333]), .B(n7903), .Z(n7905) );
  XOR U3511 ( .A(a[2336]), .B(n7891), .Z(n7893) );
  XOR U3512 ( .A(a[2339]), .B(n7878), .Z(n7880) );
  XOR U3513 ( .A(a[2342]), .B(n7866), .Z(n7868) );
  XOR U3514 ( .A(a[2345]), .B(n7854), .Z(n7856) );
  XOR U3515 ( .A(a[2348]), .B(n7842), .Z(n7844) );
  XOR U3516 ( .A(a[2351]), .B(n7829), .Z(n7831) );
  XOR U3517 ( .A(a[2354]), .B(n7817), .Z(n7819) );
  XOR U3518 ( .A(a[2357]), .B(n7805), .Z(n7807) );
  XOR U3519 ( .A(a[2360]), .B(n7792), .Z(n7794) );
  XOR U3520 ( .A(a[2363]), .B(n7780), .Z(n7782) );
  XOR U3521 ( .A(a[2366]), .B(n7768), .Z(n7770) );
  XOR U3522 ( .A(a[2369]), .B(n7755), .Z(n7757) );
  XOR U3523 ( .A(a[2372]), .B(n7743), .Z(n7745) );
  XOR U3524 ( .A(a[2375]), .B(n7731), .Z(n7733) );
  XOR U3525 ( .A(a[2378]), .B(n7719), .Z(n7721) );
  XOR U3526 ( .A(a[2381]), .B(n7706), .Z(n7708) );
  XOR U3527 ( .A(a[2384]), .B(n7694), .Z(n7696) );
  XOR U3528 ( .A(a[2387]), .B(n7682), .Z(n7684) );
  XOR U3529 ( .A(a[2390]), .B(n7669), .Z(n7671) );
  XOR U3530 ( .A(a[2393]), .B(n7657), .Z(n7659) );
  XOR U3531 ( .A(a[2396]), .B(n7645), .Z(n7647) );
  XOR U3532 ( .A(a[2399]), .B(n7631), .Z(n7633) );
  XOR U3533 ( .A(a[2402]), .B(n7619), .Z(n7621) );
  XOR U3534 ( .A(a[2405]), .B(n7607), .Z(n7609) );
  XOR U3535 ( .A(a[2408]), .B(n7595), .Z(n7597) );
  XOR U3536 ( .A(a[2411]), .B(n7582), .Z(n7584) );
  XOR U3537 ( .A(a[2414]), .B(n7570), .Z(n7572) );
  XOR U3538 ( .A(a[2417]), .B(n7558), .Z(n7560) );
  XOR U3539 ( .A(a[2420]), .B(n7545), .Z(n7547) );
  XOR U3540 ( .A(a[2423]), .B(n7533), .Z(n7535) );
  XOR U3541 ( .A(a[2426]), .B(n7521), .Z(n7523) );
  XOR U3542 ( .A(a[2429]), .B(n7508), .Z(n7510) );
  XOR U3543 ( .A(a[2432]), .B(n7496), .Z(n7498) );
  XOR U3544 ( .A(a[2435]), .B(n7484), .Z(n7486) );
  XOR U3545 ( .A(a[2438]), .B(n7472), .Z(n7474) );
  XOR U3546 ( .A(a[2441]), .B(n7459), .Z(n7461) );
  XOR U3547 ( .A(a[2444]), .B(n7447), .Z(n7449) );
  XOR U3548 ( .A(a[2447]), .B(n7435), .Z(n7437) );
  XOR U3549 ( .A(a[2450]), .B(n7422), .Z(n7424) );
  XOR U3550 ( .A(a[2453]), .B(n7410), .Z(n7412) );
  XOR U3551 ( .A(a[2456]), .B(n7398), .Z(n7400) );
  XOR U3552 ( .A(a[2459]), .B(n7385), .Z(n7387) );
  XOR U3553 ( .A(a[2462]), .B(n7373), .Z(n7375) );
  XOR U3554 ( .A(a[2465]), .B(n7361), .Z(n7363) );
  XOR U3555 ( .A(a[2468]), .B(n7349), .Z(n7351) );
  XOR U3556 ( .A(a[2471]), .B(n7336), .Z(n7338) );
  XOR U3557 ( .A(a[2474]), .B(n7324), .Z(n7326) );
  XOR U3558 ( .A(a[2477]), .B(n7312), .Z(n7314) );
  XOR U3559 ( .A(a[2480]), .B(n7299), .Z(n7301) );
  XOR U3560 ( .A(a[2483]), .B(n7287), .Z(n7289) );
  XOR U3561 ( .A(a[2486]), .B(n7275), .Z(n7277) );
  XOR U3562 ( .A(a[2489]), .B(n7262), .Z(n7264) );
  XOR U3563 ( .A(a[2492]), .B(n7250), .Z(n7252) );
  XOR U3564 ( .A(a[2495]), .B(n7238), .Z(n7240) );
  XOR U3565 ( .A(a[2498]), .B(n7226), .Z(n7228) );
  XOR U3566 ( .A(a[2501]), .B(n7212), .Z(n7214) );
  XOR U3567 ( .A(a[2504]), .B(n7200), .Z(n7202) );
  XOR U3568 ( .A(a[2507]), .B(n7188), .Z(n7190) );
  XOR U3569 ( .A(a[2510]), .B(n7175), .Z(n7177) );
  XOR U3570 ( .A(a[2513]), .B(n7163), .Z(n7165) );
  XOR U3571 ( .A(a[2516]), .B(n7151), .Z(n7153) );
  XOR U3572 ( .A(a[2519]), .B(n7138), .Z(n7140) );
  XOR U3573 ( .A(a[2522]), .B(n7126), .Z(n7128) );
  XOR U3574 ( .A(a[2525]), .B(n7114), .Z(n7116) );
  XOR U3575 ( .A(a[2528]), .B(n7102), .Z(n7104) );
  XOR U3576 ( .A(a[2531]), .B(n7089), .Z(n7091) );
  XOR U3577 ( .A(a[2534]), .B(n7077), .Z(n7079) );
  XOR U3578 ( .A(a[2537]), .B(n7065), .Z(n7067) );
  XOR U3579 ( .A(a[2540]), .B(n7052), .Z(n7054) );
  XOR U3580 ( .A(a[2543]), .B(n7040), .Z(n7042) );
  XOR U3581 ( .A(a[2546]), .B(n7028), .Z(n7030) );
  XOR U3582 ( .A(a[2549]), .B(n7015), .Z(n7017) );
  XOR U3583 ( .A(a[2552]), .B(n7003), .Z(n7005) );
  XOR U3584 ( .A(a[2555]), .B(n6991), .Z(n6993) );
  XOR U3585 ( .A(a[2558]), .B(n6979), .Z(n6981) );
  XOR U3586 ( .A(a[2561]), .B(n6966), .Z(n6968) );
  XOR U3587 ( .A(a[2564]), .B(n6954), .Z(n6956) );
  XOR U3588 ( .A(a[2567]), .B(n6942), .Z(n6944) );
  XOR U3589 ( .A(a[2570]), .B(n6929), .Z(n6931) );
  XOR U3590 ( .A(a[2573]), .B(n6917), .Z(n6919) );
  XOR U3591 ( .A(a[2576]), .B(n6905), .Z(n6907) );
  XOR U3592 ( .A(a[2579]), .B(n6892), .Z(n6894) );
  XOR U3593 ( .A(a[2582]), .B(n6880), .Z(n6882) );
  XOR U3594 ( .A(a[2585]), .B(n6868), .Z(n6870) );
  XOR U3595 ( .A(a[2588]), .B(n6856), .Z(n6858) );
  XOR U3596 ( .A(a[2591]), .B(n6843), .Z(n6845) );
  XOR U3597 ( .A(a[2594]), .B(n6831), .Z(n6833) );
  XOR U3598 ( .A(a[2597]), .B(n6819), .Z(n6821) );
  XOR U3599 ( .A(a[2600]), .B(n6805), .Z(n6807) );
  XOR U3600 ( .A(a[2603]), .B(n6793), .Z(n6795) );
  XOR U3601 ( .A(a[2606]), .B(n6781), .Z(n6783) );
  XOR U3602 ( .A(a[2609]), .B(n6768), .Z(n6770) );
  XOR U3603 ( .A(a[2612]), .B(n6756), .Z(n6758) );
  XOR U3604 ( .A(a[2615]), .B(n6744), .Z(n6746) );
  XOR U3605 ( .A(a[2618]), .B(n6732), .Z(n6734) );
  XOR U3606 ( .A(a[2621]), .B(n6719), .Z(n6721) );
  XOR U3607 ( .A(a[2624]), .B(n6707), .Z(n6709) );
  XOR U3608 ( .A(a[2627]), .B(n6695), .Z(n6697) );
  XOR U3609 ( .A(a[2630]), .B(n6682), .Z(n6684) );
  XOR U3610 ( .A(a[2633]), .B(n6670), .Z(n6672) );
  XOR U3611 ( .A(a[2636]), .B(n6658), .Z(n6660) );
  XOR U3612 ( .A(a[2639]), .B(n6645), .Z(n6647) );
  XOR U3613 ( .A(a[2642]), .B(n6633), .Z(n6635) );
  XOR U3614 ( .A(a[2645]), .B(n6621), .Z(n6623) );
  XOR U3615 ( .A(a[2648]), .B(n6609), .Z(n6611) );
  XOR U3616 ( .A(a[2651]), .B(n6596), .Z(n6598) );
  XOR U3617 ( .A(a[2654]), .B(n6584), .Z(n6586) );
  XOR U3618 ( .A(a[2657]), .B(n6572), .Z(n6574) );
  XOR U3619 ( .A(a[2660]), .B(n6559), .Z(n6561) );
  XOR U3620 ( .A(a[2663]), .B(n6547), .Z(n6549) );
  XOR U3621 ( .A(a[2666]), .B(n6535), .Z(n6537) );
  XOR U3622 ( .A(a[2669]), .B(n6522), .Z(n6524) );
  XOR U3623 ( .A(a[2672]), .B(n6510), .Z(n6512) );
  XOR U3624 ( .A(a[2675]), .B(n6498), .Z(n6500) );
  XOR U3625 ( .A(a[2678]), .B(n6486), .Z(n6488) );
  XOR U3626 ( .A(a[2681]), .B(n6473), .Z(n6475) );
  XOR U3627 ( .A(a[2684]), .B(n6461), .Z(n6463) );
  XOR U3628 ( .A(a[2687]), .B(n6449), .Z(n6451) );
  XOR U3629 ( .A(a[2690]), .B(n6436), .Z(n6438) );
  XOR U3630 ( .A(a[2693]), .B(n6424), .Z(n6426) );
  XOR U3631 ( .A(a[2696]), .B(n6412), .Z(n6414) );
  XOR U3632 ( .A(a[2699]), .B(n6398), .Z(n6400) );
  XOR U3633 ( .A(a[2702]), .B(n6386), .Z(n6388) );
  XOR U3634 ( .A(a[2705]), .B(n6374), .Z(n6376) );
  XOR U3635 ( .A(a[2708]), .B(n6362), .Z(n6364) );
  XOR U3636 ( .A(a[2711]), .B(n6349), .Z(n6351) );
  XOR U3637 ( .A(a[2714]), .B(n6337), .Z(n6339) );
  XOR U3638 ( .A(a[2717]), .B(n6325), .Z(n6327) );
  XOR U3639 ( .A(a[2720]), .B(n6312), .Z(n6314) );
  XOR U3640 ( .A(a[2723]), .B(n6300), .Z(n6302) );
  XOR U3641 ( .A(a[2726]), .B(n6288), .Z(n6290) );
  XOR U3642 ( .A(a[2729]), .B(n6275), .Z(n6277) );
  XOR U3643 ( .A(a[2732]), .B(n6263), .Z(n6265) );
  XOR U3644 ( .A(a[2735]), .B(n6251), .Z(n6253) );
  XOR U3645 ( .A(a[2738]), .B(n6239), .Z(n6241) );
  XOR U3646 ( .A(a[2741]), .B(n6226), .Z(n6228) );
  XOR U3647 ( .A(a[2744]), .B(n6214), .Z(n6216) );
  XOR U3648 ( .A(a[2747]), .B(n6202), .Z(n6204) );
  XOR U3649 ( .A(a[2750]), .B(n6189), .Z(n6191) );
  XOR U3650 ( .A(a[2753]), .B(n6177), .Z(n6179) );
  XOR U3651 ( .A(a[2756]), .B(n6165), .Z(n6167) );
  XOR U3652 ( .A(a[2759]), .B(n6152), .Z(n6154) );
  XOR U3653 ( .A(a[2762]), .B(n6140), .Z(n6142) );
  XOR U3654 ( .A(a[2765]), .B(n6128), .Z(n6130) );
  XOR U3655 ( .A(a[2768]), .B(n6116), .Z(n6118) );
  XOR U3656 ( .A(a[2771]), .B(n6103), .Z(n6105) );
  XOR U3657 ( .A(a[2774]), .B(n6091), .Z(n6093) );
  XOR U3658 ( .A(a[2777]), .B(n6079), .Z(n6081) );
  XOR U3659 ( .A(a[2780]), .B(n6066), .Z(n6068) );
  XOR U3660 ( .A(a[2783]), .B(n6054), .Z(n6056) );
  XOR U3661 ( .A(a[2786]), .B(n6042), .Z(n6044) );
  XOR U3662 ( .A(a[2789]), .B(n6029), .Z(n6031) );
  XOR U3663 ( .A(a[2792]), .B(n6017), .Z(n6019) );
  XOR U3664 ( .A(a[2795]), .B(n6005), .Z(n6007) );
  XOR U3665 ( .A(a[2798]), .B(n5993), .Z(n5995) );
  XOR U3666 ( .A(a[2801]), .B(n5979), .Z(n5981) );
  XOR U3667 ( .A(a[2804]), .B(n5967), .Z(n5969) );
  XOR U3668 ( .A(a[2807]), .B(n5955), .Z(n5957) );
  XOR U3669 ( .A(a[2810]), .B(n5942), .Z(n5944) );
  XOR U3670 ( .A(a[2813]), .B(n5930), .Z(n5932) );
  XOR U3671 ( .A(a[2816]), .B(n5918), .Z(n5920) );
  XOR U3672 ( .A(a[2819]), .B(n5905), .Z(n5907) );
  XOR U3673 ( .A(a[2822]), .B(n5893), .Z(n5895) );
  XOR U3674 ( .A(a[2825]), .B(n5881), .Z(n5883) );
  XOR U3675 ( .A(a[2828]), .B(n5869), .Z(n5871) );
  XOR U3676 ( .A(a[2831]), .B(n5856), .Z(n5858) );
  XOR U3677 ( .A(a[2834]), .B(n5844), .Z(n5846) );
  XOR U3678 ( .A(a[2837]), .B(n5832), .Z(n5834) );
  XOR U3679 ( .A(a[2840]), .B(n5819), .Z(n5821) );
  XOR U3680 ( .A(a[2843]), .B(n5807), .Z(n5809) );
  XOR U3681 ( .A(a[2846]), .B(n5795), .Z(n5797) );
  XOR U3682 ( .A(a[2849]), .B(n5782), .Z(n5784) );
  XOR U3683 ( .A(a[2852]), .B(n5770), .Z(n5772) );
  XOR U3684 ( .A(a[2855]), .B(n5758), .Z(n5760) );
  XOR U3685 ( .A(a[2858]), .B(n5746), .Z(n5748) );
  XOR U3686 ( .A(a[2861]), .B(n5733), .Z(n5735) );
  XOR U3687 ( .A(a[2864]), .B(n5721), .Z(n5723) );
  XOR U3688 ( .A(a[2867]), .B(n5709), .Z(n5711) );
  XOR U3689 ( .A(a[2870]), .B(n5696), .Z(n5698) );
  XOR U3690 ( .A(a[2873]), .B(n5684), .Z(n5686) );
  XOR U3691 ( .A(a[2876]), .B(n5672), .Z(n5674) );
  XOR U3692 ( .A(a[2879]), .B(n5659), .Z(n5661) );
  XOR U3693 ( .A(a[2882]), .B(n5647), .Z(n5649) );
  XOR U3694 ( .A(a[2885]), .B(n5635), .Z(n5637) );
  XOR U3695 ( .A(a[2888]), .B(n5623), .Z(n5625) );
  XOR U3696 ( .A(a[2891]), .B(n5610), .Z(n5612) );
  XOR U3697 ( .A(a[2894]), .B(n5598), .Z(n5600) );
  XOR U3698 ( .A(a[2897]), .B(n5586), .Z(n5588) );
  XOR U3699 ( .A(a[2900]), .B(n5572), .Z(n5574) );
  XOR U3700 ( .A(a[2903]), .B(n5560), .Z(n5562) );
  XOR U3701 ( .A(a[2906]), .B(n5548), .Z(n5550) );
  XOR U3702 ( .A(a[2909]), .B(n5535), .Z(n5537) );
  XOR U3703 ( .A(a[2912]), .B(n5523), .Z(n5525) );
  XOR U3704 ( .A(a[2915]), .B(n5511), .Z(n5513) );
  XOR U3705 ( .A(a[2918]), .B(n5499), .Z(n5501) );
  XOR U3706 ( .A(a[2921]), .B(n5486), .Z(n5488) );
  XOR U3707 ( .A(a[2924]), .B(n5474), .Z(n5476) );
  XOR U3708 ( .A(a[2927]), .B(n5462), .Z(n5464) );
  XOR U3709 ( .A(a[2930]), .B(n5449), .Z(n5451) );
  XOR U3710 ( .A(a[2933]), .B(n5437), .Z(n5439) );
  XOR U3711 ( .A(a[2936]), .B(n5425), .Z(n5427) );
  XOR U3712 ( .A(a[2939]), .B(n5412), .Z(n5414) );
  XOR U3713 ( .A(a[2942]), .B(n5400), .Z(n5402) );
  XOR U3714 ( .A(a[2945]), .B(n5388), .Z(n5390) );
  XOR U3715 ( .A(a[2948]), .B(n5376), .Z(n5378) );
  XOR U3716 ( .A(a[2951]), .B(n5363), .Z(n5365) );
  XOR U3717 ( .A(a[2954]), .B(n5351), .Z(n5353) );
  XOR U3718 ( .A(a[2957]), .B(n5339), .Z(n5341) );
  XOR U3719 ( .A(a[2960]), .B(n5326), .Z(n5328) );
  XOR U3720 ( .A(a[2963]), .B(n5314), .Z(n5316) );
  XOR U3721 ( .A(a[2966]), .B(n5302), .Z(n5304) );
  XOR U3722 ( .A(a[2969]), .B(n5289), .Z(n5291) );
  XOR U3723 ( .A(a[2972]), .B(n5277), .Z(n5279) );
  XOR U3724 ( .A(a[2975]), .B(n5265), .Z(n5267) );
  XOR U3725 ( .A(a[2978]), .B(n5253), .Z(n5255) );
  XOR U3726 ( .A(a[2981]), .B(n5240), .Z(n5242) );
  XOR U3727 ( .A(a[2984]), .B(n5228), .Z(n5230) );
  XOR U3728 ( .A(a[2987]), .B(n5216), .Z(n5218) );
  XOR U3729 ( .A(a[2990]), .B(n5203), .Z(n5205) );
  XOR U3730 ( .A(a[2993]), .B(n5191), .Z(n5193) );
  XOR U3731 ( .A(a[2996]), .B(n5179), .Z(n5181) );
  XOR U3732 ( .A(a[2999]), .B(n5164), .Z(n5166) );
  XOR U3733 ( .A(a[3002]), .B(n5152), .Z(n5154) );
  XOR U3734 ( .A(a[3005]), .B(n5140), .Z(n5142) );
  XOR U3735 ( .A(a[3008]), .B(n5128), .Z(n5130) );
  XOR U3736 ( .A(a[3011]), .B(n5115), .Z(n5117) );
  XOR U3737 ( .A(a[3014]), .B(n5103), .Z(n5105) );
  XOR U3738 ( .A(a[3017]), .B(n5091), .Z(n5093) );
  XOR U3739 ( .A(a[3020]), .B(n5078), .Z(n5080) );
  XOR U3740 ( .A(a[3023]), .B(n5066), .Z(n5068) );
  XOR U3741 ( .A(a[3026]), .B(n5054), .Z(n5056) );
  XOR U3742 ( .A(a[3029]), .B(n5041), .Z(n5043) );
  XOR U3743 ( .A(a[3032]), .B(n5029), .Z(n5031) );
  XOR U3744 ( .A(a[3035]), .B(n5017), .Z(n5019) );
  XOR U3745 ( .A(a[3038]), .B(n5005), .Z(n5007) );
  XOR U3746 ( .A(a[3041]), .B(n4992), .Z(n4994) );
  XOR U3747 ( .A(a[3044]), .B(n4980), .Z(n4982) );
  XOR U3748 ( .A(a[3047]), .B(n4968), .Z(n4970) );
  XOR U3749 ( .A(a[3050]), .B(n4955), .Z(n4957) );
  XOR U3750 ( .A(a[3053]), .B(n4943), .Z(n4945) );
  XOR U3751 ( .A(a[3056]), .B(n4931), .Z(n4933) );
  XOR U3752 ( .A(a[3059]), .B(n4918), .Z(n4920) );
  XOR U3753 ( .A(a[3062]), .B(n4906), .Z(n4908) );
  XOR U3754 ( .A(a[3065]), .B(n4894), .Z(n4896) );
  XOR U3755 ( .A(a[3068]), .B(n4882), .Z(n4884) );
  XOR U3756 ( .A(a[3071]), .B(n4869), .Z(n4871) );
  XOR U3757 ( .A(a[3074]), .B(n4857), .Z(n4859) );
  XOR U3758 ( .A(a[3077]), .B(n4845), .Z(n4847) );
  XOR U3759 ( .A(a[3080]), .B(n4832), .Z(n4834) );
  XOR U3760 ( .A(a[3083]), .B(n4820), .Z(n4822) );
  XOR U3761 ( .A(a[3086]), .B(n4808), .Z(n4810) );
  XOR U3762 ( .A(a[3089]), .B(n4795), .Z(n4797) );
  XOR U3763 ( .A(a[3092]), .B(n4783), .Z(n4785) );
  XOR U3764 ( .A(a[3095]), .B(n4771), .Z(n4773) );
  XOR U3765 ( .A(a[3098]), .B(n4759), .Z(n4761) );
  XOR U3766 ( .A(a[3101]), .B(n4745), .Z(n4747) );
  XOR U3767 ( .A(a[3104]), .B(n4733), .Z(n4735) );
  XOR U3768 ( .A(a[3107]), .B(n4721), .Z(n4723) );
  XOR U3769 ( .A(a[3110]), .B(n4708), .Z(n4710) );
  XOR U3770 ( .A(a[3113]), .B(n4696), .Z(n4698) );
  XOR U3771 ( .A(a[3116]), .B(n4684), .Z(n4686) );
  XOR U3772 ( .A(a[3119]), .B(n4671), .Z(n4673) );
  XOR U3773 ( .A(a[3122]), .B(n4659), .Z(n4661) );
  XOR U3774 ( .A(a[3125]), .B(n4647), .Z(n4649) );
  XOR U3775 ( .A(a[3128]), .B(n4635), .Z(n4637) );
  XOR U3776 ( .A(a[3131]), .B(n4622), .Z(n4624) );
  XOR U3777 ( .A(a[3134]), .B(n4610), .Z(n4612) );
  XOR U3778 ( .A(a[3137]), .B(n4598), .Z(n4600) );
  XOR U3779 ( .A(a[3140]), .B(n4585), .Z(n4587) );
  XOR U3780 ( .A(a[3143]), .B(n4573), .Z(n4575) );
  XOR U3781 ( .A(a[3146]), .B(n4561), .Z(n4563) );
  XOR U3782 ( .A(a[3149]), .B(n4548), .Z(n4550) );
  XOR U3783 ( .A(a[3152]), .B(n4536), .Z(n4538) );
  XOR U3784 ( .A(a[3155]), .B(n4524), .Z(n4526) );
  XOR U3785 ( .A(a[3158]), .B(n4512), .Z(n4514) );
  XOR U3786 ( .A(a[3161]), .B(n4499), .Z(n4501) );
  XOR U3787 ( .A(a[3164]), .B(n4487), .Z(n4489) );
  XOR U3788 ( .A(a[3167]), .B(n4475), .Z(n4477) );
  XOR U3789 ( .A(a[3170]), .B(n4462), .Z(n4464) );
  XOR U3790 ( .A(a[3173]), .B(n4450), .Z(n4452) );
  XOR U3791 ( .A(a[3176]), .B(n4438), .Z(n4440) );
  XOR U3792 ( .A(a[3179]), .B(n4425), .Z(n4427) );
  XOR U3793 ( .A(a[3182]), .B(n4413), .Z(n4415) );
  XOR U3794 ( .A(a[3185]), .B(n4401), .Z(n4403) );
  XOR U3795 ( .A(a[3188]), .B(n4389), .Z(n4391) );
  XOR U3796 ( .A(a[3191]), .B(n4376), .Z(n4378) );
  XOR U3797 ( .A(a[3194]), .B(n4364), .Z(n4366) );
  XOR U3798 ( .A(a[3197]), .B(n4352), .Z(n4354) );
  XOR U3799 ( .A(a[3200]), .B(n4338), .Z(n4340) );
  XOR U3800 ( .A(a[3203]), .B(n4326), .Z(n4328) );
  XOR U3801 ( .A(a[3206]), .B(n4314), .Z(n4316) );
  XOR U3802 ( .A(a[3209]), .B(n4301), .Z(n4303) );
  XOR U3803 ( .A(a[3212]), .B(n4289), .Z(n4291) );
  XOR U3804 ( .A(a[3215]), .B(n4277), .Z(n4279) );
  XOR U3805 ( .A(a[3218]), .B(n4265), .Z(n4267) );
  XOR U3806 ( .A(a[3221]), .B(n4252), .Z(n4254) );
  XOR U3807 ( .A(a[3224]), .B(n4240), .Z(n4242) );
  XOR U3808 ( .A(a[3227]), .B(n4228), .Z(n4230) );
  XOR U3809 ( .A(a[3230]), .B(n4215), .Z(n4217) );
  XOR U3810 ( .A(a[3233]), .B(n4203), .Z(n4205) );
  XOR U3811 ( .A(a[3236]), .B(n4191), .Z(n4193) );
  XOR U3812 ( .A(a[3239]), .B(n4178), .Z(n4180) );
  XOR U3813 ( .A(a[3242]), .B(n4166), .Z(n4168) );
  XOR U3814 ( .A(a[3245]), .B(n4154), .Z(n4156) );
  XOR U3815 ( .A(a[3248]), .B(n4142), .Z(n4144) );
  XOR U3816 ( .A(a[3251]), .B(n4129), .Z(n4131) );
  XOR U3817 ( .A(a[3254]), .B(n4117), .Z(n4119) );
  XOR U3818 ( .A(a[3257]), .B(n4105), .Z(n4107) );
  XOR U3819 ( .A(a[3260]), .B(n4092), .Z(n4094) );
  XOR U3820 ( .A(a[3263]), .B(n4080), .Z(n4082) );
  XOR U3821 ( .A(a[3266]), .B(n4068), .Z(n4070) );
  XOR U3822 ( .A(a[3269]), .B(n4055), .Z(n4057) );
  XOR U3823 ( .A(a[3272]), .B(n4043), .Z(n4045) );
  XOR U3824 ( .A(a[3275]), .B(n4031), .Z(n4033) );
  XOR U3825 ( .A(a[3278]), .B(n4019), .Z(n4021) );
  XOR U3826 ( .A(a[3281]), .B(n4006), .Z(n4008) );
  XOR U3827 ( .A(a[3284]), .B(n3994), .Z(n3996) );
  XOR U3828 ( .A(a[3287]), .B(n3982), .Z(n3984) );
  XOR U3829 ( .A(a[3290]), .B(n3969), .Z(n3971) );
  XOR U3830 ( .A(a[3293]), .B(n3957), .Z(n3959) );
  XOR U3831 ( .A(a[3296]), .B(n3945), .Z(n3947) );
  XOR U3832 ( .A(a[3299]), .B(n3931), .Z(n3933) );
  XOR U3833 ( .A(a[3302]), .B(n3919), .Z(n3921) );
  XOR U3834 ( .A(a[3305]), .B(n3907), .Z(n3909) );
  XOR U3835 ( .A(a[3308]), .B(n3895), .Z(n3897) );
  XOR U3836 ( .A(a[3311]), .B(n3882), .Z(n3884) );
  XOR U3837 ( .A(a[3314]), .B(n3870), .Z(n3872) );
  XOR U3838 ( .A(a[3317]), .B(n3858), .Z(n3860) );
  XOR U3839 ( .A(a[3320]), .B(n3845), .Z(n3847) );
  XOR U3840 ( .A(a[3323]), .B(n3833), .Z(n3835) );
  XOR U3841 ( .A(a[3326]), .B(n3821), .Z(n3823) );
  XOR U3842 ( .A(a[3329]), .B(n3808), .Z(n3810) );
  XOR U3843 ( .A(a[3332]), .B(n3796), .Z(n3798) );
  XOR U3844 ( .A(a[3335]), .B(n3784), .Z(n3786) );
  XOR U3845 ( .A(a[3338]), .B(n3772), .Z(n3774) );
  XOR U3846 ( .A(a[3341]), .B(n3759), .Z(n3761) );
  XOR U3847 ( .A(a[3344]), .B(n3747), .Z(n3749) );
  XOR U3848 ( .A(a[3347]), .B(n3735), .Z(n3737) );
  XOR U3849 ( .A(a[3350]), .B(n3722), .Z(n3724) );
  XOR U3850 ( .A(a[3353]), .B(n3710), .Z(n3712) );
  XOR U3851 ( .A(a[3356]), .B(n3698), .Z(n3700) );
  XOR U3852 ( .A(a[3359]), .B(n3685), .Z(n3687) );
  XOR U3853 ( .A(a[3362]), .B(n3673), .Z(n3675) );
  XOR U3854 ( .A(a[3365]), .B(n3661), .Z(n3663) );
  XOR U3855 ( .A(a[3368]), .B(n3649), .Z(n3651) );
  XOR U3856 ( .A(a[3371]), .B(n3636), .Z(n3638) );
  XOR U3857 ( .A(a[3374]), .B(n3624), .Z(n3626) );
  XOR U3858 ( .A(a[3377]), .B(n3612), .Z(n3614) );
  XOR U3859 ( .A(a[3380]), .B(n3599), .Z(n3601) );
  XOR U3860 ( .A(a[3383]), .B(n3587), .Z(n3589) );
  XOR U3861 ( .A(a[3386]), .B(n3575), .Z(n3577) );
  XOR U3862 ( .A(a[3389]), .B(n3562), .Z(n3564) );
  XOR U3863 ( .A(a[3392]), .B(n3550), .Z(n3552) );
  XOR U3864 ( .A(a[3395]), .B(n3538), .Z(n3540) );
  XOR U3865 ( .A(a[3398]), .B(n3526), .Z(n3528) );
  XOR U3866 ( .A(a[3401]), .B(n3512), .Z(n3514) );
  XOR U3867 ( .A(a[3404]), .B(n3500), .Z(n3502) );
  XOR U3868 ( .A(a[3407]), .B(n3488), .Z(n3490) );
  XOR U3869 ( .A(a[3410]), .B(n3475), .Z(n3477) );
  XOR U3870 ( .A(a[3413]), .B(n3463), .Z(n3465) );
  XOR U3871 ( .A(a[3416]), .B(n3451), .Z(n3453) );
  XOR U3872 ( .A(a[3419]), .B(n3438), .Z(n3440) );
  XOR U3873 ( .A(a[3422]), .B(n3426), .Z(n3428) );
  XOR U3874 ( .A(a[3425]), .B(n3414), .Z(n3416) );
  XOR U3875 ( .A(a[3428]), .B(n3402), .Z(n3404) );
  XOR U3876 ( .A(a[3431]), .B(n3389), .Z(n3391) );
  XOR U3877 ( .A(a[3434]), .B(n3377), .Z(n3379) );
  XOR U3878 ( .A(a[3437]), .B(n3365), .Z(n3367) );
  XOR U3879 ( .A(a[3440]), .B(n3352), .Z(n3354) );
  XOR U3880 ( .A(a[3443]), .B(n3340), .Z(n3342) );
  XOR U3881 ( .A(a[3446]), .B(n3328), .Z(n3330) );
  XOR U3882 ( .A(a[3449]), .B(n3315), .Z(n3317) );
  XOR U3883 ( .A(a[3452]), .B(n3303), .Z(n3305) );
  XOR U3884 ( .A(a[3455]), .B(n3291), .Z(n3293) );
  XOR U3885 ( .A(a[3458]), .B(n3279), .Z(n3281) );
  XOR U3886 ( .A(a[3461]), .B(n3266), .Z(n3268) );
  XOR U3887 ( .A(a[3464]), .B(n3254), .Z(n3256) );
  XOR U3888 ( .A(a[3467]), .B(n3242), .Z(n3244) );
  XOR U3889 ( .A(a[3470]), .B(n3229), .Z(n3231) );
  XOR U3890 ( .A(a[3473]), .B(n3217), .Z(n3219) );
  XOR U3891 ( .A(a[3476]), .B(n3205), .Z(n3207) );
  XOR U3892 ( .A(a[3479]), .B(n3192), .Z(n3194) );
  XOR U3893 ( .A(a[3482]), .B(n3180), .Z(n3182) );
  XOR U3894 ( .A(a[3485]), .B(n3168), .Z(n3170) );
  XOR U3895 ( .A(a[3488]), .B(n3156), .Z(n3158) );
  XOR U3896 ( .A(a[3491]), .B(n3143), .Z(n3145) );
  XOR U3897 ( .A(a[3494]), .B(n3131), .Z(n3133) );
  XOR U3898 ( .A(a[3497]), .B(n3119), .Z(n3121) );
  XOR U3899 ( .A(a[3500]), .B(n3105), .Z(n3107) );
  XOR U3900 ( .A(a[3503]), .B(n3093), .Z(n3095) );
  XOR U3901 ( .A(a[3506]), .B(n3081), .Z(n3083) );
  XOR U3902 ( .A(a[3509]), .B(n3068), .Z(n3070) );
  XOR U3903 ( .A(a[3512]), .B(n3056), .Z(n3058) );
  XOR U3904 ( .A(a[3515]), .B(n3044), .Z(n3046) );
  XOR U3905 ( .A(a[3518]), .B(n3032), .Z(n3034) );
  XOR U3906 ( .A(a[3521]), .B(n3019), .Z(n3021) );
  XOR U3907 ( .A(a[3524]), .B(n3007), .Z(n3009) );
  XOR U3908 ( .A(a[3527]), .B(n2995), .Z(n2997) );
  XOR U3909 ( .A(a[3530]), .B(n2982), .Z(n2984) );
  XOR U3910 ( .A(a[3533]), .B(n2970), .Z(n2972) );
  XOR U3911 ( .A(a[3536]), .B(n2958), .Z(n2960) );
  XOR U3912 ( .A(a[3539]), .B(n2945), .Z(n2947) );
  XOR U3913 ( .A(a[3542]), .B(n2933), .Z(n2935) );
  XOR U3914 ( .A(a[3545]), .B(n2921), .Z(n2923) );
  XOR U3915 ( .A(a[3548]), .B(n2909), .Z(n2911) );
  XOR U3916 ( .A(a[3551]), .B(n2896), .Z(n2898) );
  XOR U3917 ( .A(a[3554]), .B(n2884), .Z(n2886) );
  XOR U3918 ( .A(a[3557]), .B(n2872), .Z(n2874) );
  XOR U3919 ( .A(a[3560]), .B(n2859), .Z(n2861) );
  XOR U3920 ( .A(a[3563]), .B(n2847), .Z(n2849) );
  XOR U3921 ( .A(a[3566]), .B(n2835), .Z(n2837) );
  XOR U3922 ( .A(a[3569]), .B(n2822), .Z(n2824) );
  XOR U3923 ( .A(a[3572]), .B(n2810), .Z(n2812) );
  XOR U3924 ( .A(a[3575]), .B(n2798), .Z(n2800) );
  XOR U3925 ( .A(a[3578]), .B(n2786), .Z(n2788) );
  XOR U3926 ( .A(a[3581]), .B(n2773), .Z(n2775) );
  XOR U3927 ( .A(a[3584]), .B(n2761), .Z(n2763) );
  XOR U3928 ( .A(a[3587]), .B(n2749), .Z(n2751) );
  XOR U3929 ( .A(a[3590]), .B(n2736), .Z(n2738) );
  XOR U3930 ( .A(a[3593]), .B(n2724), .Z(n2726) );
  XOR U3931 ( .A(a[3596]), .B(n2712), .Z(n2714) );
  XOR U3932 ( .A(a[3599]), .B(n2698), .Z(n2700) );
  XOR U3933 ( .A(a[3602]), .B(n2686), .Z(n2688) );
  XOR U3934 ( .A(a[3605]), .B(n2674), .Z(n2676) );
  XOR U3935 ( .A(a[3608]), .B(n2662), .Z(n2664) );
  XOR U3936 ( .A(a[3611]), .B(n2649), .Z(n2651) );
  XOR U3937 ( .A(a[3614]), .B(n2637), .Z(n2639) );
  XOR U3938 ( .A(a[3617]), .B(n2625), .Z(n2627) );
  XOR U3939 ( .A(a[3620]), .B(n2612), .Z(n2614) );
  XOR U3940 ( .A(a[3623]), .B(n2600), .Z(n2602) );
  XOR U3941 ( .A(a[3626]), .B(n2588), .Z(n2590) );
  XOR U3942 ( .A(a[3629]), .B(n2575), .Z(n2577) );
  XOR U3943 ( .A(a[3632]), .B(n2563), .Z(n2565) );
  XOR U3944 ( .A(a[3635]), .B(n2551), .Z(n2553) );
  XOR U3945 ( .A(a[3638]), .B(n2539), .Z(n2541) );
  XOR U3946 ( .A(a[3641]), .B(n2526), .Z(n2528) );
  XOR U3947 ( .A(a[3644]), .B(n2514), .Z(n2516) );
  XOR U3948 ( .A(a[3647]), .B(n2502), .Z(n2504) );
  XOR U3949 ( .A(a[3650]), .B(n2489), .Z(n2491) );
  XOR U3950 ( .A(a[3653]), .B(n2477), .Z(n2479) );
  XOR U3951 ( .A(a[3656]), .B(n2465), .Z(n2467) );
  XOR U3952 ( .A(a[3659]), .B(n2452), .Z(n2454) );
  XOR U3953 ( .A(a[3662]), .B(n2440), .Z(n2442) );
  XOR U3954 ( .A(a[3665]), .B(n2428), .Z(n2430) );
  XOR U3955 ( .A(a[3668]), .B(n2416), .Z(n2418) );
  XOR U3956 ( .A(a[3671]), .B(n2403), .Z(n2405) );
  XOR U3957 ( .A(a[3674]), .B(n2391), .Z(n2393) );
  XOR U3958 ( .A(a[3677]), .B(n2379), .Z(n2381) );
  XOR U3959 ( .A(a[3680]), .B(n2366), .Z(n2368) );
  XOR U3960 ( .A(a[3683]), .B(n2354), .Z(n2356) );
  XOR U3961 ( .A(a[3686]), .B(n2342), .Z(n2344) );
  XOR U3962 ( .A(a[3689]), .B(n2329), .Z(n2331) );
  XOR U3963 ( .A(a[3692]), .B(n2317), .Z(n2319) );
  XOR U3964 ( .A(a[3695]), .B(n2305), .Z(n2307) );
  XOR U3965 ( .A(a[3698]), .B(n2293), .Z(n2295) );
  XOR U3966 ( .A(a[3701]), .B(n2279), .Z(n2281) );
  XOR U3967 ( .A(a[3704]), .B(n2267), .Z(n2269) );
  XOR U3968 ( .A(a[3707]), .B(n2255), .Z(n2257) );
  XOR U3969 ( .A(a[3710]), .B(n2242), .Z(n2244) );
  XOR U3970 ( .A(a[3713]), .B(n2230), .Z(n2232) );
  XOR U3971 ( .A(a[3716]), .B(n2218), .Z(n2220) );
  XOR U3972 ( .A(a[3719]), .B(n2205), .Z(n2207) );
  XOR U3973 ( .A(a[3722]), .B(n2193), .Z(n2195) );
  XOR U3974 ( .A(a[3725]), .B(n2181), .Z(n2183) );
  XOR U3975 ( .A(a[3728]), .B(n2169), .Z(n2171) );
  XOR U3976 ( .A(a[3731]), .B(n2156), .Z(n2158) );
  XOR U3977 ( .A(a[3734]), .B(n2144), .Z(n2146) );
  XOR U3978 ( .A(a[3737]), .B(n2132), .Z(n2134) );
  XOR U3979 ( .A(a[3740]), .B(n2119), .Z(n2121) );
  XOR U3980 ( .A(a[3743]), .B(n2107), .Z(n2109) );
  XOR U3981 ( .A(a[3746]), .B(n2095), .Z(n2097) );
  XOR U3982 ( .A(a[3749]), .B(n2082), .Z(n2084) );
  XOR U3983 ( .A(a[3752]), .B(n2070), .Z(n2072) );
  XOR U3984 ( .A(a[3755]), .B(n2058), .Z(n2060) );
  XOR U3985 ( .A(a[3758]), .B(n2046), .Z(n2048) );
  XOR U3986 ( .A(a[3761]), .B(n2033), .Z(n2035) );
  XOR U3987 ( .A(a[3764]), .B(n2021), .Z(n2023) );
  XOR U3988 ( .A(a[3767]), .B(n2009), .Z(n2011) );
  XOR U3989 ( .A(a[3770]), .B(n1996), .Z(n1998) );
  XOR U3990 ( .A(a[3773]), .B(n1984), .Z(n1986) );
  XOR U3991 ( .A(a[3776]), .B(n1972), .Z(n1974) );
  XOR U3992 ( .A(a[3779]), .B(n1959), .Z(n1961) );
  XOR U3993 ( .A(a[3782]), .B(n1947), .Z(n1949) );
  XOR U3994 ( .A(a[3785]), .B(n1935), .Z(n1937) );
  XOR U3995 ( .A(a[3788]), .B(n1923), .Z(n1925) );
  XOR U3996 ( .A(a[3791]), .B(n1910), .Z(n1912) );
  XOR U3997 ( .A(a[3794]), .B(n1898), .Z(n1900) );
  XOR U3998 ( .A(a[3797]), .B(n1886), .Z(n1888) );
  XOR U3999 ( .A(a[3800]), .B(n1872), .Z(n1874) );
  XOR U4000 ( .A(a[3803]), .B(n1860), .Z(n1862) );
  XOR U4001 ( .A(a[3806]), .B(n1848), .Z(n1850) );
  XOR U4002 ( .A(a[3809]), .B(n1835), .Z(n1837) );
  XOR U4003 ( .A(a[3812]), .B(n1823), .Z(n1825) );
  XOR U4004 ( .A(a[3815]), .B(n1811), .Z(n1813) );
  XOR U4005 ( .A(a[3818]), .B(n1799), .Z(n1801) );
  XOR U4006 ( .A(a[3821]), .B(n1786), .Z(n1788) );
  XOR U4007 ( .A(a[3824]), .B(n1774), .Z(n1776) );
  XOR U4008 ( .A(a[3827]), .B(n1762), .Z(n1764) );
  XOR U4009 ( .A(a[3830]), .B(n1749), .Z(n1751) );
  XOR U4010 ( .A(a[3833]), .B(n1737), .Z(n1739) );
  XOR U4011 ( .A(a[3836]), .B(n1725), .Z(n1727) );
  XOR U4012 ( .A(a[3839]), .B(n1712), .Z(n1714) );
  XOR U4013 ( .A(a[3842]), .B(n1700), .Z(n1702) );
  XOR U4014 ( .A(a[3845]), .B(n1688), .Z(n1690) );
  XOR U4015 ( .A(a[3848]), .B(n1676), .Z(n1678) );
  XOR U4016 ( .A(a[3851]), .B(n1663), .Z(n1665) );
  XOR U4017 ( .A(a[3854]), .B(n1651), .Z(n1653) );
  XOR U4018 ( .A(a[3857]), .B(n1639), .Z(n1641) );
  XOR U4019 ( .A(a[3860]), .B(n1626), .Z(n1628) );
  XOR U4020 ( .A(a[3863]), .B(n1614), .Z(n1616) );
  XOR U4021 ( .A(a[3866]), .B(n1602), .Z(n1604) );
  XOR U4022 ( .A(a[3869]), .B(n1589), .Z(n1591) );
  XOR U4023 ( .A(a[3872]), .B(n1577), .Z(n1579) );
  XOR U4024 ( .A(a[3875]), .B(n1565), .Z(n1567) );
  XOR U4025 ( .A(a[3878]), .B(n1553), .Z(n1555) );
  XOR U4026 ( .A(a[3881]), .B(n1540), .Z(n1542) );
  XOR U4027 ( .A(a[3884]), .B(n1528), .Z(n1530) );
  XOR U4028 ( .A(a[3887]), .B(n1516), .Z(n1518) );
  XOR U4029 ( .A(a[3890]), .B(n1503), .Z(n1505) );
  XOR U4030 ( .A(a[3893]), .B(n1491), .Z(n1493) );
  XOR U4031 ( .A(a[3896]), .B(n1479), .Z(n1481) );
  XOR U4032 ( .A(a[3899]), .B(n1465), .Z(n1467) );
  XOR U4033 ( .A(a[3902]), .B(n1453), .Z(n1455) );
  XOR U4034 ( .A(a[3905]), .B(n1441), .Z(n1443) );
  XOR U4035 ( .A(a[3908]), .B(n1429), .Z(n1431) );
  XOR U4036 ( .A(a[3911]), .B(n1416), .Z(n1418) );
  XOR U4037 ( .A(a[3914]), .B(n1404), .Z(n1406) );
  XOR U4038 ( .A(a[3917]), .B(n1392), .Z(n1394) );
  XOR U4039 ( .A(a[3920]), .B(n1379), .Z(n1381) );
  XOR U4040 ( .A(a[3923]), .B(n1367), .Z(n1369) );
  XOR U4041 ( .A(a[3926]), .B(n1355), .Z(n1357) );
  XOR U4042 ( .A(a[3929]), .B(n1342), .Z(n1344) );
  XOR U4043 ( .A(a[3932]), .B(n1330), .Z(n1332) );
  XOR U4044 ( .A(a[3935]), .B(n1318), .Z(n1320) );
  XOR U4045 ( .A(a[3938]), .B(n1306), .Z(n1308) );
  XOR U4046 ( .A(a[3941]), .B(n1293), .Z(n1295) );
  XOR U4047 ( .A(a[3944]), .B(n1281), .Z(n1283) );
  XOR U4048 ( .A(a[3947]), .B(n1269), .Z(n1271) );
  XOR U4049 ( .A(a[3950]), .B(n1256), .Z(n1258) );
  XOR U4050 ( .A(a[3953]), .B(n1244), .Z(n1246) );
  XOR U4051 ( .A(a[3956]), .B(n1232), .Z(n1234) );
  XOR U4052 ( .A(a[3959]), .B(n1219), .Z(n1221) );
  XOR U4053 ( .A(a[3962]), .B(n1207), .Z(n1209) );
  XOR U4054 ( .A(a[3965]), .B(n1195), .Z(n1197) );
  XOR U4055 ( .A(a[3968]), .B(n1183), .Z(n1185) );
  XOR U4056 ( .A(a[3971]), .B(n1170), .Z(n1172) );
  XOR U4057 ( .A(a[3974]), .B(n1158), .Z(n1160) );
  XOR U4058 ( .A(a[3977]), .B(n1146), .Z(n1148) );
  XOR U4059 ( .A(a[3980]), .B(n1133), .Z(n1135) );
  XOR U4060 ( .A(a[3983]), .B(n1121), .Z(n1123) );
  XOR U4061 ( .A(a[3986]), .B(n1109), .Z(n1111) );
  XOR U4062 ( .A(a[3989]), .B(n1096), .Z(n1098) );
  XOR U4063 ( .A(a[3992]), .B(n1084), .Z(n1086) );
  XOR U4064 ( .A(a[3995]), .B(n1072), .Z(n1074) );
  XOR U4065 ( .A(a[3998]), .B(n1060), .Z(n1062) );
  XOR U4066 ( .A(a[4001]), .B(n1045), .Z(n1047) );
  XOR U4067 ( .A(a[4004]), .B(n1033), .Z(n1035) );
  XOR U4068 ( .A(a[4007]), .B(n1021), .Z(n1023) );
  XOR U4069 ( .A(a[4010]), .B(n1008), .Z(n1010) );
  XOR U4070 ( .A(a[4013]), .B(n996), .Z(n998) );
  XOR U4071 ( .A(a[4016]), .B(n984), .Z(n986) );
  XOR U4072 ( .A(a[4019]), .B(n971), .Z(n973) );
  XOR U4073 ( .A(a[4022]), .B(n959), .Z(n961) );
  XOR U4074 ( .A(a[4025]), .B(n947), .Z(n949) );
  XOR U4075 ( .A(a[4028]), .B(n935), .Z(n937) );
  XOR U4076 ( .A(a[4031]), .B(n922), .Z(n924) );
  XOR U4077 ( .A(a[4034]), .B(n910), .Z(n912) );
  XOR U4078 ( .A(a[4037]), .B(n898), .Z(n900) );
  XOR U4079 ( .A(a[4040]), .B(n885), .Z(n887) );
  XOR U4080 ( .A(a[4043]), .B(n873), .Z(n875) );
  XOR U4081 ( .A(a[4046]), .B(n861), .Z(n863) );
  XOR U4082 ( .A(a[4049]), .B(n848), .Z(n850) );
  XOR U4083 ( .A(a[4052]), .B(n836), .Z(n838) );
  XOR U4084 ( .A(a[4055]), .B(n824), .Z(n826) );
  XOR U4085 ( .A(a[4058]), .B(n812), .Z(n814) );
  XOR U4086 ( .A(a[4061]), .B(n799), .Z(n801) );
  XOR U4087 ( .A(a[4064]), .B(n787), .Z(n789) );
  XOR U4088 ( .A(a[4067]), .B(n775), .Z(n777) );
  XOR U4089 ( .A(a[4070]), .B(n762), .Z(n764) );
  XOR U4090 ( .A(a[4073]), .B(n750), .Z(n752) );
  XOR U4091 ( .A(a[4076]), .B(n738), .Z(n740) );
  XOR U4092 ( .A(a[4079]), .B(n725), .Z(n727) );
  XOR U4093 ( .A(a[4082]), .B(n713), .Z(n715) );
  XOR U4094 ( .A(a[4085]), .B(n701), .Z(n703) );
  XOR U4095 ( .A(a[4088]), .B(n689), .Z(n691) );
  XOR U4096 ( .A(a[4091]), .B(n676), .Z(n678) );
  XOR U4097 ( .A(a[4094]), .B(n664), .Z(n666) );
  XOR U4098 ( .A(n2), .B(n3), .Z(carry_on_d) );
  ANDN U4099 ( .B(n4), .A(n5), .Z(n2) );
  XOR U4100 ( .A(b[4095]), .B(n3), .Z(n4) );
  XNOR U4101 ( .A(b[9]), .B(n6), .Z(c[9]) );
  XNOR U4102 ( .A(b[99]), .B(n7), .Z(c[99]) );
  XNOR U4103 ( .A(b[999]), .B(n8), .Z(c[999]) );
  XNOR U4104 ( .A(b[998]), .B(n9), .Z(c[998]) );
  XNOR U4105 ( .A(b[997]), .B(n10), .Z(c[997]) );
  XNOR U4106 ( .A(b[996]), .B(n11), .Z(c[996]) );
  XNOR U4107 ( .A(b[995]), .B(n12), .Z(c[995]) );
  XNOR U4108 ( .A(b[994]), .B(n13), .Z(c[994]) );
  XNOR U4109 ( .A(b[993]), .B(n14), .Z(c[993]) );
  XNOR U4110 ( .A(b[992]), .B(n15), .Z(c[992]) );
  XNOR U4111 ( .A(b[991]), .B(n16), .Z(c[991]) );
  XNOR U4112 ( .A(b[990]), .B(n17), .Z(c[990]) );
  XNOR U4113 ( .A(b[98]), .B(n18), .Z(c[98]) );
  XNOR U4114 ( .A(b[989]), .B(n19), .Z(c[989]) );
  XNOR U4115 ( .A(b[988]), .B(n20), .Z(c[988]) );
  XNOR U4116 ( .A(b[987]), .B(n21), .Z(c[987]) );
  XNOR U4117 ( .A(b[986]), .B(n22), .Z(c[986]) );
  XNOR U4118 ( .A(b[985]), .B(n23), .Z(c[985]) );
  XNOR U4119 ( .A(b[984]), .B(n24), .Z(c[984]) );
  XNOR U4120 ( .A(b[983]), .B(n25), .Z(c[983]) );
  XNOR U4121 ( .A(b[982]), .B(n26), .Z(c[982]) );
  XNOR U4122 ( .A(b[981]), .B(n27), .Z(c[981]) );
  XNOR U4123 ( .A(b[980]), .B(n28), .Z(c[980]) );
  XNOR U4124 ( .A(b[97]), .B(n29), .Z(c[97]) );
  XNOR U4125 ( .A(b[979]), .B(n30), .Z(c[979]) );
  XNOR U4126 ( .A(b[978]), .B(n31), .Z(c[978]) );
  XNOR U4127 ( .A(b[977]), .B(n32), .Z(c[977]) );
  XNOR U4128 ( .A(b[976]), .B(n33), .Z(c[976]) );
  XNOR U4129 ( .A(b[975]), .B(n34), .Z(c[975]) );
  XNOR U4130 ( .A(b[974]), .B(n35), .Z(c[974]) );
  XNOR U4131 ( .A(b[973]), .B(n36), .Z(c[973]) );
  XNOR U4132 ( .A(b[972]), .B(n37), .Z(c[972]) );
  XNOR U4133 ( .A(b[971]), .B(n38), .Z(c[971]) );
  XNOR U4134 ( .A(b[970]), .B(n39), .Z(c[970]) );
  XNOR U4135 ( .A(b[96]), .B(n40), .Z(c[96]) );
  XNOR U4136 ( .A(b[969]), .B(n41), .Z(c[969]) );
  XNOR U4137 ( .A(b[968]), .B(n42), .Z(c[968]) );
  XNOR U4138 ( .A(b[967]), .B(n43), .Z(c[967]) );
  XNOR U4139 ( .A(b[966]), .B(n44), .Z(c[966]) );
  XNOR U4140 ( .A(b[965]), .B(n45), .Z(c[965]) );
  XNOR U4141 ( .A(b[964]), .B(n46), .Z(c[964]) );
  XNOR U4142 ( .A(b[963]), .B(n47), .Z(c[963]) );
  XNOR U4143 ( .A(b[962]), .B(n48), .Z(c[962]) );
  XNOR U4144 ( .A(b[961]), .B(n49), .Z(c[961]) );
  XNOR U4145 ( .A(b[960]), .B(n50), .Z(c[960]) );
  XNOR U4146 ( .A(b[95]), .B(n51), .Z(c[95]) );
  XNOR U4147 ( .A(b[959]), .B(n52), .Z(c[959]) );
  XNOR U4148 ( .A(b[958]), .B(n53), .Z(c[958]) );
  XNOR U4149 ( .A(b[957]), .B(n54), .Z(c[957]) );
  XNOR U4150 ( .A(b[956]), .B(n55), .Z(c[956]) );
  XNOR U4151 ( .A(b[955]), .B(n56), .Z(c[955]) );
  XNOR U4152 ( .A(b[954]), .B(n57), .Z(c[954]) );
  XNOR U4153 ( .A(b[953]), .B(n58), .Z(c[953]) );
  XNOR U4154 ( .A(b[952]), .B(n59), .Z(c[952]) );
  XNOR U4155 ( .A(b[951]), .B(n60), .Z(c[951]) );
  XNOR U4156 ( .A(b[950]), .B(n61), .Z(c[950]) );
  XNOR U4157 ( .A(b[94]), .B(n62), .Z(c[94]) );
  XNOR U4158 ( .A(b[949]), .B(n63), .Z(c[949]) );
  XNOR U4159 ( .A(b[948]), .B(n64), .Z(c[948]) );
  XNOR U4160 ( .A(b[947]), .B(n65), .Z(c[947]) );
  XNOR U4161 ( .A(b[946]), .B(n66), .Z(c[946]) );
  XNOR U4162 ( .A(b[945]), .B(n67), .Z(c[945]) );
  XNOR U4163 ( .A(b[944]), .B(n68), .Z(c[944]) );
  XNOR U4164 ( .A(b[943]), .B(n69), .Z(c[943]) );
  XNOR U4165 ( .A(b[942]), .B(n70), .Z(c[942]) );
  XNOR U4166 ( .A(b[941]), .B(n71), .Z(c[941]) );
  XNOR U4167 ( .A(b[940]), .B(n72), .Z(c[940]) );
  XNOR U4168 ( .A(b[93]), .B(n73), .Z(c[93]) );
  XNOR U4169 ( .A(b[939]), .B(n74), .Z(c[939]) );
  XNOR U4170 ( .A(b[938]), .B(n75), .Z(c[938]) );
  XNOR U4171 ( .A(b[937]), .B(n76), .Z(c[937]) );
  XNOR U4172 ( .A(b[936]), .B(n77), .Z(c[936]) );
  XNOR U4173 ( .A(b[935]), .B(n78), .Z(c[935]) );
  XNOR U4174 ( .A(b[934]), .B(n79), .Z(c[934]) );
  XNOR U4175 ( .A(b[933]), .B(n80), .Z(c[933]) );
  XNOR U4176 ( .A(b[932]), .B(n81), .Z(c[932]) );
  XNOR U4177 ( .A(b[931]), .B(n82), .Z(c[931]) );
  XNOR U4178 ( .A(b[930]), .B(n83), .Z(c[930]) );
  XNOR U4179 ( .A(b[92]), .B(n84), .Z(c[92]) );
  XNOR U4180 ( .A(b[929]), .B(n85), .Z(c[929]) );
  XNOR U4181 ( .A(b[928]), .B(n86), .Z(c[928]) );
  XNOR U4182 ( .A(b[927]), .B(n87), .Z(c[927]) );
  XNOR U4183 ( .A(b[926]), .B(n88), .Z(c[926]) );
  XNOR U4184 ( .A(b[925]), .B(n89), .Z(c[925]) );
  XNOR U4185 ( .A(b[924]), .B(n90), .Z(c[924]) );
  XNOR U4186 ( .A(b[923]), .B(n91), .Z(c[923]) );
  XNOR U4187 ( .A(b[922]), .B(n92), .Z(c[922]) );
  XNOR U4188 ( .A(b[921]), .B(n93), .Z(c[921]) );
  XNOR U4189 ( .A(b[920]), .B(n94), .Z(c[920]) );
  XNOR U4190 ( .A(b[91]), .B(n95), .Z(c[91]) );
  XNOR U4191 ( .A(b[919]), .B(n96), .Z(c[919]) );
  XNOR U4192 ( .A(b[918]), .B(n97), .Z(c[918]) );
  XNOR U4193 ( .A(b[917]), .B(n98), .Z(c[917]) );
  XNOR U4194 ( .A(b[916]), .B(n99), .Z(c[916]) );
  XNOR U4195 ( .A(b[915]), .B(n100), .Z(c[915]) );
  XNOR U4196 ( .A(b[914]), .B(n101), .Z(c[914]) );
  XNOR U4197 ( .A(b[913]), .B(n102), .Z(c[913]) );
  XNOR U4198 ( .A(b[912]), .B(n103), .Z(c[912]) );
  XNOR U4199 ( .A(b[911]), .B(n104), .Z(c[911]) );
  XNOR U4200 ( .A(b[910]), .B(n105), .Z(c[910]) );
  XNOR U4201 ( .A(b[90]), .B(n106), .Z(c[90]) );
  XNOR U4202 ( .A(b[909]), .B(n107), .Z(c[909]) );
  XNOR U4203 ( .A(b[908]), .B(n108), .Z(c[908]) );
  XNOR U4204 ( .A(b[907]), .B(n109), .Z(c[907]) );
  XNOR U4205 ( .A(b[906]), .B(n110), .Z(c[906]) );
  XNOR U4206 ( .A(b[905]), .B(n111), .Z(c[905]) );
  XNOR U4207 ( .A(b[904]), .B(n112), .Z(c[904]) );
  XNOR U4208 ( .A(b[903]), .B(n113), .Z(c[903]) );
  XNOR U4209 ( .A(b[902]), .B(n114), .Z(c[902]) );
  XNOR U4210 ( .A(b[901]), .B(n115), .Z(c[901]) );
  XNOR U4211 ( .A(b[900]), .B(n116), .Z(c[900]) );
  XNOR U4212 ( .A(b[8]), .B(n117), .Z(c[8]) );
  XNOR U4213 ( .A(b[89]), .B(n118), .Z(c[89]) );
  XNOR U4214 ( .A(b[899]), .B(n119), .Z(c[899]) );
  XNOR U4215 ( .A(b[898]), .B(n120), .Z(c[898]) );
  XNOR U4216 ( .A(b[897]), .B(n121), .Z(c[897]) );
  XNOR U4217 ( .A(b[896]), .B(n122), .Z(c[896]) );
  XNOR U4218 ( .A(b[895]), .B(n123), .Z(c[895]) );
  XNOR U4219 ( .A(b[894]), .B(n124), .Z(c[894]) );
  XNOR U4220 ( .A(b[893]), .B(n125), .Z(c[893]) );
  XNOR U4221 ( .A(b[892]), .B(n126), .Z(c[892]) );
  XNOR U4222 ( .A(b[891]), .B(n127), .Z(c[891]) );
  XNOR U4223 ( .A(b[890]), .B(n128), .Z(c[890]) );
  XNOR U4224 ( .A(b[88]), .B(n129), .Z(c[88]) );
  XNOR U4225 ( .A(b[889]), .B(n130), .Z(c[889]) );
  XNOR U4226 ( .A(b[888]), .B(n131), .Z(c[888]) );
  XNOR U4227 ( .A(b[887]), .B(n132), .Z(c[887]) );
  XNOR U4228 ( .A(b[886]), .B(n133), .Z(c[886]) );
  XNOR U4229 ( .A(b[885]), .B(n134), .Z(c[885]) );
  XNOR U4230 ( .A(b[884]), .B(n135), .Z(c[884]) );
  XNOR U4231 ( .A(b[883]), .B(n136), .Z(c[883]) );
  XNOR U4232 ( .A(b[882]), .B(n137), .Z(c[882]) );
  XNOR U4233 ( .A(b[881]), .B(n138), .Z(c[881]) );
  XNOR U4234 ( .A(b[880]), .B(n139), .Z(c[880]) );
  XNOR U4235 ( .A(b[87]), .B(n140), .Z(c[87]) );
  XNOR U4236 ( .A(b[879]), .B(n141), .Z(c[879]) );
  XNOR U4237 ( .A(b[878]), .B(n142), .Z(c[878]) );
  XNOR U4238 ( .A(b[877]), .B(n143), .Z(c[877]) );
  XNOR U4239 ( .A(b[876]), .B(n144), .Z(c[876]) );
  XNOR U4240 ( .A(b[875]), .B(n145), .Z(c[875]) );
  XNOR U4241 ( .A(b[874]), .B(n146), .Z(c[874]) );
  XNOR U4242 ( .A(b[873]), .B(n147), .Z(c[873]) );
  XNOR U4243 ( .A(b[872]), .B(n148), .Z(c[872]) );
  XNOR U4244 ( .A(b[871]), .B(n149), .Z(c[871]) );
  XNOR U4245 ( .A(b[870]), .B(n150), .Z(c[870]) );
  XNOR U4246 ( .A(b[86]), .B(n151), .Z(c[86]) );
  XNOR U4247 ( .A(b[869]), .B(n152), .Z(c[869]) );
  XNOR U4248 ( .A(b[868]), .B(n153), .Z(c[868]) );
  XNOR U4249 ( .A(b[867]), .B(n154), .Z(c[867]) );
  XNOR U4250 ( .A(b[866]), .B(n155), .Z(c[866]) );
  XNOR U4251 ( .A(b[865]), .B(n156), .Z(c[865]) );
  XNOR U4252 ( .A(b[864]), .B(n157), .Z(c[864]) );
  XNOR U4253 ( .A(b[863]), .B(n158), .Z(c[863]) );
  XNOR U4254 ( .A(b[862]), .B(n159), .Z(c[862]) );
  XNOR U4255 ( .A(b[861]), .B(n160), .Z(c[861]) );
  XNOR U4256 ( .A(b[860]), .B(n161), .Z(c[860]) );
  XNOR U4257 ( .A(b[85]), .B(n162), .Z(c[85]) );
  XNOR U4258 ( .A(b[859]), .B(n163), .Z(c[859]) );
  XNOR U4259 ( .A(b[858]), .B(n164), .Z(c[858]) );
  XNOR U4260 ( .A(b[857]), .B(n165), .Z(c[857]) );
  XNOR U4261 ( .A(b[856]), .B(n166), .Z(c[856]) );
  XNOR U4262 ( .A(b[855]), .B(n167), .Z(c[855]) );
  XNOR U4263 ( .A(b[854]), .B(n168), .Z(c[854]) );
  XNOR U4264 ( .A(b[853]), .B(n169), .Z(c[853]) );
  XNOR U4265 ( .A(b[852]), .B(n170), .Z(c[852]) );
  XNOR U4266 ( .A(b[851]), .B(n171), .Z(c[851]) );
  XNOR U4267 ( .A(b[850]), .B(n172), .Z(c[850]) );
  XNOR U4268 ( .A(b[84]), .B(n173), .Z(c[84]) );
  XNOR U4269 ( .A(b[849]), .B(n174), .Z(c[849]) );
  XNOR U4270 ( .A(b[848]), .B(n175), .Z(c[848]) );
  XNOR U4271 ( .A(b[847]), .B(n176), .Z(c[847]) );
  XNOR U4272 ( .A(b[846]), .B(n177), .Z(c[846]) );
  XNOR U4273 ( .A(b[845]), .B(n178), .Z(c[845]) );
  XNOR U4274 ( .A(b[844]), .B(n179), .Z(c[844]) );
  XNOR U4275 ( .A(b[843]), .B(n180), .Z(c[843]) );
  XNOR U4276 ( .A(b[842]), .B(n181), .Z(c[842]) );
  XNOR U4277 ( .A(b[841]), .B(n182), .Z(c[841]) );
  XNOR U4278 ( .A(b[840]), .B(n183), .Z(c[840]) );
  XNOR U4279 ( .A(b[83]), .B(n184), .Z(c[83]) );
  XNOR U4280 ( .A(b[839]), .B(n185), .Z(c[839]) );
  XNOR U4281 ( .A(b[838]), .B(n186), .Z(c[838]) );
  XNOR U4282 ( .A(b[837]), .B(n187), .Z(c[837]) );
  XNOR U4283 ( .A(b[836]), .B(n188), .Z(c[836]) );
  XNOR U4284 ( .A(b[835]), .B(n189), .Z(c[835]) );
  XNOR U4285 ( .A(b[834]), .B(n190), .Z(c[834]) );
  XNOR U4286 ( .A(b[833]), .B(n191), .Z(c[833]) );
  XNOR U4287 ( .A(b[832]), .B(n192), .Z(c[832]) );
  XNOR U4288 ( .A(b[831]), .B(n193), .Z(c[831]) );
  XNOR U4289 ( .A(b[830]), .B(n194), .Z(c[830]) );
  XNOR U4290 ( .A(b[82]), .B(n195), .Z(c[82]) );
  XNOR U4291 ( .A(b[829]), .B(n196), .Z(c[829]) );
  XNOR U4292 ( .A(b[828]), .B(n197), .Z(c[828]) );
  XNOR U4293 ( .A(b[827]), .B(n198), .Z(c[827]) );
  XNOR U4294 ( .A(b[826]), .B(n199), .Z(c[826]) );
  XNOR U4295 ( .A(b[825]), .B(n200), .Z(c[825]) );
  XNOR U4296 ( .A(b[824]), .B(n201), .Z(c[824]) );
  XNOR U4297 ( .A(b[823]), .B(n202), .Z(c[823]) );
  XNOR U4298 ( .A(b[822]), .B(n203), .Z(c[822]) );
  XNOR U4299 ( .A(b[821]), .B(n204), .Z(c[821]) );
  XNOR U4300 ( .A(b[820]), .B(n205), .Z(c[820]) );
  XNOR U4301 ( .A(b[81]), .B(n206), .Z(c[81]) );
  XNOR U4302 ( .A(b[819]), .B(n207), .Z(c[819]) );
  XNOR U4303 ( .A(b[818]), .B(n208), .Z(c[818]) );
  XNOR U4304 ( .A(b[817]), .B(n209), .Z(c[817]) );
  XNOR U4305 ( .A(b[816]), .B(n210), .Z(c[816]) );
  XNOR U4306 ( .A(b[815]), .B(n211), .Z(c[815]) );
  XNOR U4307 ( .A(b[814]), .B(n212), .Z(c[814]) );
  XNOR U4308 ( .A(b[813]), .B(n213), .Z(c[813]) );
  XNOR U4309 ( .A(b[812]), .B(n214), .Z(c[812]) );
  XNOR U4310 ( .A(b[811]), .B(n215), .Z(c[811]) );
  XNOR U4311 ( .A(b[810]), .B(n216), .Z(c[810]) );
  XNOR U4312 ( .A(b[80]), .B(n217), .Z(c[80]) );
  XNOR U4313 ( .A(b[809]), .B(n218), .Z(c[809]) );
  XNOR U4314 ( .A(b[808]), .B(n219), .Z(c[808]) );
  XNOR U4315 ( .A(b[807]), .B(n220), .Z(c[807]) );
  XNOR U4316 ( .A(b[806]), .B(n221), .Z(c[806]) );
  XNOR U4317 ( .A(b[805]), .B(n222), .Z(c[805]) );
  XNOR U4318 ( .A(b[804]), .B(n223), .Z(c[804]) );
  XNOR U4319 ( .A(b[803]), .B(n224), .Z(c[803]) );
  XNOR U4320 ( .A(b[802]), .B(n225), .Z(c[802]) );
  XNOR U4321 ( .A(b[801]), .B(n226), .Z(c[801]) );
  XNOR U4322 ( .A(b[800]), .B(n227), .Z(c[800]) );
  XNOR U4323 ( .A(b[7]), .B(n228), .Z(c[7]) );
  XNOR U4324 ( .A(b[79]), .B(n229), .Z(c[79]) );
  XNOR U4325 ( .A(b[799]), .B(n230), .Z(c[799]) );
  XNOR U4326 ( .A(b[798]), .B(n231), .Z(c[798]) );
  XNOR U4327 ( .A(b[797]), .B(n232), .Z(c[797]) );
  XNOR U4328 ( .A(b[796]), .B(n233), .Z(c[796]) );
  XNOR U4329 ( .A(b[795]), .B(n234), .Z(c[795]) );
  XNOR U4330 ( .A(b[794]), .B(n235), .Z(c[794]) );
  XNOR U4331 ( .A(b[793]), .B(n236), .Z(c[793]) );
  XNOR U4332 ( .A(b[792]), .B(n237), .Z(c[792]) );
  XNOR U4333 ( .A(b[791]), .B(n238), .Z(c[791]) );
  XNOR U4334 ( .A(b[790]), .B(n239), .Z(c[790]) );
  XNOR U4335 ( .A(b[78]), .B(n240), .Z(c[78]) );
  XNOR U4336 ( .A(b[789]), .B(n241), .Z(c[789]) );
  XNOR U4337 ( .A(b[788]), .B(n242), .Z(c[788]) );
  XNOR U4338 ( .A(b[787]), .B(n243), .Z(c[787]) );
  XNOR U4339 ( .A(b[786]), .B(n244), .Z(c[786]) );
  XNOR U4340 ( .A(b[785]), .B(n245), .Z(c[785]) );
  XNOR U4341 ( .A(b[784]), .B(n246), .Z(c[784]) );
  XNOR U4342 ( .A(b[783]), .B(n247), .Z(c[783]) );
  XNOR U4343 ( .A(b[782]), .B(n248), .Z(c[782]) );
  XNOR U4344 ( .A(b[781]), .B(n249), .Z(c[781]) );
  XNOR U4345 ( .A(b[780]), .B(n250), .Z(c[780]) );
  XNOR U4346 ( .A(b[77]), .B(n251), .Z(c[77]) );
  XNOR U4347 ( .A(b[779]), .B(n252), .Z(c[779]) );
  XNOR U4348 ( .A(b[778]), .B(n253), .Z(c[778]) );
  XNOR U4349 ( .A(b[777]), .B(n254), .Z(c[777]) );
  XNOR U4350 ( .A(b[776]), .B(n255), .Z(c[776]) );
  XNOR U4351 ( .A(b[775]), .B(n256), .Z(c[775]) );
  XNOR U4352 ( .A(b[774]), .B(n257), .Z(c[774]) );
  XNOR U4353 ( .A(b[773]), .B(n258), .Z(c[773]) );
  XNOR U4354 ( .A(b[772]), .B(n259), .Z(c[772]) );
  XNOR U4355 ( .A(b[771]), .B(n260), .Z(c[771]) );
  XNOR U4356 ( .A(b[770]), .B(n261), .Z(c[770]) );
  XNOR U4357 ( .A(b[76]), .B(n262), .Z(c[76]) );
  XNOR U4358 ( .A(b[769]), .B(n263), .Z(c[769]) );
  XNOR U4359 ( .A(b[768]), .B(n264), .Z(c[768]) );
  XNOR U4360 ( .A(b[767]), .B(n265), .Z(c[767]) );
  XNOR U4361 ( .A(b[766]), .B(n266), .Z(c[766]) );
  XNOR U4362 ( .A(b[765]), .B(n267), .Z(c[765]) );
  XNOR U4363 ( .A(b[764]), .B(n268), .Z(c[764]) );
  XNOR U4364 ( .A(b[763]), .B(n269), .Z(c[763]) );
  XNOR U4365 ( .A(b[762]), .B(n270), .Z(c[762]) );
  XNOR U4366 ( .A(b[761]), .B(n271), .Z(c[761]) );
  XNOR U4367 ( .A(b[760]), .B(n272), .Z(c[760]) );
  XNOR U4368 ( .A(b[75]), .B(n273), .Z(c[75]) );
  XNOR U4369 ( .A(b[759]), .B(n274), .Z(c[759]) );
  XNOR U4370 ( .A(b[758]), .B(n275), .Z(c[758]) );
  XNOR U4371 ( .A(b[757]), .B(n276), .Z(c[757]) );
  XNOR U4372 ( .A(b[756]), .B(n277), .Z(c[756]) );
  XNOR U4373 ( .A(b[755]), .B(n278), .Z(c[755]) );
  XNOR U4374 ( .A(b[754]), .B(n279), .Z(c[754]) );
  XNOR U4375 ( .A(b[753]), .B(n280), .Z(c[753]) );
  XNOR U4376 ( .A(b[752]), .B(n281), .Z(c[752]) );
  XNOR U4377 ( .A(b[751]), .B(n282), .Z(c[751]) );
  XNOR U4378 ( .A(b[750]), .B(n283), .Z(c[750]) );
  XNOR U4379 ( .A(b[74]), .B(n284), .Z(c[74]) );
  XNOR U4380 ( .A(b[749]), .B(n285), .Z(c[749]) );
  XNOR U4381 ( .A(b[748]), .B(n286), .Z(c[748]) );
  XNOR U4382 ( .A(b[747]), .B(n287), .Z(c[747]) );
  XNOR U4383 ( .A(b[746]), .B(n288), .Z(c[746]) );
  XNOR U4384 ( .A(b[745]), .B(n289), .Z(c[745]) );
  XNOR U4385 ( .A(b[744]), .B(n290), .Z(c[744]) );
  XNOR U4386 ( .A(b[743]), .B(n291), .Z(c[743]) );
  XNOR U4387 ( .A(b[742]), .B(n292), .Z(c[742]) );
  XNOR U4388 ( .A(b[741]), .B(n293), .Z(c[741]) );
  XNOR U4389 ( .A(b[740]), .B(n294), .Z(c[740]) );
  XNOR U4390 ( .A(b[73]), .B(n295), .Z(c[73]) );
  XNOR U4391 ( .A(b[739]), .B(n296), .Z(c[739]) );
  XNOR U4392 ( .A(b[738]), .B(n297), .Z(c[738]) );
  XNOR U4393 ( .A(b[737]), .B(n298), .Z(c[737]) );
  XNOR U4394 ( .A(b[736]), .B(n299), .Z(c[736]) );
  XNOR U4395 ( .A(b[735]), .B(n300), .Z(c[735]) );
  XNOR U4396 ( .A(b[734]), .B(n301), .Z(c[734]) );
  XNOR U4397 ( .A(b[733]), .B(n302), .Z(c[733]) );
  XNOR U4398 ( .A(b[732]), .B(n303), .Z(c[732]) );
  XNOR U4399 ( .A(b[731]), .B(n304), .Z(c[731]) );
  XNOR U4400 ( .A(b[730]), .B(n305), .Z(c[730]) );
  XNOR U4401 ( .A(b[72]), .B(n306), .Z(c[72]) );
  XNOR U4402 ( .A(b[729]), .B(n307), .Z(c[729]) );
  XNOR U4403 ( .A(b[728]), .B(n308), .Z(c[728]) );
  XNOR U4404 ( .A(b[727]), .B(n309), .Z(c[727]) );
  XNOR U4405 ( .A(b[726]), .B(n310), .Z(c[726]) );
  XNOR U4406 ( .A(b[725]), .B(n311), .Z(c[725]) );
  XNOR U4407 ( .A(b[724]), .B(n312), .Z(c[724]) );
  XNOR U4408 ( .A(b[723]), .B(n313), .Z(c[723]) );
  XNOR U4409 ( .A(b[722]), .B(n314), .Z(c[722]) );
  XNOR U4410 ( .A(b[721]), .B(n315), .Z(c[721]) );
  XNOR U4411 ( .A(b[720]), .B(n316), .Z(c[720]) );
  XNOR U4412 ( .A(b[71]), .B(n317), .Z(c[71]) );
  XNOR U4413 ( .A(b[719]), .B(n318), .Z(c[719]) );
  XNOR U4414 ( .A(b[718]), .B(n319), .Z(c[718]) );
  XNOR U4415 ( .A(b[717]), .B(n320), .Z(c[717]) );
  XNOR U4416 ( .A(b[716]), .B(n321), .Z(c[716]) );
  XNOR U4417 ( .A(b[715]), .B(n322), .Z(c[715]) );
  XNOR U4418 ( .A(b[714]), .B(n323), .Z(c[714]) );
  XNOR U4419 ( .A(b[713]), .B(n324), .Z(c[713]) );
  XNOR U4420 ( .A(b[712]), .B(n325), .Z(c[712]) );
  XNOR U4421 ( .A(b[711]), .B(n326), .Z(c[711]) );
  XNOR U4422 ( .A(b[710]), .B(n327), .Z(c[710]) );
  XNOR U4423 ( .A(b[70]), .B(n328), .Z(c[70]) );
  XNOR U4424 ( .A(b[709]), .B(n329), .Z(c[709]) );
  XNOR U4425 ( .A(b[708]), .B(n330), .Z(c[708]) );
  XNOR U4426 ( .A(b[707]), .B(n331), .Z(c[707]) );
  XNOR U4427 ( .A(b[706]), .B(n332), .Z(c[706]) );
  XNOR U4428 ( .A(b[705]), .B(n333), .Z(c[705]) );
  XNOR U4429 ( .A(b[704]), .B(n334), .Z(c[704]) );
  XNOR U4430 ( .A(b[703]), .B(n335), .Z(c[703]) );
  XNOR U4431 ( .A(b[702]), .B(n336), .Z(c[702]) );
  XNOR U4432 ( .A(b[701]), .B(n337), .Z(c[701]) );
  XNOR U4433 ( .A(b[700]), .B(n338), .Z(c[700]) );
  XNOR U4434 ( .A(b[6]), .B(n339), .Z(c[6]) );
  XNOR U4435 ( .A(b[69]), .B(n340), .Z(c[69]) );
  XNOR U4436 ( .A(b[699]), .B(n341), .Z(c[699]) );
  XNOR U4437 ( .A(b[698]), .B(n342), .Z(c[698]) );
  XNOR U4438 ( .A(b[697]), .B(n343), .Z(c[697]) );
  XNOR U4439 ( .A(b[696]), .B(n344), .Z(c[696]) );
  XNOR U4440 ( .A(b[695]), .B(n345), .Z(c[695]) );
  XNOR U4441 ( .A(b[694]), .B(n346), .Z(c[694]) );
  XNOR U4442 ( .A(b[693]), .B(n347), .Z(c[693]) );
  XNOR U4443 ( .A(b[692]), .B(n348), .Z(c[692]) );
  XNOR U4444 ( .A(b[691]), .B(n349), .Z(c[691]) );
  XNOR U4445 ( .A(b[690]), .B(n350), .Z(c[690]) );
  XNOR U4446 ( .A(b[68]), .B(n351), .Z(c[68]) );
  XNOR U4447 ( .A(b[689]), .B(n352), .Z(c[689]) );
  XNOR U4448 ( .A(b[688]), .B(n353), .Z(c[688]) );
  XNOR U4449 ( .A(b[687]), .B(n354), .Z(c[687]) );
  XNOR U4450 ( .A(b[686]), .B(n355), .Z(c[686]) );
  XNOR U4451 ( .A(b[685]), .B(n356), .Z(c[685]) );
  XNOR U4452 ( .A(b[684]), .B(n357), .Z(c[684]) );
  XNOR U4453 ( .A(b[683]), .B(n358), .Z(c[683]) );
  XNOR U4454 ( .A(b[682]), .B(n359), .Z(c[682]) );
  XNOR U4455 ( .A(b[681]), .B(n360), .Z(c[681]) );
  XNOR U4456 ( .A(b[680]), .B(n361), .Z(c[680]) );
  XNOR U4457 ( .A(b[67]), .B(n362), .Z(c[67]) );
  XNOR U4458 ( .A(b[679]), .B(n363), .Z(c[679]) );
  XNOR U4459 ( .A(b[678]), .B(n364), .Z(c[678]) );
  XNOR U4460 ( .A(b[677]), .B(n365), .Z(c[677]) );
  XNOR U4461 ( .A(b[676]), .B(n366), .Z(c[676]) );
  XNOR U4462 ( .A(b[675]), .B(n367), .Z(c[675]) );
  XNOR U4463 ( .A(b[674]), .B(n368), .Z(c[674]) );
  XNOR U4464 ( .A(b[673]), .B(n369), .Z(c[673]) );
  XNOR U4465 ( .A(b[672]), .B(n370), .Z(c[672]) );
  XNOR U4466 ( .A(b[671]), .B(n371), .Z(c[671]) );
  XNOR U4467 ( .A(b[670]), .B(n372), .Z(c[670]) );
  XNOR U4468 ( .A(b[66]), .B(n373), .Z(c[66]) );
  XNOR U4469 ( .A(b[669]), .B(n374), .Z(c[669]) );
  XNOR U4470 ( .A(b[668]), .B(n375), .Z(c[668]) );
  XNOR U4471 ( .A(b[667]), .B(n376), .Z(c[667]) );
  XNOR U4472 ( .A(b[666]), .B(n377), .Z(c[666]) );
  XNOR U4473 ( .A(b[665]), .B(n378), .Z(c[665]) );
  XNOR U4474 ( .A(b[664]), .B(n379), .Z(c[664]) );
  XNOR U4475 ( .A(b[663]), .B(n380), .Z(c[663]) );
  XNOR U4476 ( .A(b[662]), .B(n381), .Z(c[662]) );
  XNOR U4477 ( .A(b[661]), .B(n382), .Z(c[661]) );
  XNOR U4478 ( .A(b[660]), .B(n383), .Z(c[660]) );
  XNOR U4479 ( .A(b[65]), .B(n384), .Z(c[65]) );
  XNOR U4480 ( .A(b[659]), .B(n385), .Z(c[659]) );
  XNOR U4481 ( .A(b[658]), .B(n386), .Z(c[658]) );
  XNOR U4482 ( .A(b[657]), .B(n387), .Z(c[657]) );
  XNOR U4483 ( .A(b[656]), .B(n388), .Z(c[656]) );
  XNOR U4484 ( .A(b[655]), .B(n389), .Z(c[655]) );
  XNOR U4485 ( .A(b[654]), .B(n390), .Z(c[654]) );
  XNOR U4486 ( .A(b[653]), .B(n391), .Z(c[653]) );
  XNOR U4487 ( .A(b[652]), .B(n392), .Z(c[652]) );
  XNOR U4488 ( .A(b[651]), .B(n393), .Z(c[651]) );
  XNOR U4489 ( .A(b[650]), .B(n394), .Z(c[650]) );
  XNOR U4490 ( .A(b[64]), .B(n395), .Z(c[64]) );
  XNOR U4491 ( .A(b[649]), .B(n396), .Z(c[649]) );
  XNOR U4492 ( .A(b[648]), .B(n397), .Z(c[648]) );
  XNOR U4493 ( .A(b[647]), .B(n398), .Z(c[647]) );
  XNOR U4494 ( .A(b[646]), .B(n399), .Z(c[646]) );
  XNOR U4495 ( .A(b[645]), .B(n400), .Z(c[645]) );
  XNOR U4496 ( .A(b[644]), .B(n401), .Z(c[644]) );
  XNOR U4497 ( .A(b[643]), .B(n402), .Z(c[643]) );
  XNOR U4498 ( .A(b[642]), .B(n403), .Z(c[642]) );
  XNOR U4499 ( .A(b[641]), .B(n404), .Z(c[641]) );
  XNOR U4500 ( .A(b[640]), .B(n405), .Z(c[640]) );
  XNOR U4501 ( .A(b[63]), .B(n406), .Z(c[63]) );
  XNOR U4502 ( .A(b[639]), .B(n407), .Z(c[639]) );
  XNOR U4503 ( .A(b[638]), .B(n408), .Z(c[638]) );
  XNOR U4504 ( .A(b[637]), .B(n409), .Z(c[637]) );
  XNOR U4505 ( .A(b[636]), .B(n410), .Z(c[636]) );
  XNOR U4506 ( .A(b[635]), .B(n411), .Z(c[635]) );
  XNOR U4507 ( .A(b[634]), .B(n412), .Z(c[634]) );
  XNOR U4508 ( .A(b[633]), .B(n413), .Z(c[633]) );
  XNOR U4509 ( .A(b[632]), .B(n414), .Z(c[632]) );
  XNOR U4510 ( .A(b[631]), .B(n415), .Z(c[631]) );
  XNOR U4511 ( .A(b[630]), .B(n416), .Z(c[630]) );
  XNOR U4512 ( .A(b[62]), .B(n417), .Z(c[62]) );
  XNOR U4513 ( .A(b[629]), .B(n418), .Z(c[629]) );
  XNOR U4514 ( .A(b[628]), .B(n419), .Z(c[628]) );
  XNOR U4515 ( .A(b[627]), .B(n420), .Z(c[627]) );
  XNOR U4516 ( .A(b[626]), .B(n421), .Z(c[626]) );
  XNOR U4517 ( .A(b[625]), .B(n422), .Z(c[625]) );
  XNOR U4518 ( .A(b[624]), .B(n423), .Z(c[624]) );
  XNOR U4519 ( .A(b[623]), .B(n424), .Z(c[623]) );
  XNOR U4520 ( .A(b[622]), .B(n425), .Z(c[622]) );
  XNOR U4521 ( .A(b[621]), .B(n426), .Z(c[621]) );
  XNOR U4522 ( .A(b[620]), .B(n427), .Z(c[620]) );
  XNOR U4523 ( .A(b[61]), .B(n428), .Z(c[61]) );
  XNOR U4524 ( .A(b[619]), .B(n429), .Z(c[619]) );
  XNOR U4525 ( .A(b[618]), .B(n430), .Z(c[618]) );
  XNOR U4526 ( .A(b[617]), .B(n431), .Z(c[617]) );
  XNOR U4527 ( .A(b[616]), .B(n432), .Z(c[616]) );
  XNOR U4528 ( .A(b[615]), .B(n433), .Z(c[615]) );
  XNOR U4529 ( .A(b[614]), .B(n434), .Z(c[614]) );
  XNOR U4530 ( .A(b[613]), .B(n435), .Z(c[613]) );
  XNOR U4531 ( .A(b[612]), .B(n436), .Z(c[612]) );
  XNOR U4532 ( .A(b[611]), .B(n437), .Z(c[611]) );
  XNOR U4533 ( .A(b[610]), .B(n438), .Z(c[610]) );
  XNOR U4534 ( .A(b[60]), .B(n439), .Z(c[60]) );
  XNOR U4535 ( .A(b[609]), .B(n440), .Z(c[609]) );
  XNOR U4536 ( .A(b[608]), .B(n441), .Z(c[608]) );
  XNOR U4537 ( .A(b[607]), .B(n442), .Z(c[607]) );
  XNOR U4538 ( .A(b[606]), .B(n443), .Z(c[606]) );
  XNOR U4539 ( .A(b[605]), .B(n444), .Z(c[605]) );
  XNOR U4540 ( .A(b[604]), .B(n445), .Z(c[604]) );
  XNOR U4541 ( .A(b[603]), .B(n446), .Z(c[603]) );
  XNOR U4542 ( .A(b[602]), .B(n447), .Z(c[602]) );
  XNOR U4543 ( .A(b[601]), .B(n448), .Z(c[601]) );
  XNOR U4544 ( .A(b[600]), .B(n449), .Z(c[600]) );
  XNOR U4545 ( .A(b[5]), .B(n450), .Z(c[5]) );
  XNOR U4546 ( .A(b[59]), .B(n451), .Z(c[59]) );
  XNOR U4547 ( .A(b[599]), .B(n452), .Z(c[599]) );
  XNOR U4548 ( .A(b[598]), .B(n453), .Z(c[598]) );
  XNOR U4549 ( .A(b[597]), .B(n454), .Z(c[597]) );
  XNOR U4550 ( .A(b[596]), .B(n455), .Z(c[596]) );
  XNOR U4551 ( .A(b[595]), .B(n456), .Z(c[595]) );
  XNOR U4552 ( .A(b[594]), .B(n457), .Z(c[594]) );
  XNOR U4553 ( .A(b[593]), .B(n458), .Z(c[593]) );
  XNOR U4554 ( .A(b[592]), .B(n459), .Z(c[592]) );
  XNOR U4555 ( .A(b[591]), .B(n460), .Z(c[591]) );
  XNOR U4556 ( .A(b[590]), .B(n461), .Z(c[590]) );
  XNOR U4557 ( .A(b[58]), .B(n462), .Z(c[58]) );
  XNOR U4558 ( .A(b[589]), .B(n463), .Z(c[589]) );
  XNOR U4559 ( .A(b[588]), .B(n464), .Z(c[588]) );
  XNOR U4560 ( .A(b[587]), .B(n465), .Z(c[587]) );
  XNOR U4561 ( .A(b[586]), .B(n466), .Z(c[586]) );
  XNOR U4562 ( .A(b[585]), .B(n467), .Z(c[585]) );
  XNOR U4563 ( .A(b[584]), .B(n468), .Z(c[584]) );
  XNOR U4564 ( .A(b[583]), .B(n469), .Z(c[583]) );
  XNOR U4565 ( .A(b[582]), .B(n470), .Z(c[582]) );
  XNOR U4566 ( .A(b[581]), .B(n471), .Z(c[581]) );
  XNOR U4567 ( .A(b[580]), .B(n472), .Z(c[580]) );
  XNOR U4568 ( .A(b[57]), .B(n473), .Z(c[57]) );
  XNOR U4569 ( .A(b[579]), .B(n474), .Z(c[579]) );
  XNOR U4570 ( .A(b[578]), .B(n475), .Z(c[578]) );
  XNOR U4571 ( .A(b[577]), .B(n476), .Z(c[577]) );
  XNOR U4572 ( .A(b[576]), .B(n477), .Z(c[576]) );
  XNOR U4573 ( .A(b[575]), .B(n478), .Z(c[575]) );
  XNOR U4574 ( .A(b[574]), .B(n479), .Z(c[574]) );
  XNOR U4575 ( .A(b[573]), .B(n480), .Z(c[573]) );
  XNOR U4576 ( .A(b[572]), .B(n481), .Z(c[572]) );
  XNOR U4577 ( .A(b[571]), .B(n482), .Z(c[571]) );
  XNOR U4578 ( .A(b[570]), .B(n483), .Z(c[570]) );
  XNOR U4579 ( .A(b[56]), .B(n484), .Z(c[56]) );
  XNOR U4580 ( .A(b[569]), .B(n485), .Z(c[569]) );
  XNOR U4581 ( .A(b[568]), .B(n486), .Z(c[568]) );
  XNOR U4582 ( .A(b[567]), .B(n487), .Z(c[567]) );
  XNOR U4583 ( .A(b[566]), .B(n488), .Z(c[566]) );
  XNOR U4584 ( .A(b[565]), .B(n489), .Z(c[565]) );
  XNOR U4585 ( .A(b[564]), .B(n490), .Z(c[564]) );
  XNOR U4586 ( .A(b[563]), .B(n491), .Z(c[563]) );
  XNOR U4587 ( .A(b[562]), .B(n492), .Z(c[562]) );
  XNOR U4588 ( .A(b[561]), .B(n493), .Z(c[561]) );
  XNOR U4589 ( .A(b[560]), .B(n494), .Z(c[560]) );
  XNOR U4590 ( .A(b[55]), .B(n495), .Z(c[55]) );
  XNOR U4591 ( .A(b[559]), .B(n496), .Z(c[559]) );
  XNOR U4592 ( .A(b[558]), .B(n497), .Z(c[558]) );
  XNOR U4593 ( .A(b[557]), .B(n498), .Z(c[557]) );
  XNOR U4594 ( .A(b[556]), .B(n499), .Z(c[556]) );
  XNOR U4595 ( .A(b[555]), .B(n500), .Z(c[555]) );
  XNOR U4596 ( .A(b[554]), .B(n501), .Z(c[554]) );
  XNOR U4597 ( .A(b[553]), .B(n502), .Z(c[553]) );
  XNOR U4598 ( .A(b[552]), .B(n503), .Z(c[552]) );
  XNOR U4599 ( .A(b[551]), .B(n504), .Z(c[551]) );
  XNOR U4600 ( .A(b[550]), .B(n505), .Z(c[550]) );
  XNOR U4601 ( .A(b[54]), .B(n506), .Z(c[54]) );
  XNOR U4602 ( .A(b[549]), .B(n507), .Z(c[549]) );
  XNOR U4603 ( .A(b[548]), .B(n508), .Z(c[548]) );
  XNOR U4604 ( .A(b[547]), .B(n509), .Z(c[547]) );
  XNOR U4605 ( .A(b[546]), .B(n510), .Z(c[546]) );
  XNOR U4606 ( .A(b[545]), .B(n511), .Z(c[545]) );
  XNOR U4607 ( .A(b[544]), .B(n512), .Z(c[544]) );
  XNOR U4608 ( .A(b[543]), .B(n513), .Z(c[543]) );
  XNOR U4609 ( .A(b[542]), .B(n514), .Z(c[542]) );
  XNOR U4610 ( .A(b[541]), .B(n515), .Z(c[541]) );
  XNOR U4611 ( .A(b[540]), .B(n516), .Z(c[540]) );
  XNOR U4612 ( .A(b[53]), .B(n517), .Z(c[53]) );
  XNOR U4613 ( .A(b[539]), .B(n518), .Z(c[539]) );
  XNOR U4614 ( .A(b[538]), .B(n519), .Z(c[538]) );
  XNOR U4615 ( .A(b[537]), .B(n520), .Z(c[537]) );
  XNOR U4616 ( .A(b[536]), .B(n521), .Z(c[536]) );
  XNOR U4617 ( .A(b[535]), .B(n522), .Z(c[535]) );
  XNOR U4618 ( .A(b[534]), .B(n523), .Z(c[534]) );
  XNOR U4619 ( .A(b[533]), .B(n524), .Z(c[533]) );
  XNOR U4620 ( .A(b[532]), .B(n525), .Z(c[532]) );
  XNOR U4621 ( .A(b[531]), .B(n526), .Z(c[531]) );
  XNOR U4622 ( .A(b[530]), .B(n527), .Z(c[530]) );
  XNOR U4623 ( .A(b[52]), .B(n528), .Z(c[52]) );
  XNOR U4624 ( .A(b[529]), .B(n529), .Z(c[529]) );
  XNOR U4625 ( .A(b[528]), .B(n530), .Z(c[528]) );
  XNOR U4626 ( .A(b[527]), .B(n531), .Z(c[527]) );
  XNOR U4627 ( .A(b[526]), .B(n532), .Z(c[526]) );
  XNOR U4628 ( .A(b[525]), .B(n533), .Z(c[525]) );
  XNOR U4629 ( .A(b[524]), .B(n534), .Z(c[524]) );
  XNOR U4630 ( .A(b[523]), .B(n535), .Z(c[523]) );
  XNOR U4631 ( .A(b[522]), .B(n536), .Z(c[522]) );
  XNOR U4632 ( .A(b[521]), .B(n537), .Z(c[521]) );
  XNOR U4633 ( .A(b[520]), .B(n538), .Z(c[520]) );
  XNOR U4634 ( .A(b[51]), .B(n539), .Z(c[51]) );
  XNOR U4635 ( .A(b[519]), .B(n540), .Z(c[519]) );
  XNOR U4636 ( .A(b[518]), .B(n541), .Z(c[518]) );
  XNOR U4637 ( .A(b[517]), .B(n542), .Z(c[517]) );
  XNOR U4638 ( .A(b[516]), .B(n543), .Z(c[516]) );
  XNOR U4639 ( .A(b[515]), .B(n544), .Z(c[515]) );
  XNOR U4640 ( .A(b[514]), .B(n545), .Z(c[514]) );
  XNOR U4641 ( .A(b[513]), .B(n546), .Z(c[513]) );
  XNOR U4642 ( .A(b[512]), .B(n547), .Z(c[512]) );
  XNOR U4643 ( .A(b[511]), .B(n548), .Z(c[511]) );
  XNOR U4644 ( .A(b[510]), .B(n549), .Z(c[510]) );
  XNOR U4645 ( .A(b[50]), .B(n550), .Z(c[50]) );
  XNOR U4646 ( .A(b[509]), .B(n551), .Z(c[509]) );
  XNOR U4647 ( .A(b[508]), .B(n552), .Z(c[508]) );
  XNOR U4648 ( .A(b[507]), .B(n553), .Z(c[507]) );
  XNOR U4649 ( .A(b[506]), .B(n554), .Z(c[506]) );
  XNOR U4650 ( .A(b[505]), .B(n555), .Z(c[505]) );
  XNOR U4651 ( .A(b[504]), .B(n556), .Z(c[504]) );
  XNOR U4652 ( .A(b[503]), .B(n557), .Z(c[503]) );
  XNOR U4653 ( .A(b[502]), .B(n558), .Z(c[502]) );
  XNOR U4654 ( .A(b[501]), .B(n559), .Z(c[501]) );
  XNOR U4655 ( .A(b[500]), .B(n560), .Z(c[500]) );
  XNOR U4656 ( .A(b[4]), .B(n561), .Z(c[4]) );
  XNOR U4657 ( .A(b[49]), .B(n562), .Z(c[49]) );
  XNOR U4658 ( .A(b[499]), .B(n563), .Z(c[499]) );
  XNOR U4659 ( .A(b[498]), .B(n564), .Z(c[498]) );
  XNOR U4660 ( .A(b[497]), .B(n565), .Z(c[497]) );
  XNOR U4661 ( .A(b[496]), .B(n566), .Z(c[496]) );
  XNOR U4662 ( .A(b[495]), .B(n567), .Z(c[495]) );
  XNOR U4663 ( .A(b[494]), .B(n568), .Z(c[494]) );
  XNOR U4664 ( .A(b[493]), .B(n569), .Z(c[493]) );
  XNOR U4665 ( .A(b[492]), .B(n570), .Z(c[492]) );
  XNOR U4666 ( .A(b[491]), .B(n571), .Z(c[491]) );
  XNOR U4667 ( .A(b[490]), .B(n572), .Z(c[490]) );
  XNOR U4668 ( .A(b[48]), .B(n573), .Z(c[48]) );
  XNOR U4669 ( .A(b[489]), .B(n574), .Z(c[489]) );
  XNOR U4670 ( .A(b[488]), .B(n575), .Z(c[488]) );
  XNOR U4671 ( .A(b[487]), .B(n576), .Z(c[487]) );
  XNOR U4672 ( .A(b[486]), .B(n577), .Z(c[486]) );
  XNOR U4673 ( .A(b[485]), .B(n578), .Z(c[485]) );
  XNOR U4674 ( .A(b[484]), .B(n579), .Z(c[484]) );
  XNOR U4675 ( .A(b[483]), .B(n580), .Z(c[483]) );
  XNOR U4676 ( .A(b[482]), .B(n581), .Z(c[482]) );
  XNOR U4677 ( .A(b[481]), .B(n582), .Z(c[481]) );
  XNOR U4678 ( .A(b[480]), .B(n583), .Z(c[480]) );
  XNOR U4679 ( .A(b[47]), .B(n584), .Z(c[47]) );
  XNOR U4680 ( .A(b[479]), .B(n585), .Z(c[479]) );
  XNOR U4681 ( .A(b[478]), .B(n586), .Z(c[478]) );
  XNOR U4682 ( .A(b[477]), .B(n587), .Z(c[477]) );
  XNOR U4683 ( .A(b[476]), .B(n588), .Z(c[476]) );
  XNOR U4684 ( .A(b[475]), .B(n589), .Z(c[475]) );
  XNOR U4685 ( .A(b[474]), .B(n590), .Z(c[474]) );
  XNOR U4686 ( .A(b[473]), .B(n591), .Z(c[473]) );
  XNOR U4687 ( .A(b[472]), .B(n592), .Z(c[472]) );
  XNOR U4688 ( .A(b[471]), .B(n593), .Z(c[471]) );
  XNOR U4689 ( .A(b[470]), .B(n594), .Z(c[470]) );
  XNOR U4690 ( .A(b[46]), .B(n595), .Z(c[46]) );
  XNOR U4691 ( .A(b[469]), .B(n596), .Z(c[469]) );
  XNOR U4692 ( .A(b[468]), .B(n597), .Z(c[468]) );
  XNOR U4693 ( .A(b[467]), .B(n598), .Z(c[467]) );
  XNOR U4694 ( .A(b[466]), .B(n599), .Z(c[466]) );
  XNOR U4695 ( .A(b[465]), .B(n600), .Z(c[465]) );
  XNOR U4696 ( .A(b[464]), .B(n601), .Z(c[464]) );
  XNOR U4697 ( .A(b[463]), .B(n602), .Z(c[463]) );
  XNOR U4698 ( .A(b[462]), .B(n603), .Z(c[462]) );
  XNOR U4699 ( .A(b[461]), .B(n604), .Z(c[461]) );
  XNOR U4700 ( .A(b[460]), .B(n605), .Z(c[460]) );
  XNOR U4701 ( .A(b[45]), .B(n606), .Z(c[45]) );
  XNOR U4702 ( .A(b[459]), .B(n607), .Z(c[459]) );
  XNOR U4703 ( .A(b[458]), .B(n608), .Z(c[458]) );
  XNOR U4704 ( .A(b[457]), .B(n609), .Z(c[457]) );
  XNOR U4705 ( .A(b[456]), .B(n610), .Z(c[456]) );
  XNOR U4706 ( .A(b[455]), .B(n611), .Z(c[455]) );
  XNOR U4707 ( .A(b[454]), .B(n612), .Z(c[454]) );
  XNOR U4708 ( .A(b[453]), .B(n613), .Z(c[453]) );
  XNOR U4709 ( .A(b[452]), .B(n614), .Z(c[452]) );
  XNOR U4710 ( .A(b[451]), .B(n615), .Z(c[451]) );
  XNOR U4711 ( .A(b[450]), .B(n616), .Z(c[450]) );
  XNOR U4712 ( .A(b[44]), .B(n617), .Z(c[44]) );
  XNOR U4713 ( .A(b[449]), .B(n618), .Z(c[449]) );
  XNOR U4714 ( .A(b[448]), .B(n619), .Z(c[448]) );
  XNOR U4715 ( .A(b[447]), .B(n620), .Z(c[447]) );
  XNOR U4716 ( .A(b[446]), .B(n621), .Z(c[446]) );
  XNOR U4717 ( .A(b[445]), .B(n622), .Z(c[445]) );
  XNOR U4718 ( .A(b[444]), .B(n623), .Z(c[444]) );
  XNOR U4719 ( .A(b[443]), .B(n624), .Z(c[443]) );
  XNOR U4720 ( .A(b[442]), .B(n625), .Z(c[442]) );
  XNOR U4721 ( .A(b[441]), .B(n626), .Z(c[441]) );
  XNOR U4722 ( .A(b[440]), .B(n627), .Z(c[440]) );
  XNOR U4723 ( .A(b[43]), .B(n628), .Z(c[43]) );
  XNOR U4724 ( .A(b[439]), .B(n629), .Z(c[439]) );
  XNOR U4725 ( .A(b[438]), .B(n630), .Z(c[438]) );
  XNOR U4726 ( .A(b[437]), .B(n631), .Z(c[437]) );
  XNOR U4727 ( .A(b[436]), .B(n632), .Z(c[436]) );
  XNOR U4728 ( .A(b[435]), .B(n633), .Z(c[435]) );
  XNOR U4729 ( .A(b[434]), .B(n634), .Z(c[434]) );
  XNOR U4730 ( .A(b[433]), .B(n635), .Z(c[433]) );
  XNOR U4731 ( .A(b[432]), .B(n636), .Z(c[432]) );
  XNOR U4732 ( .A(b[431]), .B(n637), .Z(c[431]) );
  XNOR U4733 ( .A(b[430]), .B(n638), .Z(c[430]) );
  XNOR U4734 ( .A(b[42]), .B(n639), .Z(c[42]) );
  XNOR U4735 ( .A(b[429]), .B(n640), .Z(c[429]) );
  XNOR U4736 ( .A(b[428]), .B(n641), .Z(c[428]) );
  XNOR U4737 ( .A(b[427]), .B(n642), .Z(c[427]) );
  XNOR U4738 ( .A(b[426]), .B(n643), .Z(c[426]) );
  XNOR U4739 ( .A(b[425]), .B(n644), .Z(c[425]) );
  XNOR U4740 ( .A(b[424]), .B(n645), .Z(c[424]) );
  XNOR U4741 ( .A(b[423]), .B(n646), .Z(c[423]) );
  XNOR U4742 ( .A(b[422]), .B(n647), .Z(c[422]) );
  XNOR U4743 ( .A(b[421]), .B(n648), .Z(c[421]) );
  XNOR U4744 ( .A(b[420]), .B(n649), .Z(c[420]) );
  XNOR U4745 ( .A(b[41]), .B(n650), .Z(c[41]) );
  XNOR U4746 ( .A(b[419]), .B(n651), .Z(c[419]) );
  XNOR U4747 ( .A(b[418]), .B(n652), .Z(c[418]) );
  XNOR U4748 ( .A(b[417]), .B(n653), .Z(c[417]) );
  XNOR U4749 ( .A(b[416]), .B(n654), .Z(c[416]) );
  XNOR U4750 ( .A(b[415]), .B(n655), .Z(c[415]) );
  XNOR U4751 ( .A(b[414]), .B(n656), .Z(c[414]) );
  XNOR U4752 ( .A(b[413]), .B(n657), .Z(c[413]) );
  XNOR U4753 ( .A(b[412]), .B(n658), .Z(c[412]) );
  XNOR U4754 ( .A(b[411]), .B(n659), .Z(c[411]) );
  XNOR U4755 ( .A(b[410]), .B(n660), .Z(c[410]) );
  XNOR U4756 ( .A(b[40]), .B(n661), .Z(c[40]) );
  XNOR U4757 ( .A(b[409]), .B(n662), .Z(c[409]) );
  XNOR U4758 ( .A(b[4095]), .B(n5), .Z(c[4095]) );
  XNOR U4759 ( .A(a[4095]), .B(n3), .Z(n5) );
  XNOR U4760 ( .A(n663), .B(n664), .Z(n3) );
  ANDN U4761 ( .B(n665), .A(n666), .Z(n663) );
  XNOR U4762 ( .A(b[4094]), .B(n664), .Z(n665) );
  XNOR U4763 ( .A(b[4094]), .B(n666), .Z(c[4094]) );
  XOR U4764 ( .A(n667), .B(n668), .Z(n664) );
  ANDN U4765 ( .B(n669), .A(n670), .Z(n667) );
  XNOR U4766 ( .A(b[4093]), .B(n668), .Z(n669) );
  XNOR U4767 ( .A(b[4093]), .B(n670), .Z(c[4093]) );
  XOR U4768 ( .A(n671), .B(n672), .Z(n668) );
  ANDN U4769 ( .B(n673), .A(n674), .Z(n671) );
  XNOR U4770 ( .A(b[4092]), .B(n672), .Z(n673) );
  XNOR U4771 ( .A(b[4092]), .B(n674), .Z(c[4092]) );
  XOR U4772 ( .A(n675), .B(n676), .Z(n672) );
  ANDN U4773 ( .B(n677), .A(n678), .Z(n675) );
  XNOR U4774 ( .A(b[4091]), .B(n676), .Z(n677) );
  XNOR U4775 ( .A(b[4091]), .B(n678), .Z(c[4091]) );
  XOR U4776 ( .A(n679), .B(n680), .Z(n676) );
  ANDN U4777 ( .B(n681), .A(n682), .Z(n679) );
  XNOR U4778 ( .A(b[4090]), .B(n680), .Z(n681) );
  XNOR U4779 ( .A(b[4090]), .B(n682), .Z(c[4090]) );
  XOR U4780 ( .A(n683), .B(n684), .Z(n680) );
  ANDN U4781 ( .B(n685), .A(n686), .Z(n683) );
  XNOR U4782 ( .A(b[4089]), .B(n684), .Z(n685) );
  XNOR U4783 ( .A(b[408]), .B(n687), .Z(c[408]) );
  XNOR U4784 ( .A(b[4089]), .B(n686), .Z(c[4089]) );
  XOR U4785 ( .A(n688), .B(n689), .Z(n684) );
  ANDN U4786 ( .B(n690), .A(n691), .Z(n688) );
  XNOR U4787 ( .A(b[4088]), .B(n689), .Z(n690) );
  XNOR U4788 ( .A(b[4088]), .B(n691), .Z(c[4088]) );
  XOR U4789 ( .A(n692), .B(n693), .Z(n689) );
  ANDN U4790 ( .B(n694), .A(n695), .Z(n692) );
  XNOR U4791 ( .A(b[4087]), .B(n693), .Z(n694) );
  XNOR U4792 ( .A(b[4087]), .B(n695), .Z(c[4087]) );
  XOR U4793 ( .A(n696), .B(n697), .Z(n693) );
  ANDN U4794 ( .B(n698), .A(n699), .Z(n696) );
  XNOR U4795 ( .A(b[4086]), .B(n697), .Z(n698) );
  XNOR U4796 ( .A(b[4086]), .B(n699), .Z(c[4086]) );
  XOR U4797 ( .A(n700), .B(n701), .Z(n697) );
  ANDN U4798 ( .B(n702), .A(n703), .Z(n700) );
  XNOR U4799 ( .A(b[4085]), .B(n701), .Z(n702) );
  XNOR U4800 ( .A(b[4085]), .B(n703), .Z(c[4085]) );
  XOR U4801 ( .A(n704), .B(n705), .Z(n701) );
  ANDN U4802 ( .B(n706), .A(n707), .Z(n704) );
  XNOR U4803 ( .A(b[4084]), .B(n705), .Z(n706) );
  XNOR U4804 ( .A(b[4084]), .B(n707), .Z(c[4084]) );
  XOR U4805 ( .A(n708), .B(n709), .Z(n705) );
  ANDN U4806 ( .B(n710), .A(n711), .Z(n708) );
  XNOR U4807 ( .A(b[4083]), .B(n709), .Z(n710) );
  XNOR U4808 ( .A(b[4083]), .B(n711), .Z(c[4083]) );
  XOR U4809 ( .A(n712), .B(n713), .Z(n709) );
  ANDN U4810 ( .B(n714), .A(n715), .Z(n712) );
  XNOR U4811 ( .A(b[4082]), .B(n713), .Z(n714) );
  XNOR U4812 ( .A(b[4082]), .B(n715), .Z(c[4082]) );
  XOR U4813 ( .A(n716), .B(n717), .Z(n713) );
  ANDN U4814 ( .B(n718), .A(n719), .Z(n716) );
  XNOR U4815 ( .A(b[4081]), .B(n717), .Z(n718) );
  XNOR U4816 ( .A(b[4081]), .B(n719), .Z(c[4081]) );
  XOR U4817 ( .A(n720), .B(n721), .Z(n717) );
  ANDN U4818 ( .B(n722), .A(n723), .Z(n720) );
  XNOR U4819 ( .A(b[4080]), .B(n721), .Z(n722) );
  XNOR U4820 ( .A(b[4080]), .B(n723), .Z(c[4080]) );
  XOR U4821 ( .A(n724), .B(n725), .Z(n721) );
  ANDN U4822 ( .B(n726), .A(n727), .Z(n724) );
  XNOR U4823 ( .A(b[4079]), .B(n725), .Z(n726) );
  XNOR U4824 ( .A(b[407]), .B(n728), .Z(c[407]) );
  XNOR U4825 ( .A(b[4079]), .B(n727), .Z(c[4079]) );
  XOR U4826 ( .A(n729), .B(n730), .Z(n725) );
  ANDN U4827 ( .B(n731), .A(n732), .Z(n729) );
  XNOR U4828 ( .A(b[4078]), .B(n730), .Z(n731) );
  XNOR U4829 ( .A(b[4078]), .B(n732), .Z(c[4078]) );
  XOR U4830 ( .A(n733), .B(n734), .Z(n730) );
  ANDN U4831 ( .B(n735), .A(n736), .Z(n733) );
  XNOR U4832 ( .A(b[4077]), .B(n734), .Z(n735) );
  XNOR U4833 ( .A(b[4077]), .B(n736), .Z(c[4077]) );
  XOR U4834 ( .A(n737), .B(n738), .Z(n734) );
  ANDN U4835 ( .B(n739), .A(n740), .Z(n737) );
  XNOR U4836 ( .A(b[4076]), .B(n738), .Z(n739) );
  XNOR U4837 ( .A(b[4076]), .B(n740), .Z(c[4076]) );
  XOR U4838 ( .A(n741), .B(n742), .Z(n738) );
  ANDN U4839 ( .B(n743), .A(n744), .Z(n741) );
  XNOR U4840 ( .A(b[4075]), .B(n742), .Z(n743) );
  XNOR U4841 ( .A(b[4075]), .B(n744), .Z(c[4075]) );
  XOR U4842 ( .A(n745), .B(n746), .Z(n742) );
  ANDN U4843 ( .B(n747), .A(n748), .Z(n745) );
  XNOR U4844 ( .A(b[4074]), .B(n746), .Z(n747) );
  XNOR U4845 ( .A(b[4074]), .B(n748), .Z(c[4074]) );
  XOR U4846 ( .A(n749), .B(n750), .Z(n746) );
  ANDN U4847 ( .B(n751), .A(n752), .Z(n749) );
  XNOR U4848 ( .A(b[4073]), .B(n750), .Z(n751) );
  XNOR U4849 ( .A(b[4073]), .B(n752), .Z(c[4073]) );
  XOR U4850 ( .A(n753), .B(n754), .Z(n750) );
  ANDN U4851 ( .B(n755), .A(n756), .Z(n753) );
  XNOR U4852 ( .A(b[4072]), .B(n754), .Z(n755) );
  XNOR U4853 ( .A(b[4072]), .B(n756), .Z(c[4072]) );
  XOR U4854 ( .A(n757), .B(n758), .Z(n754) );
  ANDN U4855 ( .B(n759), .A(n760), .Z(n757) );
  XNOR U4856 ( .A(b[4071]), .B(n758), .Z(n759) );
  XNOR U4857 ( .A(b[4071]), .B(n760), .Z(c[4071]) );
  XOR U4858 ( .A(n761), .B(n762), .Z(n758) );
  ANDN U4859 ( .B(n763), .A(n764), .Z(n761) );
  XNOR U4860 ( .A(b[4070]), .B(n762), .Z(n763) );
  XNOR U4861 ( .A(b[4070]), .B(n764), .Z(c[4070]) );
  XOR U4862 ( .A(n765), .B(n766), .Z(n762) );
  ANDN U4863 ( .B(n767), .A(n768), .Z(n765) );
  XNOR U4864 ( .A(b[4069]), .B(n766), .Z(n767) );
  XNOR U4865 ( .A(b[406]), .B(n769), .Z(c[406]) );
  XNOR U4866 ( .A(b[4069]), .B(n768), .Z(c[4069]) );
  XOR U4867 ( .A(n770), .B(n771), .Z(n766) );
  ANDN U4868 ( .B(n772), .A(n773), .Z(n770) );
  XNOR U4869 ( .A(b[4068]), .B(n771), .Z(n772) );
  XNOR U4870 ( .A(b[4068]), .B(n773), .Z(c[4068]) );
  XOR U4871 ( .A(n774), .B(n775), .Z(n771) );
  ANDN U4872 ( .B(n776), .A(n777), .Z(n774) );
  XNOR U4873 ( .A(b[4067]), .B(n775), .Z(n776) );
  XNOR U4874 ( .A(b[4067]), .B(n777), .Z(c[4067]) );
  XOR U4875 ( .A(n778), .B(n779), .Z(n775) );
  ANDN U4876 ( .B(n780), .A(n781), .Z(n778) );
  XNOR U4877 ( .A(b[4066]), .B(n779), .Z(n780) );
  XNOR U4878 ( .A(b[4066]), .B(n781), .Z(c[4066]) );
  XOR U4879 ( .A(n782), .B(n783), .Z(n779) );
  ANDN U4880 ( .B(n784), .A(n785), .Z(n782) );
  XNOR U4881 ( .A(b[4065]), .B(n783), .Z(n784) );
  XNOR U4882 ( .A(b[4065]), .B(n785), .Z(c[4065]) );
  XOR U4883 ( .A(n786), .B(n787), .Z(n783) );
  ANDN U4884 ( .B(n788), .A(n789), .Z(n786) );
  XNOR U4885 ( .A(b[4064]), .B(n787), .Z(n788) );
  XNOR U4886 ( .A(b[4064]), .B(n789), .Z(c[4064]) );
  XOR U4887 ( .A(n790), .B(n791), .Z(n787) );
  ANDN U4888 ( .B(n792), .A(n793), .Z(n790) );
  XNOR U4889 ( .A(b[4063]), .B(n791), .Z(n792) );
  XNOR U4890 ( .A(b[4063]), .B(n793), .Z(c[4063]) );
  XOR U4891 ( .A(n794), .B(n795), .Z(n791) );
  ANDN U4892 ( .B(n796), .A(n797), .Z(n794) );
  XNOR U4893 ( .A(b[4062]), .B(n795), .Z(n796) );
  XNOR U4894 ( .A(b[4062]), .B(n797), .Z(c[4062]) );
  XOR U4895 ( .A(n798), .B(n799), .Z(n795) );
  ANDN U4896 ( .B(n800), .A(n801), .Z(n798) );
  XNOR U4897 ( .A(b[4061]), .B(n799), .Z(n800) );
  XNOR U4898 ( .A(b[4061]), .B(n801), .Z(c[4061]) );
  XOR U4899 ( .A(n802), .B(n803), .Z(n799) );
  ANDN U4900 ( .B(n804), .A(n805), .Z(n802) );
  XNOR U4901 ( .A(b[4060]), .B(n803), .Z(n804) );
  XNOR U4902 ( .A(b[4060]), .B(n805), .Z(c[4060]) );
  XOR U4903 ( .A(n806), .B(n807), .Z(n803) );
  ANDN U4904 ( .B(n808), .A(n809), .Z(n806) );
  XNOR U4905 ( .A(b[4059]), .B(n807), .Z(n808) );
  XNOR U4906 ( .A(b[405]), .B(n810), .Z(c[405]) );
  XNOR U4907 ( .A(b[4059]), .B(n809), .Z(c[4059]) );
  XOR U4908 ( .A(n811), .B(n812), .Z(n807) );
  ANDN U4909 ( .B(n813), .A(n814), .Z(n811) );
  XNOR U4910 ( .A(b[4058]), .B(n812), .Z(n813) );
  XNOR U4911 ( .A(b[4058]), .B(n814), .Z(c[4058]) );
  XOR U4912 ( .A(n815), .B(n816), .Z(n812) );
  ANDN U4913 ( .B(n817), .A(n818), .Z(n815) );
  XNOR U4914 ( .A(b[4057]), .B(n816), .Z(n817) );
  XNOR U4915 ( .A(b[4057]), .B(n818), .Z(c[4057]) );
  XOR U4916 ( .A(n819), .B(n820), .Z(n816) );
  ANDN U4917 ( .B(n821), .A(n822), .Z(n819) );
  XNOR U4918 ( .A(b[4056]), .B(n820), .Z(n821) );
  XNOR U4919 ( .A(b[4056]), .B(n822), .Z(c[4056]) );
  XOR U4920 ( .A(n823), .B(n824), .Z(n820) );
  ANDN U4921 ( .B(n825), .A(n826), .Z(n823) );
  XNOR U4922 ( .A(b[4055]), .B(n824), .Z(n825) );
  XNOR U4923 ( .A(b[4055]), .B(n826), .Z(c[4055]) );
  XOR U4924 ( .A(n827), .B(n828), .Z(n824) );
  ANDN U4925 ( .B(n829), .A(n830), .Z(n827) );
  XNOR U4926 ( .A(b[4054]), .B(n828), .Z(n829) );
  XNOR U4927 ( .A(b[4054]), .B(n830), .Z(c[4054]) );
  XOR U4928 ( .A(n831), .B(n832), .Z(n828) );
  ANDN U4929 ( .B(n833), .A(n834), .Z(n831) );
  XNOR U4930 ( .A(b[4053]), .B(n832), .Z(n833) );
  XNOR U4931 ( .A(b[4053]), .B(n834), .Z(c[4053]) );
  XOR U4932 ( .A(n835), .B(n836), .Z(n832) );
  ANDN U4933 ( .B(n837), .A(n838), .Z(n835) );
  XNOR U4934 ( .A(b[4052]), .B(n836), .Z(n837) );
  XNOR U4935 ( .A(b[4052]), .B(n838), .Z(c[4052]) );
  XOR U4936 ( .A(n839), .B(n840), .Z(n836) );
  ANDN U4937 ( .B(n841), .A(n842), .Z(n839) );
  XNOR U4938 ( .A(b[4051]), .B(n840), .Z(n841) );
  XNOR U4939 ( .A(b[4051]), .B(n842), .Z(c[4051]) );
  XOR U4940 ( .A(n843), .B(n844), .Z(n840) );
  ANDN U4941 ( .B(n845), .A(n846), .Z(n843) );
  XNOR U4942 ( .A(b[4050]), .B(n844), .Z(n845) );
  XNOR U4943 ( .A(b[4050]), .B(n846), .Z(c[4050]) );
  XOR U4944 ( .A(n847), .B(n848), .Z(n844) );
  ANDN U4945 ( .B(n849), .A(n850), .Z(n847) );
  XNOR U4946 ( .A(b[4049]), .B(n848), .Z(n849) );
  XNOR U4947 ( .A(b[404]), .B(n851), .Z(c[404]) );
  XNOR U4948 ( .A(b[4049]), .B(n850), .Z(c[4049]) );
  XOR U4949 ( .A(n852), .B(n853), .Z(n848) );
  ANDN U4950 ( .B(n854), .A(n855), .Z(n852) );
  XNOR U4951 ( .A(b[4048]), .B(n853), .Z(n854) );
  XNOR U4952 ( .A(b[4048]), .B(n855), .Z(c[4048]) );
  XOR U4953 ( .A(n856), .B(n857), .Z(n853) );
  ANDN U4954 ( .B(n858), .A(n859), .Z(n856) );
  XNOR U4955 ( .A(b[4047]), .B(n857), .Z(n858) );
  XNOR U4956 ( .A(b[4047]), .B(n859), .Z(c[4047]) );
  XOR U4957 ( .A(n860), .B(n861), .Z(n857) );
  ANDN U4958 ( .B(n862), .A(n863), .Z(n860) );
  XNOR U4959 ( .A(b[4046]), .B(n861), .Z(n862) );
  XNOR U4960 ( .A(b[4046]), .B(n863), .Z(c[4046]) );
  XOR U4961 ( .A(n864), .B(n865), .Z(n861) );
  ANDN U4962 ( .B(n866), .A(n867), .Z(n864) );
  XNOR U4963 ( .A(b[4045]), .B(n865), .Z(n866) );
  XNOR U4964 ( .A(b[4045]), .B(n867), .Z(c[4045]) );
  XOR U4965 ( .A(n868), .B(n869), .Z(n865) );
  ANDN U4966 ( .B(n870), .A(n871), .Z(n868) );
  XNOR U4967 ( .A(b[4044]), .B(n869), .Z(n870) );
  XNOR U4968 ( .A(b[4044]), .B(n871), .Z(c[4044]) );
  XOR U4969 ( .A(n872), .B(n873), .Z(n869) );
  ANDN U4970 ( .B(n874), .A(n875), .Z(n872) );
  XNOR U4971 ( .A(b[4043]), .B(n873), .Z(n874) );
  XNOR U4972 ( .A(b[4043]), .B(n875), .Z(c[4043]) );
  XOR U4973 ( .A(n876), .B(n877), .Z(n873) );
  ANDN U4974 ( .B(n878), .A(n879), .Z(n876) );
  XNOR U4975 ( .A(b[4042]), .B(n877), .Z(n878) );
  XNOR U4976 ( .A(b[4042]), .B(n879), .Z(c[4042]) );
  XOR U4977 ( .A(n880), .B(n881), .Z(n877) );
  ANDN U4978 ( .B(n882), .A(n883), .Z(n880) );
  XNOR U4979 ( .A(b[4041]), .B(n881), .Z(n882) );
  XNOR U4980 ( .A(b[4041]), .B(n883), .Z(c[4041]) );
  XOR U4981 ( .A(n884), .B(n885), .Z(n881) );
  ANDN U4982 ( .B(n886), .A(n887), .Z(n884) );
  XNOR U4983 ( .A(b[4040]), .B(n885), .Z(n886) );
  XNOR U4984 ( .A(b[4040]), .B(n887), .Z(c[4040]) );
  XOR U4985 ( .A(n888), .B(n889), .Z(n885) );
  ANDN U4986 ( .B(n890), .A(n891), .Z(n888) );
  XNOR U4987 ( .A(b[4039]), .B(n889), .Z(n890) );
  XNOR U4988 ( .A(b[403]), .B(n892), .Z(c[403]) );
  XNOR U4989 ( .A(b[4039]), .B(n891), .Z(c[4039]) );
  XOR U4990 ( .A(n893), .B(n894), .Z(n889) );
  ANDN U4991 ( .B(n895), .A(n896), .Z(n893) );
  XNOR U4992 ( .A(b[4038]), .B(n894), .Z(n895) );
  XNOR U4993 ( .A(b[4038]), .B(n896), .Z(c[4038]) );
  XOR U4994 ( .A(n897), .B(n898), .Z(n894) );
  ANDN U4995 ( .B(n899), .A(n900), .Z(n897) );
  XNOR U4996 ( .A(b[4037]), .B(n898), .Z(n899) );
  XNOR U4997 ( .A(b[4037]), .B(n900), .Z(c[4037]) );
  XOR U4998 ( .A(n901), .B(n902), .Z(n898) );
  ANDN U4999 ( .B(n903), .A(n904), .Z(n901) );
  XNOR U5000 ( .A(b[4036]), .B(n902), .Z(n903) );
  XNOR U5001 ( .A(b[4036]), .B(n904), .Z(c[4036]) );
  XOR U5002 ( .A(n905), .B(n906), .Z(n902) );
  ANDN U5003 ( .B(n907), .A(n908), .Z(n905) );
  XNOR U5004 ( .A(b[4035]), .B(n906), .Z(n907) );
  XNOR U5005 ( .A(b[4035]), .B(n908), .Z(c[4035]) );
  XOR U5006 ( .A(n909), .B(n910), .Z(n906) );
  ANDN U5007 ( .B(n911), .A(n912), .Z(n909) );
  XNOR U5008 ( .A(b[4034]), .B(n910), .Z(n911) );
  XNOR U5009 ( .A(b[4034]), .B(n912), .Z(c[4034]) );
  XOR U5010 ( .A(n913), .B(n914), .Z(n910) );
  ANDN U5011 ( .B(n915), .A(n916), .Z(n913) );
  XNOR U5012 ( .A(b[4033]), .B(n914), .Z(n915) );
  XNOR U5013 ( .A(b[4033]), .B(n916), .Z(c[4033]) );
  XOR U5014 ( .A(n917), .B(n918), .Z(n914) );
  ANDN U5015 ( .B(n919), .A(n920), .Z(n917) );
  XNOR U5016 ( .A(b[4032]), .B(n918), .Z(n919) );
  XNOR U5017 ( .A(b[4032]), .B(n920), .Z(c[4032]) );
  XOR U5018 ( .A(n921), .B(n922), .Z(n918) );
  ANDN U5019 ( .B(n923), .A(n924), .Z(n921) );
  XNOR U5020 ( .A(b[4031]), .B(n922), .Z(n923) );
  XNOR U5021 ( .A(b[4031]), .B(n924), .Z(c[4031]) );
  XOR U5022 ( .A(n925), .B(n926), .Z(n922) );
  ANDN U5023 ( .B(n927), .A(n928), .Z(n925) );
  XNOR U5024 ( .A(b[4030]), .B(n926), .Z(n927) );
  XNOR U5025 ( .A(b[4030]), .B(n928), .Z(c[4030]) );
  XOR U5026 ( .A(n929), .B(n930), .Z(n926) );
  ANDN U5027 ( .B(n931), .A(n932), .Z(n929) );
  XNOR U5028 ( .A(b[4029]), .B(n930), .Z(n931) );
  XNOR U5029 ( .A(b[402]), .B(n933), .Z(c[402]) );
  XNOR U5030 ( .A(b[4029]), .B(n932), .Z(c[4029]) );
  XOR U5031 ( .A(n934), .B(n935), .Z(n930) );
  ANDN U5032 ( .B(n936), .A(n937), .Z(n934) );
  XNOR U5033 ( .A(b[4028]), .B(n935), .Z(n936) );
  XNOR U5034 ( .A(b[4028]), .B(n937), .Z(c[4028]) );
  XOR U5035 ( .A(n938), .B(n939), .Z(n935) );
  ANDN U5036 ( .B(n940), .A(n941), .Z(n938) );
  XNOR U5037 ( .A(b[4027]), .B(n939), .Z(n940) );
  XNOR U5038 ( .A(b[4027]), .B(n941), .Z(c[4027]) );
  XOR U5039 ( .A(n942), .B(n943), .Z(n939) );
  ANDN U5040 ( .B(n944), .A(n945), .Z(n942) );
  XNOR U5041 ( .A(b[4026]), .B(n943), .Z(n944) );
  XNOR U5042 ( .A(b[4026]), .B(n945), .Z(c[4026]) );
  XOR U5043 ( .A(n946), .B(n947), .Z(n943) );
  ANDN U5044 ( .B(n948), .A(n949), .Z(n946) );
  XNOR U5045 ( .A(b[4025]), .B(n947), .Z(n948) );
  XNOR U5046 ( .A(b[4025]), .B(n949), .Z(c[4025]) );
  XOR U5047 ( .A(n950), .B(n951), .Z(n947) );
  ANDN U5048 ( .B(n952), .A(n953), .Z(n950) );
  XNOR U5049 ( .A(b[4024]), .B(n951), .Z(n952) );
  XNOR U5050 ( .A(b[4024]), .B(n953), .Z(c[4024]) );
  XOR U5051 ( .A(n954), .B(n955), .Z(n951) );
  ANDN U5052 ( .B(n956), .A(n957), .Z(n954) );
  XNOR U5053 ( .A(b[4023]), .B(n955), .Z(n956) );
  XNOR U5054 ( .A(b[4023]), .B(n957), .Z(c[4023]) );
  XOR U5055 ( .A(n958), .B(n959), .Z(n955) );
  ANDN U5056 ( .B(n960), .A(n961), .Z(n958) );
  XNOR U5057 ( .A(b[4022]), .B(n959), .Z(n960) );
  XNOR U5058 ( .A(b[4022]), .B(n961), .Z(c[4022]) );
  XOR U5059 ( .A(n962), .B(n963), .Z(n959) );
  ANDN U5060 ( .B(n964), .A(n965), .Z(n962) );
  XNOR U5061 ( .A(b[4021]), .B(n963), .Z(n964) );
  XNOR U5062 ( .A(b[4021]), .B(n965), .Z(c[4021]) );
  XOR U5063 ( .A(n966), .B(n967), .Z(n963) );
  ANDN U5064 ( .B(n968), .A(n969), .Z(n966) );
  XNOR U5065 ( .A(b[4020]), .B(n967), .Z(n968) );
  XNOR U5066 ( .A(b[4020]), .B(n969), .Z(c[4020]) );
  XOR U5067 ( .A(n970), .B(n971), .Z(n967) );
  ANDN U5068 ( .B(n972), .A(n973), .Z(n970) );
  XNOR U5069 ( .A(b[4019]), .B(n971), .Z(n972) );
  XNOR U5070 ( .A(b[401]), .B(n974), .Z(c[401]) );
  XNOR U5071 ( .A(b[4019]), .B(n973), .Z(c[4019]) );
  XOR U5072 ( .A(n975), .B(n976), .Z(n971) );
  ANDN U5073 ( .B(n977), .A(n978), .Z(n975) );
  XNOR U5074 ( .A(b[4018]), .B(n976), .Z(n977) );
  XNOR U5075 ( .A(b[4018]), .B(n978), .Z(c[4018]) );
  XOR U5076 ( .A(n979), .B(n980), .Z(n976) );
  ANDN U5077 ( .B(n981), .A(n982), .Z(n979) );
  XNOR U5078 ( .A(b[4017]), .B(n980), .Z(n981) );
  XNOR U5079 ( .A(b[4017]), .B(n982), .Z(c[4017]) );
  XOR U5080 ( .A(n983), .B(n984), .Z(n980) );
  ANDN U5081 ( .B(n985), .A(n986), .Z(n983) );
  XNOR U5082 ( .A(b[4016]), .B(n984), .Z(n985) );
  XNOR U5083 ( .A(b[4016]), .B(n986), .Z(c[4016]) );
  XOR U5084 ( .A(n987), .B(n988), .Z(n984) );
  ANDN U5085 ( .B(n989), .A(n990), .Z(n987) );
  XNOR U5086 ( .A(b[4015]), .B(n988), .Z(n989) );
  XNOR U5087 ( .A(b[4015]), .B(n990), .Z(c[4015]) );
  XOR U5088 ( .A(n991), .B(n992), .Z(n988) );
  ANDN U5089 ( .B(n993), .A(n994), .Z(n991) );
  XNOR U5090 ( .A(b[4014]), .B(n992), .Z(n993) );
  XNOR U5091 ( .A(b[4014]), .B(n994), .Z(c[4014]) );
  XOR U5092 ( .A(n995), .B(n996), .Z(n992) );
  ANDN U5093 ( .B(n997), .A(n998), .Z(n995) );
  XNOR U5094 ( .A(b[4013]), .B(n996), .Z(n997) );
  XNOR U5095 ( .A(b[4013]), .B(n998), .Z(c[4013]) );
  XOR U5096 ( .A(n999), .B(n1000), .Z(n996) );
  ANDN U5097 ( .B(n1001), .A(n1002), .Z(n999) );
  XNOR U5098 ( .A(b[4012]), .B(n1000), .Z(n1001) );
  XNOR U5099 ( .A(b[4012]), .B(n1002), .Z(c[4012]) );
  XOR U5100 ( .A(n1003), .B(n1004), .Z(n1000) );
  ANDN U5101 ( .B(n1005), .A(n1006), .Z(n1003) );
  XNOR U5102 ( .A(b[4011]), .B(n1004), .Z(n1005) );
  XNOR U5103 ( .A(b[4011]), .B(n1006), .Z(c[4011]) );
  XOR U5104 ( .A(n1007), .B(n1008), .Z(n1004) );
  ANDN U5105 ( .B(n1009), .A(n1010), .Z(n1007) );
  XNOR U5106 ( .A(b[4010]), .B(n1008), .Z(n1009) );
  XNOR U5107 ( .A(b[4010]), .B(n1010), .Z(c[4010]) );
  XOR U5108 ( .A(n1011), .B(n1012), .Z(n1008) );
  ANDN U5109 ( .B(n1013), .A(n1014), .Z(n1011) );
  XNOR U5110 ( .A(b[4009]), .B(n1012), .Z(n1013) );
  XNOR U5111 ( .A(b[400]), .B(n1015), .Z(c[400]) );
  XNOR U5112 ( .A(b[4009]), .B(n1014), .Z(c[4009]) );
  XOR U5113 ( .A(n1016), .B(n1017), .Z(n1012) );
  ANDN U5114 ( .B(n1018), .A(n1019), .Z(n1016) );
  XNOR U5115 ( .A(b[4008]), .B(n1017), .Z(n1018) );
  XNOR U5116 ( .A(b[4008]), .B(n1019), .Z(c[4008]) );
  XOR U5117 ( .A(n1020), .B(n1021), .Z(n1017) );
  ANDN U5118 ( .B(n1022), .A(n1023), .Z(n1020) );
  XNOR U5119 ( .A(b[4007]), .B(n1021), .Z(n1022) );
  XNOR U5120 ( .A(b[4007]), .B(n1023), .Z(c[4007]) );
  XOR U5121 ( .A(n1024), .B(n1025), .Z(n1021) );
  ANDN U5122 ( .B(n1026), .A(n1027), .Z(n1024) );
  XNOR U5123 ( .A(b[4006]), .B(n1025), .Z(n1026) );
  XNOR U5124 ( .A(b[4006]), .B(n1027), .Z(c[4006]) );
  XOR U5125 ( .A(n1028), .B(n1029), .Z(n1025) );
  ANDN U5126 ( .B(n1030), .A(n1031), .Z(n1028) );
  XNOR U5127 ( .A(b[4005]), .B(n1029), .Z(n1030) );
  XNOR U5128 ( .A(b[4005]), .B(n1031), .Z(c[4005]) );
  XOR U5129 ( .A(n1032), .B(n1033), .Z(n1029) );
  ANDN U5130 ( .B(n1034), .A(n1035), .Z(n1032) );
  XNOR U5131 ( .A(b[4004]), .B(n1033), .Z(n1034) );
  XNOR U5132 ( .A(b[4004]), .B(n1035), .Z(c[4004]) );
  XOR U5133 ( .A(n1036), .B(n1037), .Z(n1033) );
  ANDN U5134 ( .B(n1038), .A(n1039), .Z(n1036) );
  XNOR U5135 ( .A(b[4003]), .B(n1037), .Z(n1038) );
  XNOR U5136 ( .A(b[4003]), .B(n1039), .Z(c[4003]) );
  XOR U5137 ( .A(n1040), .B(n1041), .Z(n1037) );
  ANDN U5138 ( .B(n1042), .A(n1043), .Z(n1040) );
  XNOR U5139 ( .A(b[4002]), .B(n1041), .Z(n1042) );
  XNOR U5140 ( .A(b[4002]), .B(n1043), .Z(c[4002]) );
  XOR U5141 ( .A(n1044), .B(n1045), .Z(n1041) );
  ANDN U5142 ( .B(n1046), .A(n1047), .Z(n1044) );
  XNOR U5143 ( .A(b[4001]), .B(n1045), .Z(n1046) );
  XNOR U5144 ( .A(b[4001]), .B(n1047), .Z(c[4001]) );
  XOR U5145 ( .A(n1048), .B(n1049), .Z(n1045) );
  ANDN U5146 ( .B(n1050), .A(n1051), .Z(n1048) );
  XNOR U5147 ( .A(b[4000]), .B(n1049), .Z(n1050) );
  XNOR U5148 ( .A(b[4000]), .B(n1051), .Z(c[4000]) );
  XOR U5149 ( .A(n1052), .B(n1053), .Z(n1049) );
  ANDN U5150 ( .B(n1054), .A(n1055), .Z(n1052) );
  XNOR U5151 ( .A(b[3999]), .B(n1053), .Z(n1054) );
  XNOR U5152 ( .A(b[3]), .B(n1056), .Z(c[3]) );
  XNOR U5153 ( .A(b[39]), .B(n1057), .Z(c[39]) );
  XNOR U5154 ( .A(b[399]), .B(n1058), .Z(c[399]) );
  XNOR U5155 ( .A(b[3999]), .B(n1055), .Z(c[3999]) );
  XOR U5156 ( .A(n1059), .B(n1060), .Z(n1053) );
  ANDN U5157 ( .B(n1061), .A(n1062), .Z(n1059) );
  XNOR U5158 ( .A(b[3998]), .B(n1060), .Z(n1061) );
  XNOR U5159 ( .A(b[3998]), .B(n1062), .Z(c[3998]) );
  XOR U5160 ( .A(n1063), .B(n1064), .Z(n1060) );
  ANDN U5161 ( .B(n1065), .A(n1066), .Z(n1063) );
  XNOR U5162 ( .A(b[3997]), .B(n1064), .Z(n1065) );
  XNOR U5163 ( .A(b[3997]), .B(n1066), .Z(c[3997]) );
  XOR U5164 ( .A(n1067), .B(n1068), .Z(n1064) );
  ANDN U5165 ( .B(n1069), .A(n1070), .Z(n1067) );
  XNOR U5166 ( .A(b[3996]), .B(n1068), .Z(n1069) );
  XNOR U5167 ( .A(b[3996]), .B(n1070), .Z(c[3996]) );
  XOR U5168 ( .A(n1071), .B(n1072), .Z(n1068) );
  ANDN U5169 ( .B(n1073), .A(n1074), .Z(n1071) );
  XNOR U5170 ( .A(b[3995]), .B(n1072), .Z(n1073) );
  XNOR U5171 ( .A(b[3995]), .B(n1074), .Z(c[3995]) );
  XOR U5172 ( .A(n1075), .B(n1076), .Z(n1072) );
  ANDN U5173 ( .B(n1077), .A(n1078), .Z(n1075) );
  XNOR U5174 ( .A(b[3994]), .B(n1076), .Z(n1077) );
  XNOR U5175 ( .A(b[3994]), .B(n1078), .Z(c[3994]) );
  XOR U5176 ( .A(n1079), .B(n1080), .Z(n1076) );
  ANDN U5177 ( .B(n1081), .A(n1082), .Z(n1079) );
  XNOR U5178 ( .A(b[3993]), .B(n1080), .Z(n1081) );
  XNOR U5179 ( .A(b[3993]), .B(n1082), .Z(c[3993]) );
  XOR U5180 ( .A(n1083), .B(n1084), .Z(n1080) );
  ANDN U5181 ( .B(n1085), .A(n1086), .Z(n1083) );
  XNOR U5182 ( .A(b[3992]), .B(n1084), .Z(n1085) );
  XNOR U5183 ( .A(b[3992]), .B(n1086), .Z(c[3992]) );
  XOR U5184 ( .A(n1087), .B(n1088), .Z(n1084) );
  ANDN U5185 ( .B(n1089), .A(n1090), .Z(n1087) );
  XNOR U5186 ( .A(b[3991]), .B(n1088), .Z(n1089) );
  XNOR U5187 ( .A(b[3991]), .B(n1090), .Z(c[3991]) );
  XOR U5188 ( .A(n1091), .B(n1092), .Z(n1088) );
  ANDN U5189 ( .B(n1093), .A(n1094), .Z(n1091) );
  XNOR U5190 ( .A(b[3990]), .B(n1092), .Z(n1093) );
  XNOR U5191 ( .A(b[3990]), .B(n1094), .Z(c[3990]) );
  XOR U5192 ( .A(n1095), .B(n1096), .Z(n1092) );
  ANDN U5193 ( .B(n1097), .A(n1098), .Z(n1095) );
  XNOR U5194 ( .A(b[3989]), .B(n1096), .Z(n1097) );
  XNOR U5195 ( .A(b[398]), .B(n1099), .Z(c[398]) );
  XNOR U5196 ( .A(b[3989]), .B(n1098), .Z(c[3989]) );
  XOR U5197 ( .A(n1100), .B(n1101), .Z(n1096) );
  ANDN U5198 ( .B(n1102), .A(n1103), .Z(n1100) );
  XNOR U5199 ( .A(b[3988]), .B(n1101), .Z(n1102) );
  XNOR U5200 ( .A(b[3988]), .B(n1103), .Z(c[3988]) );
  XOR U5201 ( .A(n1104), .B(n1105), .Z(n1101) );
  ANDN U5202 ( .B(n1106), .A(n1107), .Z(n1104) );
  XNOR U5203 ( .A(b[3987]), .B(n1105), .Z(n1106) );
  XNOR U5204 ( .A(b[3987]), .B(n1107), .Z(c[3987]) );
  XOR U5205 ( .A(n1108), .B(n1109), .Z(n1105) );
  ANDN U5206 ( .B(n1110), .A(n1111), .Z(n1108) );
  XNOR U5207 ( .A(b[3986]), .B(n1109), .Z(n1110) );
  XNOR U5208 ( .A(b[3986]), .B(n1111), .Z(c[3986]) );
  XOR U5209 ( .A(n1112), .B(n1113), .Z(n1109) );
  ANDN U5210 ( .B(n1114), .A(n1115), .Z(n1112) );
  XNOR U5211 ( .A(b[3985]), .B(n1113), .Z(n1114) );
  XNOR U5212 ( .A(b[3985]), .B(n1115), .Z(c[3985]) );
  XOR U5213 ( .A(n1116), .B(n1117), .Z(n1113) );
  ANDN U5214 ( .B(n1118), .A(n1119), .Z(n1116) );
  XNOR U5215 ( .A(b[3984]), .B(n1117), .Z(n1118) );
  XNOR U5216 ( .A(b[3984]), .B(n1119), .Z(c[3984]) );
  XOR U5217 ( .A(n1120), .B(n1121), .Z(n1117) );
  ANDN U5218 ( .B(n1122), .A(n1123), .Z(n1120) );
  XNOR U5219 ( .A(b[3983]), .B(n1121), .Z(n1122) );
  XNOR U5220 ( .A(b[3983]), .B(n1123), .Z(c[3983]) );
  XOR U5221 ( .A(n1124), .B(n1125), .Z(n1121) );
  ANDN U5222 ( .B(n1126), .A(n1127), .Z(n1124) );
  XNOR U5223 ( .A(b[3982]), .B(n1125), .Z(n1126) );
  XNOR U5224 ( .A(b[3982]), .B(n1127), .Z(c[3982]) );
  XOR U5225 ( .A(n1128), .B(n1129), .Z(n1125) );
  ANDN U5226 ( .B(n1130), .A(n1131), .Z(n1128) );
  XNOR U5227 ( .A(b[3981]), .B(n1129), .Z(n1130) );
  XNOR U5228 ( .A(b[3981]), .B(n1131), .Z(c[3981]) );
  XOR U5229 ( .A(n1132), .B(n1133), .Z(n1129) );
  ANDN U5230 ( .B(n1134), .A(n1135), .Z(n1132) );
  XNOR U5231 ( .A(b[3980]), .B(n1133), .Z(n1134) );
  XNOR U5232 ( .A(b[3980]), .B(n1135), .Z(c[3980]) );
  XOR U5233 ( .A(n1136), .B(n1137), .Z(n1133) );
  ANDN U5234 ( .B(n1138), .A(n1139), .Z(n1136) );
  XNOR U5235 ( .A(b[3979]), .B(n1137), .Z(n1138) );
  XNOR U5236 ( .A(b[397]), .B(n1140), .Z(c[397]) );
  XNOR U5237 ( .A(b[3979]), .B(n1139), .Z(c[3979]) );
  XOR U5238 ( .A(n1141), .B(n1142), .Z(n1137) );
  ANDN U5239 ( .B(n1143), .A(n1144), .Z(n1141) );
  XNOR U5240 ( .A(b[3978]), .B(n1142), .Z(n1143) );
  XNOR U5241 ( .A(b[3978]), .B(n1144), .Z(c[3978]) );
  XOR U5242 ( .A(n1145), .B(n1146), .Z(n1142) );
  ANDN U5243 ( .B(n1147), .A(n1148), .Z(n1145) );
  XNOR U5244 ( .A(b[3977]), .B(n1146), .Z(n1147) );
  XNOR U5245 ( .A(b[3977]), .B(n1148), .Z(c[3977]) );
  XOR U5246 ( .A(n1149), .B(n1150), .Z(n1146) );
  ANDN U5247 ( .B(n1151), .A(n1152), .Z(n1149) );
  XNOR U5248 ( .A(b[3976]), .B(n1150), .Z(n1151) );
  XNOR U5249 ( .A(b[3976]), .B(n1152), .Z(c[3976]) );
  XOR U5250 ( .A(n1153), .B(n1154), .Z(n1150) );
  ANDN U5251 ( .B(n1155), .A(n1156), .Z(n1153) );
  XNOR U5252 ( .A(b[3975]), .B(n1154), .Z(n1155) );
  XNOR U5253 ( .A(b[3975]), .B(n1156), .Z(c[3975]) );
  XOR U5254 ( .A(n1157), .B(n1158), .Z(n1154) );
  ANDN U5255 ( .B(n1159), .A(n1160), .Z(n1157) );
  XNOR U5256 ( .A(b[3974]), .B(n1158), .Z(n1159) );
  XNOR U5257 ( .A(b[3974]), .B(n1160), .Z(c[3974]) );
  XOR U5258 ( .A(n1161), .B(n1162), .Z(n1158) );
  ANDN U5259 ( .B(n1163), .A(n1164), .Z(n1161) );
  XNOR U5260 ( .A(b[3973]), .B(n1162), .Z(n1163) );
  XNOR U5261 ( .A(b[3973]), .B(n1164), .Z(c[3973]) );
  XOR U5262 ( .A(n1165), .B(n1166), .Z(n1162) );
  ANDN U5263 ( .B(n1167), .A(n1168), .Z(n1165) );
  XNOR U5264 ( .A(b[3972]), .B(n1166), .Z(n1167) );
  XNOR U5265 ( .A(b[3972]), .B(n1168), .Z(c[3972]) );
  XOR U5266 ( .A(n1169), .B(n1170), .Z(n1166) );
  ANDN U5267 ( .B(n1171), .A(n1172), .Z(n1169) );
  XNOR U5268 ( .A(b[3971]), .B(n1170), .Z(n1171) );
  XNOR U5269 ( .A(b[3971]), .B(n1172), .Z(c[3971]) );
  XOR U5270 ( .A(n1173), .B(n1174), .Z(n1170) );
  ANDN U5271 ( .B(n1175), .A(n1176), .Z(n1173) );
  XNOR U5272 ( .A(b[3970]), .B(n1174), .Z(n1175) );
  XNOR U5273 ( .A(b[3970]), .B(n1176), .Z(c[3970]) );
  XOR U5274 ( .A(n1177), .B(n1178), .Z(n1174) );
  ANDN U5275 ( .B(n1179), .A(n1180), .Z(n1177) );
  XNOR U5276 ( .A(b[3969]), .B(n1178), .Z(n1179) );
  XNOR U5277 ( .A(b[396]), .B(n1181), .Z(c[396]) );
  XNOR U5278 ( .A(b[3969]), .B(n1180), .Z(c[3969]) );
  XOR U5279 ( .A(n1182), .B(n1183), .Z(n1178) );
  ANDN U5280 ( .B(n1184), .A(n1185), .Z(n1182) );
  XNOR U5281 ( .A(b[3968]), .B(n1183), .Z(n1184) );
  XNOR U5282 ( .A(b[3968]), .B(n1185), .Z(c[3968]) );
  XOR U5283 ( .A(n1186), .B(n1187), .Z(n1183) );
  ANDN U5284 ( .B(n1188), .A(n1189), .Z(n1186) );
  XNOR U5285 ( .A(b[3967]), .B(n1187), .Z(n1188) );
  XNOR U5286 ( .A(b[3967]), .B(n1189), .Z(c[3967]) );
  XOR U5287 ( .A(n1190), .B(n1191), .Z(n1187) );
  ANDN U5288 ( .B(n1192), .A(n1193), .Z(n1190) );
  XNOR U5289 ( .A(b[3966]), .B(n1191), .Z(n1192) );
  XNOR U5290 ( .A(b[3966]), .B(n1193), .Z(c[3966]) );
  XOR U5291 ( .A(n1194), .B(n1195), .Z(n1191) );
  ANDN U5292 ( .B(n1196), .A(n1197), .Z(n1194) );
  XNOR U5293 ( .A(b[3965]), .B(n1195), .Z(n1196) );
  XNOR U5294 ( .A(b[3965]), .B(n1197), .Z(c[3965]) );
  XOR U5295 ( .A(n1198), .B(n1199), .Z(n1195) );
  ANDN U5296 ( .B(n1200), .A(n1201), .Z(n1198) );
  XNOR U5297 ( .A(b[3964]), .B(n1199), .Z(n1200) );
  XNOR U5298 ( .A(b[3964]), .B(n1201), .Z(c[3964]) );
  XOR U5299 ( .A(n1202), .B(n1203), .Z(n1199) );
  ANDN U5300 ( .B(n1204), .A(n1205), .Z(n1202) );
  XNOR U5301 ( .A(b[3963]), .B(n1203), .Z(n1204) );
  XNOR U5302 ( .A(b[3963]), .B(n1205), .Z(c[3963]) );
  XOR U5303 ( .A(n1206), .B(n1207), .Z(n1203) );
  ANDN U5304 ( .B(n1208), .A(n1209), .Z(n1206) );
  XNOR U5305 ( .A(b[3962]), .B(n1207), .Z(n1208) );
  XNOR U5306 ( .A(b[3962]), .B(n1209), .Z(c[3962]) );
  XOR U5307 ( .A(n1210), .B(n1211), .Z(n1207) );
  ANDN U5308 ( .B(n1212), .A(n1213), .Z(n1210) );
  XNOR U5309 ( .A(b[3961]), .B(n1211), .Z(n1212) );
  XNOR U5310 ( .A(b[3961]), .B(n1213), .Z(c[3961]) );
  XOR U5311 ( .A(n1214), .B(n1215), .Z(n1211) );
  ANDN U5312 ( .B(n1216), .A(n1217), .Z(n1214) );
  XNOR U5313 ( .A(b[3960]), .B(n1215), .Z(n1216) );
  XNOR U5314 ( .A(b[3960]), .B(n1217), .Z(c[3960]) );
  XOR U5315 ( .A(n1218), .B(n1219), .Z(n1215) );
  ANDN U5316 ( .B(n1220), .A(n1221), .Z(n1218) );
  XNOR U5317 ( .A(b[3959]), .B(n1219), .Z(n1220) );
  XNOR U5318 ( .A(b[395]), .B(n1222), .Z(c[395]) );
  XNOR U5319 ( .A(b[3959]), .B(n1221), .Z(c[3959]) );
  XOR U5320 ( .A(n1223), .B(n1224), .Z(n1219) );
  ANDN U5321 ( .B(n1225), .A(n1226), .Z(n1223) );
  XNOR U5322 ( .A(b[3958]), .B(n1224), .Z(n1225) );
  XNOR U5323 ( .A(b[3958]), .B(n1226), .Z(c[3958]) );
  XOR U5324 ( .A(n1227), .B(n1228), .Z(n1224) );
  ANDN U5325 ( .B(n1229), .A(n1230), .Z(n1227) );
  XNOR U5326 ( .A(b[3957]), .B(n1228), .Z(n1229) );
  XNOR U5327 ( .A(b[3957]), .B(n1230), .Z(c[3957]) );
  XOR U5328 ( .A(n1231), .B(n1232), .Z(n1228) );
  ANDN U5329 ( .B(n1233), .A(n1234), .Z(n1231) );
  XNOR U5330 ( .A(b[3956]), .B(n1232), .Z(n1233) );
  XNOR U5331 ( .A(b[3956]), .B(n1234), .Z(c[3956]) );
  XOR U5332 ( .A(n1235), .B(n1236), .Z(n1232) );
  ANDN U5333 ( .B(n1237), .A(n1238), .Z(n1235) );
  XNOR U5334 ( .A(b[3955]), .B(n1236), .Z(n1237) );
  XNOR U5335 ( .A(b[3955]), .B(n1238), .Z(c[3955]) );
  XOR U5336 ( .A(n1239), .B(n1240), .Z(n1236) );
  ANDN U5337 ( .B(n1241), .A(n1242), .Z(n1239) );
  XNOR U5338 ( .A(b[3954]), .B(n1240), .Z(n1241) );
  XNOR U5339 ( .A(b[3954]), .B(n1242), .Z(c[3954]) );
  XOR U5340 ( .A(n1243), .B(n1244), .Z(n1240) );
  ANDN U5341 ( .B(n1245), .A(n1246), .Z(n1243) );
  XNOR U5342 ( .A(b[3953]), .B(n1244), .Z(n1245) );
  XNOR U5343 ( .A(b[3953]), .B(n1246), .Z(c[3953]) );
  XOR U5344 ( .A(n1247), .B(n1248), .Z(n1244) );
  ANDN U5345 ( .B(n1249), .A(n1250), .Z(n1247) );
  XNOR U5346 ( .A(b[3952]), .B(n1248), .Z(n1249) );
  XNOR U5347 ( .A(b[3952]), .B(n1250), .Z(c[3952]) );
  XOR U5348 ( .A(n1251), .B(n1252), .Z(n1248) );
  ANDN U5349 ( .B(n1253), .A(n1254), .Z(n1251) );
  XNOR U5350 ( .A(b[3951]), .B(n1252), .Z(n1253) );
  XNOR U5351 ( .A(b[3951]), .B(n1254), .Z(c[3951]) );
  XOR U5352 ( .A(n1255), .B(n1256), .Z(n1252) );
  ANDN U5353 ( .B(n1257), .A(n1258), .Z(n1255) );
  XNOR U5354 ( .A(b[3950]), .B(n1256), .Z(n1257) );
  XNOR U5355 ( .A(b[3950]), .B(n1258), .Z(c[3950]) );
  XOR U5356 ( .A(n1259), .B(n1260), .Z(n1256) );
  ANDN U5357 ( .B(n1261), .A(n1262), .Z(n1259) );
  XNOR U5358 ( .A(b[3949]), .B(n1260), .Z(n1261) );
  XNOR U5359 ( .A(b[394]), .B(n1263), .Z(c[394]) );
  XNOR U5360 ( .A(b[3949]), .B(n1262), .Z(c[3949]) );
  XOR U5361 ( .A(n1264), .B(n1265), .Z(n1260) );
  ANDN U5362 ( .B(n1266), .A(n1267), .Z(n1264) );
  XNOR U5363 ( .A(b[3948]), .B(n1265), .Z(n1266) );
  XNOR U5364 ( .A(b[3948]), .B(n1267), .Z(c[3948]) );
  XOR U5365 ( .A(n1268), .B(n1269), .Z(n1265) );
  ANDN U5366 ( .B(n1270), .A(n1271), .Z(n1268) );
  XNOR U5367 ( .A(b[3947]), .B(n1269), .Z(n1270) );
  XNOR U5368 ( .A(b[3947]), .B(n1271), .Z(c[3947]) );
  XOR U5369 ( .A(n1272), .B(n1273), .Z(n1269) );
  ANDN U5370 ( .B(n1274), .A(n1275), .Z(n1272) );
  XNOR U5371 ( .A(b[3946]), .B(n1273), .Z(n1274) );
  XNOR U5372 ( .A(b[3946]), .B(n1275), .Z(c[3946]) );
  XOR U5373 ( .A(n1276), .B(n1277), .Z(n1273) );
  ANDN U5374 ( .B(n1278), .A(n1279), .Z(n1276) );
  XNOR U5375 ( .A(b[3945]), .B(n1277), .Z(n1278) );
  XNOR U5376 ( .A(b[3945]), .B(n1279), .Z(c[3945]) );
  XOR U5377 ( .A(n1280), .B(n1281), .Z(n1277) );
  ANDN U5378 ( .B(n1282), .A(n1283), .Z(n1280) );
  XNOR U5379 ( .A(b[3944]), .B(n1281), .Z(n1282) );
  XNOR U5380 ( .A(b[3944]), .B(n1283), .Z(c[3944]) );
  XOR U5381 ( .A(n1284), .B(n1285), .Z(n1281) );
  ANDN U5382 ( .B(n1286), .A(n1287), .Z(n1284) );
  XNOR U5383 ( .A(b[3943]), .B(n1285), .Z(n1286) );
  XNOR U5384 ( .A(b[3943]), .B(n1287), .Z(c[3943]) );
  XOR U5385 ( .A(n1288), .B(n1289), .Z(n1285) );
  ANDN U5386 ( .B(n1290), .A(n1291), .Z(n1288) );
  XNOR U5387 ( .A(b[3942]), .B(n1289), .Z(n1290) );
  XNOR U5388 ( .A(b[3942]), .B(n1291), .Z(c[3942]) );
  XOR U5389 ( .A(n1292), .B(n1293), .Z(n1289) );
  ANDN U5390 ( .B(n1294), .A(n1295), .Z(n1292) );
  XNOR U5391 ( .A(b[3941]), .B(n1293), .Z(n1294) );
  XNOR U5392 ( .A(b[3941]), .B(n1295), .Z(c[3941]) );
  XOR U5393 ( .A(n1296), .B(n1297), .Z(n1293) );
  ANDN U5394 ( .B(n1298), .A(n1299), .Z(n1296) );
  XNOR U5395 ( .A(b[3940]), .B(n1297), .Z(n1298) );
  XNOR U5396 ( .A(b[3940]), .B(n1299), .Z(c[3940]) );
  XOR U5397 ( .A(n1300), .B(n1301), .Z(n1297) );
  ANDN U5398 ( .B(n1302), .A(n1303), .Z(n1300) );
  XNOR U5399 ( .A(b[3939]), .B(n1301), .Z(n1302) );
  XNOR U5400 ( .A(b[393]), .B(n1304), .Z(c[393]) );
  XNOR U5401 ( .A(b[3939]), .B(n1303), .Z(c[3939]) );
  XOR U5402 ( .A(n1305), .B(n1306), .Z(n1301) );
  ANDN U5403 ( .B(n1307), .A(n1308), .Z(n1305) );
  XNOR U5404 ( .A(b[3938]), .B(n1306), .Z(n1307) );
  XNOR U5405 ( .A(b[3938]), .B(n1308), .Z(c[3938]) );
  XOR U5406 ( .A(n1309), .B(n1310), .Z(n1306) );
  ANDN U5407 ( .B(n1311), .A(n1312), .Z(n1309) );
  XNOR U5408 ( .A(b[3937]), .B(n1310), .Z(n1311) );
  XNOR U5409 ( .A(b[3937]), .B(n1312), .Z(c[3937]) );
  XOR U5410 ( .A(n1313), .B(n1314), .Z(n1310) );
  ANDN U5411 ( .B(n1315), .A(n1316), .Z(n1313) );
  XNOR U5412 ( .A(b[3936]), .B(n1314), .Z(n1315) );
  XNOR U5413 ( .A(b[3936]), .B(n1316), .Z(c[3936]) );
  XOR U5414 ( .A(n1317), .B(n1318), .Z(n1314) );
  ANDN U5415 ( .B(n1319), .A(n1320), .Z(n1317) );
  XNOR U5416 ( .A(b[3935]), .B(n1318), .Z(n1319) );
  XNOR U5417 ( .A(b[3935]), .B(n1320), .Z(c[3935]) );
  XOR U5418 ( .A(n1321), .B(n1322), .Z(n1318) );
  ANDN U5419 ( .B(n1323), .A(n1324), .Z(n1321) );
  XNOR U5420 ( .A(b[3934]), .B(n1322), .Z(n1323) );
  XNOR U5421 ( .A(b[3934]), .B(n1324), .Z(c[3934]) );
  XOR U5422 ( .A(n1325), .B(n1326), .Z(n1322) );
  ANDN U5423 ( .B(n1327), .A(n1328), .Z(n1325) );
  XNOR U5424 ( .A(b[3933]), .B(n1326), .Z(n1327) );
  XNOR U5425 ( .A(b[3933]), .B(n1328), .Z(c[3933]) );
  XOR U5426 ( .A(n1329), .B(n1330), .Z(n1326) );
  ANDN U5427 ( .B(n1331), .A(n1332), .Z(n1329) );
  XNOR U5428 ( .A(b[3932]), .B(n1330), .Z(n1331) );
  XNOR U5429 ( .A(b[3932]), .B(n1332), .Z(c[3932]) );
  XOR U5430 ( .A(n1333), .B(n1334), .Z(n1330) );
  ANDN U5431 ( .B(n1335), .A(n1336), .Z(n1333) );
  XNOR U5432 ( .A(b[3931]), .B(n1334), .Z(n1335) );
  XNOR U5433 ( .A(b[3931]), .B(n1336), .Z(c[3931]) );
  XOR U5434 ( .A(n1337), .B(n1338), .Z(n1334) );
  ANDN U5435 ( .B(n1339), .A(n1340), .Z(n1337) );
  XNOR U5436 ( .A(b[3930]), .B(n1338), .Z(n1339) );
  XNOR U5437 ( .A(b[3930]), .B(n1340), .Z(c[3930]) );
  XOR U5438 ( .A(n1341), .B(n1342), .Z(n1338) );
  ANDN U5439 ( .B(n1343), .A(n1344), .Z(n1341) );
  XNOR U5440 ( .A(b[3929]), .B(n1342), .Z(n1343) );
  XNOR U5441 ( .A(b[392]), .B(n1345), .Z(c[392]) );
  XNOR U5442 ( .A(b[3929]), .B(n1344), .Z(c[3929]) );
  XOR U5443 ( .A(n1346), .B(n1347), .Z(n1342) );
  ANDN U5444 ( .B(n1348), .A(n1349), .Z(n1346) );
  XNOR U5445 ( .A(b[3928]), .B(n1347), .Z(n1348) );
  XNOR U5446 ( .A(b[3928]), .B(n1349), .Z(c[3928]) );
  XOR U5447 ( .A(n1350), .B(n1351), .Z(n1347) );
  ANDN U5448 ( .B(n1352), .A(n1353), .Z(n1350) );
  XNOR U5449 ( .A(b[3927]), .B(n1351), .Z(n1352) );
  XNOR U5450 ( .A(b[3927]), .B(n1353), .Z(c[3927]) );
  XOR U5451 ( .A(n1354), .B(n1355), .Z(n1351) );
  ANDN U5452 ( .B(n1356), .A(n1357), .Z(n1354) );
  XNOR U5453 ( .A(b[3926]), .B(n1355), .Z(n1356) );
  XNOR U5454 ( .A(b[3926]), .B(n1357), .Z(c[3926]) );
  XOR U5455 ( .A(n1358), .B(n1359), .Z(n1355) );
  ANDN U5456 ( .B(n1360), .A(n1361), .Z(n1358) );
  XNOR U5457 ( .A(b[3925]), .B(n1359), .Z(n1360) );
  XNOR U5458 ( .A(b[3925]), .B(n1361), .Z(c[3925]) );
  XOR U5459 ( .A(n1362), .B(n1363), .Z(n1359) );
  ANDN U5460 ( .B(n1364), .A(n1365), .Z(n1362) );
  XNOR U5461 ( .A(b[3924]), .B(n1363), .Z(n1364) );
  XNOR U5462 ( .A(b[3924]), .B(n1365), .Z(c[3924]) );
  XOR U5463 ( .A(n1366), .B(n1367), .Z(n1363) );
  ANDN U5464 ( .B(n1368), .A(n1369), .Z(n1366) );
  XNOR U5465 ( .A(b[3923]), .B(n1367), .Z(n1368) );
  XNOR U5466 ( .A(b[3923]), .B(n1369), .Z(c[3923]) );
  XOR U5467 ( .A(n1370), .B(n1371), .Z(n1367) );
  ANDN U5468 ( .B(n1372), .A(n1373), .Z(n1370) );
  XNOR U5469 ( .A(b[3922]), .B(n1371), .Z(n1372) );
  XNOR U5470 ( .A(b[3922]), .B(n1373), .Z(c[3922]) );
  XOR U5471 ( .A(n1374), .B(n1375), .Z(n1371) );
  ANDN U5472 ( .B(n1376), .A(n1377), .Z(n1374) );
  XNOR U5473 ( .A(b[3921]), .B(n1375), .Z(n1376) );
  XNOR U5474 ( .A(b[3921]), .B(n1377), .Z(c[3921]) );
  XOR U5475 ( .A(n1378), .B(n1379), .Z(n1375) );
  ANDN U5476 ( .B(n1380), .A(n1381), .Z(n1378) );
  XNOR U5477 ( .A(b[3920]), .B(n1379), .Z(n1380) );
  XNOR U5478 ( .A(b[3920]), .B(n1381), .Z(c[3920]) );
  XOR U5479 ( .A(n1382), .B(n1383), .Z(n1379) );
  ANDN U5480 ( .B(n1384), .A(n1385), .Z(n1382) );
  XNOR U5481 ( .A(b[3919]), .B(n1383), .Z(n1384) );
  XNOR U5482 ( .A(b[391]), .B(n1386), .Z(c[391]) );
  XNOR U5483 ( .A(b[3919]), .B(n1385), .Z(c[3919]) );
  XOR U5484 ( .A(n1387), .B(n1388), .Z(n1383) );
  ANDN U5485 ( .B(n1389), .A(n1390), .Z(n1387) );
  XNOR U5486 ( .A(b[3918]), .B(n1388), .Z(n1389) );
  XNOR U5487 ( .A(b[3918]), .B(n1390), .Z(c[3918]) );
  XOR U5488 ( .A(n1391), .B(n1392), .Z(n1388) );
  ANDN U5489 ( .B(n1393), .A(n1394), .Z(n1391) );
  XNOR U5490 ( .A(b[3917]), .B(n1392), .Z(n1393) );
  XNOR U5491 ( .A(b[3917]), .B(n1394), .Z(c[3917]) );
  XOR U5492 ( .A(n1395), .B(n1396), .Z(n1392) );
  ANDN U5493 ( .B(n1397), .A(n1398), .Z(n1395) );
  XNOR U5494 ( .A(b[3916]), .B(n1396), .Z(n1397) );
  XNOR U5495 ( .A(b[3916]), .B(n1398), .Z(c[3916]) );
  XOR U5496 ( .A(n1399), .B(n1400), .Z(n1396) );
  ANDN U5497 ( .B(n1401), .A(n1402), .Z(n1399) );
  XNOR U5498 ( .A(b[3915]), .B(n1400), .Z(n1401) );
  XNOR U5499 ( .A(b[3915]), .B(n1402), .Z(c[3915]) );
  XOR U5500 ( .A(n1403), .B(n1404), .Z(n1400) );
  ANDN U5501 ( .B(n1405), .A(n1406), .Z(n1403) );
  XNOR U5502 ( .A(b[3914]), .B(n1404), .Z(n1405) );
  XNOR U5503 ( .A(b[3914]), .B(n1406), .Z(c[3914]) );
  XOR U5504 ( .A(n1407), .B(n1408), .Z(n1404) );
  ANDN U5505 ( .B(n1409), .A(n1410), .Z(n1407) );
  XNOR U5506 ( .A(b[3913]), .B(n1408), .Z(n1409) );
  XNOR U5507 ( .A(b[3913]), .B(n1410), .Z(c[3913]) );
  XOR U5508 ( .A(n1411), .B(n1412), .Z(n1408) );
  ANDN U5509 ( .B(n1413), .A(n1414), .Z(n1411) );
  XNOR U5510 ( .A(b[3912]), .B(n1412), .Z(n1413) );
  XNOR U5511 ( .A(b[3912]), .B(n1414), .Z(c[3912]) );
  XOR U5512 ( .A(n1415), .B(n1416), .Z(n1412) );
  ANDN U5513 ( .B(n1417), .A(n1418), .Z(n1415) );
  XNOR U5514 ( .A(b[3911]), .B(n1416), .Z(n1417) );
  XNOR U5515 ( .A(b[3911]), .B(n1418), .Z(c[3911]) );
  XOR U5516 ( .A(n1419), .B(n1420), .Z(n1416) );
  ANDN U5517 ( .B(n1421), .A(n1422), .Z(n1419) );
  XNOR U5518 ( .A(b[3910]), .B(n1420), .Z(n1421) );
  XNOR U5519 ( .A(b[3910]), .B(n1422), .Z(c[3910]) );
  XOR U5520 ( .A(n1423), .B(n1424), .Z(n1420) );
  ANDN U5521 ( .B(n1425), .A(n1426), .Z(n1423) );
  XNOR U5522 ( .A(b[3909]), .B(n1424), .Z(n1425) );
  XNOR U5523 ( .A(b[390]), .B(n1427), .Z(c[390]) );
  XNOR U5524 ( .A(b[3909]), .B(n1426), .Z(c[3909]) );
  XOR U5525 ( .A(n1428), .B(n1429), .Z(n1424) );
  ANDN U5526 ( .B(n1430), .A(n1431), .Z(n1428) );
  XNOR U5527 ( .A(b[3908]), .B(n1429), .Z(n1430) );
  XNOR U5528 ( .A(b[3908]), .B(n1431), .Z(c[3908]) );
  XOR U5529 ( .A(n1432), .B(n1433), .Z(n1429) );
  ANDN U5530 ( .B(n1434), .A(n1435), .Z(n1432) );
  XNOR U5531 ( .A(b[3907]), .B(n1433), .Z(n1434) );
  XNOR U5532 ( .A(b[3907]), .B(n1435), .Z(c[3907]) );
  XOR U5533 ( .A(n1436), .B(n1437), .Z(n1433) );
  ANDN U5534 ( .B(n1438), .A(n1439), .Z(n1436) );
  XNOR U5535 ( .A(b[3906]), .B(n1437), .Z(n1438) );
  XNOR U5536 ( .A(b[3906]), .B(n1439), .Z(c[3906]) );
  XOR U5537 ( .A(n1440), .B(n1441), .Z(n1437) );
  ANDN U5538 ( .B(n1442), .A(n1443), .Z(n1440) );
  XNOR U5539 ( .A(b[3905]), .B(n1441), .Z(n1442) );
  XNOR U5540 ( .A(b[3905]), .B(n1443), .Z(c[3905]) );
  XOR U5541 ( .A(n1444), .B(n1445), .Z(n1441) );
  ANDN U5542 ( .B(n1446), .A(n1447), .Z(n1444) );
  XNOR U5543 ( .A(b[3904]), .B(n1445), .Z(n1446) );
  XNOR U5544 ( .A(b[3904]), .B(n1447), .Z(c[3904]) );
  XOR U5545 ( .A(n1448), .B(n1449), .Z(n1445) );
  ANDN U5546 ( .B(n1450), .A(n1451), .Z(n1448) );
  XNOR U5547 ( .A(b[3903]), .B(n1449), .Z(n1450) );
  XNOR U5548 ( .A(b[3903]), .B(n1451), .Z(c[3903]) );
  XOR U5549 ( .A(n1452), .B(n1453), .Z(n1449) );
  ANDN U5550 ( .B(n1454), .A(n1455), .Z(n1452) );
  XNOR U5551 ( .A(b[3902]), .B(n1453), .Z(n1454) );
  XNOR U5552 ( .A(b[3902]), .B(n1455), .Z(c[3902]) );
  XOR U5553 ( .A(n1456), .B(n1457), .Z(n1453) );
  ANDN U5554 ( .B(n1458), .A(n1459), .Z(n1456) );
  XNOR U5555 ( .A(b[3901]), .B(n1457), .Z(n1458) );
  XNOR U5556 ( .A(b[3901]), .B(n1459), .Z(c[3901]) );
  XOR U5557 ( .A(n1460), .B(n1461), .Z(n1457) );
  ANDN U5558 ( .B(n1462), .A(n1463), .Z(n1460) );
  XNOR U5559 ( .A(b[3900]), .B(n1461), .Z(n1462) );
  XNOR U5560 ( .A(b[3900]), .B(n1463), .Z(c[3900]) );
  XOR U5561 ( .A(n1464), .B(n1465), .Z(n1461) );
  ANDN U5562 ( .B(n1466), .A(n1467), .Z(n1464) );
  XNOR U5563 ( .A(b[3899]), .B(n1465), .Z(n1466) );
  XNOR U5564 ( .A(b[38]), .B(n1468), .Z(c[38]) );
  XNOR U5565 ( .A(b[389]), .B(n1469), .Z(c[389]) );
  XNOR U5566 ( .A(b[3899]), .B(n1467), .Z(c[3899]) );
  XOR U5567 ( .A(n1470), .B(n1471), .Z(n1465) );
  ANDN U5568 ( .B(n1472), .A(n1473), .Z(n1470) );
  XNOR U5569 ( .A(b[3898]), .B(n1471), .Z(n1472) );
  XNOR U5570 ( .A(b[3898]), .B(n1473), .Z(c[3898]) );
  XOR U5571 ( .A(n1474), .B(n1475), .Z(n1471) );
  ANDN U5572 ( .B(n1476), .A(n1477), .Z(n1474) );
  XNOR U5573 ( .A(b[3897]), .B(n1475), .Z(n1476) );
  XNOR U5574 ( .A(b[3897]), .B(n1477), .Z(c[3897]) );
  XOR U5575 ( .A(n1478), .B(n1479), .Z(n1475) );
  ANDN U5576 ( .B(n1480), .A(n1481), .Z(n1478) );
  XNOR U5577 ( .A(b[3896]), .B(n1479), .Z(n1480) );
  XNOR U5578 ( .A(b[3896]), .B(n1481), .Z(c[3896]) );
  XOR U5579 ( .A(n1482), .B(n1483), .Z(n1479) );
  ANDN U5580 ( .B(n1484), .A(n1485), .Z(n1482) );
  XNOR U5581 ( .A(b[3895]), .B(n1483), .Z(n1484) );
  XNOR U5582 ( .A(b[3895]), .B(n1485), .Z(c[3895]) );
  XOR U5583 ( .A(n1486), .B(n1487), .Z(n1483) );
  ANDN U5584 ( .B(n1488), .A(n1489), .Z(n1486) );
  XNOR U5585 ( .A(b[3894]), .B(n1487), .Z(n1488) );
  XNOR U5586 ( .A(b[3894]), .B(n1489), .Z(c[3894]) );
  XOR U5587 ( .A(n1490), .B(n1491), .Z(n1487) );
  ANDN U5588 ( .B(n1492), .A(n1493), .Z(n1490) );
  XNOR U5589 ( .A(b[3893]), .B(n1491), .Z(n1492) );
  XNOR U5590 ( .A(b[3893]), .B(n1493), .Z(c[3893]) );
  XOR U5591 ( .A(n1494), .B(n1495), .Z(n1491) );
  ANDN U5592 ( .B(n1496), .A(n1497), .Z(n1494) );
  XNOR U5593 ( .A(b[3892]), .B(n1495), .Z(n1496) );
  XNOR U5594 ( .A(b[3892]), .B(n1497), .Z(c[3892]) );
  XOR U5595 ( .A(n1498), .B(n1499), .Z(n1495) );
  ANDN U5596 ( .B(n1500), .A(n1501), .Z(n1498) );
  XNOR U5597 ( .A(b[3891]), .B(n1499), .Z(n1500) );
  XNOR U5598 ( .A(b[3891]), .B(n1501), .Z(c[3891]) );
  XOR U5599 ( .A(n1502), .B(n1503), .Z(n1499) );
  ANDN U5600 ( .B(n1504), .A(n1505), .Z(n1502) );
  XNOR U5601 ( .A(b[3890]), .B(n1503), .Z(n1504) );
  XNOR U5602 ( .A(b[3890]), .B(n1505), .Z(c[3890]) );
  XOR U5603 ( .A(n1506), .B(n1507), .Z(n1503) );
  ANDN U5604 ( .B(n1508), .A(n1509), .Z(n1506) );
  XNOR U5605 ( .A(b[3889]), .B(n1507), .Z(n1508) );
  XNOR U5606 ( .A(b[388]), .B(n1510), .Z(c[388]) );
  XNOR U5607 ( .A(b[3889]), .B(n1509), .Z(c[3889]) );
  XOR U5608 ( .A(n1511), .B(n1512), .Z(n1507) );
  ANDN U5609 ( .B(n1513), .A(n1514), .Z(n1511) );
  XNOR U5610 ( .A(b[3888]), .B(n1512), .Z(n1513) );
  XNOR U5611 ( .A(b[3888]), .B(n1514), .Z(c[3888]) );
  XOR U5612 ( .A(n1515), .B(n1516), .Z(n1512) );
  ANDN U5613 ( .B(n1517), .A(n1518), .Z(n1515) );
  XNOR U5614 ( .A(b[3887]), .B(n1516), .Z(n1517) );
  XNOR U5615 ( .A(b[3887]), .B(n1518), .Z(c[3887]) );
  XOR U5616 ( .A(n1519), .B(n1520), .Z(n1516) );
  ANDN U5617 ( .B(n1521), .A(n1522), .Z(n1519) );
  XNOR U5618 ( .A(b[3886]), .B(n1520), .Z(n1521) );
  XNOR U5619 ( .A(b[3886]), .B(n1522), .Z(c[3886]) );
  XOR U5620 ( .A(n1523), .B(n1524), .Z(n1520) );
  ANDN U5621 ( .B(n1525), .A(n1526), .Z(n1523) );
  XNOR U5622 ( .A(b[3885]), .B(n1524), .Z(n1525) );
  XNOR U5623 ( .A(b[3885]), .B(n1526), .Z(c[3885]) );
  XOR U5624 ( .A(n1527), .B(n1528), .Z(n1524) );
  ANDN U5625 ( .B(n1529), .A(n1530), .Z(n1527) );
  XNOR U5626 ( .A(b[3884]), .B(n1528), .Z(n1529) );
  XNOR U5627 ( .A(b[3884]), .B(n1530), .Z(c[3884]) );
  XOR U5628 ( .A(n1531), .B(n1532), .Z(n1528) );
  ANDN U5629 ( .B(n1533), .A(n1534), .Z(n1531) );
  XNOR U5630 ( .A(b[3883]), .B(n1532), .Z(n1533) );
  XNOR U5631 ( .A(b[3883]), .B(n1534), .Z(c[3883]) );
  XOR U5632 ( .A(n1535), .B(n1536), .Z(n1532) );
  ANDN U5633 ( .B(n1537), .A(n1538), .Z(n1535) );
  XNOR U5634 ( .A(b[3882]), .B(n1536), .Z(n1537) );
  XNOR U5635 ( .A(b[3882]), .B(n1538), .Z(c[3882]) );
  XOR U5636 ( .A(n1539), .B(n1540), .Z(n1536) );
  ANDN U5637 ( .B(n1541), .A(n1542), .Z(n1539) );
  XNOR U5638 ( .A(b[3881]), .B(n1540), .Z(n1541) );
  XNOR U5639 ( .A(b[3881]), .B(n1542), .Z(c[3881]) );
  XOR U5640 ( .A(n1543), .B(n1544), .Z(n1540) );
  ANDN U5641 ( .B(n1545), .A(n1546), .Z(n1543) );
  XNOR U5642 ( .A(b[3880]), .B(n1544), .Z(n1545) );
  XNOR U5643 ( .A(b[3880]), .B(n1546), .Z(c[3880]) );
  XOR U5644 ( .A(n1547), .B(n1548), .Z(n1544) );
  ANDN U5645 ( .B(n1549), .A(n1550), .Z(n1547) );
  XNOR U5646 ( .A(b[3879]), .B(n1548), .Z(n1549) );
  XNOR U5647 ( .A(b[387]), .B(n1551), .Z(c[387]) );
  XNOR U5648 ( .A(b[3879]), .B(n1550), .Z(c[3879]) );
  XOR U5649 ( .A(n1552), .B(n1553), .Z(n1548) );
  ANDN U5650 ( .B(n1554), .A(n1555), .Z(n1552) );
  XNOR U5651 ( .A(b[3878]), .B(n1553), .Z(n1554) );
  XNOR U5652 ( .A(b[3878]), .B(n1555), .Z(c[3878]) );
  XOR U5653 ( .A(n1556), .B(n1557), .Z(n1553) );
  ANDN U5654 ( .B(n1558), .A(n1559), .Z(n1556) );
  XNOR U5655 ( .A(b[3877]), .B(n1557), .Z(n1558) );
  XNOR U5656 ( .A(b[3877]), .B(n1559), .Z(c[3877]) );
  XOR U5657 ( .A(n1560), .B(n1561), .Z(n1557) );
  ANDN U5658 ( .B(n1562), .A(n1563), .Z(n1560) );
  XNOR U5659 ( .A(b[3876]), .B(n1561), .Z(n1562) );
  XNOR U5660 ( .A(b[3876]), .B(n1563), .Z(c[3876]) );
  XOR U5661 ( .A(n1564), .B(n1565), .Z(n1561) );
  ANDN U5662 ( .B(n1566), .A(n1567), .Z(n1564) );
  XNOR U5663 ( .A(b[3875]), .B(n1565), .Z(n1566) );
  XNOR U5664 ( .A(b[3875]), .B(n1567), .Z(c[3875]) );
  XOR U5665 ( .A(n1568), .B(n1569), .Z(n1565) );
  ANDN U5666 ( .B(n1570), .A(n1571), .Z(n1568) );
  XNOR U5667 ( .A(b[3874]), .B(n1569), .Z(n1570) );
  XNOR U5668 ( .A(b[3874]), .B(n1571), .Z(c[3874]) );
  XOR U5669 ( .A(n1572), .B(n1573), .Z(n1569) );
  ANDN U5670 ( .B(n1574), .A(n1575), .Z(n1572) );
  XNOR U5671 ( .A(b[3873]), .B(n1573), .Z(n1574) );
  XNOR U5672 ( .A(b[3873]), .B(n1575), .Z(c[3873]) );
  XOR U5673 ( .A(n1576), .B(n1577), .Z(n1573) );
  ANDN U5674 ( .B(n1578), .A(n1579), .Z(n1576) );
  XNOR U5675 ( .A(b[3872]), .B(n1577), .Z(n1578) );
  XNOR U5676 ( .A(b[3872]), .B(n1579), .Z(c[3872]) );
  XOR U5677 ( .A(n1580), .B(n1581), .Z(n1577) );
  ANDN U5678 ( .B(n1582), .A(n1583), .Z(n1580) );
  XNOR U5679 ( .A(b[3871]), .B(n1581), .Z(n1582) );
  XNOR U5680 ( .A(b[3871]), .B(n1583), .Z(c[3871]) );
  XOR U5681 ( .A(n1584), .B(n1585), .Z(n1581) );
  ANDN U5682 ( .B(n1586), .A(n1587), .Z(n1584) );
  XNOR U5683 ( .A(b[3870]), .B(n1585), .Z(n1586) );
  XNOR U5684 ( .A(b[3870]), .B(n1587), .Z(c[3870]) );
  XOR U5685 ( .A(n1588), .B(n1589), .Z(n1585) );
  ANDN U5686 ( .B(n1590), .A(n1591), .Z(n1588) );
  XNOR U5687 ( .A(b[3869]), .B(n1589), .Z(n1590) );
  XNOR U5688 ( .A(b[386]), .B(n1592), .Z(c[386]) );
  XNOR U5689 ( .A(b[3869]), .B(n1591), .Z(c[3869]) );
  XOR U5690 ( .A(n1593), .B(n1594), .Z(n1589) );
  ANDN U5691 ( .B(n1595), .A(n1596), .Z(n1593) );
  XNOR U5692 ( .A(b[3868]), .B(n1594), .Z(n1595) );
  XNOR U5693 ( .A(b[3868]), .B(n1596), .Z(c[3868]) );
  XOR U5694 ( .A(n1597), .B(n1598), .Z(n1594) );
  ANDN U5695 ( .B(n1599), .A(n1600), .Z(n1597) );
  XNOR U5696 ( .A(b[3867]), .B(n1598), .Z(n1599) );
  XNOR U5697 ( .A(b[3867]), .B(n1600), .Z(c[3867]) );
  XOR U5698 ( .A(n1601), .B(n1602), .Z(n1598) );
  ANDN U5699 ( .B(n1603), .A(n1604), .Z(n1601) );
  XNOR U5700 ( .A(b[3866]), .B(n1602), .Z(n1603) );
  XNOR U5701 ( .A(b[3866]), .B(n1604), .Z(c[3866]) );
  XOR U5702 ( .A(n1605), .B(n1606), .Z(n1602) );
  ANDN U5703 ( .B(n1607), .A(n1608), .Z(n1605) );
  XNOR U5704 ( .A(b[3865]), .B(n1606), .Z(n1607) );
  XNOR U5705 ( .A(b[3865]), .B(n1608), .Z(c[3865]) );
  XOR U5706 ( .A(n1609), .B(n1610), .Z(n1606) );
  ANDN U5707 ( .B(n1611), .A(n1612), .Z(n1609) );
  XNOR U5708 ( .A(b[3864]), .B(n1610), .Z(n1611) );
  XNOR U5709 ( .A(b[3864]), .B(n1612), .Z(c[3864]) );
  XOR U5710 ( .A(n1613), .B(n1614), .Z(n1610) );
  ANDN U5711 ( .B(n1615), .A(n1616), .Z(n1613) );
  XNOR U5712 ( .A(b[3863]), .B(n1614), .Z(n1615) );
  XNOR U5713 ( .A(b[3863]), .B(n1616), .Z(c[3863]) );
  XOR U5714 ( .A(n1617), .B(n1618), .Z(n1614) );
  ANDN U5715 ( .B(n1619), .A(n1620), .Z(n1617) );
  XNOR U5716 ( .A(b[3862]), .B(n1618), .Z(n1619) );
  XNOR U5717 ( .A(b[3862]), .B(n1620), .Z(c[3862]) );
  XOR U5718 ( .A(n1621), .B(n1622), .Z(n1618) );
  ANDN U5719 ( .B(n1623), .A(n1624), .Z(n1621) );
  XNOR U5720 ( .A(b[3861]), .B(n1622), .Z(n1623) );
  XNOR U5721 ( .A(b[3861]), .B(n1624), .Z(c[3861]) );
  XOR U5722 ( .A(n1625), .B(n1626), .Z(n1622) );
  ANDN U5723 ( .B(n1627), .A(n1628), .Z(n1625) );
  XNOR U5724 ( .A(b[3860]), .B(n1626), .Z(n1627) );
  XNOR U5725 ( .A(b[3860]), .B(n1628), .Z(c[3860]) );
  XOR U5726 ( .A(n1629), .B(n1630), .Z(n1626) );
  ANDN U5727 ( .B(n1631), .A(n1632), .Z(n1629) );
  XNOR U5728 ( .A(b[3859]), .B(n1630), .Z(n1631) );
  XNOR U5729 ( .A(b[385]), .B(n1633), .Z(c[385]) );
  XNOR U5730 ( .A(b[3859]), .B(n1632), .Z(c[3859]) );
  XOR U5731 ( .A(n1634), .B(n1635), .Z(n1630) );
  ANDN U5732 ( .B(n1636), .A(n1637), .Z(n1634) );
  XNOR U5733 ( .A(b[3858]), .B(n1635), .Z(n1636) );
  XNOR U5734 ( .A(b[3858]), .B(n1637), .Z(c[3858]) );
  XOR U5735 ( .A(n1638), .B(n1639), .Z(n1635) );
  ANDN U5736 ( .B(n1640), .A(n1641), .Z(n1638) );
  XNOR U5737 ( .A(b[3857]), .B(n1639), .Z(n1640) );
  XNOR U5738 ( .A(b[3857]), .B(n1641), .Z(c[3857]) );
  XOR U5739 ( .A(n1642), .B(n1643), .Z(n1639) );
  ANDN U5740 ( .B(n1644), .A(n1645), .Z(n1642) );
  XNOR U5741 ( .A(b[3856]), .B(n1643), .Z(n1644) );
  XNOR U5742 ( .A(b[3856]), .B(n1645), .Z(c[3856]) );
  XOR U5743 ( .A(n1646), .B(n1647), .Z(n1643) );
  ANDN U5744 ( .B(n1648), .A(n1649), .Z(n1646) );
  XNOR U5745 ( .A(b[3855]), .B(n1647), .Z(n1648) );
  XNOR U5746 ( .A(b[3855]), .B(n1649), .Z(c[3855]) );
  XOR U5747 ( .A(n1650), .B(n1651), .Z(n1647) );
  ANDN U5748 ( .B(n1652), .A(n1653), .Z(n1650) );
  XNOR U5749 ( .A(b[3854]), .B(n1651), .Z(n1652) );
  XNOR U5750 ( .A(b[3854]), .B(n1653), .Z(c[3854]) );
  XOR U5751 ( .A(n1654), .B(n1655), .Z(n1651) );
  ANDN U5752 ( .B(n1656), .A(n1657), .Z(n1654) );
  XNOR U5753 ( .A(b[3853]), .B(n1655), .Z(n1656) );
  XNOR U5754 ( .A(b[3853]), .B(n1657), .Z(c[3853]) );
  XOR U5755 ( .A(n1658), .B(n1659), .Z(n1655) );
  ANDN U5756 ( .B(n1660), .A(n1661), .Z(n1658) );
  XNOR U5757 ( .A(b[3852]), .B(n1659), .Z(n1660) );
  XNOR U5758 ( .A(b[3852]), .B(n1661), .Z(c[3852]) );
  XOR U5759 ( .A(n1662), .B(n1663), .Z(n1659) );
  ANDN U5760 ( .B(n1664), .A(n1665), .Z(n1662) );
  XNOR U5761 ( .A(b[3851]), .B(n1663), .Z(n1664) );
  XNOR U5762 ( .A(b[3851]), .B(n1665), .Z(c[3851]) );
  XOR U5763 ( .A(n1666), .B(n1667), .Z(n1663) );
  ANDN U5764 ( .B(n1668), .A(n1669), .Z(n1666) );
  XNOR U5765 ( .A(b[3850]), .B(n1667), .Z(n1668) );
  XNOR U5766 ( .A(b[3850]), .B(n1669), .Z(c[3850]) );
  XOR U5767 ( .A(n1670), .B(n1671), .Z(n1667) );
  ANDN U5768 ( .B(n1672), .A(n1673), .Z(n1670) );
  XNOR U5769 ( .A(b[3849]), .B(n1671), .Z(n1672) );
  XNOR U5770 ( .A(b[384]), .B(n1674), .Z(c[384]) );
  XNOR U5771 ( .A(b[3849]), .B(n1673), .Z(c[3849]) );
  XOR U5772 ( .A(n1675), .B(n1676), .Z(n1671) );
  ANDN U5773 ( .B(n1677), .A(n1678), .Z(n1675) );
  XNOR U5774 ( .A(b[3848]), .B(n1676), .Z(n1677) );
  XNOR U5775 ( .A(b[3848]), .B(n1678), .Z(c[3848]) );
  XOR U5776 ( .A(n1679), .B(n1680), .Z(n1676) );
  ANDN U5777 ( .B(n1681), .A(n1682), .Z(n1679) );
  XNOR U5778 ( .A(b[3847]), .B(n1680), .Z(n1681) );
  XNOR U5779 ( .A(b[3847]), .B(n1682), .Z(c[3847]) );
  XOR U5780 ( .A(n1683), .B(n1684), .Z(n1680) );
  ANDN U5781 ( .B(n1685), .A(n1686), .Z(n1683) );
  XNOR U5782 ( .A(b[3846]), .B(n1684), .Z(n1685) );
  XNOR U5783 ( .A(b[3846]), .B(n1686), .Z(c[3846]) );
  XOR U5784 ( .A(n1687), .B(n1688), .Z(n1684) );
  ANDN U5785 ( .B(n1689), .A(n1690), .Z(n1687) );
  XNOR U5786 ( .A(b[3845]), .B(n1688), .Z(n1689) );
  XNOR U5787 ( .A(b[3845]), .B(n1690), .Z(c[3845]) );
  XOR U5788 ( .A(n1691), .B(n1692), .Z(n1688) );
  ANDN U5789 ( .B(n1693), .A(n1694), .Z(n1691) );
  XNOR U5790 ( .A(b[3844]), .B(n1692), .Z(n1693) );
  XNOR U5791 ( .A(b[3844]), .B(n1694), .Z(c[3844]) );
  XOR U5792 ( .A(n1695), .B(n1696), .Z(n1692) );
  ANDN U5793 ( .B(n1697), .A(n1698), .Z(n1695) );
  XNOR U5794 ( .A(b[3843]), .B(n1696), .Z(n1697) );
  XNOR U5795 ( .A(b[3843]), .B(n1698), .Z(c[3843]) );
  XOR U5796 ( .A(n1699), .B(n1700), .Z(n1696) );
  ANDN U5797 ( .B(n1701), .A(n1702), .Z(n1699) );
  XNOR U5798 ( .A(b[3842]), .B(n1700), .Z(n1701) );
  XNOR U5799 ( .A(b[3842]), .B(n1702), .Z(c[3842]) );
  XOR U5800 ( .A(n1703), .B(n1704), .Z(n1700) );
  ANDN U5801 ( .B(n1705), .A(n1706), .Z(n1703) );
  XNOR U5802 ( .A(b[3841]), .B(n1704), .Z(n1705) );
  XNOR U5803 ( .A(b[3841]), .B(n1706), .Z(c[3841]) );
  XOR U5804 ( .A(n1707), .B(n1708), .Z(n1704) );
  ANDN U5805 ( .B(n1709), .A(n1710), .Z(n1707) );
  XNOR U5806 ( .A(b[3840]), .B(n1708), .Z(n1709) );
  XNOR U5807 ( .A(b[3840]), .B(n1710), .Z(c[3840]) );
  XOR U5808 ( .A(n1711), .B(n1712), .Z(n1708) );
  ANDN U5809 ( .B(n1713), .A(n1714), .Z(n1711) );
  XNOR U5810 ( .A(b[3839]), .B(n1712), .Z(n1713) );
  XNOR U5811 ( .A(b[383]), .B(n1715), .Z(c[383]) );
  XNOR U5812 ( .A(b[3839]), .B(n1714), .Z(c[3839]) );
  XOR U5813 ( .A(n1716), .B(n1717), .Z(n1712) );
  ANDN U5814 ( .B(n1718), .A(n1719), .Z(n1716) );
  XNOR U5815 ( .A(b[3838]), .B(n1717), .Z(n1718) );
  XNOR U5816 ( .A(b[3838]), .B(n1719), .Z(c[3838]) );
  XOR U5817 ( .A(n1720), .B(n1721), .Z(n1717) );
  ANDN U5818 ( .B(n1722), .A(n1723), .Z(n1720) );
  XNOR U5819 ( .A(b[3837]), .B(n1721), .Z(n1722) );
  XNOR U5820 ( .A(b[3837]), .B(n1723), .Z(c[3837]) );
  XOR U5821 ( .A(n1724), .B(n1725), .Z(n1721) );
  ANDN U5822 ( .B(n1726), .A(n1727), .Z(n1724) );
  XNOR U5823 ( .A(b[3836]), .B(n1725), .Z(n1726) );
  XNOR U5824 ( .A(b[3836]), .B(n1727), .Z(c[3836]) );
  XOR U5825 ( .A(n1728), .B(n1729), .Z(n1725) );
  ANDN U5826 ( .B(n1730), .A(n1731), .Z(n1728) );
  XNOR U5827 ( .A(b[3835]), .B(n1729), .Z(n1730) );
  XNOR U5828 ( .A(b[3835]), .B(n1731), .Z(c[3835]) );
  XOR U5829 ( .A(n1732), .B(n1733), .Z(n1729) );
  ANDN U5830 ( .B(n1734), .A(n1735), .Z(n1732) );
  XNOR U5831 ( .A(b[3834]), .B(n1733), .Z(n1734) );
  XNOR U5832 ( .A(b[3834]), .B(n1735), .Z(c[3834]) );
  XOR U5833 ( .A(n1736), .B(n1737), .Z(n1733) );
  ANDN U5834 ( .B(n1738), .A(n1739), .Z(n1736) );
  XNOR U5835 ( .A(b[3833]), .B(n1737), .Z(n1738) );
  XNOR U5836 ( .A(b[3833]), .B(n1739), .Z(c[3833]) );
  XOR U5837 ( .A(n1740), .B(n1741), .Z(n1737) );
  ANDN U5838 ( .B(n1742), .A(n1743), .Z(n1740) );
  XNOR U5839 ( .A(b[3832]), .B(n1741), .Z(n1742) );
  XNOR U5840 ( .A(b[3832]), .B(n1743), .Z(c[3832]) );
  XOR U5841 ( .A(n1744), .B(n1745), .Z(n1741) );
  ANDN U5842 ( .B(n1746), .A(n1747), .Z(n1744) );
  XNOR U5843 ( .A(b[3831]), .B(n1745), .Z(n1746) );
  XNOR U5844 ( .A(b[3831]), .B(n1747), .Z(c[3831]) );
  XOR U5845 ( .A(n1748), .B(n1749), .Z(n1745) );
  ANDN U5846 ( .B(n1750), .A(n1751), .Z(n1748) );
  XNOR U5847 ( .A(b[3830]), .B(n1749), .Z(n1750) );
  XNOR U5848 ( .A(b[3830]), .B(n1751), .Z(c[3830]) );
  XOR U5849 ( .A(n1752), .B(n1753), .Z(n1749) );
  ANDN U5850 ( .B(n1754), .A(n1755), .Z(n1752) );
  XNOR U5851 ( .A(b[3829]), .B(n1753), .Z(n1754) );
  XNOR U5852 ( .A(b[382]), .B(n1756), .Z(c[382]) );
  XNOR U5853 ( .A(b[3829]), .B(n1755), .Z(c[3829]) );
  XOR U5854 ( .A(n1757), .B(n1758), .Z(n1753) );
  ANDN U5855 ( .B(n1759), .A(n1760), .Z(n1757) );
  XNOR U5856 ( .A(b[3828]), .B(n1758), .Z(n1759) );
  XNOR U5857 ( .A(b[3828]), .B(n1760), .Z(c[3828]) );
  XOR U5858 ( .A(n1761), .B(n1762), .Z(n1758) );
  ANDN U5859 ( .B(n1763), .A(n1764), .Z(n1761) );
  XNOR U5860 ( .A(b[3827]), .B(n1762), .Z(n1763) );
  XNOR U5861 ( .A(b[3827]), .B(n1764), .Z(c[3827]) );
  XOR U5862 ( .A(n1765), .B(n1766), .Z(n1762) );
  ANDN U5863 ( .B(n1767), .A(n1768), .Z(n1765) );
  XNOR U5864 ( .A(b[3826]), .B(n1766), .Z(n1767) );
  XNOR U5865 ( .A(b[3826]), .B(n1768), .Z(c[3826]) );
  XOR U5866 ( .A(n1769), .B(n1770), .Z(n1766) );
  ANDN U5867 ( .B(n1771), .A(n1772), .Z(n1769) );
  XNOR U5868 ( .A(b[3825]), .B(n1770), .Z(n1771) );
  XNOR U5869 ( .A(b[3825]), .B(n1772), .Z(c[3825]) );
  XOR U5870 ( .A(n1773), .B(n1774), .Z(n1770) );
  ANDN U5871 ( .B(n1775), .A(n1776), .Z(n1773) );
  XNOR U5872 ( .A(b[3824]), .B(n1774), .Z(n1775) );
  XNOR U5873 ( .A(b[3824]), .B(n1776), .Z(c[3824]) );
  XOR U5874 ( .A(n1777), .B(n1778), .Z(n1774) );
  ANDN U5875 ( .B(n1779), .A(n1780), .Z(n1777) );
  XNOR U5876 ( .A(b[3823]), .B(n1778), .Z(n1779) );
  XNOR U5877 ( .A(b[3823]), .B(n1780), .Z(c[3823]) );
  XOR U5878 ( .A(n1781), .B(n1782), .Z(n1778) );
  ANDN U5879 ( .B(n1783), .A(n1784), .Z(n1781) );
  XNOR U5880 ( .A(b[3822]), .B(n1782), .Z(n1783) );
  XNOR U5881 ( .A(b[3822]), .B(n1784), .Z(c[3822]) );
  XOR U5882 ( .A(n1785), .B(n1786), .Z(n1782) );
  ANDN U5883 ( .B(n1787), .A(n1788), .Z(n1785) );
  XNOR U5884 ( .A(b[3821]), .B(n1786), .Z(n1787) );
  XNOR U5885 ( .A(b[3821]), .B(n1788), .Z(c[3821]) );
  XOR U5886 ( .A(n1789), .B(n1790), .Z(n1786) );
  ANDN U5887 ( .B(n1791), .A(n1792), .Z(n1789) );
  XNOR U5888 ( .A(b[3820]), .B(n1790), .Z(n1791) );
  XNOR U5889 ( .A(b[3820]), .B(n1792), .Z(c[3820]) );
  XOR U5890 ( .A(n1793), .B(n1794), .Z(n1790) );
  ANDN U5891 ( .B(n1795), .A(n1796), .Z(n1793) );
  XNOR U5892 ( .A(b[3819]), .B(n1794), .Z(n1795) );
  XNOR U5893 ( .A(b[381]), .B(n1797), .Z(c[381]) );
  XNOR U5894 ( .A(b[3819]), .B(n1796), .Z(c[3819]) );
  XOR U5895 ( .A(n1798), .B(n1799), .Z(n1794) );
  ANDN U5896 ( .B(n1800), .A(n1801), .Z(n1798) );
  XNOR U5897 ( .A(b[3818]), .B(n1799), .Z(n1800) );
  XNOR U5898 ( .A(b[3818]), .B(n1801), .Z(c[3818]) );
  XOR U5899 ( .A(n1802), .B(n1803), .Z(n1799) );
  ANDN U5900 ( .B(n1804), .A(n1805), .Z(n1802) );
  XNOR U5901 ( .A(b[3817]), .B(n1803), .Z(n1804) );
  XNOR U5902 ( .A(b[3817]), .B(n1805), .Z(c[3817]) );
  XOR U5903 ( .A(n1806), .B(n1807), .Z(n1803) );
  ANDN U5904 ( .B(n1808), .A(n1809), .Z(n1806) );
  XNOR U5905 ( .A(b[3816]), .B(n1807), .Z(n1808) );
  XNOR U5906 ( .A(b[3816]), .B(n1809), .Z(c[3816]) );
  XOR U5907 ( .A(n1810), .B(n1811), .Z(n1807) );
  ANDN U5908 ( .B(n1812), .A(n1813), .Z(n1810) );
  XNOR U5909 ( .A(b[3815]), .B(n1811), .Z(n1812) );
  XNOR U5910 ( .A(b[3815]), .B(n1813), .Z(c[3815]) );
  XOR U5911 ( .A(n1814), .B(n1815), .Z(n1811) );
  ANDN U5912 ( .B(n1816), .A(n1817), .Z(n1814) );
  XNOR U5913 ( .A(b[3814]), .B(n1815), .Z(n1816) );
  XNOR U5914 ( .A(b[3814]), .B(n1817), .Z(c[3814]) );
  XOR U5915 ( .A(n1818), .B(n1819), .Z(n1815) );
  ANDN U5916 ( .B(n1820), .A(n1821), .Z(n1818) );
  XNOR U5917 ( .A(b[3813]), .B(n1819), .Z(n1820) );
  XNOR U5918 ( .A(b[3813]), .B(n1821), .Z(c[3813]) );
  XOR U5919 ( .A(n1822), .B(n1823), .Z(n1819) );
  ANDN U5920 ( .B(n1824), .A(n1825), .Z(n1822) );
  XNOR U5921 ( .A(b[3812]), .B(n1823), .Z(n1824) );
  XNOR U5922 ( .A(b[3812]), .B(n1825), .Z(c[3812]) );
  XOR U5923 ( .A(n1826), .B(n1827), .Z(n1823) );
  ANDN U5924 ( .B(n1828), .A(n1829), .Z(n1826) );
  XNOR U5925 ( .A(b[3811]), .B(n1827), .Z(n1828) );
  XNOR U5926 ( .A(b[3811]), .B(n1829), .Z(c[3811]) );
  XOR U5927 ( .A(n1830), .B(n1831), .Z(n1827) );
  ANDN U5928 ( .B(n1832), .A(n1833), .Z(n1830) );
  XNOR U5929 ( .A(b[3810]), .B(n1831), .Z(n1832) );
  XNOR U5930 ( .A(b[3810]), .B(n1833), .Z(c[3810]) );
  XOR U5931 ( .A(n1834), .B(n1835), .Z(n1831) );
  ANDN U5932 ( .B(n1836), .A(n1837), .Z(n1834) );
  XNOR U5933 ( .A(b[3809]), .B(n1835), .Z(n1836) );
  XNOR U5934 ( .A(b[380]), .B(n1838), .Z(c[380]) );
  XNOR U5935 ( .A(b[3809]), .B(n1837), .Z(c[3809]) );
  XOR U5936 ( .A(n1839), .B(n1840), .Z(n1835) );
  ANDN U5937 ( .B(n1841), .A(n1842), .Z(n1839) );
  XNOR U5938 ( .A(b[3808]), .B(n1840), .Z(n1841) );
  XNOR U5939 ( .A(b[3808]), .B(n1842), .Z(c[3808]) );
  XOR U5940 ( .A(n1843), .B(n1844), .Z(n1840) );
  ANDN U5941 ( .B(n1845), .A(n1846), .Z(n1843) );
  XNOR U5942 ( .A(b[3807]), .B(n1844), .Z(n1845) );
  XNOR U5943 ( .A(b[3807]), .B(n1846), .Z(c[3807]) );
  XOR U5944 ( .A(n1847), .B(n1848), .Z(n1844) );
  ANDN U5945 ( .B(n1849), .A(n1850), .Z(n1847) );
  XNOR U5946 ( .A(b[3806]), .B(n1848), .Z(n1849) );
  XNOR U5947 ( .A(b[3806]), .B(n1850), .Z(c[3806]) );
  XOR U5948 ( .A(n1851), .B(n1852), .Z(n1848) );
  ANDN U5949 ( .B(n1853), .A(n1854), .Z(n1851) );
  XNOR U5950 ( .A(b[3805]), .B(n1852), .Z(n1853) );
  XNOR U5951 ( .A(b[3805]), .B(n1854), .Z(c[3805]) );
  XOR U5952 ( .A(n1855), .B(n1856), .Z(n1852) );
  ANDN U5953 ( .B(n1857), .A(n1858), .Z(n1855) );
  XNOR U5954 ( .A(b[3804]), .B(n1856), .Z(n1857) );
  XNOR U5955 ( .A(b[3804]), .B(n1858), .Z(c[3804]) );
  XOR U5956 ( .A(n1859), .B(n1860), .Z(n1856) );
  ANDN U5957 ( .B(n1861), .A(n1862), .Z(n1859) );
  XNOR U5958 ( .A(b[3803]), .B(n1860), .Z(n1861) );
  XNOR U5959 ( .A(b[3803]), .B(n1862), .Z(c[3803]) );
  XOR U5960 ( .A(n1863), .B(n1864), .Z(n1860) );
  ANDN U5961 ( .B(n1865), .A(n1866), .Z(n1863) );
  XNOR U5962 ( .A(b[3802]), .B(n1864), .Z(n1865) );
  XNOR U5963 ( .A(b[3802]), .B(n1866), .Z(c[3802]) );
  XOR U5964 ( .A(n1867), .B(n1868), .Z(n1864) );
  ANDN U5965 ( .B(n1869), .A(n1870), .Z(n1867) );
  XNOR U5966 ( .A(b[3801]), .B(n1868), .Z(n1869) );
  XNOR U5967 ( .A(b[3801]), .B(n1870), .Z(c[3801]) );
  XOR U5968 ( .A(n1871), .B(n1872), .Z(n1868) );
  ANDN U5969 ( .B(n1873), .A(n1874), .Z(n1871) );
  XNOR U5970 ( .A(b[3800]), .B(n1872), .Z(n1873) );
  XNOR U5971 ( .A(b[3800]), .B(n1874), .Z(c[3800]) );
  XOR U5972 ( .A(n1875), .B(n1876), .Z(n1872) );
  ANDN U5973 ( .B(n1877), .A(n1878), .Z(n1875) );
  XNOR U5974 ( .A(b[3799]), .B(n1876), .Z(n1877) );
  XNOR U5975 ( .A(b[37]), .B(n1879), .Z(c[37]) );
  XNOR U5976 ( .A(b[379]), .B(n1880), .Z(c[379]) );
  XNOR U5977 ( .A(b[3799]), .B(n1878), .Z(c[3799]) );
  XOR U5978 ( .A(n1881), .B(n1882), .Z(n1876) );
  ANDN U5979 ( .B(n1883), .A(n1884), .Z(n1881) );
  XNOR U5980 ( .A(b[3798]), .B(n1882), .Z(n1883) );
  XNOR U5981 ( .A(b[3798]), .B(n1884), .Z(c[3798]) );
  XOR U5982 ( .A(n1885), .B(n1886), .Z(n1882) );
  ANDN U5983 ( .B(n1887), .A(n1888), .Z(n1885) );
  XNOR U5984 ( .A(b[3797]), .B(n1886), .Z(n1887) );
  XNOR U5985 ( .A(b[3797]), .B(n1888), .Z(c[3797]) );
  XOR U5986 ( .A(n1889), .B(n1890), .Z(n1886) );
  ANDN U5987 ( .B(n1891), .A(n1892), .Z(n1889) );
  XNOR U5988 ( .A(b[3796]), .B(n1890), .Z(n1891) );
  XNOR U5989 ( .A(b[3796]), .B(n1892), .Z(c[3796]) );
  XOR U5990 ( .A(n1893), .B(n1894), .Z(n1890) );
  ANDN U5991 ( .B(n1895), .A(n1896), .Z(n1893) );
  XNOR U5992 ( .A(b[3795]), .B(n1894), .Z(n1895) );
  XNOR U5993 ( .A(b[3795]), .B(n1896), .Z(c[3795]) );
  XOR U5994 ( .A(n1897), .B(n1898), .Z(n1894) );
  ANDN U5995 ( .B(n1899), .A(n1900), .Z(n1897) );
  XNOR U5996 ( .A(b[3794]), .B(n1898), .Z(n1899) );
  XNOR U5997 ( .A(b[3794]), .B(n1900), .Z(c[3794]) );
  XOR U5998 ( .A(n1901), .B(n1902), .Z(n1898) );
  ANDN U5999 ( .B(n1903), .A(n1904), .Z(n1901) );
  XNOR U6000 ( .A(b[3793]), .B(n1902), .Z(n1903) );
  XNOR U6001 ( .A(b[3793]), .B(n1904), .Z(c[3793]) );
  XOR U6002 ( .A(n1905), .B(n1906), .Z(n1902) );
  ANDN U6003 ( .B(n1907), .A(n1908), .Z(n1905) );
  XNOR U6004 ( .A(b[3792]), .B(n1906), .Z(n1907) );
  XNOR U6005 ( .A(b[3792]), .B(n1908), .Z(c[3792]) );
  XOR U6006 ( .A(n1909), .B(n1910), .Z(n1906) );
  ANDN U6007 ( .B(n1911), .A(n1912), .Z(n1909) );
  XNOR U6008 ( .A(b[3791]), .B(n1910), .Z(n1911) );
  XNOR U6009 ( .A(b[3791]), .B(n1912), .Z(c[3791]) );
  XOR U6010 ( .A(n1913), .B(n1914), .Z(n1910) );
  ANDN U6011 ( .B(n1915), .A(n1916), .Z(n1913) );
  XNOR U6012 ( .A(b[3790]), .B(n1914), .Z(n1915) );
  XNOR U6013 ( .A(b[3790]), .B(n1916), .Z(c[3790]) );
  XOR U6014 ( .A(n1917), .B(n1918), .Z(n1914) );
  ANDN U6015 ( .B(n1919), .A(n1920), .Z(n1917) );
  XNOR U6016 ( .A(b[3789]), .B(n1918), .Z(n1919) );
  XNOR U6017 ( .A(b[378]), .B(n1921), .Z(c[378]) );
  XNOR U6018 ( .A(b[3789]), .B(n1920), .Z(c[3789]) );
  XOR U6019 ( .A(n1922), .B(n1923), .Z(n1918) );
  ANDN U6020 ( .B(n1924), .A(n1925), .Z(n1922) );
  XNOR U6021 ( .A(b[3788]), .B(n1923), .Z(n1924) );
  XNOR U6022 ( .A(b[3788]), .B(n1925), .Z(c[3788]) );
  XOR U6023 ( .A(n1926), .B(n1927), .Z(n1923) );
  ANDN U6024 ( .B(n1928), .A(n1929), .Z(n1926) );
  XNOR U6025 ( .A(b[3787]), .B(n1927), .Z(n1928) );
  XNOR U6026 ( .A(b[3787]), .B(n1929), .Z(c[3787]) );
  XOR U6027 ( .A(n1930), .B(n1931), .Z(n1927) );
  ANDN U6028 ( .B(n1932), .A(n1933), .Z(n1930) );
  XNOR U6029 ( .A(b[3786]), .B(n1931), .Z(n1932) );
  XNOR U6030 ( .A(b[3786]), .B(n1933), .Z(c[3786]) );
  XOR U6031 ( .A(n1934), .B(n1935), .Z(n1931) );
  ANDN U6032 ( .B(n1936), .A(n1937), .Z(n1934) );
  XNOR U6033 ( .A(b[3785]), .B(n1935), .Z(n1936) );
  XNOR U6034 ( .A(b[3785]), .B(n1937), .Z(c[3785]) );
  XOR U6035 ( .A(n1938), .B(n1939), .Z(n1935) );
  ANDN U6036 ( .B(n1940), .A(n1941), .Z(n1938) );
  XNOR U6037 ( .A(b[3784]), .B(n1939), .Z(n1940) );
  XNOR U6038 ( .A(b[3784]), .B(n1941), .Z(c[3784]) );
  XOR U6039 ( .A(n1942), .B(n1943), .Z(n1939) );
  ANDN U6040 ( .B(n1944), .A(n1945), .Z(n1942) );
  XNOR U6041 ( .A(b[3783]), .B(n1943), .Z(n1944) );
  XNOR U6042 ( .A(b[3783]), .B(n1945), .Z(c[3783]) );
  XOR U6043 ( .A(n1946), .B(n1947), .Z(n1943) );
  ANDN U6044 ( .B(n1948), .A(n1949), .Z(n1946) );
  XNOR U6045 ( .A(b[3782]), .B(n1947), .Z(n1948) );
  XNOR U6046 ( .A(b[3782]), .B(n1949), .Z(c[3782]) );
  XOR U6047 ( .A(n1950), .B(n1951), .Z(n1947) );
  ANDN U6048 ( .B(n1952), .A(n1953), .Z(n1950) );
  XNOR U6049 ( .A(b[3781]), .B(n1951), .Z(n1952) );
  XNOR U6050 ( .A(b[3781]), .B(n1953), .Z(c[3781]) );
  XOR U6051 ( .A(n1954), .B(n1955), .Z(n1951) );
  ANDN U6052 ( .B(n1956), .A(n1957), .Z(n1954) );
  XNOR U6053 ( .A(b[3780]), .B(n1955), .Z(n1956) );
  XNOR U6054 ( .A(b[3780]), .B(n1957), .Z(c[3780]) );
  XOR U6055 ( .A(n1958), .B(n1959), .Z(n1955) );
  ANDN U6056 ( .B(n1960), .A(n1961), .Z(n1958) );
  XNOR U6057 ( .A(b[3779]), .B(n1959), .Z(n1960) );
  XNOR U6058 ( .A(b[377]), .B(n1962), .Z(c[377]) );
  XNOR U6059 ( .A(b[3779]), .B(n1961), .Z(c[3779]) );
  XOR U6060 ( .A(n1963), .B(n1964), .Z(n1959) );
  ANDN U6061 ( .B(n1965), .A(n1966), .Z(n1963) );
  XNOR U6062 ( .A(b[3778]), .B(n1964), .Z(n1965) );
  XNOR U6063 ( .A(b[3778]), .B(n1966), .Z(c[3778]) );
  XOR U6064 ( .A(n1967), .B(n1968), .Z(n1964) );
  ANDN U6065 ( .B(n1969), .A(n1970), .Z(n1967) );
  XNOR U6066 ( .A(b[3777]), .B(n1968), .Z(n1969) );
  XNOR U6067 ( .A(b[3777]), .B(n1970), .Z(c[3777]) );
  XOR U6068 ( .A(n1971), .B(n1972), .Z(n1968) );
  ANDN U6069 ( .B(n1973), .A(n1974), .Z(n1971) );
  XNOR U6070 ( .A(b[3776]), .B(n1972), .Z(n1973) );
  XNOR U6071 ( .A(b[3776]), .B(n1974), .Z(c[3776]) );
  XOR U6072 ( .A(n1975), .B(n1976), .Z(n1972) );
  ANDN U6073 ( .B(n1977), .A(n1978), .Z(n1975) );
  XNOR U6074 ( .A(b[3775]), .B(n1976), .Z(n1977) );
  XNOR U6075 ( .A(b[3775]), .B(n1978), .Z(c[3775]) );
  XOR U6076 ( .A(n1979), .B(n1980), .Z(n1976) );
  ANDN U6077 ( .B(n1981), .A(n1982), .Z(n1979) );
  XNOR U6078 ( .A(b[3774]), .B(n1980), .Z(n1981) );
  XNOR U6079 ( .A(b[3774]), .B(n1982), .Z(c[3774]) );
  XOR U6080 ( .A(n1983), .B(n1984), .Z(n1980) );
  ANDN U6081 ( .B(n1985), .A(n1986), .Z(n1983) );
  XNOR U6082 ( .A(b[3773]), .B(n1984), .Z(n1985) );
  XNOR U6083 ( .A(b[3773]), .B(n1986), .Z(c[3773]) );
  XOR U6084 ( .A(n1987), .B(n1988), .Z(n1984) );
  ANDN U6085 ( .B(n1989), .A(n1990), .Z(n1987) );
  XNOR U6086 ( .A(b[3772]), .B(n1988), .Z(n1989) );
  XNOR U6087 ( .A(b[3772]), .B(n1990), .Z(c[3772]) );
  XOR U6088 ( .A(n1991), .B(n1992), .Z(n1988) );
  ANDN U6089 ( .B(n1993), .A(n1994), .Z(n1991) );
  XNOR U6090 ( .A(b[3771]), .B(n1992), .Z(n1993) );
  XNOR U6091 ( .A(b[3771]), .B(n1994), .Z(c[3771]) );
  XOR U6092 ( .A(n1995), .B(n1996), .Z(n1992) );
  ANDN U6093 ( .B(n1997), .A(n1998), .Z(n1995) );
  XNOR U6094 ( .A(b[3770]), .B(n1996), .Z(n1997) );
  XNOR U6095 ( .A(b[3770]), .B(n1998), .Z(c[3770]) );
  XOR U6096 ( .A(n1999), .B(n2000), .Z(n1996) );
  ANDN U6097 ( .B(n2001), .A(n2002), .Z(n1999) );
  XNOR U6098 ( .A(b[3769]), .B(n2000), .Z(n2001) );
  XNOR U6099 ( .A(b[376]), .B(n2003), .Z(c[376]) );
  XNOR U6100 ( .A(b[3769]), .B(n2002), .Z(c[3769]) );
  XOR U6101 ( .A(n2004), .B(n2005), .Z(n2000) );
  ANDN U6102 ( .B(n2006), .A(n2007), .Z(n2004) );
  XNOR U6103 ( .A(b[3768]), .B(n2005), .Z(n2006) );
  XNOR U6104 ( .A(b[3768]), .B(n2007), .Z(c[3768]) );
  XOR U6105 ( .A(n2008), .B(n2009), .Z(n2005) );
  ANDN U6106 ( .B(n2010), .A(n2011), .Z(n2008) );
  XNOR U6107 ( .A(b[3767]), .B(n2009), .Z(n2010) );
  XNOR U6108 ( .A(b[3767]), .B(n2011), .Z(c[3767]) );
  XOR U6109 ( .A(n2012), .B(n2013), .Z(n2009) );
  ANDN U6110 ( .B(n2014), .A(n2015), .Z(n2012) );
  XNOR U6111 ( .A(b[3766]), .B(n2013), .Z(n2014) );
  XNOR U6112 ( .A(b[3766]), .B(n2015), .Z(c[3766]) );
  XOR U6113 ( .A(n2016), .B(n2017), .Z(n2013) );
  ANDN U6114 ( .B(n2018), .A(n2019), .Z(n2016) );
  XNOR U6115 ( .A(b[3765]), .B(n2017), .Z(n2018) );
  XNOR U6116 ( .A(b[3765]), .B(n2019), .Z(c[3765]) );
  XOR U6117 ( .A(n2020), .B(n2021), .Z(n2017) );
  ANDN U6118 ( .B(n2022), .A(n2023), .Z(n2020) );
  XNOR U6119 ( .A(b[3764]), .B(n2021), .Z(n2022) );
  XNOR U6120 ( .A(b[3764]), .B(n2023), .Z(c[3764]) );
  XOR U6121 ( .A(n2024), .B(n2025), .Z(n2021) );
  ANDN U6122 ( .B(n2026), .A(n2027), .Z(n2024) );
  XNOR U6123 ( .A(b[3763]), .B(n2025), .Z(n2026) );
  XNOR U6124 ( .A(b[3763]), .B(n2027), .Z(c[3763]) );
  XOR U6125 ( .A(n2028), .B(n2029), .Z(n2025) );
  ANDN U6126 ( .B(n2030), .A(n2031), .Z(n2028) );
  XNOR U6127 ( .A(b[3762]), .B(n2029), .Z(n2030) );
  XNOR U6128 ( .A(b[3762]), .B(n2031), .Z(c[3762]) );
  XOR U6129 ( .A(n2032), .B(n2033), .Z(n2029) );
  ANDN U6130 ( .B(n2034), .A(n2035), .Z(n2032) );
  XNOR U6131 ( .A(b[3761]), .B(n2033), .Z(n2034) );
  XNOR U6132 ( .A(b[3761]), .B(n2035), .Z(c[3761]) );
  XOR U6133 ( .A(n2036), .B(n2037), .Z(n2033) );
  ANDN U6134 ( .B(n2038), .A(n2039), .Z(n2036) );
  XNOR U6135 ( .A(b[3760]), .B(n2037), .Z(n2038) );
  XNOR U6136 ( .A(b[3760]), .B(n2039), .Z(c[3760]) );
  XOR U6137 ( .A(n2040), .B(n2041), .Z(n2037) );
  ANDN U6138 ( .B(n2042), .A(n2043), .Z(n2040) );
  XNOR U6139 ( .A(b[3759]), .B(n2041), .Z(n2042) );
  XNOR U6140 ( .A(b[375]), .B(n2044), .Z(c[375]) );
  XNOR U6141 ( .A(b[3759]), .B(n2043), .Z(c[3759]) );
  XOR U6142 ( .A(n2045), .B(n2046), .Z(n2041) );
  ANDN U6143 ( .B(n2047), .A(n2048), .Z(n2045) );
  XNOR U6144 ( .A(b[3758]), .B(n2046), .Z(n2047) );
  XNOR U6145 ( .A(b[3758]), .B(n2048), .Z(c[3758]) );
  XOR U6146 ( .A(n2049), .B(n2050), .Z(n2046) );
  ANDN U6147 ( .B(n2051), .A(n2052), .Z(n2049) );
  XNOR U6148 ( .A(b[3757]), .B(n2050), .Z(n2051) );
  XNOR U6149 ( .A(b[3757]), .B(n2052), .Z(c[3757]) );
  XOR U6150 ( .A(n2053), .B(n2054), .Z(n2050) );
  ANDN U6151 ( .B(n2055), .A(n2056), .Z(n2053) );
  XNOR U6152 ( .A(b[3756]), .B(n2054), .Z(n2055) );
  XNOR U6153 ( .A(b[3756]), .B(n2056), .Z(c[3756]) );
  XOR U6154 ( .A(n2057), .B(n2058), .Z(n2054) );
  ANDN U6155 ( .B(n2059), .A(n2060), .Z(n2057) );
  XNOR U6156 ( .A(b[3755]), .B(n2058), .Z(n2059) );
  XNOR U6157 ( .A(b[3755]), .B(n2060), .Z(c[3755]) );
  XOR U6158 ( .A(n2061), .B(n2062), .Z(n2058) );
  ANDN U6159 ( .B(n2063), .A(n2064), .Z(n2061) );
  XNOR U6160 ( .A(b[3754]), .B(n2062), .Z(n2063) );
  XNOR U6161 ( .A(b[3754]), .B(n2064), .Z(c[3754]) );
  XOR U6162 ( .A(n2065), .B(n2066), .Z(n2062) );
  ANDN U6163 ( .B(n2067), .A(n2068), .Z(n2065) );
  XNOR U6164 ( .A(b[3753]), .B(n2066), .Z(n2067) );
  XNOR U6165 ( .A(b[3753]), .B(n2068), .Z(c[3753]) );
  XOR U6166 ( .A(n2069), .B(n2070), .Z(n2066) );
  ANDN U6167 ( .B(n2071), .A(n2072), .Z(n2069) );
  XNOR U6168 ( .A(b[3752]), .B(n2070), .Z(n2071) );
  XNOR U6169 ( .A(b[3752]), .B(n2072), .Z(c[3752]) );
  XOR U6170 ( .A(n2073), .B(n2074), .Z(n2070) );
  ANDN U6171 ( .B(n2075), .A(n2076), .Z(n2073) );
  XNOR U6172 ( .A(b[3751]), .B(n2074), .Z(n2075) );
  XNOR U6173 ( .A(b[3751]), .B(n2076), .Z(c[3751]) );
  XOR U6174 ( .A(n2077), .B(n2078), .Z(n2074) );
  ANDN U6175 ( .B(n2079), .A(n2080), .Z(n2077) );
  XNOR U6176 ( .A(b[3750]), .B(n2078), .Z(n2079) );
  XNOR U6177 ( .A(b[3750]), .B(n2080), .Z(c[3750]) );
  XOR U6178 ( .A(n2081), .B(n2082), .Z(n2078) );
  ANDN U6179 ( .B(n2083), .A(n2084), .Z(n2081) );
  XNOR U6180 ( .A(b[3749]), .B(n2082), .Z(n2083) );
  XNOR U6181 ( .A(b[374]), .B(n2085), .Z(c[374]) );
  XNOR U6182 ( .A(b[3749]), .B(n2084), .Z(c[3749]) );
  XOR U6183 ( .A(n2086), .B(n2087), .Z(n2082) );
  ANDN U6184 ( .B(n2088), .A(n2089), .Z(n2086) );
  XNOR U6185 ( .A(b[3748]), .B(n2087), .Z(n2088) );
  XNOR U6186 ( .A(b[3748]), .B(n2089), .Z(c[3748]) );
  XOR U6187 ( .A(n2090), .B(n2091), .Z(n2087) );
  ANDN U6188 ( .B(n2092), .A(n2093), .Z(n2090) );
  XNOR U6189 ( .A(b[3747]), .B(n2091), .Z(n2092) );
  XNOR U6190 ( .A(b[3747]), .B(n2093), .Z(c[3747]) );
  XOR U6191 ( .A(n2094), .B(n2095), .Z(n2091) );
  ANDN U6192 ( .B(n2096), .A(n2097), .Z(n2094) );
  XNOR U6193 ( .A(b[3746]), .B(n2095), .Z(n2096) );
  XNOR U6194 ( .A(b[3746]), .B(n2097), .Z(c[3746]) );
  XOR U6195 ( .A(n2098), .B(n2099), .Z(n2095) );
  ANDN U6196 ( .B(n2100), .A(n2101), .Z(n2098) );
  XNOR U6197 ( .A(b[3745]), .B(n2099), .Z(n2100) );
  XNOR U6198 ( .A(b[3745]), .B(n2101), .Z(c[3745]) );
  XOR U6199 ( .A(n2102), .B(n2103), .Z(n2099) );
  ANDN U6200 ( .B(n2104), .A(n2105), .Z(n2102) );
  XNOR U6201 ( .A(b[3744]), .B(n2103), .Z(n2104) );
  XNOR U6202 ( .A(b[3744]), .B(n2105), .Z(c[3744]) );
  XOR U6203 ( .A(n2106), .B(n2107), .Z(n2103) );
  ANDN U6204 ( .B(n2108), .A(n2109), .Z(n2106) );
  XNOR U6205 ( .A(b[3743]), .B(n2107), .Z(n2108) );
  XNOR U6206 ( .A(b[3743]), .B(n2109), .Z(c[3743]) );
  XOR U6207 ( .A(n2110), .B(n2111), .Z(n2107) );
  ANDN U6208 ( .B(n2112), .A(n2113), .Z(n2110) );
  XNOR U6209 ( .A(b[3742]), .B(n2111), .Z(n2112) );
  XNOR U6210 ( .A(b[3742]), .B(n2113), .Z(c[3742]) );
  XOR U6211 ( .A(n2114), .B(n2115), .Z(n2111) );
  ANDN U6212 ( .B(n2116), .A(n2117), .Z(n2114) );
  XNOR U6213 ( .A(b[3741]), .B(n2115), .Z(n2116) );
  XNOR U6214 ( .A(b[3741]), .B(n2117), .Z(c[3741]) );
  XOR U6215 ( .A(n2118), .B(n2119), .Z(n2115) );
  ANDN U6216 ( .B(n2120), .A(n2121), .Z(n2118) );
  XNOR U6217 ( .A(b[3740]), .B(n2119), .Z(n2120) );
  XNOR U6218 ( .A(b[3740]), .B(n2121), .Z(c[3740]) );
  XOR U6219 ( .A(n2122), .B(n2123), .Z(n2119) );
  ANDN U6220 ( .B(n2124), .A(n2125), .Z(n2122) );
  XNOR U6221 ( .A(b[3739]), .B(n2123), .Z(n2124) );
  XNOR U6222 ( .A(b[373]), .B(n2126), .Z(c[373]) );
  XNOR U6223 ( .A(b[3739]), .B(n2125), .Z(c[3739]) );
  XOR U6224 ( .A(n2127), .B(n2128), .Z(n2123) );
  ANDN U6225 ( .B(n2129), .A(n2130), .Z(n2127) );
  XNOR U6226 ( .A(b[3738]), .B(n2128), .Z(n2129) );
  XNOR U6227 ( .A(b[3738]), .B(n2130), .Z(c[3738]) );
  XOR U6228 ( .A(n2131), .B(n2132), .Z(n2128) );
  ANDN U6229 ( .B(n2133), .A(n2134), .Z(n2131) );
  XNOR U6230 ( .A(b[3737]), .B(n2132), .Z(n2133) );
  XNOR U6231 ( .A(b[3737]), .B(n2134), .Z(c[3737]) );
  XOR U6232 ( .A(n2135), .B(n2136), .Z(n2132) );
  ANDN U6233 ( .B(n2137), .A(n2138), .Z(n2135) );
  XNOR U6234 ( .A(b[3736]), .B(n2136), .Z(n2137) );
  XNOR U6235 ( .A(b[3736]), .B(n2138), .Z(c[3736]) );
  XOR U6236 ( .A(n2139), .B(n2140), .Z(n2136) );
  ANDN U6237 ( .B(n2141), .A(n2142), .Z(n2139) );
  XNOR U6238 ( .A(b[3735]), .B(n2140), .Z(n2141) );
  XNOR U6239 ( .A(b[3735]), .B(n2142), .Z(c[3735]) );
  XOR U6240 ( .A(n2143), .B(n2144), .Z(n2140) );
  ANDN U6241 ( .B(n2145), .A(n2146), .Z(n2143) );
  XNOR U6242 ( .A(b[3734]), .B(n2144), .Z(n2145) );
  XNOR U6243 ( .A(b[3734]), .B(n2146), .Z(c[3734]) );
  XOR U6244 ( .A(n2147), .B(n2148), .Z(n2144) );
  ANDN U6245 ( .B(n2149), .A(n2150), .Z(n2147) );
  XNOR U6246 ( .A(b[3733]), .B(n2148), .Z(n2149) );
  XNOR U6247 ( .A(b[3733]), .B(n2150), .Z(c[3733]) );
  XOR U6248 ( .A(n2151), .B(n2152), .Z(n2148) );
  ANDN U6249 ( .B(n2153), .A(n2154), .Z(n2151) );
  XNOR U6250 ( .A(b[3732]), .B(n2152), .Z(n2153) );
  XNOR U6251 ( .A(b[3732]), .B(n2154), .Z(c[3732]) );
  XOR U6252 ( .A(n2155), .B(n2156), .Z(n2152) );
  ANDN U6253 ( .B(n2157), .A(n2158), .Z(n2155) );
  XNOR U6254 ( .A(b[3731]), .B(n2156), .Z(n2157) );
  XNOR U6255 ( .A(b[3731]), .B(n2158), .Z(c[3731]) );
  XOR U6256 ( .A(n2159), .B(n2160), .Z(n2156) );
  ANDN U6257 ( .B(n2161), .A(n2162), .Z(n2159) );
  XNOR U6258 ( .A(b[3730]), .B(n2160), .Z(n2161) );
  XNOR U6259 ( .A(b[3730]), .B(n2162), .Z(c[3730]) );
  XOR U6260 ( .A(n2163), .B(n2164), .Z(n2160) );
  ANDN U6261 ( .B(n2165), .A(n2166), .Z(n2163) );
  XNOR U6262 ( .A(b[3729]), .B(n2164), .Z(n2165) );
  XNOR U6263 ( .A(b[372]), .B(n2167), .Z(c[372]) );
  XNOR U6264 ( .A(b[3729]), .B(n2166), .Z(c[3729]) );
  XOR U6265 ( .A(n2168), .B(n2169), .Z(n2164) );
  ANDN U6266 ( .B(n2170), .A(n2171), .Z(n2168) );
  XNOR U6267 ( .A(b[3728]), .B(n2169), .Z(n2170) );
  XNOR U6268 ( .A(b[3728]), .B(n2171), .Z(c[3728]) );
  XOR U6269 ( .A(n2172), .B(n2173), .Z(n2169) );
  ANDN U6270 ( .B(n2174), .A(n2175), .Z(n2172) );
  XNOR U6271 ( .A(b[3727]), .B(n2173), .Z(n2174) );
  XNOR U6272 ( .A(b[3727]), .B(n2175), .Z(c[3727]) );
  XOR U6273 ( .A(n2176), .B(n2177), .Z(n2173) );
  ANDN U6274 ( .B(n2178), .A(n2179), .Z(n2176) );
  XNOR U6275 ( .A(b[3726]), .B(n2177), .Z(n2178) );
  XNOR U6276 ( .A(b[3726]), .B(n2179), .Z(c[3726]) );
  XOR U6277 ( .A(n2180), .B(n2181), .Z(n2177) );
  ANDN U6278 ( .B(n2182), .A(n2183), .Z(n2180) );
  XNOR U6279 ( .A(b[3725]), .B(n2181), .Z(n2182) );
  XNOR U6280 ( .A(b[3725]), .B(n2183), .Z(c[3725]) );
  XOR U6281 ( .A(n2184), .B(n2185), .Z(n2181) );
  ANDN U6282 ( .B(n2186), .A(n2187), .Z(n2184) );
  XNOR U6283 ( .A(b[3724]), .B(n2185), .Z(n2186) );
  XNOR U6284 ( .A(b[3724]), .B(n2187), .Z(c[3724]) );
  XOR U6285 ( .A(n2188), .B(n2189), .Z(n2185) );
  ANDN U6286 ( .B(n2190), .A(n2191), .Z(n2188) );
  XNOR U6287 ( .A(b[3723]), .B(n2189), .Z(n2190) );
  XNOR U6288 ( .A(b[3723]), .B(n2191), .Z(c[3723]) );
  XOR U6289 ( .A(n2192), .B(n2193), .Z(n2189) );
  ANDN U6290 ( .B(n2194), .A(n2195), .Z(n2192) );
  XNOR U6291 ( .A(b[3722]), .B(n2193), .Z(n2194) );
  XNOR U6292 ( .A(b[3722]), .B(n2195), .Z(c[3722]) );
  XOR U6293 ( .A(n2196), .B(n2197), .Z(n2193) );
  ANDN U6294 ( .B(n2198), .A(n2199), .Z(n2196) );
  XNOR U6295 ( .A(b[3721]), .B(n2197), .Z(n2198) );
  XNOR U6296 ( .A(b[3721]), .B(n2199), .Z(c[3721]) );
  XOR U6297 ( .A(n2200), .B(n2201), .Z(n2197) );
  ANDN U6298 ( .B(n2202), .A(n2203), .Z(n2200) );
  XNOR U6299 ( .A(b[3720]), .B(n2201), .Z(n2202) );
  XNOR U6300 ( .A(b[3720]), .B(n2203), .Z(c[3720]) );
  XOR U6301 ( .A(n2204), .B(n2205), .Z(n2201) );
  ANDN U6302 ( .B(n2206), .A(n2207), .Z(n2204) );
  XNOR U6303 ( .A(b[3719]), .B(n2205), .Z(n2206) );
  XNOR U6304 ( .A(b[371]), .B(n2208), .Z(c[371]) );
  XNOR U6305 ( .A(b[3719]), .B(n2207), .Z(c[3719]) );
  XOR U6306 ( .A(n2209), .B(n2210), .Z(n2205) );
  ANDN U6307 ( .B(n2211), .A(n2212), .Z(n2209) );
  XNOR U6308 ( .A(b[3718]), .B(n2210), .Z(n2211) );
  XNOR U6309 ( .A(b[3718]), .B(n2212), .Z(c[3718]) );
  XOR U6310 ( .A(n2213), .B(n2214), .Z(n2210) );
  ANDN U6311 ( .B(n2215), .A(n2216), .Z(n2213) );
  XNOR U6312 ( .A(b[3717]), .B(n2214), .Z(n2215) );
  XNOR U6313 ( .A(b[3717]), .B(n2216), .Z(c[3717]) );
  XOR U6314 ( .A(n2217), .B(n2218), .Z(n2214) );
  ANDN U6315 ( .B(n2219), .A(n2220), .Z(n2217) );
  XNOR U6316 ( .A(b[3716]), .B(n2218), .Z(n2219) );
  XNOR U6317 ( .A(b[3716]), .B(n2220), .Z(c[3716]) );
  XOR U6318 ( .A(n2221), .B(n2222), .Z(n2218) );
  ANDN U6319 ( .B(n2223), .A(n2224), .Z(n2221) );
  XNOR U6320 ( .A(b[3715]), .B(n2222), .Z(n2223) );
  XNOR U6321 ( .A(b[3715]), .B(n2224), .Z(c[3715]) );
  XOR U6322 ( .A(n2225), .B(n2226), .Z(n2222) );
  ANDN U6323 ( .B(n2227), .A(n2228), .Z(n2225) );
  XNOR U6324 ( .A(b[3714]), .B(n2226), .Z(n2227) );
  XNOR U6325 ( .A(b[3714]), .B(n2228), .Z(c[3714]) );
  XOR U6326 ( .A(n2229), .B(n2230), .Z(n2226) );
  ANDN U6327 ( .B(n2231), .A(n2232), .Z(n2229) );
  XNOR U6328 ( .A(b[3713]), .B(n2230), .Z(n2231) );
  XNOR U6329 ( .A(b[3713]), .B(n2232), .Z(c[3713]) );
  XOR U6330 ( .A(n2233), .B(n2234), .Z(n2230) );
  ANDN U6331 ( .B(n2235), .A(n2236), .Z(n2233) );
  XNOR U6332 ( .A(b[3712]), .B(n2234), .Z(n2235) );
  XNOR U6333 ( .A(b[3712]), .B(n2236), .Z(c[3712]) );
  XOR U6334 ( .A(n2237), .B(n2238), .Z(n2234) );
  ANDN U6335 ( .B(n2239), .A(n2240), .Z(n2237) );
  XNOR U6336 ( .A(b[3711]), .B(n2238), .Z(n2239) );
  XNOR U6337 ( .A(b[3711]), .B(n2240), .Z(c[3711]) );
  XOR U6338 ( .A(n2241), .B(n2242), .Z(n2238) );
  ANDN U6339 ( .B(n2243), .A(n2244), .Z(n2241) );
  XNOR U6340 ( .A(b[3710]), .B(n2242), .Z(n2243) );
  XNOR U6341 ( .A(b[3710]), .B(n2244), .Z(c[3710]) );
  XOR U6342 ( .A(n2245), .B(n2246), .Z(n2242) );
  ANDN U6343 ( .B(n2247), .A(n2248), .Z(n2245) );
  XNOR U6344 ( .A(b[3709]), .B(n2246), .Z(n2247) );
  XNOR U6345 ( .A(b[370]), .B(n2249), .Z(c[370]) );
  XNOR U6346 ( .A(b[3709]), .B(n2248), .Z(c[3709]) );
  XOR U6347 ( .A(n2250), .B(n2251), .Z(n2246) );
  ANDN U6348 ( .B(n2252), .A(n2253), .Z(n2250) );
  XNOR U6349 ( .A(b[3708]), .B(n2251), .Z(n2252) );
  XNOR U6350 ( .A(b[3708]), .B(n2253), .Z(c[3708]) );
  XOR U6351 ( .A(n2254), .B(n2255), .Z(n2251) );
  ANDN U6352 ( .B(n2256), .A(n2257), .Z(n2254) );
  XNOR U6353 ( .A(b[3707]), .B(n2255), .Z(n2256) );
  XNOR U6354 ( .A(b[3707]), .B(n2257), .Z(c[3707]) );
  XOR U6355 ( .A(n2258), .B(n2259), .Z(n2255) );
  ANDN U6356 ( .B(n2260), .A(n2261), .Z(n2258) );
  XNOR U6357 ( .A(b[3706]), .B(n2259), .Z(n2260) );
  XNOR U6358 ( .A(b[3706]), .B(n2261), .Z(c[3706]) );
  XOR U6359 ( .A(n2262), .B(n2263), .Z(n2259) );
  ANDN U6360 ( .B(n2264), .A(n2265), .Z(n2262) );
  XNOR U6361 ( .A(b[3705]), .B(n2263), .Z(n2264) );
  XNOR U6362 ( .A(b[3705]), .B(n2265), .Z(c[3705]) );
  XOR U6363 ( .A(n2266), .B(n2267), .Z(n2263) );
  ANDN U6364 ( .B(n2268), .A(n2269), .Z(n2266) );
  XNOR U6365 ( .A(b[3704]), .B(n2267), .Z(n2268) );
  XNOR U6366 ( .A(b[3704]), .B(n2269), .Z(c[3704]) );
  XOR U6367 ( .A(n2270), .B(n2271), .Z(n2267) );
  ANDN U6368 ( .B(n2272), .A(n2273), .Z(n2270) );
  XNOR U6369 ( .A(b[3703]), .B(n2271), .Z(n2272) );
  XNOR U6370 ( .A(b[3703]), .B(n2273), .Z(c[3703]) );
  XOR U6371 ( .A(n2274), .B(n2275), .Z(n2271) );
  ANDN U6372 ( .B(n2276), .A(n2277), .Z(n2274) );
  XNOR U6373 ( .A(b[3702]), .B(n2275), .Z(n2276) );
  XNOR U6374 ( .A(b[3702]), .B(n2277), .Z(c[3702]) );
  XOR U6375 ( .A(n2278), .B(n2279), .Z(n2275) );
  ANDN U6376 ( .B(n2280), .A(n2281), .Z(n2278) );
  XNOR U6377 ( .A(b[3701]), .B(n2279), .Z(n2280) );
  XNOR U6378 ( .A(b[3701]), .B(n2281), .Z(c[3701]) );
  XOR U6379 ( .A(n2282), .B(n2283), .Z(n2279) );
  ANDN U6380 ( .B(n2284), .A(n2285), .Z(n2282) );
  XNOR U6381 ( .A(b[3700]), .B(n2283), .Z(n2284) );
  XNOR U6382 ( .A(b[3700]), .B(n2285), .Z(c[3700]) );
  XOR U6383 ( .A(n2286), .B(n2287), .Z(n2283) );
  ANDN U6384 ( .B(n2288), .A(n2289), .Z(n2286) );
  XNOR U6385 ( .A(b[3699]), .B(n2287), .Z(n2288) );
  XNOR U6386 ( .A(b[36]), .B(n2290), .Z(c[36]) );
  XNOR U6387 ( .A(b[369]), .B(n2291), .Z(c[369]) );
  XNOR U6388 ( .A(b[3699]), .B(n2289), .Z(c[3699]) );
  XOR U6389 ( .A(n2292), .B(n2293), .Z(n2287) );
  ANDN U6390 ( .B(n2294), .A(n2295), .Z(n2292) );
  XNOR U6391 ( .A(b[3698]), .B(n2293), .Z(n2294) );
  XNOR U6392 ( .A(b[3698]), .B(n2295), .Z(c[3698]) );
  XOR U6393 ( .A(n2296), .B(n2297), .Z(n2293) );
  ANDN U6394 ( .B(n2298), .A(n2299), .Z(n2296) );
  XNOR U6395 ( .A(b[3697]), .B(n2297), .Z(n2298) );
  XNOR U6396 ( .A(b[3697]), .B(n2299), .Z(c[3697]) );
  XOR U6397 ( .A(n2300), .B(n2301), .Z(n2297) );
  ANDN U6398 ( .B(n2302), .A(n2303), .Z(n2300) );
  XNOR U6399 ( .A(b[3696]), .B(n2301), .Z(n2302) );
  XNOR U6400 ( .A(b[3696]), .B(n2303), .Z(c[3696]) );
  XOR U6401 ( .A(n2304), .B(n2305), .Z(n2301) );
  ANDN U6402 ( .B(n2306), .A(n2307), .Z(n2304) );
  XNOR U6403 ( .A(b[3695]), .B(n2305), .Z(n2306) );
  XNOR U6404 ( .A(b[3695]), .B(n2307), .Z(c[3695]) );
  XOR U6405 ( .A(n2308), .B(n2309), .Z(n2305) );
  ANDN U6406 ( .B(n2310), .A(n2311), .Z(n2308) );
  XNOR U6407 ( .A(b[3694]), .B(n2309), .Z(n2310) );
  XNOR U6408 ( .A(b[3694]), .B(n2311), .Z(c[3694]) );
  XOR U6409 ( .A(n2312), .B(n2313), .Z(n2309) );
  ANDN U6410 ( .B(n2314), .A(n2315), .Z(n2312) );
  XNOR U6411 ( .A(b[3693]), .B(n2313), .Z(n2314) );
  XNOR U6412 ( .A(b[3693]), .B(n2315), .Z(c[3693]) );
  XOR U6413 ( .A(n2316), .B(n2317), .Z(n2313) );
  ANDN U6414 ( .B(n2318), .A(n2319), .Z(n2316) );
  XNOR U6415 ( .A(b[3692]), .B(n2317), .Z(n2318) );
  XNOR U6416 ( .A(b[3692]), .B(n2319), .Z(c[3692]) );
  XOR U6417 ( .A(n2320), .B(n2321), .Z(n2317) );
  ANDN U6418 ( .B(n2322), .A(n2323), .Z(n2320) );
  XNOR U6419 ( .A(b[3691]), .B(n2321), .Z(n2322) );
  XNOR U6420 ( .A(b[3691]), .B(n2323), .Z(c[3691]) );
  XOR U6421 ( .A(n2324), .B(n2325), .Z(n2321) );
  ANDN U6422 ( .B(n2326), .A(n2327), .Z(n2324) );
  XNOR U6423 ( .A(b[3690]), .B(n2325), .Z(n2326) );
  XNOR U6424 ( .A(b[3690]), .B(n2327), .Z(c[3690]) );
  XOR U6425 ( .A(n2328), .B(n2329), .Z(n2325) );
  ANDN U6426 ( .B(n2330), .A(n2331), .Z(n2328) );
  XNOR U6427 ( .A(b[3689]), .B(n2329), .Z(n2330) );
  XNOR U6428 ( .A(b[368]), .B(n2332), .Z(c[368]) );
  XNOR U6429 ( .A(b[3689]), .B(n2331), .Z(c[3689]) );
  XOR U6430 ( .A(n2333), .B(n2334), .Z(n2329) );
  ANDN U6431 ( .B(n2335), .A(n2336), .Z(n2333) );
  XNOR U6432 ( .A(b[3688]), .B(n2334), .Z(n2335) );
  XNOR U6433 ( .A(b[3688]), .B(n2336), .Z(c[3688]) );
  XOR U6434 ( .A(n2337), .B(n2338), .Z(n2334) );
  ANDN U6435 ( .B(n2339), .A(n2340), .Z(n2337) );
  XNOR U6436 ( .A(b[3687]), .B(n2338), .Z(n2339) );
  XNOR U6437 ( .A(b[3687]), .B(n2340), .Z(c[3687]) );
  XOR U6438 ( .A(n2341), .B(n2342), .Z(n2338) );
  ANDN U6439 ( .B(n2343), .A(n2344), .Z(n2341) );
  XNOR U6440 ( .A(b[3686]), .B(n2342), .Z(n2343) );
  XNOR U6441 ( .A(b[3686]), .B(n2344), .Z(c[3686]) );
  XOR U6442 ( .A(n2345), .B(n2346), .Z(n2342) );
  ANDN U6443 ( .B(n2347), .A(n2348), .Z(n2345) );
  XNOR U6444 ( .A(b[3685]), .B(n2346), .Z(n2347) );
  XNOR U6445 ( .A(b[3685]), .B(n2348), .Z(c[3685]) );
  XOR U6446 ( .A(n2349), .B(n2350), .Z(n2346) );
  ANDN U6447 ( .B(n2351), .A(n2352), .Z(n2349) );
  XNOR U6448 ( .A(b[3684]), .B(n2350), .Z(n2351) );
  XNOR U6449 ( .A(b[3684]), .B(n2352), .Z(c[3684]) );
  XOR U6450 ( .A(n2353), .B(n2354), .Z(n2350) );
  ANDN U6451 ( .B(n2355), .A(n2356), .Z(n2353) );
  XNOR U6452 ( .A(b[3683]), .B(n2354), .Z(n2355) );
  XNOR U6453 ( .A(b[3683]), .B(n2356), .Z(c[3683]) );
  XOR U6454 ( .A(n2357), .B(n2358), .Z(n2354) );
  ANDN U6455 ( .B(n2359), .A(n2360), .Z(n2357) );
  XNOR U6456 ( .A(b[3682]), .B(n2358), .Z(n2359) );
  XNOR U6457 ( .A(b[3682]), .B(n2360), .Z(c[3682]) );
  XOR U6458 ( .A(n2361), .B(n2362), .Z(n2358) );
  ANDN U6459 ( .B(n2363), .A(n2364), .Z(n2361) );
  XNOR U6460 ( .A(b[3681]), .B(n2362), .Z(n2363) );
  XNOR U6461 ( .A(b[3681]), .B(n2364), .Z(c[3681]) );
  XOR U6462 ( .A(n2365), .B(n2366), .Z(n2362) );
  ANDN U6463 ( .B(n2367), .A(n2368), .Z(n2365) );
  XNOR U6464 ( .A(b[3680]), .B(n2366), .Z(n2367) );
  XNOR U6465 ( .A(b[3680]), .B(n2368), .Z(c[3680]) );
  XOR U6466 ( .A(n2369), .B(n2370), .Z(n2366) );
  ANDN U6467 ( .B(n2371), .A(n2372), .Z(n2369) );
  XNOR U6468 ( .A(b[3679]), .B(n2370), .Z(n2371) );
  XNOR U6469 ( .A(b[367]), .B(n2373), .Z(c[367]) );
  XNOR U6470 ( .A(b[3679]), .B(n2372), .Z(c[3679]) );
  XOR U6471 ( .A(n2374), .B(n2375), .Z(n2370) );
  ANDN U6472 ( .B(n2376), .A(n2377), .Z(n2374) );
  XNOR U6473 ( .A(b[3678]), .B(n2375), .Z(n2376) );
  XNOR U6474 ( .A(b[3678]), .B(n2377), .Z(c[3678]) );
  XOR U6475 ( .A(n2378), .B(n2379), .Z(n2375) );
  ANDN U6476 ( .B(n2380), .A(n2381), .Z(n2378) );
  XNOR U6477 ( .A(b[3677]), .B(n2379), .Z(n2380) );
  XNOR U6478 ( .A(b[3677]), .B(n2381), .Z(c[3677]) );
  XOR U6479 ( .A(n2382), .B(n2383), .Z(n2379) );
  ANDN U6480 ( .B(n2384), .A(n2385), .Z(n2382) );
  XNOR U6481 ( .A(b[3676]), .B(n2383), .Z(n2384) );
  XNOR U6482 ( .A(b[3676]), .B(n2385), .Z(c[3676]) );
  XOR U6483 ( .A(n2386), .B(n2387), .Z(n2383) );
  ANDN U6484 ( .B(n2388), .A(n2389), .Z(n2386) );
  XNOR U6485 ( .A(b[3675]), .B(n2387), .Z(n2388) );
  XNOR U6486 ( .A(b[3675]), .B(n2389), .Z(c[3675]) );
  XOR U6487 ( .A(n2390), .B(n2391), .Z(n2387) );
  ANDN U6488 ( .B(n2392), .A(n2393), .Z(n2390) );
  XNOR U6489 ( .A(b[3674]), .B(n2391), .Z(n2392) );
  XNOR U6490 ( .A(b[3674]), .B(n2393), .Z(c[3674]) );
  XOR U6491 ( .A(n2394), .B(n2395), .Z(n2391) );
  ANDN U6492 ( .B(n2396), .A(n2397), .Z(n2394) );
  XNOR U6493 ( .A(b[3673]), .B(n2395), .Z(n2396) );
  XNOR U6494 ( .A(b[3673]), .B(n2397), .Z(c[3673]) );
  XOR U6495 ( .A(n2398), .B(n2399), .Z(n2395) );
  ANDN U6496 ( .B(n2400), .A(n2401), .Z(n2398) );
  XNOR U6497 ( .A(b[3672]), .B(n2399), .Z(n2400) );
  XNOR U6498 ( .A(b[3672]), .B(n2401), .Z(c[3672]) );
  XOR U6499 ( .A(n2402), .B(n2403), .Z(n2399) );
  ANDN U6500 ( .B(n2404), .A(n2405), .Z(n2402) );
  XNOR U6501 ( .A(b[3671]), .B(n2403), .Z(n2404) );
  XNOR U6502 ( .A(b[3671]), .B(n2405), .Z(c[3671]) );
  XOR U6503 ( .A(n2406), .B(n2407), .Z(n2403) );
  ANDN U6504 ( .B(n2408), .A(n2409), .Z(n2406) );
  XNOR U6505 ( .A(b[3670]), .B(n2407), .Z(n2408) );
  XNOR U6506 ( .A(b[3670]), .B(n2409), .Z(c[3670]) );
  XOR U6507 ( .A(n2410), .B(n2411), .Z(n2407) );
  ANDN U6508 ( .B(n2412), .A(n2413), .Z(n2410) );
  XNOR U6509 ( .A(b[3669]), .B(n2411), .Z(n2412) );
  XNOR U6510 ( .A(b[366]), .B(n2414), .Z(c[366]) );
  XNOR U6511 ( .A(b[3669]), .B(n2413), .Z(c[3669]) );
  XOR U6512 ( .A(n2415), .B(n2416), .Z(n2411) );
  ANDN U6513 ( .B(n2417), .A(n2418), .Z(n2415) );
  XNOR U6514 ( .A(b[3668]), .B(n2416), .Z(n2417) );
  XNOR U6515 ( .A(b[3668]), .B(n2418), .Z(c[3668]) );
  XOR U6516 ( .A(n2419), .B(n2420), .Z(n2416) );
  ANDN U6517 ( .B(n2421), .A(n2422), .Z(n2419) );
  XNOR U6518 ( .A(b[3667]), .B(n2420), .Z(n2421) );
  XNOR U6519 ( .A(b[3667]), .B(n2422), .Z(c[3667]) );
  XOR U6520 ( .A(n2423), .B(n2424), .Z(n2420) );
  ANDN U6521 ( .B(n2425), .A(n2426), .Z(n2423) );
  XNOR U6522 ( .A(b[3666]), .B(n2424), .Z(n2425) );
  XNOR U6523 ( .A(b[3666]), .B(n2426), .Z(c[3666]) );
  XOR U6524 ( .A(n2427), .B(n2428), .Z(n2424) );
  ANDN U6525 ( .B(n2429), .A(n2430), .Z(n2427) );
  XNOR U6526 ( .A(b[3665]), .B(n2428), .Z(n2429) );
  XNOR U6527 ( .A(b[3665]), .B(n2430), .Z(c[3665]) );
  XOR U6528 ( .A(n2431), .B(n2432), .Z(n2428) );
  ANDN U6529 ( .B(n2433), .A(n2434), .Z(n2431) );
  XNOR U6530 ( .A(b[3664]), .B(n2432), .Z(n2433) );
  XNOR U6531 ( .A(b[3664]), .B(n2434), .Z(c[3664]) );
  XOR U6532 ( .A(n2435), .B(n2436), .Z(n2432) );
  ANDN U6533 ( .B(n2437), .A(n2438), .Z(n2435) );
  XNOR U6534 ( .A(b[3663]), .B(n2436), .Z(n2437) );
  XNOR U6535 ( .A(b[3663]), .B(n2438), .Z(c[3663]) );
  XOR U6536 ( .A(n2439), .B(n2440), .Z(n2436) );
  ANDN U6537 ( .B(n2441), .A(n2442), .Z(n2439) );
  XNOR U6538 ( .A(b[3662]), .B(n2440), .Z(n2441) );
  XNOR U6539 ( .A(b[3662]), .B(n2442), .Z(c[3662]) );
  XOR U6540 ( .A(n2443), .B(n2444), .Z(n2440) );
  ANDN U6541 ( .B(n2445), .A(n2446), .Z(n2443) );
  XNOR U6542 ( .A(b[3661]), .B(n2444), .Z(n2445) );
  XNOR U6543 ( .A(b[3661]), .B(n2446), .Z(c[3661]) );
  XOR U6544 ( .A(n2447), .B(n2448), .Z(n2444) );
  ANDN U6545 ( .B(n2449), .A(n2450), .Z(n2447) );
  XNOR U6546 ( .A(b[3660]), .B(n2448), .Z(n2449) );
  XNOR U6547 ( .A(b[3660]), .B(n2450), .Z(c[3660]) );
  XOR U6548 ( .A(n2451), .B(n2452), .Z(n2448) );
  ANDN U6549 ( .B(n2453), .A(n2454), .Z(n2451) );
  XNOR U6550 ( .A(b[3659]), .B(n2452), .Z(n2453) );
  XNOR U6551 ( .A(b[365]), .B(n2455), .Z(c[365]) );
  XNOR U6552 ( .A(b[3659]), .B(n2454), .Z(c[3659]) );
  XOR U6553 ( .A(n2456), .B(n2457), .Z(n2452) );
  ANDN U6554 ( .B(n2458), .A(n2459), .Z(n2456) );
  XNOR U6555 ( .A(b[3658]), .B(n2457), .Z(n2458) );
  XNOR U6556 ( .A(b[3658]), .B(n2459), .Z(c[3658]) );
  XOR U6557 ( .A(n2460), .B(n2461), .Z(n2457) );
  ANDN U6558 ( .B(n2462), .A(n2463), .Z(n2460) );
  XNOR U6559 ( .A(b[3657]), .B(n2461), .Z(n2462) );
  XNOR U6560 ( .A(b[3657]), .B(n2463), .Z(c[3657]) );
  XOR U6561 ( .A(n2464), .B(n2465), .Z(n2461) );
  ANDN U6562 ( .B(n2466), .A(n2467), .Z(n2464) );
  XNOR U6563 ( .A(b[3656]), .B(n2465), .Z(n2466) );
  XNOR U6564 ( .A(b[3656]), .B(n2467), .Z(c[3656]) );
  XOR U6565 ( .A(n2468), .B(n2469), .Z(n2465) );
  ANDN U6566 ( .B(n2470), .A(n2471), .Z(n2468) );
  XNOR U6567 ( .A(b[3655]), .B(n2469), .Z(n2470) );
  XNOR U6568 ( .A(b[3655]), .B(n2471), .Z(c[3655]) );
  XOR U6569 ( .A(n2472), .B(n2473), .Z(n2469) );
  ANDN U6570 ( .B(n2474), .A(n2475), .Z(n2472) );
  XNOR U6571 ( .A(b[3654]), .B(n2473), .Z(n2474) );
  XNOR U6572 ( .A(b[3654]), .B(n2475), .Z(c[3654]) );
  XOR U6573 ( .A(n2476), .B(n2477), .Z(n2473) );
  ANDN U6574 ( .B(n2478), .A(n2479), .Z(n2476) );
  XNOR U6575 ( .A(b[3653]), .B(n2477), .Z(n2478) );
  XNOR U6576 ( .A(b[3653]), .B(n2479), .Z(c[3653]) );
  XOR U6577 ( .A(n2480), .B(n2481), .Z(n2477) );
  ANDN U6578 ( .B(n2482), .A(n2483), .Z(n2480) );
  XNOR U6579 ( .A(b[3652]), .B(n2481), .Z(n2482) );
  XNOR U6580 ( .A(b[3652]), .B(n2483), .Z(c[3652]) );
  XOR U6581 ( .A(n2484), .B(n2485), .Z(n2481) );
  ANDN U6582 ( .B(n2486), .A(n2487), .Z(n2484) );
  XNOR U6583 ( .A(b[3651]), .B(n2485), .Z(n2486) );
  XNOR U6584 ( .A(b[3651]), .B(n2487), .Z(c[3651]) );
  XOR U6585 ( .A(n2488), .B(n2489), .Z(n2485) );
  ANDN U6586 ( .B(n2490), .A(n2491), .Z(n2488) );
  XNOR U6587 ( .A(b[3650]), .B(n2489), .Z(n2490) );
  XNOR U6588 ( .A(b[3650]), .B(n2491), .Z(c[3650]) );
  XOR U6589 ( .A(n2492), .B(n2493), .Z(n2489) );
  ANDN U6590 ( .B(n2494), .A(n2495), .Z(n2492) );
  XNOR U6591 ( .A(b[3649]), .B(n2493), .Z(n2494) );
  XNOR U6592 ( .A(b[364]), .B(n2496), .Z(c[364]) );
  XNOR U6593 ( .A(b[3649]), .B(n2495), .Z(c[3649]) );
  XOR U6594 ( .A(n2497), .B(n2498), .Z(n2493) );
  ANDN U6595 ( .B(n2499), .A(n2500), .Z(n2497) );
  XNOR U6596 ( .A(b[3648]), .B(n2498), .Z(n2499) );
  XNOR U6597 ( .A(b[3648]), .B(n2500), .Z(c[3648]) );
  XOR U6598 ( .A(n2501), .B(n2502), .Z(n2498) );
  ANDN U6599 ( .B(n2503), .A(n2504), .Z(n2501) );
  XNOR U6600 ( .A(b[3647]), .B(n2502), .Z(n2503) );
  XNOR U6601 ( .A(b[3647]), .B(n2504), .Z(c[3647]) );
  XOR U6602 ( .A(n2505), .B(n2506), .Z(n2502) );
  ANDN U6603 ( .B(n2507), .A(n2508), .Z(n2505) );
  XNOR U6604 ( .A(b[3646]), .B(n2506), .Z(n2507) );
  XNOR U6605 ( .A(b[3646]), .B(n2508), .Z(c[3646]) );
  XOR U6606 ( .A(n2509), .B(n2510), .Z(n2506) );
  ANDN U6607 ( .B(n2511), .A(n2512), .Z(n2509) );
  XNOR U6608 ( .A(b[3645]), .B(n2510), .Z(n2511) );
  XNOR U6609 ( .A(b[3645]), .B(n2512), .Z(c[3645]) );
  XOR U6610 ( .A(n2513), .B(n2514), .Z(n2510) );
  ANDN U6611 ( .B(n2515), .A(n2516), .Z(n2513) );
  XNOR U6612 ( .A(b[3644]), .B(n2514), .Z(n2515) );
  XNOR U6613 ( .A(b[3644]), .B(n2516), .Z(c[3644]) );
  XOR U6614 ( .A(n2517), .B(n2518), .Z(n2514) );
  ANDN U6615 ( .B(n2519), .A(n2520), .Z(n2517) );
  XNOR U6616 ( .A(b[3643]), .B(n2518), .Z(n2519) );
  XNOR U6617 ( .A(b[3643]), .B(n2520), .Z(c[3643]) );
  XOR U6618 ( .A(n2521), .B(n2522), .Z(n2518) );
  ANDN U6619 ( .B(n2523), .A(n2524), .Z(n2521) );
  XNOR U6620 ( .A(b[3642]), .B(n2522), .Z(n2523) );
  XNOR U6621 ( .A(b[3642]), .B(n2524), .Z(c[3642]) );
  XOR U6622 ( .A(n2525), .B(n2526), .Z(n2522) );
  ANDN U6623 ( .B(n2527), .A(n2528), .Z(n2525) );
  XNOR U6624 ( .A(b[3641]), .B(n2526), .Z(n2527) );
  XNOR U6625 ( .A(b[3641]), .B(n2528), .Z(c[3641]) );
  XOR U6626 ( .A(n2529), .B(n2530), .Z(n2526) );
  ANDN U6627 ( .B(n2531), .A(n2532), .Z(n2529) );
  XNOR U6628 ( .A(b[3640]), .B(n2530), .Z(n2531) );
  XNOR U6629 ( .A(b[3640]), .B(n2532), .Z(c[3640]) );
  XOR U6630 ( .A(n2533), .B(n2534), .Z(n2530) );
  ANDN U6631 ( .B(n2535), .A(n2536), .Z(n2533) );
  XNOR U6632 ( .A(b[3639]), .B(n2534), .Z(n2535) );
  XNOR U6633 ( .A(b[363]), .B(n2537), .Z(c[363]) );
  XNOR U6634 ( .A(b[3639]), .B(n2536), .Z(c[3639]) );
  XOR U6635 ( .A(n2538), .B(n2539), .Z(n2534) );
  ANDN U6636 ( .B(n2540), .A(n2541), .Z(n2538) );
  XNOR U6637 ( .A(b[3638]), .B(n2539), .Z(n2540) );
  XNOR U6638 ( .A(b[3638]), .B(n2541), .Z(c[3638]) );
  XOR U6639 ( .A(n2542), .B(n2543), .Z(n2539) );
  ANDN U6640 ( .B(n2544), .A(n2545), .Z(n2542) );
  XNOR U6641 ( .A(b[3637]), .B(n2543), .Z(n2544) );
  XNOR U6642 ( .A(b[3637]), .B(n2545), .Z(c[3637]) );
  XOR U6643 ( .A(n2546), .B(n2547), .Z(n2543) );
  ANDN U6644 ( .B(n2548), .A(n2549), .Z(n2546) );
  XNOR U6645 ( .A(b[3636]), .B(n2547), .Z(n2548) );
  XNOR U6646 ( .A(b[3636]), .B(n2549), .Z(c[3636]) );
  XOR U6647 ( .A(n2550), .B(n2551), .Z(n2547) );
  ANDN U6648 ( .B(n2552), .A(n2553), .Z(n2550) );
  XNOR U6649 ( .A(b[3635]), .B(n2551), .Z(n2552) );
  XNOR U6650 ( .A(b[3635]), .B(n2553), .Z(c[3635]) );
  XOR U6651 ( .A(n2554), .B(n2555), .Z(n2551) );
  ANDN U6652 ( .B(n2556), .A(n2557), .Z(n2554) );
  XNOR U6653 ( .A(b[3634]), .B(n2555), .Z(n2556) );
  XNOR U6654 ( .A(b[3634]), .B(n2557), .Z(c[3634]) );
  XOR U6655 ( .A(n2558), .B(n2559), .Z(n2555) );
  ANDN U6656 ( .B(n2560), .A(n2561), .Z(n2558) );
  XNOR U6657 ( .A(b[3633]), .B(n2559), .Z(n2560) );
  XNOR U6658 ( .A(b[3633]), .B(n2561), .Z(c[3633]) );
  XOR U6659 ( .A(n2562), .B(n2563), .Z(n2559) );
  ANDN U6660 ( .B(n2564), .A(n2565), .Z(n2562) );
  XNOR U6661 ( .A(b[3632]), .B(n2563), .Z(n2564) );
  XNOR U6662 ( .A(b[3632]), .B(n2565), .Z(c[3632]) );
  XOR U6663 ( .A(n2566), .B(n2567), .Z(n2563) );
  ANDN U6664 ( .B(n2568), .A(n2569), .Z(n2566) );
  XNOR U6665 ( .A(b[3631]), .B(n2567), .Z(n2568) );
  XNOR U6666 ( .A(b[3631]), .B(n2569), .Z(c[3631]) );
  XOR U6667 ( .A(n2570), .B(n2571), .Z(n2567) );
  ANDN U6668 ( .B(n2572), .A(n2573), .Z(n2570) );
  XNOR U6669 ( .A(b[3630]), .B(n2571), .Z(n2572) );
  XNOR U6670 ( .A(b[3630]), .B(n2573), .Z(c[3630]) );
  XOR U6671 ( .A(n2574), .B(n2575), .Z(n2571) );
  ANDN U6672 ( .B(n2576), .A(n2577), .Z(n2574) );
  XNOR U6673 ( .A(b[3629]), .B(n2575), .Z(n2576) );
  XNOR U6674 ( .A(b[362]), .B(n2578), .Z(c[362]) );
  XNOR U6675 ( .A(b[3629]), .B(n2577), .Z(c[3629]) );
  XOR U6676 ( .A(n2579), .B(n2580), .Z(n2575) );
  ANDN U6677 ( .B(n2581), .A(n2582), .Z(n2579) );
  XNOR U6678 ( .A(b[3628]), .B(n2580), .Z(n2581) );
  XNOR U6679 ( .A(b[3628]), .B(n2582), .Z(c[3628]) );
  XOR U6680 ( .A(n2583), .B(n2584), .Z(n2580) );
  ANDN U6681 ( .B(n2585), .A(n2586), .Z(n2583) );
  XNOR U6682 ( .A(b[3627]), .B(n2584), .Z(n2585) );
  XNOR U6683 ( .A(b[3627]), .B(n2586), .Z(c[3627]) );
  XOR U6684 ( .A(n2587), .B(n2588), .Z(n2584) );
  ANDN U6685 ( .B(n2589), .A(n2590), .Z(n2587) );
  XNOR U6686 ( .A(b[3626]), .B(n2588), .Z(n2589) );
  XNOR U6687 ( .A(b[3626]), .B(n2590), .Z(c[3626]) );
  XOR U6688 ( .A(n2591), .B(n2592), .Z(n2588) );
  ANDN U6689 ( .B(n2593), .A(n2594), .Z(n2591) );
  XNOR U6690 ( .A(b[3625]), .B(n2592), .Z(n2593) );
  XNOR U6691 ( .A(b[3625]), .B(n2594), .Z(c[3625]) );
  XOR U6692 ( .A(n2595), .B(n2596), .Z(n2592) );
  ANDN U6693 ( .B(n2597), .A(n2598), .Z(n2595) );
  XNOR U6694 ( .A(b[3624]), .B(n2596), .Z(n2597) );
  XNOR U6695 ( .A(b[3624]), .B(n2598), .Z(c[3624]) );
  XOR U6696 ( .A(n2599), .B(n2600), .Z(n2596) );
  ANDN U6697 ( .B(n2601), .A(n2602), .Z(n2599) );
  XNOR U6698 ( .A(b[3623]), .B(n2600), .Z(n2601) );
  XNOR U6699 ( .A(b[3623]), .B(n2602), .Z(c[3623]) );
  XOR U6700 ( .A(n2603), .B(n2604), .Z(n2600) );
  ANDN U6701 ( .B(n2605), .A(n2606), .Z(n2603) );
  XNOR U6702 ( .A(b[3622]), .B(n2604), .Z(n2605) );
  XNOR U6703 ( .A(b[3622]), .B(n2606), .Z(c[3622]) );
  XOR U6704 ( .A(n2607), .B(n2608), .Z(n2604) );
  ANDN U6705 ( .B(n2609), .A(n2610), .Z(n2607) );
  XNOR U6706 ( .A(b[3621]), .B(n2608), .Z(n2609) );
  XNOR U6707 ( .A(b[3621]), .B(n2610), .Z(c[3621]) );
  XOR U6708 ( .A(n2611), .B(n2612), .Z(n2608) );
  ANDN U6709 ( .B(n2613), .A(n2614), .Z(n2611) );
  XNOR U6710 ( .A(b[3620]), .B(n2612), .Z(n2613) );
  XNOR U6711 ( .A(b[3620]), .B(n2614), .Z(c[3620]) );
  XOR U6712 ( .A(n2615), .B(n2616), .Z(n2612) );
  ANDN U6713 ( .B(n2617), .A(n2618), .Z(n2615) );
  XNOR U6714 ( .A(b[3619]), .B(n2616), .Z(n2617) );
  XNOR U6715 ( .A(b[361]), .B(n2619), .Z(c[361]) );
  XNOR U6716 ( .A(b[3619]), .B(n2618), .Z(c[3619]) );
  XOR U6717 ( .A(n2620), .B(n2621), .Z(n2616) );
  ANDN U6718 ( .B(n2622), .A(n2623), .Z(n2620) );
  XNOR U6719 ( .A(b[3618]), .B(n2621), .Z(n2622) );
  XNOR U6720 ( .A(b[3618]), .B(n2623), .Z(c[3618]) );
  XOR U6721 ( .A(n2624), .B(n2625), .Z(n2621) );
  ANDN U6722 ( .B(n2626), .A(n2627), .Z(n2624) );
  XNOR U6723 ( .A(b[3617]), .B(n2625), .Z(n2626) );
  XNOR U6724 ( .A(b[3617]), .B(n2627), .Z(c[3617]) );
  XOR U6725 ( .A(n2628), .B(n2629), .Z(n2625) );
  ANDN U6726 ( .B(n2630), .A(n2631), .Z(n2628) );
  XNOR U6727 ( .A(b[3616]), .B(n2629), .Z(n2630) );
  XNOR U6728 ( .A(b[3616]), .B(n2631), .Z(c[3616]) );
  XOR U6729 ( .A(n2632), .B(n2633), .Z(n2629) );
  ANDN U6730 ( .B(n2634), .A(n2635), .Z(n2632) );
  XNOR U6731 ( .A(b[3615]), .B(n2633), .Z(n2634) );
  XNOR U6732 ( .A(b[3615]), .B(n2635), .Z(c[3615]) );
  XOR U6733 ( .A(n2636), .B(n2637), .Z(n2633) );
  ANDN U6734 ( .B(n2638), .A(n2639), .Z(n2636) );
  XNOR U6735 ( .A(b[3614]), .B(n2637), .Z(n2638) );
  XNOR U6736 ( .A(b[3614]), .B(n2639), .Z(c[3614]) );
  XOR U6737 ( .A(n2640), .B(n2641), .Z(n2637) );
  ANDN U6738 ( .B(n2642), .A(n2643), .Z(n2640) );
  XNOR U6739 ( .A(b[3613]), .B(n2641), .Z(n2642) );
  XNOR U6740 ( .A(b[3613]), .B(n2643), .Z(c[3613]) );
  XOR U6741 ( .A(n2644), .B(n2645), .Z(n2641) );
  ANDN U6742 ( .B(n2646), .A(n2647), .Z(n2644) );
  XNOR U6743 ( .A(b[3612]), .B(n2645), .Z(n2646) );
  XNOR U6744 ( .A(b[3612]), .B(n2647), .Z(c[3612]) );
  XOR U6745 ( .A(n2648), .B(n2649), .Z(n2645) );
  ANDN U6746 ( .B(n2650), .A(n2651), .Z(n2648) );
  XNOR U6747 ( .A(b[3611]), .B(n2649), .Z(n2650) );
  XNOR U6748 ( .A(b[3611]), .B(n2651), .Z(c[3611]) );
  XOR U6749 ( .A(n2652), .B(n2653), .Z(n2649) );
  ANDN U6750 ( .B(n2654), .A(n2655), .Z(n2652) );
  XNOR U6751 ( .A(b[3610]), .B(n2653), .Z(n2654) );
  XNOR U6752 ( .A(b[3610]), .B(n2655), .Z(c[3610]) );
  XOR U6753 ( .A(n2656), .B(n2657), .Z(n2653) );
  ANDN U6754 ( .B(n2658), .A(n2659), .Z(n2656) );
  XNOR U6755 ( .A(b[3609]), .B(n2657), .Z(n2658) );
  XNOR U6756 ( .A(b[360]), .B(n2660), .Z(c[360]) );
  XNOR U6757 ( .A(b[3609]), .B(n2659), .Z(c[3609]) );
  XOR U6758 ( .A(n2661), .B(n2662), .Z(n2657) );
  ANDN U6759 ( .B(n2663), .A(n2664), .Z(n2661) );
  XNOR U6760 ( .A(b[3608]), .B(n2662), .Z(n2663) );
  XNOR U6761 ( .A(b[3608]), .B(n2664), .Z(c[3608]) );
  XOR U6762 ( .A(n2665), .B(n2666), .Z(n2662) );
  ANDN U6763 ( .B(n2667), .A(n2668), .Z(n2665) );
  XNOR U6764 ( .A(b[3607]), .B(n2666), .Z(n2667) );
  XNOR U6765 ( .A(b[3607]), .B(n2668), .Z(c[3607]) );
  XOR U6766 ( .A(n2669), .B(n2670), .Z(n2666) );
  ANDN U6767 ( .B(n2671), .A(n2672), .Z(n2669) );
  XNOR U6768 ( .A(b[3606]), .B(n2670), .Z(n2671) );
  XNOR U6769 ( .A(b[3606]), .B(n2672), .Z(c[3606]) );
  XOR U6770 ( .A(n2673), .B(n2674), .Z(n2670) );
  ANDN U6771 ( .B(n2675), .A(n2676), .Z(n2673) );
  XNOR U6772 ( .A(b[3605]), .B(n2674), .Z(n2675) );
  XNOR U6773 ( .A(b[3605]), .B(n2676), .Z(c[3605]) );
  XOR U6774 ( .A(n2677), .B(n2678), .Z(n2674) );
  ANDN U6775 ( .B(n2679), .A(n2680), .Z(n2677) );
  XNOR U6776 ( .A(b[3604]), .B(n2678), .Z(n2679) );
  XNOR U6777 ( .A(b[3604]), .B(n2680), .Z(c[3604]) );
  XOR U6778 ( .A(n2681), .B(n2682), .Z(n2678) );
  ANDN U6779 ( .B(n2683), .A(n2684), .Z(n2681) );
  XNOR U6780 ( .A(b[3603]), .B(n2682), .Z(n2683) );
  XNOR U6781 ( .A(b[3603]), .B(n2684), .Z(c[3603]) );
  XOR U6782 ( .A(n2685), .B(n2686), .Z(n2682) );
  ANDN U6783 ( .B(n2687), .A(n2688), .Z(n2685) );
  XNOR U6784 ( .A(b[3602]), .B(n2686), .Z(n2687) );
  XNOR U6785 ( .A(b[3602]), .B(n2688), .Z(c[3602]) );
  XOR U6786 ( .A(n2689), .B(n2690), .Z(n2686) );
  ANDN U6787 ( .B(n2691), .A(n2692), .Z(n2689) );
  XNOR U6788 ( .A(b[3601]), .B(n2690), .Z(n2691) );
  XNOR U6789 ( .A(b[3601]), .B(n2692), .Z(c[3601]) );
  XOR U6790 ( .A(n2693), .B(n2694), .Z(n2690) );
  ANDN U6791 ( .B(n2695), .A(n2696), .Z(n2693) );
  XNOR U6792 ( .A(b[3600]), .B(n2694), .Z(n2695) );
  XNOR U6793 ( .A(b[3600]), .B(n2696), .Z(c[3600]) );
  XOR U6794 ( .A(n2697), .B(n2698), .Z(n2694) );
  ANDN U6795 ( .B(n2699), .A(n2700), .Z(n2697) );
  XNOR U6796 ( .A(b[3599]), .B(n2698), .Z(n2699) );
  XNOR U6797 ( .A(b[35]), .B(n2701), .Z(c[35]) );
  XNOR U6798 ( .A(b[359]), .B(n2702), .Z(c[359]) );
  XNOR U6799 ( .A(b[3599]), .B(n2700), .Z(c[3599]) );
  XOR U6800 ( .A(n2703), .B(n2704), .Z(n2698) );
  ANDN U6801 ( .B(n2705), .A(n2706), .Z(n2703) );
  XNOR U6802 ( .A(b[3598]), .B(n2704), .Z(n2705) );
  XNOR U6803 ( .A(b[3598]), .B(n2706), .Z(c[3598]) );
  XOR U6804 ( .A(n2707), .B(n2708), .Z(n2704) );
  ANDN U6805 ( .B(n2709), .A(n2710), .Z(n2707) );
  XNOR U6806 ( .A(b[3597]), .B(n2708), .Z(n2709) );
  XNOR U6807 ( .A(b[3597]), .B(n2710), .Z(c[3597]) );
  XOR U6808 ( .A(n2711), .B(n2712), .Z(n2708) );
  ANDN U6809 ( .B(n2713), .A(n2714), .Z(n2711) );
  XNOR U6810 ( .A(b[3596]), .B(n2712), .Z(n2713) );
  XNOR U6811 ( .A(b[3596]), .B(n2714), .Z(c[3596]) );
  XOR U6812 ( .A(n2715), .B(n2716), .Z(n2712) );
  ANDN U6813 ( .B(n2717), .A(n2718), .Z(n2715) );
  XNOR U6814 ( .A(b[3595]), .B(n2716), .Z(n2717) );
  XNOR U6815 ( .A(b[3595]), .B(n2718), .Z(c[3595]) );
  XOR U6816 ( .A(n2719), .B(n2720), .Z(n2716) );
  ANDN U6817 ( .B(n2721), .A(n2722), .Z(n2719) );
  XNOR U6818 ( .A(b[3594]), .B(n2720), .Z(n2721) );
  XNOR U6819 ( .A(b[3594]), .B(n2722), .Z(c[3594]) );
  XOR U6820 ( .A(n2723), .B(n2724), .Z(n2720) );
  ANDN U6821 ( .B(n2725), .A(n2726), .Z(n2723) );
  XNOR U6822 ( .A(b[3593]), .B(n2724), .Z(n2725) );
  XNOR U6823 ( .A(b[3593]), .B(n2726), .Z(c[3593]) );
  XOR U6824 ( .A(n2727), .B(n2728), .Z(n2724) );
  ANDN U6825 ( .B(n2729), .A(n2730), .Z(n2727) );
  XNOR U6826 ( .A(b[3592]), .B(n2728), .Z(n2729) );
  XNOR U6827 ( .A(b[3592]), .B(n2730), .Z(c[3592]) );
  XOR U6828 ( .A(n2731), .B(n2732), .Z(n2728) );
  ANDN U6829 ( .B(n2733), .A(n2734), .Z(n2731) );
  XNOR U6830 ( .A(b[3591]), .B(n2732), .Z(n2733) );
  XNOR U6831 ( .A(b[3591]), .B(n2734), .Z(c[3591]) );
  XOR U6832 ( .A(n2735), .B(n2736), .Z(n2732) );
  ANDN U6833 ( .B(n2737), .A(n2738), .Z(n2735) );
  XNOR U6834 ( .A(b[3590]), .B(n2736), .Z(n2737) );
  XNOR U6835 ( .A(b[3590]), .B(n2738), .Z(c[3590]) );
  XOR U6836 ( .A(n2739), .B(n2740), .Z(n2736) );
  ANDN U6837 ( .B(n2741), .A(n2742), .Z(n2739) );
  XNOR U6838 ( .A(b[3589]), .B(n2740), .Z(n2741) );
  XNOR U6839 ( .A(b[358]), .B(n2743), .Z(c[358]) );
  XNOR U6840 ( .A(b[3589]), .B(n2742), .Z(c[3589]) );
  XOR U6841 ( .A(n2744), .B(n2745), .Z(n2740) );
  ANDN U6842 ( .B(n2746), .A(n2747), .Z(n2744) );
  XNOR U6843 ( .A(b[3588]), .B(n2745), .Z(n2746) );
  XNOR U6844 ( .A(b[3588]), .B(n2747), .Z(c[3588]) );
  XOR U6845 ( .A(n2748), .B(n2749), .Z(n2745) );
  ANDN U6846 ( .B(n2750), .A(n2751), .Z(n2748) );
  XNOR U6847 ( .A(b[3587]), .B(n2749), .Z(n2750) );
  XNOR U6848 ( .A(b[3587]), .B(n2751), .Z(c[3587]) );
  XOR U6849 ( .A(n2752), .B(n2753), .Z(n2749) );
  ANDN U6850 ( .B(n2754), .A(n2755), .Z(n2752) );
  XNOR U6851 ( .A(b[3586]), .B(n2753), .Z(n2754) );
  XNOR U6852 ( .A(b[3586]), .B(n2755), .Z(c[3586]) );
  XOR U6853 ( .A(n2756), .B(n2757), .Z(n2753) );
  ANDN U6854 ( .B(n2758), .A(n2759), .Z(n2756) );
  XNOR U6855 ( .A(b[3585]), .B(n2757), .Z(n2758) );
  XNOR U6856 ( .A(b[3585]), .B(n2759), .Z(c[3585]) );
  XOR U6857 ( .A(n2760), .B(n2761), .Z(n2757) );
  ANDN U6858 ( .B(n2762), .A(n2763), .Z(n2760) );
  XNOR U6859 ( .A(b[3584]), .B(n2761), .Z(n2762) );
  XNOR U6860 ( .A(b[3584]), .B(n2763), .Z(c[3584]) );
  XOR U6861 ( .A(n2764), .B(n2765), .Z(n2761) );
  ANDN U6862 ( .B(n2766), .A(n2767), .Z(n2764) );
  XNOR U6863 ( .A(b[3583]), .B(n2765), .Z(n2766) );
  XNOR U6864 ( .A(b[3583]), .B(n2767), .Z(c[3583]) );
  XOR U6865 ( .A(n2768), .B(n2769), .Z(n2765) );
  ANDN U6866 ( .B(n2770), .A(n2771), .Z(n2768) );
  XNOR U6867 ( .A(b[3582]), .B(n2769), .Z(n2770) );
  XNOR U6868 ( .A(b[3582]), .B(n2771), .Z(c[3582]) );
  XOR U6869 ( .A(n2772), .B(n2773), .Z(n2769) );
  ANDN U6870 ( .B(n2774), .A(n2775), .Z(n2772) );
  XNOR U6871 ( .A(b[3581]), .B(n2773), .Z(n2774) );
  XNOR U6872 ( .A(b[3581]), .B(n2775), .Z(c[3581]) );
  XOR U6873 ( .A(n2776), .B(n2777), .Z(n2773) );
  ANDN U6874 ( .B(n2778), .A(n2779), .Z(n2776) );
  XNOR U6875 ( .A(b[3580]), .B(n2777), .Z(n2778) );
  XNOR U6876 ( .A(b[3580]), .B(n2779), .Z(c[3580]) );
  XOR U6877 ( .A(n2780), .B(n2781), .Z(n2777) );
  ANDN U6878 ( .B(n2782), .A(n2783), .Z(n2780) );
  XNOR U6879 ( .A(b[3579]), .B(n2781), .Z(n2782) );
  XNOR U6880 ( .A(b[357]), .B(n2784), .Z(c[357]) );
  XNOR U6881 ( .A(b[3579]), .B(n2783), .Z(c[3579]) );
  XOR U6882 ( .A(n2785), .B(n2786), .Z(n2781) );
  ANDN U6883 ( .B(n2787), .A(n2788), .Z(n2785) );
  XNOR U6884 ( .A(b[3578]), .B(n2786), .Z(n2787) );
  XNOR U6885 ( .A(b[3578]), .B(n2788), .Z(c[3578]) );
  XOR U6886 ( .A(n2789), .B(n2790), .Z(n2786) );
  ANDN U6887 ( .B(n2791), .A(n2792), .Z(n2789) );
  XNOR U6888 ( .A(b[3577]), .B(n2790), .Z(n2791) );
  XNOR U6889 ( .A(b[3577]), .B(n2792), .Z(c[3577]) );
  XOR U6890 ( .A(n2793), .B(n2794), .Z(n2790) );
  ANDN U6891 ( .B(n2795), .A(n2796), .Z(n2793) );
  XNOR U6892 ( .A(b[3576]), .B(n2794), .Z(n2795) );
  XNOR U6893 ( .A(b[3576]), .B(n2796), .Z(c[3576]) );
  XOR U6894 ( .A(n2797), .B(n2798), .Z(n2794) );
  ANDN U6895 ( .B(n2799), .A(n2800), .Z(n2797) );
  XNOR U6896 ( .A(b[3575]), .B(n2798), .Z(n2799) );
  XNOR U6897 ( .A(b[3575]), .B(n2800), .Z(c[3575]) );
  XOR U6898 ( .A(n2801), .B(n2802), .Z(n2798) );
  ANDN U6899 ( .B(n2803), .A(n2804), .Z(n2801) );
  XNOR U6900 ( .A(b[3574]), .B(n2802), .Z(n2803) );
  XNOR U6901 ( .A(b[3574]), .B(n2804), .Z(c[3574]) );
  XOR U6902 ( .A(n2805), .B(n2806), .Z(n2802) );
  ANDN U6903 ( .B(n2807), .A(n2808), .Z(n2805) );
  XNOR U6904 ( .A(b[3573]), .B(n2806), .Z(n2807) );
  XNOR U6905 ( .A(b[3573]), .B(n2808), .Z(c[3573]) );
  XOR U6906 ( .A(n2809), .B(n2810), .Z(n2806) );
  ANDN U6907 ( .B(n2811), .A(n2812), .Z(n2809) );
  XNOR U6908 ( .A(b[3572]), .B(n2810), .Z(n2811) );
  XNOR U6909 ( .A(b[3572]), .B(n2812), .Z(c[3572]) );
  XOR U6910 ( .A(n2813), .B(n2814), .Z(n2810) );
  ANDN U6911 ( .B(n2815), .A(n2816), .Z(n2813) );
  XNOR U6912 ( .A(b[3571]), .B(n2814), .Z(n2815) );
  XNOR U6913 ( .A(b[3571]), .B(n2816), .Z(c[3571]) );
  XOR U6914 ( .A(n2817), .B(n2818), .Z(n2814) );
  ANDN U6915 ( .B(n2819), .A(n2820), .Z(n2817) );
  XNOR U6916 ( .A(b[3570]), .B(n2818), .Z(n2819) );
  XNOR U6917 ( .A(b[3570]), .B(n2820), .Z(c[3570]) );
  XOR U6918 ( .A(n2821), .B(n2822), .Z(n2818) );
  ANDN U6919 ( .B(n2823), .A(n2824), .Z(n2821) );
  XNOR U6920 ( .A(b[3569]), .B(n2822), .Z(n2823) );
  XNOR U6921 ( .A(b[356]), .B(n2825), .Z(c[356]) );
  XNOR U6922 ( .A(b[3569]), .B(n2824), .Z(c[3569]) );
  XOR U6923 ( .A(n2826), .B(n2827), .Z(n2822) );
  ANDN U6924 ( .B(n2828), .A(n2829), .Z(n2826) );
  XNOR U6925 ( .A(b[3568]), .B(n2827), .Z(n2828) );
  XNOR U6926 ( .A(b[3568]), .B(n2829), .Z(c[3568]) );
  XOR U6927 ( .A(n2830), .B(n2831), .Z(n2827) );
  ANDN U6928 ( .B(n2832), .A(n2833), .Z(n2830) );
  XNOR U6929 ( .A(b[3567]), .B(n2831), .Z(n2832) );
  XNOR U6930 ( .A(b[3567]), .B(n2833), .Z(c[3567]) );
  XOR U6931 ( .A(n2834), .B(n2835), .Z(n2831) );
  ANDN U6932 ( .B(n2836), .A(n2837), .Z(n2834) );
  XNOR U6933 ( .A(b[3566]), .B(n2835), .Z(n2836) );
  XNOR U6934 ( .A(b[3566]), .B(n2837), .Z(c[3566]) );
  XOR U6935 ( .A(n2838), .B(n2839), .Z(n2835) );
  ANDN U6936 ( .B(n2840), .A(n2841), .Z(n2838) );
  XNOR U6937 ( .A(b[3565]), .B(n2839), .Z(n2840) );
  XNOR U6938 ( .A(b[3565]), .B(n2841), .Z(c[3565]) );
  XOR U6939 ( .A(n2842), .B(n2843), .Z(n2839) );
  ANDN U6940 ( .B(n2844), .A(n2845), .Z(n2842) );
  XNOR U6941 ( .A(b[3564]), .B(n2843), .Z(n2844) );
  XNOR U6942 ( .A(b[3564]), .B(n2845), .Z(c[3564]) );
  XOR U6943 ( .A(n2846), .B(n2847), .Z(n2843) );
  ANDN U6944 ( .B(n2848), .A(n2849), .Z(n2846) );
  XNOR U6945 ( .A(b[3563]), .B(n2847), .Z(n2848) );
  XNOR U6946 ( .A(b[3563]), .B(n2849), .Z(c[3563]) );
  XOR U6947 ( .A(n2850), .B(n2851), .Z(n2847) );
  ANDN U6948 ( .B(n2852), .A(n2853), .Z(n2850) );
  XNOR U6949 ( .A(b[3562]), .B(n2851), .Z(n2852) );
  XNOR U6950 ( .A(b[3562]), .B(n2853), .Z(c[3562]) );
  XOR U6951 ( .A(n2854), .B(n2855), .Z(n2851) );
  ANDN U6952 ( .B(n2856), .A(n2857), .Z(n2854) );
  XNOR U6953 ( .A(b[3561]), .B(n2855), .Z(n2856) );
  XNOR U6954 ( .A(b[3561]), .B(n2857), .Z(c[3561]) );
  XOR U6955 ( .A(n2858), .B(n2859), .Z(n2855) );
  ANDN U6956 ( .B(n2860), .A(n2861), .Z(n2858) );
  XNOR U6957 ( .A(b[3560]), .B(n2859), .Z(n2860) );
  XNOR U6958 ( .A(b[3560]), .B(n2861), .Z(c[3560]) );
  XOR U6959 ( .A(n2862), .B(n2863), .Z(n2859) );
  ANDN U6960 ( .B(n2864), .A(n2865), .Z(n2862) );
  XNOR U6961 ( .A(b[3559]), .B(n2863), .Z(n2864) );
  XNOR U6962 ( .A(b[355]), .B(n2866), .Z(c[355]) );
  XNOR U6963 ( .A(b[3559]), .B(n2865), .Z(c[3559]) );
  XOR U6964 ( .A(n2867), .B(n2868), .Z(n2863) );
  ANDN U6965 ( .B(n2869), .A(n2870), .Z(n2867) );
  XNOR U6966 ( .A(b[3558]), .B(n2868), .Z(n2869) );
  XNOR U6967 ( .A(b[3558]), .B(n2870), .Z(c[3558]) );
  XOR U6968 ( .A(n2871), .B(n2872), .Z(n2868) );
  ANDN U6969 ( .B(n2873), .A(n2874), .Z(n2871) );
  XNOR U6970 ( .A(b[3557]), .B(n2872), .Z(n2873) );
  XNOR U6971 ( .A(b[3557]), .B(n2874), .Z(c[3557]) );
  XOR U6972 ( .A(n2875), .B(n2876), .Z(n2872) );
  ANDN U6973 ( .B(n2877), .A(n2878), .Z(n2875) );
  XNOR U6974 ( .A(b[3556]), .B(n2876), .Z(n2877) );
  XNOR U6975 ( .A(b[3556]), .B(n2878), .Z(c[3556]) );
  XOR U6976 ( .A(n2879), .B(n2880), .Z(n2876) );
  ANDN U6977 ( .B(n2881), .A(n2882), .Z(n2879) );
  XNOR U6978 ( .A(b[3555]), .B(n2880), .Z(n2881) );
  XNOR U6979 ( .A(b[3555]), .B(n2882), .Z(c[3555]) );
  XOR U6980 ( .A(n2883), .B(n2884), .Z(n2880) );
  ANDN U6981 ( .B(n2885), .A(n2886), .Z(n2883) );
  XNOR U6982 ( .A(b[3554]), .B(n2884), .Z(n2885) );
  XNOR U6983 ( .A(b[3554]), .B(n2886), .Z(c[3554]) );
  XOR U6984 ( .A(n2887), .B(n2888), .Z(n2884) );
  ANDN U6985 ( .B(n2889), .A(n2890), .Z(n2887) );
  XNOR U6986 ( .A(b[3553]), .B(n2888), .Z(n2889) );
  XNOR U6987 ( .A(b[3553]), .B(n2890), .Z(c[3553]) );
  XOR U6988 ( .A(n2891), .B(n2892), .Z(n2888) );
  ANDN U6989 ( .B(n2893), .A(n2894), .Z(n2891) );
  XNOR U6990 ( .A(b[3552]), .B(n2892), .Z(n2893) );
  XNOR U6991 ( .A(b[3552]), .B(n2894), .Z(c[3552]) );
  XOR U6992 ( .A(n2895), .B(n2896), .Z(n2892) );
  ANDN U6993 ( .B(n2897), .A(n2898), .Z(n2895) );
  XNOR U6994 ( .A(b[3551]), .B(n2896), .Z(n2897) );
  XNOR U6995 ( .A(b[3551]), .B(n2898), .Z(c[3551]) );
  XOR U6996 ( .A(n2899), .B(n2900), .Z(n2896) );
  ANDN U6997 ( .B(n2901), .A(n2902), .Z(n2899) );
  XNOR U6998 ( .A(b[3550]), .B(n2900), .Z(n2901) );
  XNOR U6999 ( .A(b[3550]), .B(n2902), .Z(c[3550]) );
  XOR U7000 ( .A(n2903), .B(n2904), .Z(n2900) );
  ANDN U7001 ( .B(n2905), .A(n2906), .Z(n2903) );
  XNOR U7002 ( .A(b[3549]), .B(n2904), .Z(n2905) );
  XNOR U7003 ( .A(b[354]), .B(n2907), .Z(c[354]) );
  XNOR U7004 ( .A(b[3549]), .B(n2906), .Z(c[3549]) );
  XOR U7005 ( .A(n2908), .B(n2909), .Z(n2904) );
  ANDN U7006 ( .B(n2910), .A(n2911), .Z(n2908) );
  XNOR U7007 ( .A(b[3548]), .B(n2909), .Z(n2910) );
  XNOR U7008 ( .A(b[3548]), .B(n2911), .Z(c[3548]) );
  XOR U7009 ( .A(n2912), .B(n2913), .Z(n2909) );
  ANDN U7010 ( .B(n2914), .A(n2915), .Z(n2912) );
  XNOR U7011 ( .A(b[3547]), .B(n2913), .Z(n2914) );
  XNOR U7012 ( .A(b[3547]), .B(n2915), .Z(c[3547]) );
  XOR U7013 ( .A(n2916), .B(n2917), .Z(n2913) );
  ANDN U7014 ( .B(n2918), .A(n2919), .Z(n2916) );
  XNOR U7015 ( .A(b[3546]), .B(n2917), .Z(n2918) );
  XNOR U7016 ( .A(b[3546]), .B(n2919), .Z(c[3546]) );
  XOR U7017 ( .A(n2920), .B(n2921), .Z(n2917) );
  ANDN U7018 ( .B(n2922), .A(n2923), .Z(n2920) );
  XNOR U7019 ( .A(b[3545]), .B(n2921), .Z(n2922) );
  XNOR U7020 ( .A(b[3545]), .B(n2923), .Z(c[3545]) );
  XOR U7021 ( .A(n2924), .B(n2925), .Z(n2921) );
  ANDN U7022 ( .B(n2926), .A(n2927), .Z(n2924) );
  XNOR U7023 ( .A(b[3544]), .B(n2925), .Z(n2926) );
  XNOR U7024 ( .A(b[3544]), .B(n2927), .Z(c[3544]) );
  XOR U7025 ( .A(n2928), .B(n2929), .Z(n2925) );
  ANDN U7026 ( .B(n2930), .A(n2931), .Z(n2928) );
  XNOR U7027 ( .A(b[3543]), .B(n2929), .Z(n2930) );
  XNOR U7028 ( .A(b[3543]), .B(n2931), .Z(c[3543]) );
  XOR U7029 ( .A(n2932), .B(n2933), .Z(n2929) );
  ANDN U7030 ( .B(n2934), .A(n2935), .Z(n2932) );
  XNOR U7031 ( .A(b[3542]), .B(n2933), .Z(n2934) );
  XNOR U7032 ( .A(b[3542]), .B(n2935), .Z(c[3542]) );
  XOR U7033 ( .A(n2936), .B(n2937), .Z(n2933) );
  ANDN U7034 ( .B(n2938), .A(n2939), .Z(n2936) );
  XNOR U7035 ( .A(b[3541]), .B(n2937), .Z(n2938) );
  XNOR U7036 ( .A(b[3541]), .B(n2939), .Z(c[3541]) );
  XOR U7037 ( .A(n2940), .B(n2941), .Z(n2937) );
  ANDN U7038 ( .B(n2942), .A(n2943), .Z(n2940) );
  XNOR U7039 ( .A(b[3540]), .B(n2941), .Z(n2942) );
  XNOR U7040 ( .A(b[3540]), .B(n2943), .Z(c[3540]) );
  XOR U7041 ( .A(n2944), .B(n2945), .Z(n2941) );
  ANDN U7042 ( .B(n2946), .A(n2947), .Z(n2944) );
  XNOR U7043 ( .A(b[3539]), .B(n2945), .Z(n2946) );
  XNOR U7044 ( .A(b[353]), .B(n2948), .Z(c[353]) );
  XNOR U7045 ( .A(b[3539]), .B(n2947), .Z(c[3539]) );
  XOR U7046 ( .A(n2949), .B(n2950), .Z(n2945) );
  ANDN U7047 ( .B(n2951), .A(n2952), .Z(n2949) );
  XNOR U7048 ( .A(b[3538]), .B(n2950), .Z(n2951) );
  XNOR U7049 ( .A(b[3538]), .B(n2952), .Z(c[3538]) );
  XOR U7050 ( .A(n2953), .B(n2954), .Z(n2950) );
  ANDN U7051 ( .B(n2955), .A(n2956), .Z(n2953) );
  XNOR U7052 ( .A(b[3537]), .B(n2954), .Z(n2955) );
  XNOR U7053 ( .A(b[3537]), .B(n2956), .Z(c[3537]) );
  XOR U7054 ( .A(n2957), .B(n2958), .Z(n2954) );
  ANDN U7055 ( .B(n2959), .A(n2960), .Z(n2957) );
  XNOR U7056 ( .A(b[3536]), .B(n2958), .Z(n2959) );
  XNOR U7057 ( .A(b[3536]), .B(n2960), .Z(c[3536]) );
  XOR U7058 ( .A(n2961), .B(n2962), .Z(n2958) );
  ANDN U7059 ( .B(n2963), .A(n2964), .Z(n2961) );
  XNOR U7060 ( .A(b[3535]), .B(n2962), .Z(n2963) );
  XNOR U7061 ( .A(b[3535]), .B(n2964), .Z(c[3535]) );
  XOR U7062 ( .A(n2965), .B(n2966), .Z(n2962) );
  ANDN U7063 ( .B(n2967), .A(n2968), .Z(n2965) );
  XNOR U7064 ( .A(b[3534]), .B(n2966), .Z(n2967) );
  XNOR U7065 ( .A(b[3534]), .B(n2968), .Z(c[3534]) );
  XOR U7066 ( .A(n2969), .B(n2970), .Z(n2966) );
  ANDN U7067 ( .B(n2971), .A(n2972), .Z(n2969) );
  XNOR U7068 ( .A(b[3533]), .B(n2970), .Z(n2971) );
  XNOR U7069 ( .A(b[3533]), .B(n2972), .Z(c[3533]) );
  XOR U7070 ( .A(n2973), .B(n2974), .Z(n2970) );
  ANDN U7071 ( .B(n2975), .A(n2976), .Z(n2973) );
  XNOR U7072 ( .A(b[3532]), .B(n2974), .Z(n2975) );
  XNOR U7073 ( .A(b[3532]), .B(n2976), .Z(c[3532]) );
  XOR U7074 ( .A(n2977), .B(n2978), .Z(n2974) );
  ANDN U7075 ( .B(n2979), .A(n2980), .Z(n2977) );
  XNOR U7076 ( .A(b[3531]), .B(n2978), .Z(n2979) );
  XNOR U7077 ( .A(b[3531]), .B(n2980), .Z(c[3531]) );
  XOR U7078 ( .A(n2981), .B(n2982), .Z(n2978) );
  ANDN U7079 ( .B(n2983), .A(n2984), .Z(n2981) );
  XNOR U7080 ( .A(b[3530]), .B(n2982), .Z(n2983) );
  XNOR U7081 ( .A(b[3530]), .B(n2984), .Z(c[3530]) );
  XOR U7082 ( .A(n2985), .B(n2986), .Z(n2982) );
  ANDN U7083 ( .B(n2987), .A(n2988), .Z(n2985) );
  XNOR U7084 ( .A(b[3529]), .B(n2986), .Z(n2987) );
  XNOR U7085 ( .A(b[352]), .B(n2989), .Z(c[352]) );
  XNOR U7086 ( .A(b[3529]), .B(n2988), .Z(c[3529]) );
  XOR U7087 ( .A(n2990), .B(n2991), .Z(n2986) );
  ANDN U7088 ( .B(n2992), .A(n2993), .Z(n2990) );
  XNOR U7089 ( .A(b[3528]), .B(n2991), .Z(n2992) );
  XNOR U7090 ( .A(b[3528]), .B(n2993), .Z(c[3528]) );
  XOR U7091 ( .A(n2994), .B(n2995), .Z(n2991) );
  ANDN U7092 ( .B(n2996), .A(n2997), .Z(n2994) );
  XNOR U7093 ( .A(b[3527]), .B(n2995), .Z(n2996) );
  XNOR U7094 ( .A(b[3527]), .B(n2997), .Z(c[3527]) );
  XOR U7095 ( .A(n2998), .B(n2999), .Z(n2995) );
  ANDN U7096 ( .B(n3000), .A(n3001), .Z(n2998) );
  XNOR U7097 ( .A(b[3526]), .B(n2999), .Z(n3000) );
  XNOR U7098 ( .A(b[3526]), .B(n3001), .Z(c[3526]) );
  XOR U7099 ( .A(n3002), .B(n3003), .Z(n2999) );
  ANDN U7100 ( .B(n3004), .A(n3005), .Z(n3002) );
  XNOR U7101 ( .A(b[3525]), .B(n3003), .Z(n3004) );
  XNOR U7102 ( .A(b[3525]), .B(n3005), .Z(c[3525]) );
  XOR U7103 ( .A(n3006), .B(n3007), .Z(n3003) );
  ANDN U7104 ( .B(n3008), .A(n3009), .Z(n3006) );
  XNOR U7105 ( .A(b[3524]), .B(n3007), .Z(n3008) );
  XNOR U7106 ( .A(b[3524]), .B(n3009), .Z(c[3524]) );
  XOR U7107 ( .A(n3010), .B(n3011), .Z(n3007) );
  ANDN U7108 ( .B(n3012), .A(n3013), .Z(n3010) );
  XNOR U7109 ( .A(b[3523]), .B(n3011), .Z(n3012) );
  XNOR U7110 ( .A(b[3523]), .B(n3013), .Z(c[3523]) );
  XOR U7111 ( .A(n3014), .B(n3015), .Z(n3011) );
  ANDN U7112 ( .B(n3016), .A(n3017), .Z(n3014) );
  XNOR U7113 ( .A(b[3522]), .B(n3015), .Z(n3016) );
  XNOR U7114 ( .A(b[3522]), .B(n3017), .Z(c[3522]) );
  XOR U7115 ( .A(n3018), .B(n3019), .Z(n3015) );
  ANDN U7116 ( .B(n3020), .A(n3021), .Z(n3018) );
  XNOR U7117 ( .A(b[3521]), .B(n3019), .Z(n3020) );
  XNOR U7118 ( .A(b[3521]), .B(n3021), .Z(c[3521]) );
  XOR U7119 ( .A(n3022), .B(n3023), .Z(n3019) );
  ANDN U7120 ( .B(n3024), .A(n3025), .Z(n3022) );
  XNOR U7121 ( .A(b[3520]), .B(n3023), .Z(n3024) );
  XNOR U7122 ( .A(b[3520]), .B(n3025), .Z(c[3520]) );
  XOR U7123 ( .A(n3026), .B(n3027), .Z(n3023) );
  ANDN U7124 ( .B(n3028), .A(n3029), .Z(n3026) );
  XNOR U7125 ( .A(b[3519]), .B(n3027), .Z(n3028) );
  XNOR U7126 ( .A(b[351]), .B(n3030), .Z(c[351]) );
  XNOR U7127 ( .A(b[3519]), .B(n3029), .Z(c[3519]) );
  XOR U7128 ( .A(n3031), .B(n3032), .Z(n3027) );
  ANDN U7129 ( .B(n3033), .A(n3034), .Z(n3031) );
  XNOR U7130 ( .A(b[3518]), .B(n3032), .Z(n3033) );
  XNOR U7131 ( .A(b[3518]), .B(n3034), .Z(c[3518]) );
  XOR U7132 ( .A(n3035), .B(n3036), .Z(n3032) );
  ANDN U7133 ( .B(n3037), .A(n3038), .Z(n3035) );
  XNOR U7134 ( .A(b[3517]), .B(n3036), .Z(n3037) );
  XNOR U7135 ( .A(b[3517]), .B(n3038), .Z(c[3517]) );
  XOR U7136 ( .A(n3039), .B(n3040), .Z(n3036) );
  ANDN U7137 ( .B(n3041), .A(n3042), .Z(n3039) );
  XNOR U7138 ( .A(b[3516]), .B(n3040), .Z(n3041) );
  XNOR U7139 ( .A(b[3516]), .B(n3042), .Z(c[3516]) );
  XOR U7140 ( .A(n3043), .B(n3044), .Z(n3040) );
  ANDN U7141 ( .B(n3045), .A(n3046), .Z(n3043) );
  XNOR U7142 ( .A(b[3515]), .B(n3044), .Z(n3045) );
  XNOR U7143 ( .A(b[3515]), .B(n3046), .Z(c[3515]) );
  XOR U7144 ( .A(n3047), .B(n3048), .Z(n3044) );
  ANDN U7145 ( .B(n3049), .A(n3050), .Z(n3047) );
  XNOR U7146 ( .A(b[3514]), .B(n3048), .Z(n3049) );
  XNOR U7147 ( .A(b[3514]), .B(n3050), .Z(c[3514]) );
  XOR U7148 ( .A(n3051), .B(n3052), .Z(n3048) );
  ANDN U7149 ( .B(n3053), .A(n3054), .Z(n3051) );
  XNOR U7150 ( .A(b[3513]), .B(n3052), .Z(n3053) );
  XNOR U7151 ( .A(b[3513]), .B(n3054), .Z(c[3513]) );
  XOR U7152 ( .A(n3055), .B(n3056), .Z(n3052) );
  ANDN U7153 ( .B(n3057), .A(n3058), .Z(n3055) );
  XNOR U7154 ( .A(b[3512]), .B(n3056), .Z(n3057) );
  XNOR U7155 ( .A(b[3512]), .B(n3058), .Z(c[3512]) );
  XOR U7156 ( .A(n3059), .B(n3060), .Z(n3056) );
  ANDN U7157 ( .B(n3061), .A(n3062), .Z(n3059) );
  XNOR U7158 ( .A(b[3511]), .B(n3060), .Z(n3061) );
  XNOR U7159 ( .A(b[3511]), .B(n3062), .Z(c[3511]) );
  XOR U7160 ( .A(n3063), .B(n3064), .Z(n3060) );
  ANDN U7161 ( .B(n3065), .A(n3066), .Z(n3063) );
  XNOR U7162 ( .A(b[3510]), .B(n3064), .Z(n3065) );
  XNOR U7163 ( .A(b[3510]), .B(n3066), .Z(c[3510]) );
  XOR U7164 ( .A(n3067), .B(n3068), .Z(n3064) );
  ANDN U7165 ( .B(n3069), .A(n3070), .Z(n3067) );
  XNOR U7166 ( .A(b[3509]), .B(n3068), .Z(n3069) );
  XNOR U7167 ( .A(b[350]), .B(n3071), .Z(c[350]) );
  XNOR U7168 ( .A(b[3509]), .B(n3070), .Z(c[3509]) );
  XOR U7169 ( .A(n3072), .B(n3073), .Z(n3068) );
  ANDN U7170 ( .B(n3074), .A(n3075), .Z(n3072) );
  XNOR U7171 ( .A(b[3508]), .B(n3073), .Z(n3074) );
  XNOR U7172 ( .A(b[3508]), .B(n3075), .Z(c[3508]) );
  XOR U7173 ( .A(n3076), .B(n3077), .Z(n3073) );
  ANDN U7174 ( .B(n3078), .A(n3079), .Z(n3076) );
  XNOR U7175 ( .A(b[3507]), .B(n3077), .Z(n3078) );
  XNOR U7176 ( .A(b[3507]), .B(n3079), .Z(c[3507]) );
  XOR U7177 ( .A(n3080), .B(n3081), .Z(n3077) );
  ANDN U7178 ( .B(n3082), .A(n3083), .Z(n3080) );
  XNOR U7179 ( .A(b[3506]), .B(n3081), .Z(n3082) );
  XNOR U7180 ( .A(b[3506]), .B(n3083), .Z(c[3506]) );
  XOR U7181 ( .A(n3084), .B(n3085), .Z(n3081) );
  ANDN U7182 ( .B(n3086), .A(n3087), .Z(n3084) );
  XNOR U7183 ( .A(b[3505]), .B(n3085), .Z(n3086) );
  XNOR U7184 ( .A(b[3505]), .B(n3087), .Z(c[3505]) );
  XOR U7185 ( .A(n3088), .B(n3089), .Z(n3085) );
  ANDN U7186 ( .B(n3090), .A(n3091), .Z(n3088) );
  XNOR U7187 ( .A(b[3504]), .B(n3089), .Z(n3090) );
  XNOR U7188 ( .A(b[3504]), .B(n3091), .Z(c[3504]) );
  XOR U7189 ( .A(n3092), .B(n3093), .Z(n3089) );
  ANDN U7190 ( .B(n3094), .A(n3095), .Z(n3092) );
  XNOR U7191 ( .A(b[3503]), .B(n3093), .Z(n3094) );
  XNOR U7192 ( .A(b[3503]), .B(n3095), .Z(c[3503]) );
  XOR U7193 ( .A(n3096), .B(n3097), .Z(n3093) );
  ANDN U7194 ( .B(n3098), .A(n3099), .Z(n3096) );
  XNOR U7195 ( .A(b[3502]), .B(n3097), .Z(n3098) );
  XNOR U7196 ( .A(b[3502]), .B(n3099), .Z(c[3502]) );
  XOR U7197 ( .A(n3100), .B(n3101), .Z(n3097) );
  ANDN U7198 ( .B(n3102), .A(n3103), .Z(n3100) );
  XNOR U7199 ( .A(b[3501]), .B(n3101), .Z(n3102) );
  XNOR U7200 ( .A(b[3501]), .B(n3103), .Z(c[3501]) );
  XOR U7201 ( .A(n3104), .B(n3105), .Z(n3101) );
  ANDN U7202 ( .B(n3106), .A(n3107), .Z(n3104) );
  XNOR U7203 ( .A(b[3500]), .B(n3105), .Z(n3106) );
  XNOR U7204 ( .A(b[3500]), .B(n3107), .Z(c[3500]) );
  XOR U7205 ( .A(n3108), .B(n3109), .Z(n3105) );
  ANDN U7206 ( .B(n3110), .A(n3111), .Z(n3108) );
  XNOR U7207 ( .A(b[3499]), .B(n3109), .Z(n3110) );
  XNOR U7208 ( .A(b[34]), .B(n3112), .Z(c[34]) );
  XNOR U7209 ( .A(b[349]), .B(n3113), .Z(c[349]) );
  XNOR U7210 ( .A(b[3499]), .B(n3111), .Z(c[3499]) );
  XOR U7211 ( .A(n3114), .B(n3115), .Z(n3109) );
  ANDN U7212 ( .B(n3116), .A(n3117), .Z(n3114) );
  XNOR U7213 ( .A(b[3498]), .B(n3115), .Z(n3116) );
  XNOR U7214 ( .A(b[3498]), .B(n3117), .Z(c[3498]) );
  XOR U7215 ( .A(n3118), .B(n3119), .Z(n3115) );
  ANDN U7216 ( .B(n3120), .A(n3121), .Z(n3118) );
  XNOR U7217 ( .A(b[3497]), .B(n3119), .Z(n3120) );
  XNOR U7218 ( .A(b[3497]), .B(n3121), .Z(c[3497]) );
  XOR U7219 ( .A(n3122), .B(n3123), .Z(n3119) );
  ANDN U7220 ( .B(n3124), .A(n3125), .Z(n3122) );
  XNOR U7221 ( .A(b[3496]), .B(n3123), .Z(n3124) );
  XNOR U7222 ( .A(b[3496]), .B(n3125), .Z(c[3496]) );
  XOR U7223 ( .A(n3126), .B(n3127), .Z(n3123) );
  ANDN U7224 ( .B(n3128), .A(n3129), .Z(n3126) );
  XNOR U7225 ( .A(b[3495]), .B(n3127), .Z(n3128) );
  XNOR U7226 ( .A(b[3495]), .B(n3129), .Z(c[3495]) );
  XOR U7227 ( .A(n3130), .B(n3131), .Z(n3127) );
  ANDN U7228 ( .B(n3132), .A(n3133), .Z(n3130) );
  XNOR U7229 ( .A(b[3494]), .B(n3131), .Z(n3132) );
  XNOR U7230 ( .A(b[3494]), .B(n3133), .Z(c[3494]) );
  XOR U7231 ( .A(n3134), .B(n3135), .Z(n3131) );
  ANDN U7232 ( .B(n3136), .A(n3137), .Z(n3134) );
  XNOR U7233 ( .A(b[3493]), .B(n3135), .Z(n3136) );
  XNOR U7234 ( .A(b[3493]), .B(n3137), .Z(c[3493]) );
  XOR U7235 ( .A(n3138), .B(n3139), .Z(n3135) );
  ANDN U7236 ( .B(n3140), .A(n3141), .Z(n3138) );
  XNOR U7237 ( .A(b[3492]), .B(n3139), .Z(n3140) );
  XNOR U7238 ( .A(b[3492]), .B(n3141), .Z(c[3492]) );
  XOR U7239 ( .A(n3142), .B(n3143), .Z(n3139) );
  ANDN U7240 ( .B(n3144), .A(n3145), .Z(n3142) );
  XNOR U7241 ( .A(b[3491]), .B(n3143), .Z(n3144) );
  XNOR U7242 ( .A(b[3491]), .B(n3145), .Z(c[3491]) );
  XOR U7243 ( .A(n3146), .B(n3147), .Z(n3143) );
  ANDN U7244 ( .B(n3148), .A(n3149), .Z(n3146) );
  XNOR U7245 ( .A(b[3490]), .B(n3147), .Z(n3148) );
  XNOR U7246 ( .A(b[3490]), .B(n3149), .Z(c[3490]) );
  XOR U7247 ( .A(n3150), .B(n3151), .Z(n3147) );
  ANDN U7248 ( .B(n3152), .A(n3153), .Z(n3150) );
  XNOR U7249 ( .A(b[3489]), .B(n3151), .Z(n3152) );
  XNOR U7250 ( .A(b[348]), .B(n3154), .Z(c[348]) );
  XNOR U7251 ( .A(b[3489]), .B(n3153), .Z(c[3489]) );
  XOR U7252 ( .A(n3155), .B(n3156), .Z(n3151) );
  ANDN U7253 ( .B(n3157), .A(n3158), .Z(n3155) );
  XNOR U7254 ( .A(b[3488]), .B(n3156), .Z(n3157) );
  XNOR U7255 ( .A(b[3488]), .B(n3158), .Z(c[3488]) );
  XOR U7256 ( .A(n3159), .B(n3160), .Z(n3156) );
  ANDN U7257 ( .B(n3161), .A(n3162), .Z(n3159) );
  XNOR U7258 ( .A(b[3487]), .B(n3160), .Z(n3161) );
  XNOR U7259 ( .A(b[3487]), .B(n3162), .Z(c[3487]) );
  XOR U7260 ( .A(n3163), .B(n3164), .Z(n3160) );
  ANDN U7261 ( .B(n3165), .A(n3166), .Z(n3163) );
  XNOR U7262 ( .A(b[3486]), .B(n3164), .Z(n3165) );
  XNOR U7263 ( .A(b[3486]), .B(n3166), .Z(c[3486]) );
  XOR U7264 ( .A(n3167), .B(n3168), .Z(n3164) );
  ANDN U7265 ( .B(n3169), .A(n3170), .Z(n3167) );
  XNOR U7266 ( .A(b[3485]), .B(n3168), .Z(n3169) );
  XNOR U7267 ( .A(b[3485]), .B(n3170), .Z(c[3485]) );
  XOR U7268 ( .A(n3171), .B(n3172), .Z(n3168) );
  ANDN U7269 ( .B(n3173), .A(n3174), .Z(n3171) );
  XNOR U7270 ( .A(b[3484]), .B(n3172), .Z(n3173) );
  XNOR U7271 ( .A(b[3484]), .B(n3174), .Z(c[3484]) );
  XOR U7272 ( .A(n3175), .B(n3176), .Z(n3172) );
  ANDN U7273 ( .B(n3177), .A(n3178), .Z(n3175) );
  XNOR U7274 ( .A(b[3483]), .B(n3176), .Z(n3177) );
  XNOR U7275 ( .A(b[3483]), .B(n3178), .Z(c[3483]) );
  XOR U7276 ( .A(n3179), .B(n3180), .Z(n3176) );
  ANDN U7277 ( .B(n3181), .A(n3182), .Z(n3179) );
  XNOR U7278 ( .A(b[3482]), .B(n3180), .Z(n3181) );
  XNOR U7279 ( .A(b[3482]), .B(n3182), .Z(c[3482]) );
  XOR U7280 ( .A(n3183), .B(n3184), .Z(n3180) );
  ANDN U7281 ( .B(n3185), .A(n3186), .Z(n3183) );
  XNOR U7282 ( .A(b[3481]), .B(n3184), .Z(n3185) );
  XNOR U7283 ( .A(b[3481]), .B(n3186), .Z(c[3481]) );
  XOR U7284 ( .A(n3187), .B(n3188), .Z(n3184) );
  ANDN U7285 ( .B(n3189), .A(n3190), .Z(n3187) );
  XNOR U7286 ( .A(b[3480]), .B(n3188), .Z(n3189) );
  XNOR U7287 ( .A(b[3480]), .B(n3190), .Z(c[3480]) );
  XOR U7288 ( .A(n3191), .B(n3192), .Z(n3188) );
  ANDN U7289 ( .B(n3193), .A(n3194), .Z(n3191) );
  XNOR U7290 ( .A(b[3479]), .B(n3192), .Z(n3193) );
  XNOR U7291 ( .A(b[347]), .B(n3195), .Z(c[347]) );
  XNOR U7292 ( .A(b[3479]), .B(n3194), .Z(c[3479]) );
  XOR U7293 ( .A(n3196), .B(n3197), .Z(n3192) );
  ANDN U7294 ( .B(n3198), .A(n3199), .Z(n3196) );
  XNOR U7295 ( .A(b[3478]), .B(n3197), .Z(n3198) );
  XNOR U7296 ( .A(b[3478]), .B(n3199), .Z(c[3478]) );
  XOR U7297 ( .A(n3200), .B(n3201), .Z(n3197) );
  ANDN U7298 ( .B(n3202), .A(n3203), .Z(n3200) );
  XNOR U7299 ( .A(b[3477]), .B(n3201), .Z(n3202) );
  XNOR U7300 ( .A(b[3477]), .B(n3203), .Z(c[3477]) );
  XOR U7301 ( .A(n3204), .B(n3205), .Z(n3201) );
  ANDN U7302 ( .B(n3206), .A(n3207), .Z(n3204) );
  XNOR U7303 ( .A(b[3476]), .B(n3205), .Z(n3206) );
  XNOR U7304 ( .A(b[3476]), .B(n3207), .Z(c[3476]) );
  XOR U7305 ( .A(n3208), .B(n3209), .Z(n3205) );
  ANDN U7306 ( .B(n3210), .A(n3211), .Z(n3208) );
  XNOR U7307 ( .A(b[3475]), .B(n3209), .Z(n3210) );
  XNOR U7308 ( .A(b[3475]), .B(n3211), .Z(c[3475]) );
  XOR U7309 ( .A(n3212), .B(n3213), .Z(n3209) );
  ANDN U7310 ( .B(n3214), .A(n3215), .Z(n3212) );
  XNOR U7311 ( .A(b[3474]), .B(n3213), .Z(n3214) );
  XNOR U7312 ( .A(b[3474]), .B(n3215), .Z(c[3474]) );
  XOR U7313 ( .A(n3216), .B(n3217), .Z(n3213) );
  ANDN U7314 ( .B(n3218), .A(n3219), .Z(n3216) );
  XNOR U7315 ( .A(b[3473]), .B(n3217), .Z(n3218) );
  XNOR U7316 ( .A(b[3473]), .B(n3219), .Z(c[3473]) );
  XOR U7317 ( .A(n3220), .B(n3221), .Z(n3217) );
  ANDN U7318 ( .B(n3222), .A(n3223), .Z(n3220) );
  XNOR U7319 ( .A(b[3472]), .B(n3221), .Z(n3222) );
  XNOR U7320 ( .A(b[3472]), .B(n3223), .Z(c[3472]) );
  XOR U7321 ( .A(n3224), .B(n3225), .Z(n3221) );
  ANDN U7322 ( .B(n3226), .A(n3227), .Z(n3224) );
  XNOR U7323 ( .A(b[3471]), .B(n3225), .Z(n3226) );
  XNOR U7324 ( .A(b[3471]), .B(n3227), .Z(c[3471]) );
  XOR U7325 ( .A(n3228), .B(n3229), .Z(n3225) );
  ANDN U7326 ( .B(n3230), .A(n3231), .Z(n3228) );
  XNOR U7327 ( .A(b[3470]), .B(n3229), .Z(n3230) );
  XNOR U7328 ( .A(b[3470]), .B(n3231), .Z(c[3470]) );
  XOR U7329 ( .A(n3232), .B(n3233), .Z(n3229) );
  ANDN U7330 ( .B(n3234), .A(n3235), .Z(n3232) );
  XNOR U7331 ( .A(b[3469]), .B(n3233), .Z(n3234) );
  XNOR U7332 ( .A(b[346]), .B(n3236), .Z(c[346]) );
  XNOR U7333 ( .A(b[3469]), .B(n3235), .Z(c[3469]) );
  XOR U7334 ( .A(n3237), .B(n3238), .Z(n3233) );
  ANDN U7335 ( .B(n3239), .A(n3240), .Z(n3237) );
  XNOR U7336 ( .A(b[3468]), .B(n3238), .Z(n3239) );
  XNOR U7337 ( .A(b[3468]), .B(n3240), .Z(c[3468]) );
  XOR U7338 ( .A(n3241), .B(n3242), .Z(n3238) );
  ANDN U7339 ( .B(n3243), .A(n3244), .Z(n3241) );
  XNOR U7340 ( .A(b[3467]), .B(n3242), .Z(n3243) );
  XNOR U7341 ( .A(b[3467]), .B(n3244), .Z(c[3467]) );
  XOR U7342 ( .A(n3245), .B(n3246), .Z(n3242) );
  ANDN U7343 ( .B(n3247), .A(n3248), .Z(n3245) );
  XNOR U7344 ( .A(b[3466]), .B(n3246), .Z(n3247) );
  XNOR U7345 ( .A(b[3466]), .B(n3248), .Z(c[3466]) );
  XOR U7346 ( .A(n3249), .B(n3250), .Z(n3246) );
  ANDN U7347 ( .B(n3251), .A(n3252), .Z(n3249) );
  XNOR U7348 ( .A(b[3465]), .B(n3250), .Z(n3251) );
  XNOR U7349 ( .A(b[3465]), .B(n3252), .Z(c[3465]) );
  XOR U7350 ( .A(n3253), .B(n3254), .Z(n3250) );
  ANDN U7351 ( .B(n3255), .A(n3256), .Z(n3253) );
  XNOR U7352 ( .A(b[3464]), .B(n3254), .Z(n3255) );
  XNOR U7353 ( .A(b[3464]), .B(n3256), .Z(c[3464]) );
  XOR U7354 ( .A(n3257), .B(n3258), .Z(n3254) );
  ANDN U7355 ( .B(n3259), .A(n3260), .Z(n3257) );
  XNOR U7356 ( .A(b[3463]), .B(n3258), .Z(n3259) );
  XNOR U7357 ( .A(b[3463]), .B(n3260), .Z(c[3463]) );
  XOR U7358 ( .A(n3261), .B(n3262), .Z(n3258) );
  ANDN U7359 ( .B(n3263), .A(n3264), .Z(n3261) );
  XNOR U7360 ( .A(b[3462]), .B(n3262), .Z(n3263) );
  XNOR U7361 ( .A(b[3462]), .B(n3264), .Z(c[3462]) );
  XOR U7362 ( .A(n3265), .B(n3266), .Z(n3262) );
  ANDN U7363 ( .B(n3267), .A(n3268), .Z(n3265) );
  XNOR U7364 ( .A(b[3461]), .B(n3266), .Z(n3267) );
  XNOR U7365 ( .A(b[3461]), .B(n3268), .Z(c[3461]) );
  XOR U7366 ( .A(n3269), .B(n3270), .Z(n3266) );
  ANDN U7367 ( .B(n3271), .A(n3272), .Z(n3269) );
  XNOR U7368 ( .A(b[3460]), .B(n3270), .Z(n3271) );
  XNOR U7369 ( .A(b[3460]), .B(n3272), .Z(c[3460]) );
  XOR U7370 ( .A(n3273), .B(n3274), .Z(n3270) );
  ANDN U7371 ( .B(n3275), .A(n3276), .Z(n3273) );
  XNOR U7372 ( .A(b[3459]), .B(n3274), .Z(n3275) );
  XNOR U7373 ( .A(b[345]), .B(n3277), .Z(c[345]) );
  XNOR U7374 ( .A(b[3459]), .B(n3276), .Z(c[3459]) );
  XOR U7375 ( .A(n3278), .B(n3279), .Z(n3274) );
  ANDN U7376 ( .B(n3280), .A(n3281), .Z(n3278) );
  XNOR U7377 ( .A(b[3458]), .B(n3279), .Z(n3280) );
  XNOR U7378 ( .A(b[3458]), .B(n3281), .Z(c[3458]) );
  XOR U7379 ( .A(n3282), .B(n3283), .Z(n3279) );
  ANDN U7380 ( .B(n3284), .A(n3285), .Z(n3282) );
  XNOR U7381 ( .A(b[3457]), .B(n3283), .Z(n3284) );
  XNOR U7382 ( .A(b[3457]), .B(n3285), .Z(c[3457]) );
  XOR U7383 ( .A(n3286), .B(n3287), .Z(n3283) );
  ANDN U7384 ( .B(n3288), .A(n3289), .Z(n3286) );
  XNOR U7385 ( .A(b[3456]), .B(n3287), .Z(n3288) );
  XNOR U7386 ( .A(b[3456]), .B(n3289), .Z(c[3456]) );
  XOR U7387 ( .A(n3290), .B(n3291), .Z(n3287) );
  ANDN U7388 ( .B(n3292), .A(n3293), .Z(n3290) );
  XNOR U7389 ( .A(b[3455]), .B(n3291), .Z(n3292) );
  XNOR U7390 ( .A(b[3455]), .B(n3293), .Z(c[3455]) );
  XOR U7391 ( .A(n3294), .B(n3295), .Z(n3291) );
  ANDN U7392 ( .B(n3296), .A(n3297), .Z(n3294) );
  XNOR U7393 ( .A(b[3454]), .B(n3295), .Z(n3296) );
  XNOR U7394 ( .A(b[3454]), .B(n3297), .Z(c[3454]) );
  XOR U7395 ( .A(n3298), .B(n3299), .Z(n3295) );
  ANDN U7396 ( .B(n3300), .A(n3301), .Z(n3298) );
  XNOR U7397 ( .A(b[3453]), .B(n3299), .Z(n3300) );
  XNOR U7398 ( .A(b[3453]), .B(n3301), .Z(c[3453]) );
  XOR U7399 ( .A(n3302), .B(n3303), .Z(n3299) );
  ANDN U7400 ( .B(n3304), .A(n3305), .Z(n3302) );
  XNOR U7401 ( .A(b[3452]), .B(n3303), .Z(n3304) );
  XNOR U7402 ( .A(b[3452]), .B(n3305), .Z(c[3452]) );
  XOR U7403 ( .A(n3306), .B(n3307), .Z(n3303) );
  ANDN U7404 ( .B(n3308), .A(n3309), .Z(n3306) );
  XNOR U7405 ( .A(b[3451]), .B(n3307), .Z(n3308) );
  XNOR U7406 ( .A(b[3451]), .B(n3309), .Z(c[3451]) );
  XOR U7407 ( .A(n3310), .B(n3311), .Z(n3307) );
  ANDN U7408 ( .B(n3312), .A(n3313), .Z(n3310) );
  XNOR U7409 ( .A(b[3450]), .B(n3311), .Z(n3312) );
  XNOR U7410 ( .A(b[3450]), .B(n3313), .Z(c[3450]) );
  XOR U7411 ( .A(n3314), .B(n3315), .Z(n3311) );
  ANDN U7412 ( .B(n3316), .A(n3317), .Z(n3314) );
  XNOR U7413 ( .A(b[3449]), .B(n3315), .Z(n3316) );
  XNOR U7414 ( .A(b[344]), .B(n3318), .Z(c[344]) );
  XNOR U7415 ( .A(b[3449]), .B(n3317), .Z(c[3449]) );
  XOR U7416 ( .A(n3319), .B(n3320), .Z(n3315) );
  ANDN U7417 ( .B(n3321), .A(n3322), .Z(n3319) );
  XNOR U7418 ( .A(b[3448]), .B(n3320), .Z(n3321) );
  XNOR U7419 ( .A(b[3448]), .B(n3322), .Z(c[3448]) );
  XOR U7420 ( .A(n3323), .B(n3324), .Z(n3320) );
  ANDN U7421 ( .B(n3325), .A(n3326), .Z(n3323) );
  XNOR U7422 ( .A(b[3447]), .B(n3324), .Z(n3325) );
  XNOR U7423 ( .A(b[3447]), .B(n3326), .Z(c[3447]) );
  XOR U7424 ( .A(n3327), .B(n3328), .Z(n3324) );
  ANDN U7425 ( .B(n3329), .A(n3330), .Z(n3327) );
  XNOR U7426 ( .A(b[3446]), .B(n3328), .Z(n3329) );
  XNOR U7427 ( .A(b[3446]), .B(n3330), .Z(c[3446]) );
  XOR U7428 ( .A(n3331), .B(n3332), .Z(n3328) );
  ANDN U7429 ( .B(n3333), .A(n3334), .Z(n3331) );
  XNOR U7430 ( .A(b[3445]), .B(n3332), .Z(n3333) );
  XNOR U7431 ( .A(b[3445]), .B(n3334), .Z(c[3445]) );
  XOR U7432 ( .A(n3335), .B(n3336), .Z(n3332) );
  ANDN U7433 ( .B(n3337), .A(n3338), .Z(n3335) );
  XNOR U7434 ( .A(b[3444]), .B(n3336), .Z(n3337) );
  XNOR U7435 ( .A(b[3444]), .B(n3338), .Z(c[3444]) );
  XOR U7436 ( .A(n3339), .B(n3340), .Z(n3336) );
  ANDN U7437 ( .B(n3341), .A(n3342), .Z(n3339) );
  XNOR U7438 ( .A(b[3443]), .B(n3340), .Z(n3341) );
  XNOR U7439 ( .A(b[3443]), .B(n3342), .Z(c[3443]) );
  XOR U7440 ( .A(n3343), .B(n3344), .Z(n3340) );
  ANDN U7441 ( .B(n3345), .A(n3346), .Z(n3343) );
  XNOR U7442 ( .A(b[3442]), .B(n3344), .Z(n3345) );
  XNOR U7443 ( .A(b[3442]), .B(n3346), .Z(c[3442]) );
  XOR U7444 ( .A(n3347), .B(n3348), .Z(n3344) );
  ANDN U7445 ( .B(n3349), .A(n3350), .Z(n3347) );
  XNOR U7446 ( .A(b[3441]), .B(n3348), .Z(n3349) );
  XNOR U7447 ( .A(b[3441]), .B(n3350), .Z(c[3441]) );
  XOR U7448 ( .A(n3351), .B(n3352), .Z(n3348) );
  ANDN U7449 ( .B(n3353), .A(n3354), .Z(n3351) );
  XNOR U7450 ( .A(b[3440]), .B(n3352), .Z(n3353) );
  XNOR U7451 ( .A(b[3440]), .B(n3354), .Z(c[3440]) );
  XOR U7452 ( .A(n3355), .B(n3356), .Z(n3352) );
  ANDN U7453 ( .B(n3357), .A(n3358), .Z(n3355) );
  XNOR U7454 ( .A(b[3439]), .B(n3356), .Z(n3357) );
  XNOR U7455 ( .A(b[343]), .B(n3359), .Z(c[343]) );
  XNOR U7456 ( .A(b[3439]), .B(n3358), .Z(c[3439]) );
  XOR U7457 ( .A(n3360), .B(n3361), .Z(n3356) );
  ANDN U7458 ( .B(n3362), .A(n3363), .Z(n3360) );
  XNOR U7459 ( .A(b[3438]), .B(n3361), .Z(n3362) );
  XNOR U7460 ( .A(b[3438]), .B(n3363), .Z(c[3438]) );
  XOR U7461 ( .A(n3364), .B(n3365), .Z(n3361) );
  ANDN U7462 ( .B(n3366), .A(n3367), .Z(n3364) );
  XNOR U7463 ( .A(b[3437]), .B(n3365), .Z(n3366) );
  XNOR U7464 ( .A(b[3437]), .B(n3367), .Z(c[3437]) );
  XOR U7465 ( .A(n3368), .B(n3369), .Z(n3365) );
  ANDN U7466 ( .B(n3370), .A(n3371), .Z(n3368) );
  XNOR U7467 ( .A(b[3436]), .B(n3369), .Z(n3370) );
  XNOR U7468 ( .A(b[3436]), .B(n3371), .Z(c[3436]) );
  XOR U7469 ( .A(n3372), .B(n3373), .Z(n3369) );
  ANDN U7470 ( .B(n3374), .A(n3375), .Z(n3372) );
  XNOR U7471 ( .A(b[3435]), .B(n3373), .Z(n3374) );
  XNOR U7472 ( .A(b[3435]), .B(n3375), .Z(c[3435]) );
  XOR U7473 ( .A(n3376), .B(n3377), .Z(n3373) );
  ANDN U7474 ( .B(n3378), .A(n3379), .Z(n3376) );
  XNOR U7475 ( .A(b[3434]), .B(n3377), .Z(n3378) );
  XNOR U7476 ( .A(b[3434]), .B(n3379), .Z(c[3434]) );
  XOR U7477 ( .A(n3380), .B(n3381), .Z(n3377) );
  ANDN U7478 ( .B(n3382), .A(n3383), .Z(n3380) );
  XNOR U7479 ( .A(b[3433]), .B(n3381), .Z(n3382) );
  XNOR U7480 ( .A(b[3433]), .B(n3383), .Z(c[3433]) );
  XOR U7481 ( .A(n3384), .B(n3385), .Z(n3381) );
  ANDN U7482 ( .B(n3386), .A(n3387), .Z(n3384) );
  XNOR U7483 ( .A(b[3432]), .B(n3385), .Z(n3386) );
  XNOR U7484 ( .A(b[3432]), .B(n3387), .Z(c[3432]) );
  XOR U7485 ( .A(n3388), .B(n3389), .Z(n3385) );
  ANDN U7486 ( .B(n3390), .A(n3391), .Z(n3388) );
  XNOR U7487 ( .A(b[3431]), .B(n3389), .Z(n3390) );
  XNOR U7488 ( .A(b[3431]), .B(n3391), .Z(c[3431]) );
  XOR U7489 ( .A(n3392), .B(n3393), .Z(n3389) );
  ANDN U7490 ( .B(n3394), .A(n3395), .Z(n3392) );
  XNOR U7491 ( .A(b[3430]), .B(n3393), .Z(n3394) );
  XNOR U7492 ( .A(b[3430]), .B(n3395), .Z(c[3430]) );
  XOR U7493 ( .A(n3396), .B(n3397), .Z(n3393) );
  ANDN U7494 ( .B(n3398), .A(n3399), .Z(n3396) );
  XNOR U7495 ( .A(b[3429]), .B(n3397), .Z(n3398) );
  XNOR U7496 ( .A(b[342]), .B(n3400), .Z(c[342]) );
  XNOR U7497 ( .A(b[3429]), .B(n3399), .Z(c[3429]) );
  XOR U7498 ( .A(n3401), .B(n3402), .Z(n3397) );
  ANDN U7499 ( .B(n3403), .A(n3404), .Z(n3401) );
  XNOR U7500 ( .A(b[3428]), .B(n3402), .Z(n3403) );
  XNOR U7501 ( .A(b[3428]), .B(n3404), .Z(c[3428]) );
  XOR U7502 ( .A(n3405), .B(n3406), .Z(n3402) );
  ANDN U7503 ( .B(n3407), .A(n3408), .Z(n3405) );
  XNOR U7504 ( .A(b[3427]), .B(n3406), .Z(n3407) );
  XNOR U7505 ( .A(b[3427]), .B(n3408), .Z(c[3427]) );
  XOR U7506 ( .A(n3409), .B(n3410), .Z(n3406) );
  ANDN U7507 ( .B(n3411), .A(n3412), .Z(n3409) );
  XNOR U7508 ( .A(b[3426]), .B(n3410), .Z(n3411) );
  XNOR U7509 ( .A(b[3426]), .B(n3412), .Z(c[3426]) );
  XOR U7510 ( .A(n3413), .B(n3414), .Z(n3410) );
  ANDN U7511 ( .B(n3415), .A(n3416), .Z(n3413) );
  XNOR U7512 ( .A(b[3425]), .B(n3414), .Z(n3415) );
  XNOR U7513 ( .A(b[3425]), .B(n3416), .Z(c[3425]) );
  XOR U7514 ( .A(n3417), .B(n3418), .Z(n3414) );
  ANDN U7515 ( .B(n3419), .A(n3420), .Z(n3417) );
  XNOR U7516 ( .A(b[3424]), .B(n3418), .Z(n3419) );
  XNOR U7517 ( .A(b[3424]), .B(n3420), .Z(c[3424]) );
  XOR U7518 ( .A(n3421), .B(n3422), .Z(n3418) );
  ANDN U7519 ( .B(n3423), .A(n3424), .Z(n3421) );
  XNOR U7520 ( .A(b[3423]), .B(n3422), .Z(n3423) );
  XNOR U7521 ( .A(b[3423]), .B(n3424), .Z(c[3423]) );
  XOR U7522 ( .A(n3425), .B(n3426), .Z(n3422) );
  ANDN U7523 ( .B(n3427), .A(n3428), .Z(n3425) );
  XNOR U7524 ( .A(b[3422]), .B(n3426), .Z(n3427) );
  XNOR U7525 ( .A(b[3422]), .B(n3428), .Z(c[3422]) );
  XOR U7526 ( .A(n3429), .B(n3430), .Z(n3426) );
  ANDN U7527 ( .B(n3431), .A(n3432), .Z(n3429) );
  XNOR U7528 ( .A(b[3421]), .B(n3430), .Z(n3431) );
  XNOR U7529 ( .A(b[3421]), .B(n3432), .Z(c[3421]) );
  XOR U7530 ( .A(n3433), .B(n3434), .Z(n3430) );
  ANDN U7531 ( .B(n3435), .A(n3436), .Z(n3433) );
  XNOR U7532 ( .A(b[3420]), .B(n3434), .Z(n3435) );
  XNOR U7533 ( .A(b[3420]), .B(n3436), .Z(c[3420]) );
  XOR U7534 ( .A(n3437), .B(n3438), .Z(n3434) );
  ANDN U7535 ( .B(n3439), .A(n3440), .Z(n3437) );
  XNOR U7536 ( .A(b[3419]), .B(n3438), .Z(n3439) );
  XNOR U7537 ( .A(b[341]), .B(n3441), .Z(c[341]) );
  XNOR U7538 ( .A(b[3419]), .B(n3440), .Z(c[3419]) );
  XOR U7539 ( .A(n3442), .B(n3443), .Z(n3438) );
  ANDN U7540 ( .B(n3444), .A(n3445), .Z(n3442) );
  XNOR U7541 ( .A(b[3418]), .B(n3443), .Z(n3444) );
  XNOR U7542 ( .A(b[3418]), .B(n3445), .Z(c[3418]) );
  XOR U7543 ( .A(n3446), .B(n3447), .Z(n3443) );
  ANDN U7544 ( .B(n3448), .A(n3449), .Z(n3446) );
  XNOR U7545 ( .A(b[3417]), .B(n3447), .Z(n3448) );
  XNOR U7546 ( .A(b[3417]), .B(n3449), .Z(c[3417]) );
  XOR U7547 ( .A(n3450), .B(n3451), .Z(n3447) );
  ANDN U7548 ( .B(n3452), .A(n3453), .Z(n3450) );
  XNOR U7549 ( .A(b[3416]), .B(n3451), .Z(n3452) );
  XNOR U7550 ( .A(b[3416]), .B(n3453), .Z(c[3416]) );
  XOR U7551 ( .A(n3454), .B(n3455), .Z(n3451) );
  ANDN U7552 ( .B(n3456), .A(n3457), .Z(n3454) );
  XNOR U7553 ( .A(b[3415]), .B(n3455), .Z(n3456) );
  XNOR U7554 ( .A(b[3415]), .B(n3457), .Z(c[3415]) );
  XOR U7555 ( .A(n3458), .B(n3459), .Z(n3455) );
  ANDN U7556 ( .B(n3460), .A(n3461), .Z(n3458) );
  XNOR U7557 ( .A(b[3414]), .B(n3459), .Z(n3460) );
  XNOR U7558 ( .A(b[3414]), .B(n3461), .Z(c[3414]) );
  XOR U7559 ( .A(n3462), .B(n3463), .Z(n3459) );
  ANDN U7560 ( .B(n3464), .A(n3465), .Z(n3462) );
  XNOR U7561 ( .A(b[3413]), .B(n3463), .Z(n3464) );
  XNOR U7562 ( .A(b[3413]), .B(n3465), .Z(c[3413]) );
  XOR U7563 ( .A(n3466), .B(n3467), .Z(n3463) );
  ANDN U7564 ( .B(n3468), .A(n3469), .Z(n3466) );
  XNOR U7565 ( .A(b[3412]), .B(n3467), .Z(n3468) );
  XNOR U7566 ( .A(b[3412]), .B(n3469), .Z(c[3412]) );
  XOR U7567 ( .A(n3470), .B(n3471), .Z(n3467) );
  ANDN U7568 ( .B(n3472), .A(n3473), .Z(n3470) );
  XNOR U7569 ( .A(b[3411]), .B(n3471), .Z(n3472) );
  XNOR U7570 ( .A(b[3411]), .B(n3473), .Z(c[3411]) );
  XOR U7571 ( .A(n3474), .B(n3475), .Z(n3471) );
  ANDN U7572 ( .B(n3476), .A(n3477), .Z(n3474) );
  XNOR U7573 ( .A(b[3410]), .B(n3475), .Z(n3476) );
  XNOR U7574 ( .A(b[3410]), .B(n3477), .Z(c[3410]) );
  XOR U7575 ( .A(n3478), .B(n3479), .Z(n3475) );
  ANDN U7576 ( .B(n3480), .A(n3481), .Z(n3478) );
  XNOR U7577 ( .A(b[3409]), .B(n3479), .Z(n3480) );
  XNOR U7578 ( .A(b[340]), .B(n3482), .Z(c[340]) );
  XNOR U7579 ( .A(b[3409]), .B(n3481), .Z(c[3409]) );
  XOR U7580 ( .A(n3483), .B(n3484), .Z(n3479) );
  ANDN U7581 ( .B(n3485), .A(n3486), .Z(n3483) );
  XNOR U7582 ( .A(b[3408]), .B(n3484), .Z(n3485) );
  XNOR U7583 ( .A(b[3408]), .B(n3486), .Z(c[3408]) );
  XOR U7584 ( .A(n3487), .B(n3488), .Z(n3484) );
  ANDN U7585 ( .B(n3489), .A(n3490), .Z(n3487) );
  XNOR U7586 ( .A(b[3407]), .B(n3488), .Z(n3489) );
  XNOR U7587 ( .A(b[3407]), .B(n3490), .Z(c[3407]) );
  XOR U7588 ( .A(n3491), .B(n3492), .Z(n3488) );
  ANDN U7589 ( .B(n3493), .A(n3494), .Z(n3491) );
  XNOR U7590 ( .A(b[3406]), .B(n3492), .Z(n3493) );
  XNOR U7591 ( .A(b[3406]), .B(n3494), .Z(c[3406]) );
  XOR U7592 ( .A(n3495), .B(n3496), .Z(n3492) );
  ANDN U7593 ( .B(n3497), .A(n3498), .Z(n3495) );
  XNOR U7594 ( .A(b[3405]), .B(n3496), .Z(n3497) );
  XNOR U7595 ( .A(b[3405]), .B(n3498), .Z(c[3405]) );
  XOR U7596 ( .A(n3499), .B(n3500), .Z(n3496) );
  ANDN U7597 ( .B(n3501), .A(n3502), .Z(n3499) );
  XNOR U7598 ( .A(b[3404]), .B(n3500), .Z(n3501) );
  XNOR U7599 ( .A(b[3404]), .B(n3502), .Z(c[3404]) );
  XOR U7600 ( .A(n3503), .B(n3504), .Z(n3500) );
  ANDN U7601 ( .B(n3505), .A(n3506), .Z(n3503) );
  XNOR U7602 ( .A(b[3403]), .B(n3504), .Z(n3505) );
  XNOR U7603 ( .A(b[3403]), .B(n3506), .Z(c[3403]) );
  XOR U7604 ( .A(n3507), .B(n3508), .Z(n3504) );
  ANDN U7605 ( .B(n3509), .A(n3510), .Z(n3507) );
  XNOR U7606 ( .A(b[3402]), .B(n3508), .Z(n3509) );
  XNOR U7607 ( .A(b[3402]), .B(n3510), .Z(c[3402]) );
  XOR U7608 ( .A(n3511), .B(n3512), .Z(n3508) );
  ANDN U7609 ( .B(n3513), .A(n3514), .Z(n3511) );
  XNOR U7610 ( .A(b[3401]), .B(n3512), .Z(n3513) );
  XNOR U7611 ( .A(b[3401]), .B(n3514), .Z(c[3401]) );
  XOR U7612 ( .A(n3515), .B(n3516), .Z(n3512) );
  ANDN U7613 ( .B(n3517), .A(n3518), .Z(n3515) );
  XNOR U7614 ( .A(b[3400]), .B(n3516), .Z(n3517) );
  XNOR U7615 ( .A(b[3400]), .B(n3518), .Z(c[3400]) );
  XOR U7616 ( .A(n3519), .B(n3520), .Z(n3516) );
  ANDN U7617 ( .B(n3521), .A(n3522), .Z(n3519) );
  XNOR U7618 ( .A(b[3399]), .B(n3520), .Z(n3521) );
  XNOR U7619 ( .A(b[33]), .B(n3523), .Z(c[33]) );
  XNOR U7620 ( .A(b[339]), .B(n3524), .Z(c[339]) );
  XNOR U7621 ( .A(b[3399]), .B(n3522), .Z(c[3399]) );
  XOR U7622 ( .A(n3525), .B(n3526), .Z(n3520) );
  ANDN U7623 ( .B(n3527), .A(n3528), .Z(n3525) );
  XNOR U7624 ( .A(b[3398]), .B(n3526), .Z(n3527) );
  XNOR U7625 ( .A(b[3398]), .B(n3528), .Z(c[3398]) );
  XOR U7626 ( .A(n3529), .B(n3530), .Z(n3526) );
  ANDN U7627 ( .B(n3531), .A(n3532), .Z(n3529) );
  XNOR U7628 ( .A(b[3397]), .B(n3530), .Z(n3531) );
  XNOR U7629 ( .A(b[3397]), .B(n3532), .Z(c[3397]) );
  XOR U7630 ( .A(n3533), .B(n3534), .Z(n3530) );
  ANDN U7631 ( .B(n3535), .A(n3536), .Z(n3533) );
  XNOR U7632 ( .A(b[3396]), .B(n3534), .Z(n3535) );
  XNOR U7633 ( .A(b[3396]), .B(n3536), .Z(c[3396]) );
  XOR U7634 ( .A(n3537), .B(n3538), .Z(n3534) );
  ANDN U7635 ( .B(n3539), .A(n3540), .Z(n3537) );
  XNOR U7636 ( .A(b[3395]), .B(n3538), .Z(n3539) );
  XNOR U7637 ( .A(b[3395]), .B(n3540), .Z(c[3395]) );
  XOR U7638 ( .A(n3541), .B(n3542), .Z(n3538) );
  ANDN U7639 ( .B(n3543), .A(n3544), .Z(n3541) );
  XNOR U7640 ( .A(b[3394]), .B(n3542), .Z(n3543) );
  XNOR U7641 ( .A(b[3394]), .B(n3544), .Z(c[3394]) );
  XOR U7642 ( .A(n3545), .B(n3546), .Z(n3542) );
  ANDN U7643 ( .B(n3547), .A(n3548), .Z(n3545) );
  XNOR U7644 ( .A(b[3393]), .B(n3546), .Z(n3547) );
  XNOR U7645 ( .A(b[3393]), .B(n3548), .Z(c[3393]) );
  XOR U7646 ( .A(n3549), .B(n3550), .Z(n3546) );
  ANDN U7647 ( .B(n3551), .A(n3552), .Z(n3549) );
  XNOR U7648 ( .A(b[3392]), .B(n3550), .Z(n3551) );
  XNOR U7649 ( .A(b[3392]), .B(n3552), .Z(c[3392]) );
  XOR U7650 ( .A(n3553), .B(n3554), .Z(n3550) );
  ANDN U7651 ( .B(n3555), .A(n3556), .Z(n3553) );
  XNOR U7652 ( .A(b[3391]), .B(n3554), .Z(n3555) );
  XNOR U7653 ( .A(b[3391]), .B(n3556), .Z(c[3391]) );
  XOR U7654 ( .A(n3557), .B(n3558), .Z(n3554) );
  ANDN U7655 ( .B(n3559), .A(n3560), .Z(n3557) );
  XNOR U7656 ( .A(b[3390]), .B(n3558), .Z(n3559) );
  XNOR U7657 ( .A(b[3390]), .B(n3560), .Z(c[3390]) );
  XOR U7658 ( .A(n3561), .B(n3562), .Z(n3558) );
  ANDN U7659 ( .B(n3563), .A(n3564), .Z(n3561) );
  XNOR U7660 ( .A(b[3389]), .B(n3562), .Z(n3563) );
  XNOR U7661 ( .A(b[338]), .B(n3565), .Z(c[338]) );
  XNOR U7662 ( .A(b[3389]), .B(n3564), .Z(c[3389]) );
  XOR U7663 ( .A(n3566), .B(n3567), .Z(n3562) );
  ANDN U7664 ( .B(n3568), .A(n3569), .Z(n3566) );
  XNOR U7665 ( .A(b[3388]), .B(n3567), .Z(n3568) );
  XNOR U7666 ( .A(b[3388]), .B(n3569), .Z(c[3388]) );
  XOR U7667 ( .A(n3570), .B(n3571), .Z(n3567) );
  ANDN U7668 ( .B(n3572), .A(n3573), .Z(n3570) );
  XNOR U7669 ( .A(b[3387]), .B(n3571), .Z(n3572) );
  XNOR U7670 ( .A(b[3387]), .B(n3573), .Z(c[3387]) );
  XOR U7671 ( .A(n3574), .B(n3575), .Z(n3571) );
  ANDN U7672 ( .B(n3576), .A(n3577), .Z(n3574) );
  XNOR U7673 ( .A(b[3386]), .B(n3575), .Z(n3576) );
  XNOR U7674 ( .A(b[3386]), .B(n3577), .Z(c[3386]) );
  XOR U7675 ( .A(n3578), .B(n3579), .Z(n3575) );
  ANDN U7676 ( .B(n3580), .A(n3581), .Z(n3578) );
  XNOR U7677 ( .A(b[3385]), .B(n3579), .Z(n3580) );
  XNOR U7678 ( .A(b[3385]), .B(n3581), .Z(c[3385]) );
  XOR U7679 ( .A(n3582), .B(n3583), .Z(n3579) );
  ANDN U7680 ( .B(n3584), .A(n3585), .Z(n3582) );
  XNOR U7681 ( .A(b[3384]), .B(n3583), .Z(n3584) );
  XNOR U7682 ( .A(b[3384]), .B(n3585), .Z(c[3384]) );
  XOR U7683 ( .A(n3586), .B(n3587), .Z(n3583) );
  ANDN U7684 ( .B(n3588), .A(n3589), .Z(n3586) );
  XNOR U7685 ( .A(b[3383]), .B(n3587), .Z(n3588) );
  XNOR U7686 ( .A(b[3383]), .B(n3589), .Z(c[3383]) );
  XOR U7687 ( .A(n3590), .B(n3591), .Z(n3587) );
  ANDN U7688 ( .B(n3592), .A(n3593), .Z(n3590) );
  XNOR U7689 ( .A(b[3382]), .B(n3591), .Z(n3592) );
  XNOR U7690 ( .A(b[3382]), .B(n3593), .Z(c[3382]) );
  XOR U7691 ( .A(n3594), .B(n3595), .Z(n3591) );
  ANDN U7692 ( .B(n3596), .A(n3597), .Z(n3594) );
  XNOR U7693 ( .A(b[3381]), .B(n3595), .Z(n3596) );
  XNOR U7694 ( .A(b[3381]), .B(n3597), .Z(c[3381]) );
  XOR U7695 ( .A(n3598), .B(n3599), .Z(n3595) );
  ANDN U7696 ( .B(n3600), .A(n3601), .Z(n3598) );
  XNOR U7697 ( .A(b[3380]), .B(n3599), .Z(n3600) );
  XNOR U7698 ( .A(b[3380]), .B(n3601), .Z(c[3380]) );
  XOR U7699 ( .A(n3602), .B(n3603), .Z(n3599) );
  ANDN U7700 ( .B(n3604), .A(n3605), .Z(n3602) );
  XNOR U7701 ( .A(b[3379]), .B(n3603), .Z(n3604) );
  XNOR U7702 ( .A(b[337]), .B(n3606), .Z(c[337]) );
  XNOR U7703 ( .A(b[3379]), .B(n3605), .Z(c[3379]) );
  XOR U7704 ( .A(n3607), .B(n3608), .Z(n3603) );
  ANDN U7705 ( .B(n3609), .A(n3610), .Z(n3607) );
  XNOR U7706 ( .A(b[3378]), .B(n3608), .Z(n3609) );
  XNOR U7707 ( .A(b[3378]), .B(n3610), .Z(c[3378]) );
  XOR U7708 ( .A(n3611), .B(n3612), .Z(n3608) );
  ANDN U7709 ( .B(n3613), .A(n3614), .Z(n3611) );
  XNOR U7710 ( .A(b[3377]), .B(n3612), .Z(n3613) );
  XNOR U7711 ( .A(b[3377]), .B(n3614), .Z(c[3377]) );
  XOR U7712 ( .A(n3615), .B(n3616), .Z(n3612) );
  ANDN U7713 ( .B(n3617), .A(n3618), .Z(n3615) );
  XNOR U7714 ( .A(b[3376]), .B(n3616), .Z(n3617) );
  XNOR U7715 ( .A(b[3376]), .B(n3618), .Z(c[3376]) );
  XOR U7716 ( .A(n3619), .B(n3620), .Z(n3616) );
  ANDN U7717 ( .B(n3621), .A(n3622), .Z(n3619) );
  XNOR U7718 ( .A(b[3375]), .B(n3620), .Z(n3621) );
  XNOR U7719 ( .A(b[3375]), .B(n3622), .Z(c[3375]) );
  XOR U7720 ( .A(n3623), .B(n3624), .Z(n3620) );
  ANDN U7721 ( .B(n3625), .A(n3626), .Z(n3623) );
  XNOR U7722 ( .A(b[3374]), .B(n3624), .Z(n3625) );
  XNOR U7723 ( .A(b[3374]), .B(n3626), .Z(c[3374]) );
  XOR U7724 ( .A(n3627), .B(n3628), .Z(n3624) );
  ANDN U7725 ( .B(n3629), .A(n3630), .Z(n3627) );
  XNOR U7726 ( .A(b[3373]), .B(n3628), .Z(n3629) );
  XNOR U7727 ( .A(b[3373]), .B(n3630), .Z(c[3373]) );
  XOR U7728 ( .A(n3631), .B(n3632), .Z(n3628) );
  ANDN U7729 ( .B(n3633), .A(n3634), .Z(n3631) );
  XNOR U7730 ( .A(b[3372]), .B(n3632), .Z(n3633) );
  XNOR U7731 ( .A(b[3372]), .B(n3634), .Z(c[3372]) );
  XOR U7732 ( .A(n3635), .B(n3636), .Z(n3632) );
  ANDN U7733 ( .B(n3637), .A(n3638), .Z(n3635) );
  XNOR U7734 ( .A(b[3371]), .B(n3636), .Z(n3637) );
  XNOR U7735 ( .A(b[3371]), .B(n3638), .Z(c[3371]) );
  XOR U7736 ( .A(n3639), .B(n3640), .Z(n3636) );
  ANDN U7737 ( .B(n3641), .A(n3642), .Z(n3639) );
  XNOR U7738 ( .A(b[3370]), .B(n3640), .Z(n3641) );
  XNOR U7739 ( .A(b[3370]), .B(n3642), .Z(c[3370]) );
  XOR U7740 ( .A(n3643), .B(n3644), .Z(n3640) );
  ANDN U7741 ( .B(n3645), .A(n3646), .Z(n3643) );
  XNOR U7742 ( .A(b[3369]), .B(n3644), .Z(n3645) );
  XNOR U7743 ( .A(b[336]), .B(n3647), .Z(c[336]) );
  XNOR U7744 ( .A(b[3369]), .B(n3646), .Z(c[3369]) );
  XOR U7745 ( .A(n3648), .B(n3649), .Z(n3644) );
  ANDN U7746 ( .B(n3650), .A(n3651), .Z(n3648) );
  XNOR U7747 ( .A(b[3368]), .B(n3649), .Z(n3650) );
  XNOR U7748 ( .A(b[3368]), .B(n3651), .Z(c[3368]) );
  XOR U7749 ( .A(n3652), .B(n3653), .Z(n3649) );
  ANDN U7750 ( .B(n3654), .A(n3655), .Z(n3652) );
  XNOR U7751 ( .A(b[3367]), .B(n3653), .Z(n3654) );
  XNOR U7752 ( .A(b[3367]), .B(n3655), .Z(c[3367]) );
  XOR U7753 ( .A(n3656), .B(n3657), .Z(n3653) );
  ANDN U7754 ( .B(n3658), .A(n3659), .Z(n3656) );
  XNOR U7755 ( .A(b[3366]), .B(n3657), .Z(n3658) );
  XNOR U7756 ( .A(b[3366]), .B(n3659), .Z(c[3366]) );
  XOR U7757 ( .A(n3660), .B(n3661), .Z(n3657) );
  ANDN U7758 ( .B(n3662), .A(n3663), .Z(n3660) );
  XNOR U7759 ( .A(b[3365]), .B(n3661), .Z(n3662) );
  XNOR U7760 ( .A(b[3365]), .B(n3663), .Z(c[3365]) );
  XOR U7761 ( .A(n3664), .B(n3665), .Z(n3661) );
  ANDN U7762 ( .B(n3666), .A(n3667), .Z(n3664) );
  XNOR U7763 ( .A(b[3364]), .B(n3665), .Z(n3666) );
  XNOR U7764 ( .A(b[3364]), .B(n3667), .Z(c[3364]) );
  XOR U7765 ( .A(n3668), .B(n3669), .Z(n3665) );
  ANDN U7766 ( .B(n3670), .A(n3671), .Z(n3668) );
  XNOR U7767 ( .A(b[3363]), .B(n3669), .Z(n3670) );
  XNOR U7768 ( .A(b[3363]), .B(n3671), .Z(c[3363]) );
  XOR U7769 ( .A(n3672), .B(n3673), .Z(n3669) );
  ANDN U7770 ( .B(n3674), .A(n3675), .Z(n3672) );
  XNOR U7771 ( .A(b[3362]), .B(n3673), .Z(n3674) );
  XNOR U7772 ( .A(b[3362]), .B(n3675), .Z(c[3362]) );
  XOR U7773 ( .A(n3676), .B(n3677), .Z(n3673) );
  ANDN U7774 ( .B(n3678), .A(n3679), .Z(n3676) );
  XNOR U7775 ( .A(b[3361]), .B(n3677), .Z(n3678) );
  XNOR U7776 ( .A(b[3361]), .B(n3679), .Z(c[3361]) );
  XOR U7777 ( .A(n3680), .B(n3681), .Z(n3677) );
  ANDN U7778 ( .B(n3682), .A(n3683), .Z(n3680) );
  XNOR U7779 ( .A(b[3360]), .B(n3681), .Z(n3682) );
  XNOR U7780 ( .A(b[3360]), .B(n3683), .Z(c[3360]) );
  XOR U7781 ( .A(n3684), .B(n3685), .Z(n3681) );
  ANDN U7782 ( .B(n3686), .A(n3687), .Z(n3684) );
  XNOR U7783 ( .A(b[3359]), .B(n3685), .Z(n3686) );
  XNOR U7784 ( .A(b[335]), .B(n3688), .Z(c[335]) );
  XNOR U7785 ( .A(b[3359]), .B(n3687), .Z(c[3359]) );
  XOR U7786 ( .A(n3689), .B(n3690), .Z(n3685) );
  ANDN U7787 ( .B(n3691), .A(n3692), .Z(n3689) );
  XNOR U7788 ( .A(b[3358]), .B(n3690), .Z(n3691) );
  XNOR U7789 ( .A(b[3358]), .B(n3692), .Z(c[3358]) );
  XOR U7790 ( .A(n3693), .B(n3694), .Z(n3690) );
  ANDN U7791 ( .B(n3695), .A(n3696), .Z(n3693) );
  XNOR U7792 ( .A(b[3357]), .B(n3694), .Z(n3695) );
  XNOR U7793 ( .A(b[3357]), .B(n3696), .Z(c[3357]) );
  XOR U7794 ( .A(n3697), .B(n3698), .Z(n3694) );
  ANDN U7795 ( .B(n3699), .A(n3700), .Z(n3697) );
  XNOR U7796 ( .A(b[3356]), .B(n3698), .Z(n3699) );
  XNOR U7797 ( .A(b[3356]), .B(n3700), .Z(c[3356]) );
  XOR U7798 ( .A(n3701), .B(n3702), .Z(n3698) );
  ANDN U7799 ( .B(n3703), .A(n3704), .Z(n3701) );
  XNOR U7800 ( .A(b[3355]), .B(n3702), .Z(n3703) );
  XNOR U7801 ( .A(b[3355]), .B(n3704), .Z(c[3355]) );
  XOR U7802 ( .A(n3705), .B(n3706), .Z(n3702) );
  ANDN U7803 ( .B(n3707), .A(n3708), .Z(n3705) );
  XNOR U7804 ( .A(b[3354]), .B(n3706), .Z(n3707) );
  XNOR U7805 ( .A(b[3354]), .B(n3708), .Z(c[3354]) );
  XOR U7806 ( .A(n3709), .B(n3710), .Z(n3706) );
  ANDN U7807 ( .B(n3711), .A(n3712), .Z(n3709) );
  XNOR U7808 ( .A(b[3353]), .B(n3710), .Z(n3711) );
  XNOR U7809 ( .A(b[3353]), .B(n3712), .Z(c[3353]) );
  XOR U7810 ( .A(n3713), .B(n3714), .Z(n3710) );
  ANDN U7811 ( .B(n3715), .A(n3716), .Z(n3713) );
  XNOR U7812 ( .A(b[3352]), .B(n3714), .Z(n3715) );
  XNOR U7813 ( .A(b[3352]), .B(n3716), .Z(c[3352]) );
  XOR U7814 ( .A(n3717), .B(n3718), .Z(n3714) );
  ANDN U7815 ( .B(n3719), .A(n3720), .Z(n3717) );
  XNOR U7816 ( .A(b[3351]), .B(n3718), .Z(n3719) );
  XNOR U7817 ( .A(b[3351]), .B(n3720), .Z(c[3351]) );
  XOR U7818 ( .A(n3721), .B(n3722), .Z(n3718) );
  ANDN U7819 ( .B(n3723), .A(n3724), .Z(n3721) );
  XNOR U7820 ( .A(b[3350]), .B(n3722), .Z(n3723) );
  XNOR U7821 ( .A(b[3350]), .B(n3724), .Z(c[3350]) );
  XOR U7822 ( .A(n3725), .B(n3726), .Z(n3722) );
  ANDN U7823 ( .B(n3727), .A(n3728), .Z(n3725) );
  XNOR U7824 ( .A(b[3349]), .B(n3726), .Z(n3727) );
  XNOR U7825 ( .A(b[334]), .B(n3729), .Z(c[334]) );
  XNOR U7826 ( .A(b[3349]), .B(n3728), .Z(c[3349]) );
  XOR U7827 ( .A(n3730), .B(n3731), .Z(n3726) );
  ANDN U7828 ( .B(n3732), .A(n3733), .Z(n3730) );
  XNOR U7829 ( .A(b[3348]), .B(n3731), .Z(n3732) );
  XNOR U7830 ( .A(b[3348]), .B(n3733), .Z(c[3348]) );
  XOR U7831 ( .A(n3734), .B(n3735), .Z(n3731) );
  ANDN U7832 ( .B(n3736), .A(n3737), .Z(n3734) );
  XNOR U7833 ( .A(b[3347]), .B(n3735), .Z(n3736) );
  XNOR U7834 ( .A(b[3347]), .B(n3737), .Z(c[3347]) );
  XOR U7835 ( .A(n3738), .B(n3739), .Z(n3735) );
  ANDN U7836 ( .B(n3740), .A(n3741), .Z(n3738) );
  XNOR U7837 ( .A(b[3346]), .B(n3739), .Z(n3740) );
  XNOR U7838 ( .A(b[3346]), .B(n3741), .Z(c[3346]) );
  XOR U7839 ( .A(n3742), .B(n3743), .Z(n3739) );
  ANDN U7840 ( .B(n3744), .A(n3745), .Z(n3742) );
  XNOR U7841 ( .A(b[3345]), .B(n3743), .Z(n3744) );
  XNOR U7842 ( .A(b[3345]), .B(n3745), .Z(c[3345]) );
  XOR U7843 ( .A(n3746), .B(n3747), .Z(n3743) );
  ANDN U7844 ( .B(n3748), .A(n3749), .Z(n3746) );
  XNOR U7845 ( .A(b[3344]), .B(n3747), .Z(n3748) );
  XNOR U7846 ( .A(b[3344]), .B(n3749), .Z(c[3344]) );
  XOR U7847 ( .A(n3750), .B(n3751), .Z(n3747) );
  ANDN U7848 ( .B(n3752), .A(n3753), .Z(n3750) );
  XNOR U7849 ( .A(b[3343]), .B(n3751), .Z(n3752) );
  XNOR U7850 ( .A(b[3343]), .B(n3753), .Z(c[3343]) );
  XOR U7851 ( .A(n3754), .B(n3755), .Z(n3751) );
  ANDN U7852 ( .B(n3756), .A(n3757), .Z(n3754) );
  XNOR U7853 ( .A(b[3342]), .B(n3755), .Z(n3756) );
  XNOR U7854 ( .A(b[3342]), .B(n3757), .Z(c[3342]) );
  XOR U7855 ( .A(n3758), .B(n3759), .Z(n3755) );
  ANDN U7856 ( .B(n3760), .A(n3761), .Z(n3758) );
  XNOR U7857 ( .A(b[3341]), .B(n3759), .Z(n3760) );
  XNOR U7858 ( .A(b[3341]), .B(n3761), .Z(c[3341]) );
  XOR U7859 ( .A(n3762), .B(n3763), .Z(n3759) );
  ANDN U7860 ( .B(n3764), .A(n3765), .Z(n3762) );
  XNOR U7861 ( .A(b[3340]), .B(n3763), .Z(n3764) );
  XNOR U7862 ( .A(b[3340]), .B(n3765), .Z(c[3340]) );
  XOR U7863 ( .A(n3766), .B(n3767), .Z(n3763) );
  ANDN U7864 ( .B(n3768), .A(n3769), .Z(n3766) );
  XNOR U7865 ( .A(b[3339]), .B(n3767), .Z(n3768) );
  XNOR U7866 ( .A(b[333]), .B(n3770), .Z(c[333]) );
  XNOR U7867 ( .A(b[3339]), .B(n3769), .Z(c[3339]) );
  XOR U7868 ( .A(n3771), .B(n3772), .Z(n3767) );
  ANDN U7869 ( .B(n3773), .A(n3774), .Z(n3771) );
  XNOR U7870 ( .A(b[3338]), .B(n3772), .Z(n3773) );
  XNOR U7871 ( .A(b[3338]), .B(n3774), .Z(c[3338]) );
  XOR U7872 ( .A(n3775), .B(n3776), .Z(n3772) );
  ANDN U7873 ( .B(n3777), .A(n3778), .Z(n3775) );
  XNOR U7874 ( .A(b[3337]), .B(n3776), .Z(n3777) );
  XNOR U7875 ( .A(b[3337]), .B(n3778), .Z(c[3337]) );
  XOR U7876 ( .A(n3779), .B(n3780), .Z(n3776) );
  ANDN U7877 ( .B(n3781), .A(n3782), .Z(n3779) );
  XNOR U7878 ( .A(b[3336]), .B(n3780), .Z(n3781) );
  XNOR U7879 ( .A(b[3336]), .B(n3782), .Z(c[3336]) );
  XOR U7880 ( .A(n3783), .B(n3784), .Z(n3780) );
  ANDN U7881 ( .B(n3785), .A(n3786), .Z(n3783) );
  XNOR U7882 ( .A(b[3335]), .B(n3784), .Z(n3785) );
  XNOR U7883 ( .A(b[3335]), .B(n3786), .Z(c[3335]) );
  XOR U7884 ( .A(n3787), .B(n3788), .Z(n3784) );
  ANDN U7885 ( .B(n3789), .A(n3790), .Z(n3787) );
  XNOR U7886 ( .A(b[3334]), .B(n3788), .Z(n3789) );
  XNOR U7887 ( .A(b[3334]), .B(n3790), .Z(c[3334]) );
  XOR U7888 ( .A(n3791), .B(n3792), .Z(n3788) );
  ANDN U7889 ( .B(n3793), .A(n3794), .Z(n3791) );
  XNOR U7890 ( .A(b[3333]), .B(n3792), .Z(n3793) );
  XNOR U7891 ( .A(b[3333]), .B(n3794), .Z(c[3333]) );
  XOR U7892 ( .A(n3795), .B(n3796), .Z(n3792) );
  ANDN U7893 ( .B(n3797), .A(n3798), .Z(n3795) );
  XNOR U7894 ( .A(b[3332]), .B(n3796), .Z(n3797) );
  XNOR U7895 ( .A(b[3332]), .B(n3798), .Z(c[3332]) );
  XOR U7896 ( .A(n3799), .B(n3800), .Z(n3796) );
  ANDN U7897 ( .B(n3801), .A(n3802), .Z(n3799) );
  XNOR U7898 ( .A(b[3331]), .B(n3800), .Z(n3801) );
  XNOR U7899 ( .A(b[3331]), .B(n3802), .Z(c[3331]) );
  XOR U7900 ( .A(n3803), .B(n3804), .Z(n3800) );
  ANDN U7901 ( .B(n3805), .A(n3806), .Z(n3803) );
  XNOR U7902 ( .A(b[3330]), .B(n3804), .Z(n3805) );
  XNOR U7903 ( .A(b[3330]), .B(n3806), .Z(c[3330]) );
  XOR U7904 ( .A(n3807), .B(n3808), .Z(n3804) );
  ANDN U7905 ( .B(n3809), .A(n3810), .Z(n3807) );
  XNOR U7906 ( .A(b[3329]), .B(n3808), .Z(n3809) );
  XNOR U7907 ( .A(b[332]), .B(n3811), .Z(c[332]) );
  XNOR U7908 ( .A(b[3329]), .B(n3810), .Z(c[3329]) );
  XOR U7909 ( .A(n3812), .B(n3813), .Z(n3808) );
  ANDN U7910 ( .B(n3814), .A(n3815), .Z(n3812) );
  XNOR U7911 ( .A(b[3328]), .B(n3813), .Z(n3814) );
  XNOR U7912 ( .A(b[3328]), .B(n3815), .Z(c[3328]) );
  XOR U7913 ( .A(n3816), .B(n3817), .Z(n3813) );
  ANDN U7914 ( .B(n3818), .A(n3819), .Z(n3816) );
  XNOR U7915 ( .A(b[3327]), .B(n3817), .Z(n3818) );
  XNOR U7916 ( .A(b[3327]), .B(n3819), .Z(c[3327]) );
  XOR U7917 ( .A(n3820), .B(n3821), .Z(n3817) );
  ANDN U7918 ( .B(n3822), .A(n3823), .Z(n3820) );
  XNOR U7919 ( .A(b[3326]), .B(n3821), .Z(n3822) );
  XNOR U7920 ( .A(b[3326]), .B(n3823), .Z(c[3326]) );
  XOR U7921 ( .A(n3824), .B(n3825), .Z(n3821) );
  ANDN U7922 ( .B(n3826), .A(n3827), .Z(n3824) );
  XNOR U7923 ( .A(b[3325]), .B(n3825), .Z(n3826) );
  XNOR U7924 ( .A(b[3325]), .B(n3827), .Z(c[3325]) );
  XOR U7925 ( .A(n3828), .B(n3829), .Z(n3825) );
  ANDN U7926 ( .B(n3830), .A(n3831), .Z(n3828) );
  XNOR U7927 ( .A(b[3324]), .B(n3829), .Z(n3830) );
  XNOR U7928 ( .A(b[3324]), .B(n3831), .Z(c[3324]) );
  XOR U7929 ( .A(n3832), .B(n3833), .Z(n3829) );
  ANDN U7930 ( .B(n3834), .A(n3835), .Z(n3832) );
  XNOR U7931 ( .A(b[3323]), .B(n3833), .Z(n3834) );
  XNOR U7932 ( .A(b[3323]), .B(n3835), .Z(c[3323]) );
  XOR U7933 ( .A(n3836), .B(n3837), .Z(n3833) );
  ANDN U7934 ( .B(n3838), .A(n3839), .Z(n3836) );
  XNOR U7935 ( .A(b[3322]), .B(n3837), .Z(n3838) );
  XNOR U7936 ( .A(b[3322]), .B(n3839), .Z(c[3322]) );
  XOR U7937 ( .A(n3840), .B(n3841), .Z(n3837) );
  ANDN U7938 ( .B(n3842), .A(n3843), .Z(n3840) );
  XNOR U7939 ( .A(b[3321]), .B(n3841), .Z(n3842) );
  XNOR U7940 ( .A(b[3321]), .B(n3843), .Z(c[3321]) );
  XOR U7941 ( .A(n3844), .B(n3845), .Z(n3841) );
  ANDN U7942 ( .B(n3846), .A(n3847), .Z(n3844) );
  XNOR U7943 ( .A(b[3320]), .B(n3845), .Z(n3846) );
  XNOR U7944 ( .A(b[3320]), .B(n3847), .Z(c[3320]) );
  XOR U7945 ( .A(n3848), .B(n3849), .Z(n3845) );
  ANDN U7946 ( .B(n3850), .A(n3851), .Z(n3848) );
  XNOR U7947 ( .A(b[3319]), .B(n3849), .Z(n3850) );
  XNOR U7948 ( .A(b[331]), .B(n3852), .Z(c[331]) );
  XNOR U7949 ( .A(b[3319]), .B(n3851), .Z(c[3319]) );
  XOR U7950 ( .A(n3853), .B(n3854), .Z(n3849) );
  ANDN U7951 ( .B(n3855), .A(n3856), .Z(n3853) );
  XNOR U7952 ( .A(b[3318]), .B(n3854), .Z(n3855) );
  XNOR U7953 ( .A(b[3318]), .B(n3856), .Z(c[3318]) );
  XOR U7954 ( .A(n3857), .B(n3858), .Z(n3854) );
  ANDN U7955 ( .B(n3859), .A(n3860), .Z(n3857) );
  XNOR U7956 ( .A(b[3317]), .B(n3858), .Z(n3859) );
  XNOR U7957 ( .A(b[3317]), .B(n3860), .Z(c[3317]) );
  XOR U7958 ( .A(n3861), .B(n3862), .Z(n3858) );
  ANDN U7959 ( .B(n3863), .A(n3864), .Z(n3861) );
  XNOR U7960 ( .A(b[3316]), .B(n3862), .Z(n3863) );
  XNOR U7961 ( .A(b[3316]), .B(n3864), .Z(c[3316]) );
  XOR U7962 ( .A(n3865), .B(n3866), .Z(n3862) );
  ANDN U7963 ( .B(n3867), .A(n3868), .Z(n3865) );
  XNOR U7964 ( .A(b[3315]), .B(n3866), .Z(n3867) );
  XNOR U7965 ( .A(b[3315]), .B(n3868), .Z(c[3315]) );
  XOR U7966 ( .A(n3869), .B(n3870), .Z(n3866) );
  ANDN U7967 ( .B(n3871), .A(n3872), .Z(n3869) );
  XNOR U7968 ( .A(b[3314]), .B(n3870), .Z(n3871) );
  XNOR U7969 ( .A(b[3314]), .B(n3872), .Z(c[3314]) );
  XOR U7970 ( .A(n3873), .B(n3874), .Z(n3870) );
  ANDN U7971 ( .B(n3875), .A(n3876), .Z(n3873) );
  XNOR U7972 ( .A(b[3313]), .B(n3874), .Z(n3875) );
  XNOR U7973 ( .A(b[3313]), .B(n3876), .Z(c[3313]) );
  XOR U7974 ( .A(n3877), .B(n3878), .Z(n3874) );
  ANDN U7975 ( .B(n3879), .A(n3880), .Z(n3877) );
  XNOR U7976 ( .A(b[3312]), .B(n3878), .Z(n3879) );
  XNOR U7977 ( .A(b[3312]), .B(n3880), .Z(c[3312]) );
  XOR U7978 ( .A(n3881), .B(n3882), .Z(n3878) );
  ANDN U7979 ( .B(n3883), .A(n3884), .Z(n3881) );
  XNOR U7980 ( .A(b[3311]), .B(n3882), .Z(n3883) );
  XNOR U7981 ( .A(b[3311]), .B(n3884), .Z(c[3311]) );
  XOR U7982 ( .A(n3885), .B(n3886), .Z(n3882) );
  ANDN U7983 ( .B(n3887), .A(n3888), .Z(n3885) );
  XNOR U7984 ( .A(b[3310]), .B(n3886), .Z(n3887) );
  XNOR U7985 ( .A(b[3310]), .B(n3888), .Z(c[3310]) );
  XOR U7986 ( .A(n3889), .B(n3890), .Z(n3886) );
  ANDN U7987 ( .B(n3891), .A(n3892), .Z(n3889) );
  XNOR U7988 ( .A(b[3309]), .B(n3890), .Z(n3891) );
  XNOR U7989 ( .A(b[330]), .B(n3893), .Z(c[330]) );
  XNOR U7990 ( .A(b[3309]), .B(n3892), .Z(c[3309]) );
  XOR U7991 ( .A(n3894), .B(n3895), .Z(n3890) );
  ANDN U7992 ( .B(n3896), .A(n3897), .Z(n3894) );
  XNOR U7993 ( .A(b[3308]), .B(n3895), .Z(n3896) );
  XNOR U7994 ( .A(b[3308]), .B(n3897), .Z(c[3308]) );
  XOR U7995 ( .A(n3898), .B(n3899), .Z(n3895) );
  ANDN U7996 ( .B(n3900), .A(n3901), .Z(n3898) );
  XNOR U7997 ( .A(b[3307]), .B(n3899), .Z(n3900) );
  XNOR U7998 ( .A(b[3307]), .B(n3901), .Z(c[3307]) );
  XOR U7999 ( .A(n3902), .B(n3903), .Z(n3899) );
  ANDN U8000 ( .B(n3904), .A(n3905), .Z(n3902) );
  XNOR U8001 ( .A(b[3306]), .B(n3903), .Z(n3904) );
  XNOR U8002 ( .A(b[3306]), .B(n3905), .Z(c[3306]) );
  XOR U8003 ( .A(n3906), .B(n3907), .Z(n3903) );
  ANDN U8004 ( .B(n3908), .A(n3909), .Z(n3906) );
  XNOR U8005 ( .A(b[3305]), .B(n3907), .Z(n3908) );
  XNOR U8006 ( .A(b[3305]), .B(n3909), .Z(c[3305]) );
  XOR U8007 ( .A(n3910), .B(n3911), .Z(n3907) );
  ANDN U8008 ( .B(n3912), .A(n3913), .Z(n3910) );
  XNOR U8009 ( .A(b[3304]), .B(n3911), .Z(n3912) );
  XNOR U8010 ( .A(b[3304]), .B(n3913), .Z(c[3304]) );
  XOR U8011 ( .A(n3914), .B(n3915), .Z(n3911) );
  ANDN U8012 ( .B(n3916), .A(n3917), .Z(n3914) );
  XNOR U8013 ( .A(b[3303]), .B(n3915), .Z(n3916) );
  XNOR U8014 ( .A(b[3303]), .B(n3917), .Z(c[3303]) );
  XOR U8015 ( .A(n3918), .B(n3919), .Z(n3915) );
  ANDN U8016 ( .B(n3920), .A(n3921), .Z(n3918) );
  XNOR U8017 ( .A(b[3302]), .B(n3919), .Z(n3920) );
  XNOR U8018 ( .A(b[3302]), .B(n3921), .Z(c[3302]) );
  XOR U8019 ( .A(n3922), .B(n3923), .Z(n3919) );
  ANDN U8020 ( .B(n3924), .A(n3925), .Z(n3922) );
  XNOR U8021 ( .A(b[3301]), .B(n3923), .Z(n3924) );
  XNOR U8022 ( .A(b[3301]), .B(n3925), .Z(c[3301]) );
  XOR U8023 ( .A(n3926), .B(n3927), .Z(n3923) );
  ANDN U8024 ( .B(n3928), .A(n3929), .Z(n3926) );
  XNOR U8025 ( .A(b[3300]), .B(n3927), .Z(n3928) );
  XNOR U8026 ( .A(b[3300]), .B(n3929), .Z(c[3300]) );
  XOR U8027 ( .A(n3930), .B(n3931), .Z(n3927) );
  ANDN U8028 ( .B(n3932), .A(n3933), .Z(n3930) );
  XNOR U8029 ( .A(b[3299]), .B(n3931), .Z(n3932) );
  XNOR U8030 ( .A(b[32]), .B(n3934), .Z(c[32]) );
  XNOR U8031 ( .A(b[329]), .B(n3935), .Z(c[329]) );
  XNOR U8032 ( .A(b[3299]), .B(n3933), .Z(c[3299]) );
  XOR U8033 ( .A(n3936), .B(n3937), .Z(n3931) );
  ANDN U8034 ( .B(n3938), .A(n3939), .Z(n3936) );
  XNOR U8035 ( .A(b[3298]), .B(n3937), .Z(n3938) );
  XNOR U8036 ( .A(b[3298]), .B(n3939), .Z(c[3298]) );
  XOR U8037 ( .A(n3940), .B(n3941), .Z(n3937) );
  ANDN U8038 ( .B(n3942), .A(n3943), .Z(n3940) );
  XNOR U8039 ( .A(b[3297]), .B(n3941), .Z(n3942) );
  XNOR U8040 ( .A(b[3297]), .B(n3943), .Z(c[3297]) );
  XOR U8041 ( .A(n3944), .B(n3945), .Z(n3941) );
  ANDN U8042 ( .B(n3946), .A(n3947), .Z(n3944) );
  XNOR U8043 ( .A(b[3296]), .B(n3945), .Z(n3946) );
  XNOR U8044 ( .A(b[3296]), .B(n3947), .Z(c[3296]) );
  XOR U8045 ( .A(n3948), .B(n3949), .Z(n3945) );
  ANDN U8046 ( .B(n3950), .A(n3951), .Z(n3948) );
  XNOR U8047 ( .A(b[3295]), .B(n3949), .Z(n3950) );
  XNOR U8048 ( .A(b[3295]), .B(n3951), .Z(c[3295]) );
  XOR U8049 ( .A(n3952), .B(n3953), .Z(n3949) );
  ANDN U8050 ( .B(n3954), .A(n3955), .Z(n3952) );
  XNOR U8051 ( .A(b[3294]), .B(n3953), .Z(n3954) );
  XNOR U8052 ( .A(b[3294]), .B(n3955), .Z(c[3294]) );
  XOR U8053 ( .A(n3956), .B(n3957), .Z(n3953) );
  ANDN U8054 ( .B(n3958), .A(n3959), .Z(n3956) );
  XNOR U8055 ( .A(b[3293]), .B(n3957), .Z(n3958) );
  XNOR U8056 ( .A(b[3293]), .B(n3959), .Z(c[3293]) );
  XOR U8057 ( .A(n3960), .B(n3961), .Z(n3957) );
  ANDN U8058 ( .B(n3962), .A(n3963), .Z(n3960) );
  XNOR U8059 ( .A(b[3292]), .B(n3961), .Z(n3962) );
  XNOR U8060 ( .A(b[3292]), .B(n3963), .Z(c[3292]) );
  XOR U8061 ( .A(n3964), .B(n3965), .Z(n3961) );
  ANDN U8062 ( .B(n3966), .A(n3967), .Z(n3964) );
  XNOR U8063 ( .A(b[3291]), .B(n3965), .Z(n3966) );
  XNOR U8064 ( .A(b[3291]), .B(n3967), .Z(c[3291]) );
  XOR U8065 ( .A(n3968), .B(n3969), .Z(n3965) );
  ANDN U8066 ( .B(n3970), .A(n3971), .Z(n3968) );
  XNOR U8067 ( .A(b[3290]), .B(n3969), .Z(n3970) );
  XNOR U8068 ( .A(b[3290]), .B(n3971), .Z(c[3290]) );
  XOR U8069 ( .A(n3972), .B(n3973), .Z(n3969) );
  ANDN U8070 ( .B(n3974), .A(n3975), .Z(n3972) );
  XNOR U8071 ( .A(b[3289]), .B(n3973), .Z(n3974) );
  XNOR U8072 ( .A(b[328]), .B(n3976), .Z(c[328]) );
  XNOR U8073 ( .A(b[3289]), .B(n3975), .Z(c[3289]) );
  XOR U8074 ( .A(n3977), .B(n3978), .Z(n3973) );
  ANDN U8075 ( .B(n3979), .A(n3980), .Z(n3977) );
  XNOR U8076 ( .A(b[3288]), .B(n3978), .Z(n3979) );
  XNOR U8077 ( .A(b[3288]), .B(n3980), .Z(c[3288]) );
  XOR U8078 ( .A(n3981), .B(n3982), .Z(n3978) );
  ANDN U8079 ( .B(n3983), .A(n3984), .Z(n3981) );
  XNOR U8080 ( .A(b[3287]), .B(n3982), .Z(n3983) );
  XNOR U8081 ( .A(b[3287]), .B(n3984), .Z(c[3287]) );
  XOR U8082 ( .A(n3985), .B(n3986), .Z(n3982) );
  ANDN U8083 ( .B(n3987), .A(n3988), .Z(n3985) );
  XNOR U8084 ( .A(b[3286]), .B(n3986), .Z(n3987) );
  XNOR U8085 ( .A(b[3286]), .B(n3988), .Z(c[3286]) );
  XOR U8086 ( .A(n3989), .B(n3990), .Z(n3986) );
  ANDN U8087 ( .B(n3991), .A(n3992), .Z(n3989) );
  XNOR U8088 ( .A(b[3285]), .B(n3990), .Z(n3991) );
  XNOR U8089 ( .A(b[3285]), .B(n3992), .Z(c[3285]) );
  XOR U8090 ( .A(n3993), .B(n3994), .Z(n3990) );
  ANDN U8091 ( .B(n3995), .A(n3996), .Z(n3993) );
  XNOR U8092 ( .A(b[3284]), .B(n3994), .Z(n3995) );
  XNOR U8093 ( .A(b[3284]), .B(n3996), .Z(c[3284]) );
  XOR U8094 ( .A(n3997), .B(n3998), .Z(n3994) );
  ANDN U8095 ( .B(n3999), .A(n4000), .Z(n3997) );
  XNOR U8096 ( .A(b[3283]), .B(n3998), .Z(n3999) );
  XNOR U8097 ( .A(b[3283]), .B(n4000), .Z(c[3283]) );
  XOR U8098 ( .A(n4001), .B(n4002), .Z(n3998) );
  ANDN U8099 ( .B(n4003), .A(n4004), .Z(n4001) );
  XNOR U8100 ( .A(b[3282]), .B(n4002), .Z(n4003) );
  XNOR U8101 ( .A(b[3282]), .B(n4004), .Z(c[3282]) );
  XOR U8102 ( .A(n4005), .B(n4006), .Z(n4002) );
  ANDN U8103 ( .B(n4007), .A(n4008), .Z(n4005) );
  XNOR U8104 ( .A(b[3281]), .B(n4006), .Z(n4007) );
  XNOR U8105 ( .A(b[3281]), .B(n4008), .Z(c[3281]) );
  XOR U8106 ( .A(n4009), .B(n4010), .Z(n4006) );
  ANDN U8107 ( .B(n4011), .A(n4012), .Z(n4009) );
  XNOR U8108 ( .A(b[3280]), .B(n4010), .Z(n4011) );
  XNOR U8109 ( .A(b[3280]), .B(n4012), .Z(c[3280]) );
  XOR U8110 ( .A(n4013), .B(n4014), .Z(n4010) );
  ANDN U8111 ( .B(n4015), .A(n4016), .Z(n4013) );
  XNOR U8112 ( .A(b[3279]), .B(n4014), .Z(n4015) );
  XNOR U8113 ( .A(b[327]), .B(n4017), .Z(c[327]) );
  XNOR U8114 ( .A(b[3279]), .B(n4016), .Z(c[3279]) );
  XOR U8115 ( .A(n4018), .B(n4019), .Z(n4014) );
  ANDN U8116 ( .B(n4020), .A(n4021), .Z(n4018) );
  XNOR U8117 ( .A(b[3278]), .B(n4019), .Z(n4020) );
  XNOR U8118 ( .A(b[3278]), .B(n4021), .Z(c[3278]) );
  XOR U8119 ( .A(n4022), .B(n4023), .Z(n4019) );
  ANDN U8120 ( .B(n4024), .A(n4025), .Z(n4022) );
  XNOR U8121 ( .A(b[3277]), .B(n4023), .Z(n4024) );
  XNOR U8122 ( .A(b[3277]), .B(n4025), .Z(c[3277]) );
  XOR U8123 ( .A(n4026), .B(n4027), .Z(n4023) );
  ANDN U8124 ( .B(n4028), .A(n4029), .Z(n4026) );
  XNOR U8125 ( .A(b[3276]), .B(n4027), .Z(n4028) );
  XNOR U8126 ( .A(b[3276]), .B(n4029), .Z(c[3276]) );
  XOR U8127 ( .A(n4030), .B(n4031), .Z(n4027) );
  ANDN U8128 ( .B(n4032), .A(n4033), .Z(n4030) );
  XNOR U8129 ( .A(b[3275]), .B(n4031), .Z(n4032) );
  XNOR U8130 ( .A(b[3275]), .B(n4033), .Z(c[3275]) );
  XOR U8131 ( .A(n4034), .B(n4035), .Z(n4031) );
  ANDN U8132 ( .B(n4036), .A(n4037), .Z(n4034) );
  XNOR U8133 ( .A(b[3274]), .B(n4035), .Z(n4036) );
  XNOR U8134 ( .A(b[3274]), .B(n4037), .Z(c[3274]) );
  XOR U8135 ( .A(n4038), .B(n4039), .Z(n4035) );
  ANDN U8136 ( .B(n4040), .A(n4041), .Z(n4038) );
  XNOR U8137 ( .A(b[3273]), .B(n4039), .Z(n4040) );
  XNOR U8138 ( .A(b[3273]), .B(n4041), .Z(c[3273]) );
  XOR U8139 ( .A(n4042), .B(n4043), .Z(n4039) );
  ANDN U8140 ( .B(n4044), .A(n4045), .Z(n4042) );
  XNOR U8141 ( .A(b[3272]), .B(n4043), .Z(n4044) );
  XNOR U8142 ( .A(b[3272]), .B(n4045), .Z(c[3272]) );
  XOR U8143 ( .A(n4046), .B(n4047), .Z(n4043) );
  ANDN U8144 ( .B(n4048), .A(n4049), .Z(n4046) );
  XNOR U8145 ( .A(b[3271]), .B(n4047), .Z(n4048) );
  XNOR U8146 ( .A(b[3271]), .B(n4049), .Z(c[3271]) );
  XOR U8147 ( .A(n4050), .B(n4051), .Z(n4047) );
  ANDN U8148 ( .B(n4052), .A(n4053), .Z(n4050) );
  XNOR U8149 ( .A(b[3270]), .B(n4051), .Z(n4052) );
  XNOR U8150 ( .A(b[3270]), .B(n4053), .Z(c[3270]) );
  XOR U8151 ( .A(n4054), .B(n4055), .Z(n4051) );
  ANDN U8152 ( .B(n4056), .A(n4057), .Z(n4054) );
  XNOR U8153 ( .A(b[3269]), .B(n4055), .Z(n4056) );
  XNOR U8154 ( .A(b[326]), .B(n4058), .Z(c[326]) );
  XNOR U8155 ( .A(b[3269]), .B(n4057), .Z(c[3269]) );
  XOR U8156 ( .A(n4059), .B(n4060), .Z(n4055) );
  ANDN U8157 ( .B(n4061), .A(n4062), .Z(n4059) );
  XNOR U8158 ( .A(b[3268]), .B(n4060), .Z(n4061) );
  XNOR U8159 ( .A(b[3268]), .B(n4062), .Z(c[3268]) );
  XOR U8160 ( .A(n4063), .B(n4064), .Z(n4060) );
  ANDN U8161 ( .B(n4065), .A(n4066), .Z(n4063) );
  XNOR U8162 ( .A(b[3267]), .B(n4064), .Z(n4065) );
  XNOR U8163 ( .A(b[3267]), .B(n4066), .Z(c[3267]) );
  XOR U8164 ( .A(n4067), .B(n4068), .Z(n4064) );
  ANDN U8165 ( .B(n4069), .A(n4070), .Z(n4067) );
  XNOR U8166 ( .A(b[3266]), .B(n4068), .Z(n4069) );
  XNOR U8167 ( .A(b[3266]), .B(n4070), .Z(c[3266]) );
  XOR U8168 ( .A(n4071), .B(n4072), .Z(n4068) );
  ANDN U8169 ( .B(n4073), .A(n4074), .Z(n4071) );
  XNOR U8170 ( .A(b[3265]), .B(n4072), .Z(n4073) );
  XNOR U8171 ( .A(b[3265]), .B(n4074), .Z(c[3265]) );
  XOR U8172 ( .A(n4075), .B(n4076), .Z(n4072) );
  ANDN U8173 ( .B(n4077), .A(n4078), .Z(n4075) );
  XNOR U8174 ( .A(b[3264]), .B(n4076), .Z(n4077) );
  XNOR U8175 ( .A(b[3264]), .B(n4078), .Z(c[3264]) );
  XOR U8176 ( .A(n4079), .B(n4080), .Z(n4076) );
  ANDN U8177 ( .B(n4081), .A(n4082), .Z(n4079) );
  XNOR U8178 ( .A(b[3263]), .B(n4080), .Z(n4081) );
  XNOR U8179 ( .A(b[3263]), .B(n4082), .Z(c[3263]) );
  XOR U8180 ( .A(n4083), .B(n4084), .Z(n4080) );
  ANDN U8181 ( .B(n4085), .A(n4086), .Z(n4083) );
  XNOR U8182 ( .A(b[3262]), .B(n4084), .Z(n4085) );
  XNOR U8183 ( .A(b[3262]), .B(n4086), .Z(c[3262]) );
  XOR U8184 ( .A(n4087), .B(n4088), .Z(n4084) );
  ANDN U8185 ( .B(n4089), .A(n4090), .Z(n4087) );
  XNOR U8186 ( .A(b[3261]), .B(n4088), .Z(n4089) );
  XNOR U8187 ( .A(b[3261]), .B(n4090), .Z(c[3261]) );
  XOR U8188 ( .A(n4091), .B(n4092), .Z(n4088) );
  ANDN U8189 ( .B(n4093), .A(n4094), .Z(n4091) );
  XNOR U8190 ( .A(b[3260]), .B(n4092), .Z(n4093) );
  XNOR U8191 ( .A(b[3260]), .B(n4094), .Z(c[3260]) );
  XOR U8192 ( .A(n4095), .B(n4096), .Z(n4092) );
  ANDN U8193 ( .B(n4097), .A(n4098), .Z(n4095) );
  XNOR U8194 ( .A(b[3259]), .B(n4096), .Z(n4097) );
  XNOR U8195 ( .A(b[325]), .B(n4099), .Z(c[325]) );
  XNOR U8196 ( .A(b[3259]), .B(n4098), .Z(c[3259]) );
  XOR U8197 ( .A(n4100), .B(n4101), .Z(n4096) );
  ANDN U8198 ( .B(n4102), .A(n4103), .Z(n4100) );
  XNOR U8199 ( .A(b[3258]), .B(n4101), .Z(n4102) );
  XNOR U8200 ( .A(b[3258]), .B(n4103), .Z(c[3258]) );
  XOR U8201 ( .A(n4104), .B(n4105), .Z(n4101) );
  ANDN U8202 ( .B(n4106), .A(n4107), .Z(n4104) );
  XNOR U8203 ( .A(b[3257]), .B(n4105), .Z(n4106) );
  XNOR U8204 ( .A(b[3257]), .B(n4107), .Z(c[3257]) );
  XOR U8205 ( .A(n4108), .B(n4109), .Z(n4105) );
  ANDN U8206 ( .B(n4110), .A(n4111), .Z(n4108) );
  XNOR U8207 ( .A(b[3256]), .B(n4109), .Z(n4110) );
  XNOR U8208 ( .A(b[3256]), .B(n4111), .Z(c[3256]) );
  XOR U8209 ( .A(n4112), .B(n4113), .Z(n4109) );
  ANDN U8210 ( .B(n4114), .A(n4115), .Z(n4112) );
  XNOR U8211 ( .A(b[3255]), .B(n4113), .Z(n4114) );
  XNOR U8212 ( .A(b[3255]), .B(n4115), .Z(c[3255]) );
  XOR U8213 ( .A(n4116), .B(n4117), .Z(n4113) );
  ANDN U8214 ( .B(n4118), .A(n4119), .Z(n4116) );
  XNOR U8215 ( .A(b[3254]), .B(n4117), .Z(n4118) );
  XNOR U8216 ( .A(b[3254]), .B(n4119), .Z(c[3254]) );
  XOR U8217 ( .A(n4120), .B(n4121), .Z(n4117) );
  ANDN U8218 ( .B(n4122), .A(n4123), .Z(n4120) );
  XNOR U8219 ( .A(b[3253]), .B(n4121), .Z(n4122) );
  XNOR U8220 ( .A(b[3253]), .B(n4123), .Z(c[3253]) );
  XOR U8221 ( .A(n4124), .B(n4125), .Z(n4121) );
  ANDN U8222 ( .B(n4126), .A(n4127), .Z(n4124) );
  XNOR U8223 ( .A(b[3252]), .B(n4125), .Z(n4126) );
  XNOR U8224 ( .A(b[3252]), .B(n4127), .Z(c[3252]) );
  XOR U8225 ( .A(n4128), .B(n4129), .Z(n4125) );
  ANDN U8226 ( .B(n4130), .A(n4131), .Z(n4128) );
  XNOR U8227 ( .A(b[3251]), .B(n4129), .Z(n4130) );
  XNOR U8228 ( .A(b[3251]), .B(n4131), .Z(c[3251]) );
  XOR U8229 ( .A(n4132), .B(n4133), .Z(n4129) );
  ANDN U8230 ( .B(n4134), .A(n4135), .Z(n4132) );
  XNOR U8231 ( .A(b[3250]), .B(n4133), .Z(n4134) );
  XNOR U8232 ( .A(b[3250]), .B(n4135), .Z(c[3250]) );
  XOR U8233 ( .A(n4136), .B(n4137), .Z(n4133) );
  ANDN U8234 ( .B(n4138), .A(n4139), .Z(n4136) );
  XNOR U8235 ( .A(b[3249]), .B(n4137), .Z(n4138) );
  XNOR U8236 ( .A(b[324]), .B(n4140), .Z(c[324]) );
  XNOR U8237 ( .A(b[3249]), .B(n4139), .Z(c[3249]) );
  XOR U8238 ( .A(n4141), .B(n4142), .Z(n4137) );
  ANDN U8239 ( .B(n4143), .A(n4144), .Z(n4141) );
  XNOR U8240 ( .A(b[3248]), .B(n4142), .Z(n4143) );
  XNOR U8241 ( .A(b[3248]), .B(n4144), .Z(c[3248]) );
  XOR U8242 ( .A(n4145), .B(n4146), .Z(n4142) );
  ANDN U8243 ( .B(n4147), .A(n4148), .Z(n4145) );
  XNOR U8244 ( .A(b[3247]), .B(n4146), .Z(n4147) );
  XNOR U8245 ( .A(b[3247]), .B(n4148), .Z(c[3247]) );
  XOR U8246 ( .A(n4149), .B(n4150), .Z(n4146) );
  ANDN U8247 ( .B(n4151), .A(n4152), .Z(n4149) );
  XNOR U8248 ( .A(b[3246]), .B(n4150), .Z(n4151) );
  XNOR U8249 ( .A(b[3246]), .B(n4152), .Z(c[3246]) );
  XOR U8250 ( .A(n4153), .B(n4154), .Z(n4150) );
  ANDN U8251 ( .B(n4155), .A(n4156), .Z(n4153) );
  XNOR U8252 ( .A(b[3245]), .B(n4154), .Z(n4155) );
  XNOR U8253 ( .A(b[3245]), .B(n4156), .Z(c[3245]) );
  XOR U8254 ( .A(n4157), .B(n4158), .Z(n4154) );
  ANDN U8255 ( .B(n4159), .A(n4160), .Z(n4157) );
  XNOR U8256 ( .A(b[3244]), .B(n4158), .Z(n4159) );
  XNOR U8257 ( .A(b[3244]), .B(n4160), .Z(c[3244]) );
  XOR U8258 ( .A(n4161), .B(n4162), .Z(n4158) );
  ANDN U8259 ( .B(n4163), .A(n4164), .Z(n4161) );
  XNOR U8260 ( .A(b[3243]), .B(n4162), .Z(n4163) );
  XNOR U8261 ( .A(b[3243]), .B(n4164), .Z(c[3243]) );
  XOR U8262 ( .A(n4165), .B(n4166), .Z(n4162) );
  ANDN U8263 ( .B(n4167), .A(n4168), .Z(n4165) );
  XNOR U8264 ( .A(b[3242]), .B(n4166), .Z(n4167) );
  XNOR U8265 ( .A(b[3242]), .B(n4168), .Z(c[3242]) );
  XOR U8266 ( .A(n4169), .B(n4170), .Z(n4166) );
  ANDN U8267 ( .B(n4171), .A(n4172), .Z(n4169) );
  XNOR U8268 ( .A(b[3241]), .B(n4170), .Z(n4171) );
  XNOR U8269 ( .A(b[3241]), .B(n4172), .Z(c[3241]) );
  XOR U8270 ( .A(n4173), .B(n4174), .Z(n4170) );
  ANDN U8271 ( .B(n4175), .A(n4176), .Z(n4173) );
  XNOR U8272 ( .A(b[3240]), .B(n4174), .Z(n4175) );
  XNOR U8273 ( .A(b[3240]), .B(n4176), .Z(c[3240]) );
  XOR U8274 ( .A(n4177), .B(n4178), .Z(n4174) );
  ANDN U8275 ( .B(n4179), .A(n4180), .Z(n4177) );
  XNOR U8276 ( .A(b[3239]), .B(n4178), .Z(n4179) );
  XNOR U8277 ( .A(b[323]), .B(n4181), .Z(c[323]) );
  XNOR U8278 ( .A(b[3239]), .B(n4180), .Z(c[3239]) );
  XOR U8279 ( .A(n4182), .B(n4183), .Z(n4178) );
  ANDN U8280 ( .B(n4184), .A(n4185), .Z(n4182) );
  XNOR U8281 ( .A(b[3238]), .B(n4183), .Z(n4184) );
  XNOR U8282 ( .A(b[3238]), .B(n4185), .Z(c[3238]) );
  XOR U8283 ( .A(n4186), .B(n4187), .Z(n4183) );
  ANDN U8284 ( .B(n4188), .A(n4189), .Z(n4186) );
  XNOR U8285 ( .A(b[3237]), .B(n4187), .Z(n4188) );
  XNOR U8286 ( .A(b[3237]), .B(n4189), .Z(c[3237]) );
  XOR U8287 ( .A(n4190), .B(n4191), .Z(n4187) );
  ANDN U8288 ( .B(n4192), .A(n4193), .Z(n4190) );
  XNOR U8289 ( .A(b[3236]), .B(n4191), .Z(n4192) );
  XNOR U8290 ( .A(b[3236]), .B(n4193), .Z(c[3236]) );
  XOR U8291 ( .A(n4194), .B(n4195), .Z(n4191) );
  ANDN U8292 ( .B(n4196), .A(n4197), .Z(n4194) );
  XNOR U8293 ( .A(b[3235]), .B(n4195), .Z(n4196) );
  XNOR U8294 ( .A(b[3235]), .B(n4197), .Z(c[3235]) );
  XOR U8295 ( .A(n4198), .B(n4199), .Z(n4195) );
  ANDN U8296 ( .B(n4200), .A(n4201), .Z(n4198) );
  XNOR U8297 ( .A(b[3234]), .B(n4199), .Z(n4200) );
  XNOR U8298 ( .A(b[3234]), .B(n4201), .Z(c[3234]) );
  XOR U8299 ( .A(n4202), .B(n4203), .Z(n4199) );
  ANDN U8300 ( .B(n4204), .A(n4205), .Z(n4202) );
  XNOR U8301 ( .A(b[3233]), .B(n4203), .Z(n4204) );
  XNOR U8302 ( .A(b[3233]), .B(n4205), .Z(c[3233]) );
  XOR U8303 ( .A(n4206), .B(n4207), .Z(n4203) );
  ANDN U8304 ( .B(n4208), .A(n4209), .Z(n4206) );
  XNOR U8305 ( .A(b[3232]), .B(n4207), .Z(n4208) );
  XNOR U8306 ( .A(b[3232]), .B(n4209), .Z(c[3232]) );
  XOR U8307 ( .A(n4210), .B(n4211), .Z(n4207) );
  ANDN U8308 ( .B(n4212), .A(n4213), .Z(n4210) );
  XNOR U8309 ( .A(b[3231]), .B(n4211), .Z(n4212) );
  XNOR U8310 ( .A(b[3231]), .B(n4213), .Z(c[3231]) );
  XOR U8311 ( .A(n4214), .B(n4215), .Z(n4211) );
  ANDN U8312 ( .B(n4216), .A(n4217), .Z(n4214) );
  XNOR U8313 ( .A(b[3230]), .B(n4215), .Z(n4216) );
  XNOR U8314 ( .A(b[3230]), .B(n4217), .Z(c[3230]) );
  XOR U8315 ( .A(n4218), .B(n4219), .Z(n4215) );
  ANDN U8316 ( .B(n4220), .A(n4221), .Z(n4218) );
  XNOR U8317 ( .A(b[3229]), .B(n4219), .Z(n4220) );
  XNOR U8318 ( .A(b[322]), .B(n4222), .Z(c[322]) );
  XNOR U8319 ( .A(b[3229]), .B(n4221), .Z(c[3229]) );
  XOR U8320 ( .A(n4223), .B(n4224), .Z(n4219) );
  ANDN U8321 ( .B(n4225), .A(n4226), .Z(n4223) );
  XNOR U8322 ( .A(b[3228]), .B(n4224), .Z(n4225) );
  XNOR U8323 ( .A(b[3228]), .B(n4226), .Z(c[3228]) );
  XOR U8324 ( .A(n4227), .B(n4228), .Z(n4224) );
  ANDN U8325 ( .B(n4229), .A(n4230), .Z(n4227) );
  XNOR U8326 ( .A(b[3227]), .B(n4228), .Z(n4229) );
  XNOR U8327 ( .A(b[3227]), .B(n4230), .Z(c[3227]) );
  XOR U8328 ( .A(n4231), .B(n4232), .Z(n4228) );
  ANDN U8329 ( .B(n4233), .A(n4234), .Z(n4231) );
  XNOR U8330 ( .A(b[3226]), .B(n4232), .Z(n4233) );
  XNOR U8331 ( .A(b[3226]), .B(n4234), .Z(c[3226]) );
  XOR U8332 ( .A(n4235), .B(n4236), .Z(n4232) );
  ANDN U8333 ( .B(n4237), .A(n4238), .Z(n4235) );
  XNOR U8334 ( .A(b[3225]), .B(n4236), .Z(n4237) );
  XNOR U8335 ( .A(b[3225]), .B(n4238), .Z(c[3225]) );
  XOR U8336 ( .A(n4239), .B(n4240), .Z(n4236) );
  ANDN U8337 ( .B(n4241), .A(n4242), .Z(n4239) );
  XNOR U8338 ( .A(b[3224]), .B(n4240), .Z(n4241) );
  XNOR U8339 ( .A(b[3224]), .B(n4242), .Z(c[3224]) );
  XOR U8340 ( .A(n4243), .B(n4244), .Z(n4240) );
  ANDN U8341 ( .B(n4245), .A(n4246), .Z(n4243) );
  XNOR U8342 ( .A(b[3223]), .B(n4244), .Z(n4245) );
  XNOR U8343 ( .A(b[3223]), .B(n4246), .Z(c[3223]) );
  XOR U8344 ( .A(n4247), .B(n4248), .Z(n4244) );
  ANDN U8345 ( .B(n4249), .A(n4250), .Z(n4247) );
  XNOR U8346 ( .A(b[3222]), .B(n4248), .Z(n4249) );
  XNOR U8347 ( .A(b[3222]), .B(n4250), .Z(c[3222]) );
  XOR U8348 ( .A(n4251), .B(n4252), .Z(n4248) );
  ANDN U8349 ( .B(n4253), .A(n4254), .Z(n4251) );
  XNOR U8350 ( .A(b[3221]), .B(n4252), .Z(n4253) );
  XNOR U8351 ( .A(b[3221]), .B(n4254), .Z(c[3221]) );
  XOR U8352 ( .A(n4255), .B(n4256), .Z(n4252) );
  ANDN U8353 ( .B(n4257), .A(n4258), .Z(n4255) );
  XNOR U8354 ( .A(b[3220]), .B(n4256), .Z(n4257) );
  XNOR U8355 ( .A(b[3220]), .B(n4258), .Z(c[3220]) );
  XOR U8356 ( .A(n4259), .B(n4260), .Z(n4256) );
  ANDN U8357 ( .B(n4261), .A(n4262), .Z(n4259) );
  XNOR U8358 ( .A(b[3219]), .B(n4260), .Z(n4261) );
  XNOR U8359 ( .A(b[321]), .B(n4263), .Z(c[321]) );
  XNOR U8360 ( .A(b[3219]), .B(n4262), .Z(c[3219]) );
  XOR U8361 ( .A(n4264), .B(n4265), .Z(n4260) );
  ANDN U8362 ( .B(n4266), .A(n4267), .Z(n4264) );
  XNOR U8363 ( .A(b[3218]), .B(n4265), .Z(n4266) );
  XNOR U8364 ( .A(b[3218]), .B(n4267), .Z(c[3218]) );
  XOR U8365 ( .A(n4268), .B(n4269), .Z(n4265) );
  ANDN U8366 ( .B(n4270), .A(n4271), .Z(n4268) );
  XNOR U8367 ( .A(b[3217]), .B(n4269), .Z(n4270) );
  XNOR U8368 ( .A(b[3217]), .B(n4271), .Z(c[3217]) );
  XOR U8369 ( .A(n4272), .B(n4273), .Z(n4269) );
  ANDN U8370 ( .B(n4274), .A(n4275), .Z(n4272) );
  XNOR U8371 ( .A(b[3216]), .B(n4273), .Z(n4274) );
  XNOR U8372 ( .A(b[3216]), .B(n4275), .Z(c[3216]) );
  XOR U8373 ( .A(n4276), .B(n4277), .Z(n4273) );
  ANDN U8374 ( .B(n4278), .A(n4279), .Z(n4276) );
  XNOR U8375 ( .A(b[3215]), .B(n4277), .Z(n4278) );
  XNOR U8376 ( .A(b[3215]), .B(n4279), .Z(c[3215]) );
  XOR U8377 ( .A(n4280), .B(n4281), .Z(n4277) );
  ANDN U8378 ( .B(n4282), .A(n4283), .Z(n4280) );
  XNOR U8379 ( .A(b[3214]), .B(n4281), .Z(n4282) );
  XNOR U8380 ( .A(b[3214]), .B(n4283), .Z(c[3214]) );
  XOR U8381 ( .A(n4284), .B(n4285), .Z(n4281) );
  ANDN U8382 ( .B(n4286), .A(n4287), .Z(n4284) );
  XNOR U8383 ( .A(b[3213]), .B(n4285), .Z(n4286) );
  XNOR U8384 ( .A(b[3213]), .B(n4287), .Z(c[3213]) );
  XOR U8385 ( .A(n4288), .B(n4289), .Z(n4285) );
  ANDN U8386 ( .B(n4290), .A(n4291), .Z(n4288) );
  XNOR U8387 ( .A(b[3212]), .B(n4289), .Z(n4290) );
  XNOR U8388 ( .A(b[3212]), .B(n4291), .Z(c[3212]) );
  XOR U8389 ( .A(n4292), .B(n4293), .Z(n4289) );
  ANDN U8390 ( .B(n4294), .A(n4295), .Z(n4292) );
  XNOR U8391 ( .A(b[3211]), .B(n4293), .Z(n4294) );
  XNOR U8392 ( .A(b[3211]), .B(n4295), .Z(c[3211]) );
  XOR U8393 ( .A(n4296), .B(n4297), .Z(n4293) );
  ANDN U8394 ( .B(n4298), .A(n4299), .Z(n4296) );
  XNOR U8395 ( .A(b[3210]), .B(n4297), .Z(n4298) );
  XNOR U8396 ( .A(b[3210]), .B(n4299), .Z(c[3210]) );
  XOR U8397 ( .A(n4300), .B(n4301), .Z(n4297) );
  ANDN U8398 ( .B(n4302), .A(n4303), .Z(n4300) );
  XNOR U8399 ( .A(b[3209]), .B(n4301), .Z(n4302) );
  XNOR U8400 ( .A(b[320]), .B(n4304), .Z(c[320]) );
  XNOR U8401 ( .A(b[3209]), .B(n4303), .Z(c[3209]) );
  XOR U8402 ( .A(n4305), .B(n4306), .Z(n4301) );
  ANDN U8403 ( .B(n4307), .A(n4308), .Z(n4305) );
  XNOR U8404 ( .A(b[3208]), .B(n4306), .Z(n4307) );
  XNOR U8405 ( .A(b[3208]), .B(n4308), .Z(c[3208]) );
  XOR U8406 ( .A(n4309), .B(n4310), .Z(n4306) );
  ANDN U8407 ( .B(n4311), .A(n4312), .Z(n4309) );
  XNOR U8408 ( .A(b[3207]), .B(n4310), .Z(n4311) );
  XNOR U8409 ( .A(b[3207]), .B(n4312), .Z(c[3207]) );
  XOR U8410 ( .A(n4313), .B(n4314), .Z(n4310) );
  ANDN U8411 ( .B(n4315), .A(n4316), .Z(n4313) );
  XNOR U8412 ( .A(b[3206]), .B(n4314), .Z(n4315) );
  XNOR U8413 ( .A(b[3206]), .B(n4316), .Z(c[3206]) );
  XOR U8414 ( .A(n4317), .B(n4318), .Z(n4314) );
  ANDN U8415 ( .B(n4319), .A(n4320), .Z(n4317) );
  XNOR U8416 ( .A(b[3205]), .B(n4318), .Z(n4319) );
  XNOR U8417 ( .A(b[3205]), .B(n4320), .Z(c[3205]) );
  XOR U8418 ( .A(n4321), .B(n4322), .Z(n4318) );
  ANDN U8419 ( .B(n4323), .A(n4324), .Z(n4321) );
  XNOR U8420 ( .A(b[3204]), .B(n4322), .Z(n4323) );
  XNOR U8421 ( .A(b[3204]), .B(n4324), .Z(c[3204]) );
  XOR U8422 ( .A(n4325), .B(n4326), .Z(n4322) );
  ANDN U8423 ( .B(n4327), .A(n4328), .Z(n4325) );
  XNOR U8424 ( .A(b[3203]), .B(n4326), .Z(n4327) );
  XNOR U8425 ( .A(b[3203]), .B(n4328), .Z(c[3203]) );
  XOR U8426 ( .A(n4329), .B(n4330), .Z(n4326) );
  ANDN U8427 ( .B(n4331), .A(n4332), .Z(n4329) );
  XNOR U8428 ( .A(b[3202]), .B(n4330), .Z(n4331) );
  XNOR U8429 ( .A(b[3202]), .B(n4332), .Z(c[3202]) );
  XOR U8430 ( .A(n4333), .B(n4334), .Z(n4330) );
  ANDN U8431 ( .B(n4335), .A(n4336), .Z(n4333) );
  XNOR U8432 ( .A(b[3201]), .B(n4334), .Z(n4335) );
  XNOR U8433 ( .A(b[3201]), .B(n4336), .Z(c[3201]) );
  XOR U8434 ( .A(n4337), .B(n4338), .Z(n4334) );
  ANDN U8435 ( .B(n4339), .A(n4340), .Z(n4337) );
  XNOR U8436 ( .A(b[3200]), .B(n4338), .Z(n4339) );
  XNOR U8437 ( .A(b[3200]), .B(n4340), .Z(c[3200]) );
  XOR U8438 ( .A(n4341), .B(n4342), .Z(n4338) );
  ANDN U8439 ( .B(n4343), .A(n4344), .Z(n4341) );
  XNOR U8440 ( .A(b[3199]), .B(n4342), .Z(n4343) );
  XNOR U8441 ( .A(b[31]), .B(n4345), .Z(c[31]) );
  XNOR U8442 ( .A(b[319]), .B(n4346), .Z(c[319]) );
  XNOR U8443 ( .A(b[3199]), .B(n4344), .Z(c[3199]) );
  XOR U8444 ( .A(n4347), .B(n4348), .Z(n4342) );
  ANDN U8445 ( .B(n4349), .A(n4350), .Z(n4347) );
  XNOR U8446 ( .A(b[3198]), .B(n4348), .Z(n4349) );
  XNOR U8447 ( .A(b[3198]), .B(n4350), .Z(c[3198]) );
  XOR U8448 ( .A(n4351), .B(n4352), .Z(n4348) );
  ANDN U8449 ( .B(n4353), .A(n4354), .Z(n4351) );
  XNOR U8450 ( .A(b[3197]), .B(n4352), .Z(n4353) );
  XNOR U8451 ( .A(b[3197]), .B(n4354), .Z(c[3197]) );
  XOR U8452 ( .A(n4355), .B(n4356), .Z(n4352) );
  ANDN U8453 ( .B(n4357), .A(n4358), .Z(n4355) );
  XNOR U8454 ( .A(b[3196]), .B(n4356), .Z(n4357) );
  XNOR U8455 ( .A(b[3196]), .B(n4358), .Z(c[3196]) );
  XOR U8456 ( .A(n4359), .B(n4360), .Z(n4356) );
  ANDN U8457 ( .B(n4361), .A(n4362), .Z(n4359) );
  XNOR U8458 ( .A(b[3195]), .B(n4360), .Z(n4361) );
  XNOR U8459 ( .A(b[3195]), .B(n4362), .Z(c[3195]) );
  XOR U8460 ( .A(n4363), .B(n4364), .Z(n4360) );
  ANDN U8461 ( .B(n4365), .A(n4366), .Z(n4363) );
  XNOR U8462 ( .A(b[3194]), .B(n4364), .Z(n4365) );
  XNOR U8463 ( .A(b[3194]), .B(n4366), .Z(c[3194]) );
  XOR U8464 ( .A(n4367), .B(n4368), .Z(n4364) );
  ANDN U8465 ( .B(n4369), .A(n4370), .Z(n4367) );
  XNOR U8466 ( .A(b[3193]), .B(n4368), .Z(n4369) );
  XNOR U8467 ( .A(b[3193]), .B(n4370), .Z(c[3193]) );
  XOR U8468 ( .A(n4371), .B(n4372), .Z(n4368) );
  ANDN U8469 ( .B(n4373), .A(n4374), .Z(n4371) );
  XNOR U8470 ( .A(b[3192]), .B(n4372), .Z(n4373) );
  XNOR U8471 ( .A(b[3192]), .B(n4374), .Z(c[3192]) );
  XOR U8472 ( .A(n4375), .B(n4376), .Z(n4372) );
  ANDN U8473 ( .B(n4377), .A(n4378), .Z(n4375) );
  XNOR U8474 ( .A(b[3191]), .B(n4376), .Z(n4377) );
  XNOR U8475 ( .A(b[3191]), .B(n4378), .Z(c[3191]) );
  XOR U8476 ( .A(n4379), .B(n4380), .Z(n4376) );
  ANDN U8477 ( .B(n4381), .A(n4382), .Z(n4379) );
  XNOR U8478 ( .A(b[3190]), .B(n4380), .Z(n4381) );
  XNOR U8479 ( .A(b[3190]), .B(n4382), .Z(c[3190]) );
  XOR U8480 ( .A(n4383), .B(n4384), .Z(n4380) );
  ANDN U8481 ( .B(n4385), .A(n4386), .Z(n4383) );
  XNOR U8482 ( .A(b[3189]), .B(n4384), .Z(n4385) );
  XNOR U8483 ( .A(b[318]), .B(n4387), .Z(c[318]) );
  XNOR U8484 ( .A(b[3189]), .B(n4386), .Z(c[3189]) );
  XOR U8485 ( .A(n4388), .B(n4389), .Z(n4384) );
  ANDN U8486 ( .B(n4390), .A(n4391), .Z(n4388) );
  XNOR U8487 ( .A(b[3188]), .B(n4389), .Z(n4390) );
  XNOR U8488 ( .A(b[3188]), .B(n4391), .Z(c[3188]) );
  XOR U8489 ( .A(n4392), .B(n4393), .Z(n4389) );
  ANDN U8490 ( .B(n4394), .A(n4395), .Z(n4392) );
  XNOR U8491 ( .A(b[3187]), .B(n4393), .Z(n4394) );
  XNOR U8492 ( .A(b[3187]), .B(n4395), .Z(c[3187]) );
  XOR U8493 ( .A(n4396), .B(n4397), .Z(n4393) );
  ANDN U8494 ( .B(n4398), .A(n4399), .Z(n4396) );
  XNOR U8495 ( .A(b[3186]), .B(n4397), .Z(n4398) );
  XNOR U8496 ( .A(b[3186]), .B(n4399), .Z(c[3186]) );
  XOR U8497 ( .A(n4400), .B(n4401), .Z(n4397) );
  ANDN U8498 ( .B(n4402), .A(n4403), .Z(n4400) );
  XNOR U8499 ( .A(b[3185]), .B(n4401), .Z(n4402) );
  XNOR U8500 ( .A(b[3185]), .B(n4403), .Z(c[3185]) );
  XOR U8501 ( .A(n4404), .B(n4405), .Z(n4401) );
  ANDN U8502 ( .B(n4406), .A(n4407), .Z(n4404) );
  XNOR U8503 ( .A(b[3184]), .B(n4405), .Z(n4406) );
  XNOR U8504 ( .A(b[3184]), .B(n4407), .Z(c[3184]) );
  XOR U8505 ( .A(n4408), .B(n4409), .Z(n4405) );
  ANDN U8506 ( .B(n4410), .A(n4411), .Z(n4408) );
  XNOR U8507 ( .A(b[3183]), .B(n4409), .Z(n4410) );
  XNOR U8508 ( .A(b[3183]), .B(n4411), .Z(c[3183]) );
  XOR U8509 ( .A(n4412), .B(n4413), .Z(n4409) );
  ANDN U8510 ( .B(n4414), .A(n4415), .Z(n4412) );
  XNOR U8511 ( .A(b[3182]), .B(n4413), .Z(n4414) );
  XNOR U8512 ( .A(b[3182]), .B(n4415), .Z(c[3182]) );
  XOR U8513 ( .A(n4416), .B(n4417), .Z(n4413) );
  ANDN U8514 ( .B(n4418), .A(n4419), .Z(n4416) );
  XNOR U8515 ( .A(b[3181]), .B(n4417), .Z(n4418) );
  XNOR U8516 ( .A(b[3181]), .B(n4419), .Z(c[3181]) );
  XOR U8517 ( .A(n4420), .B(n4421), .Z(n4417) );
  ANDN U8518 ( .B(n4422), .A(n4423), .Z(n4420) );
  XNOR U8519 ( .A(b[3180]), .B(n4421), .Z(n4422) );
  XNOR U8520 ( .A(b[3180]), .B(n4423), .Z(c[3180]) );
  XOR U8521 ( .A(n4424), .B(n4425), .Z(n4421) );
  ANDN U8522 ( .B(n4426), .A(n4427), .Z(n4424) );
  XNOR U8523 ( .A(b[3179]), .B(n4425), .Z(n4426) );
  XNOR U8524 ( .A(b[317]), .B(n4428), .Z(c[317]) );
  XNOR U8525 ( .A(b[3179]), .B(n4427), .Z(c[3179]) );
  XOR U8526 ( .A(n4429), .B(n4430), .Z(n4425) );
  ANDN U8527 ( .B(n4431), .A(n4432), .Z(n4429) );
  XNOR U8528 ( .A(b[3178]), .B(n4430), .Z(n4431) );
  XNOR U8529 ( .A(b[3178]), .B(n4432), .Z(c[3178]) );
  XOR U8530 ( .A(n4433), .B(n4434), .Z(n4430) );
  ANDN U8531 ( .B(n4435), .A(n4436), .Z(n4433) );
  XNOR U8532 ( .A(b[3177]), .B(n4434), .Z(n4435) );
  XNOR U8533 ( .A(b[3177]), .B(n4436), .Z(c[3177]) );
  XOR U8534 ( .A(n4437), .B(n4438), .Z(n4434) );
  ANDN U8535 ( .B(n4439), .A(n4440), .Z(n4437) );
  XNOR U8536 ( .A(b[3176]), .B(n4438), .Z(n4439) );
  XNOR U8537 ( .A(b[3176]), .B(n4440), .Z(c[3176]) );
  XOR U8538 ( .A(n4441), .B(n4442), .Z(n4438) );
  ANDN U8539 ( .B(n4443), .A(n4444), .Z(n4441) );
  XNOR U8540 ( .A(b[3175]), .B(n4442), .Z(n4443) );
  XNOR U8541 ( .A(b[3175]), .B(n4444), .Z(c[3175]) );
  XOR U8542 ( .A(n4445), .B(n4446), .Z(n4442) );
  ANDN U8543 ( .B(n4447), .A(n4448), .Z(n4445) );
  XNOR U8544 ( .A(b[3174]), .B(n4446), .Z(n4447) );
  XNOR U8545 ( .A(b[3174]), .B(n4448), .Z(c[3174]) );
  XOR U8546 ( .A(n4449), .B(n4450), .Z(n4446) );
  ANDN U8547 ( .B(n4451), .A(n4452), .Z(n4449) );
  XNOR U8548 ( .A(b[3173]), .B(n4450), .Z(n4451) );
  XNOR U8549 ( .A(b[3173]), .B(n4452), .Z(c[3173]) );
  XOR U8550 ( .A(n4453), .B(n4454), .Z(n4450) );
  ANDN U8551 ( .B(n4455), .A(n4456), .Z(n4453) );
  XNOR U8552 ( .A(b[3172]), .B(n4454), .Z(n4455) );
  XNOR U8553 ( .A(b[3172]), .B(n4456), .Z(c[3172]) );
  XOR U8554 ( .A(n4457), .B(n4458), .Z(n4454) );
  ANDN U8555 ( .B(n4459), .A(n4460), .Z(n4457) );
  XNOR U8556 ( .A(b[3171]), .B(n4458), .Z(n4459) );
  XNOR U8557 ( .A(b[3171]), .B(n4460), .Z(c[3171]) );
  XOR U8558 ( .A(n4461), .B(n4462), .Z(n4458) );
  ANDN U8559 ( .B(n4463), .A(n4464), .Z(n4461) );
  XNOR U8560 ( .A(b[3170]), .B(n4462), .Z(n4463) );
  XNOR U8561 ( .A(b[3170]), .B(n4464), .Z(c[3170]) );
  XOR U8562 ( .A(n4465), .B(n4466), .Z(n4462) );
  ANDN U8563 ( .B(n4467), .A(n4468), .Z(n4465) );
  XNOR U8564 ( .A(b[3169]), .B(n4466), .Z(n4467) );
  XNOR U8565 ( .A(b[316]), .B(n4469), .Z(c[316]) );
  XNOR U8566 ( .A(b[3169]), .B(n4468), .Z(c[3169]) );
  XOR U8567 ( .A(n4470), .B(n4471), .Z(n4466) );
  ANDN U8568 ( .B(n4472), .A(n4473), .Z(n4470) );
  XNOR U8569 ( .A(b[3168]), .B(n4471), .Z(n4472) );
  XNOR U8570 ( .A(b[3168]), .B(n4473), .Z(c[3168]) );
  XOR U8571 ( .A(n4474), .B(n4475), .Z(n4471) );
  ANDN U8572 ( .B(n4476), .A(n4477), .Z(n4474) );
  XNOR U8573 ( .A(b[3167]), .B(n4475), .Z(n4476) );
  XNOR U8574 ( .A(b[3167]), .B(n4477), .Z(c[3167]) );
  XOR U8575 ( .A(n4478), .B(n4479), .Z(n4475) );
  ANDN U8576 ( .B(n4480), .A(n4481), .Z(n4478) );
  XNOR U8577 ( .A(b[3166]), .B(n4479), .Z(n4480) );
  XNOR U8578 ( .A(b[3166]), .B(n4481), .Z(c[3166]) );
  XOR U8579 ( .A(n4482), .B(n4483), .Z(n4479) );
  ANDN U8580 ( .B(n4484), .A(n4485), .Z(n4482) );
  XNOR U8581 ( .A(b[3165]), .B(n4483), .Z(n4484) );
  XNOR U8582 ( .A(b[3165]), .B(n4485), .Z(c[3165]) );
  XOR U8583 ( .A(n4486), .B(n4487), .Z(n4483) );
  ANDN U8584 ( .B(n4488), .A(n4489), .Z(n4486) );
  XNOR U8585 ( .A(b[3164]), .B(n4487), .Z(n4488) );
  XNOR U8586 ( .A(b[3164]), .B(n4489), .Z(c[3164]) );
  XOR U8587 ( .A(n4490), .B(n4491), .Z(n4487) );
  ANDN U8588 ( .B(n4492), .A(n4493), .Z(n4490) );
  XNOR U8589 ( .A(b[3163]), .B(n4491), .Z(n4492) );
  XNOR U8590 ( .A(b[3163]), .B(n4493), .Z(c[3163]) );
  XOR U8591 ( .A(n4494), .B(n4495), .Z(n4491) );
  ANDN U8592 ( .B(n4496), .A(n4497), .Z(n4494) );
  XNOR U8593 ( .A(b[3162]), .B(n4495), .Z(n4496) );
  XNOR U8594 ( .A(b[3162]), .B(n4497), .Z(c[3162]) );
  XOR U8595 ( .A(n4498), .B(n4499), .Z(n4495) );
  ANDN U8596 ( .B(n4500), .A(n4501), .Z(n4498) );
  XNOR U8597 ( .A(b[3161]), .B(n4499), .Z(n4500) );
  XNOR U8598 ( .A(b[3161]), .B(n4501), .Z(c[3161]) );
  XOR U8599 ( .A(n4502), .B(n4503), .Z(n4499) );
  ANDN U8600 ( .B(n4504), .A(n4505), .Z(n4502) );
  XNOR U8601 ( .A(b[3160]), .B(n4503), .Z(n4504) );
  XNOR U8602 ( .A(b[3160]), .B(n4505), .Z(c[3160]) );
  XOR U8603 ( .A(n4506), .B(n4507), .Z(n4503) );
  ANDN U8604 ( .B(n4508), .A(n4509), .Z(n4506) );
  XNOR U8605 ( .A(b[3159]), .B(n4507), .Z(n4508) );
  XNOR U8606 ( .A(b[315]), .B(n4510), .Z(c[315]) );
  XNOR U8607 ( .A(b[3159]), .B(n4509), .Z(c[3159]) );
  XOR U8608 ( .A(n4511), .B(n4512), .Z(n4507) );
  ANDN U8609 ( .B(n4513), .A(n4514), .Z(n4511) );
  XNOR U8610 ( .A(b[3158]), .B(n4512), .Z(n4513) );
  XNOR U8611 ( .A(b[3158]), .B(n4514), .Z(c[3158]) );
  XOR U8612 ( .A(n4515), .B(n4516), .Z(n4512) );
  ANDN U8613 ( .B(n4517), .A(n4518), .Z(n4515) );
  XNOR U8614 ( .A(b[3157]), .B(n4516), .Z(n4517) );
  XNOR U8615 ( .A(b[3157]), .B(n4518), .Z(c[3157]) );
  XOR U8616 ( .A(n4519), .B(n4520), .Z(n4516) );
  ANDN U8617 ( .B(n4521), .A(n4522), .Z(n4519) );
  XNOR U8618 ( .A(b[3156]), .B(n4520), .Z(n4521) );
  XNOR U8619 ( .A(b[3156]), .B(n4522), .Z(c[3156]) );
  XOR U8620 ( .A(n4523), .B(n4524), .Z(n4520) );
  ANDN U8621 ( .B(n4525), .A(n4526), .Z(n4523) );
  XNOR U8622 ( .A(b[3155]), .B(n4524), .Z(n4525) );
  XNOR U8623 ( .A(b[3155]), .B(n4526), .Z(c[3155]) );
  XOR U8624 ( .A(n4527), .B(n4528), .Z(n4524) );
  ANDN U8625 ( .B(n4529), .A(n4530), .Z(n4527) );
  XNOR U8626 ( .A(b[3154]), .B(n4528), .Z(n4529) );
  XNOR U8627 ( .A(b[3154]), .B(n4530), .Z(c[3154]) );
  XOR U8628 ( .A(n4531), .B(n4532), .Z(n4528) );
  ANDN U8629 ( .B(n4533), .A(n4534), .Z(n4531) );
  XNOR U8630 ( .A(b[3153]), .B(n4532), .Z(n4533) );
  XNOR U8631 ( .A(b[3153]), .B(n4534), .Z(c[3153]) );
  XOR U8632 ( .A(n4535), .B(n4536), .Z(n4532) );
  ANDN U8633 ( .B(n4537), .A(n4538), .Z(n4535) );
  XNOR U8634 ( .A(b[3152]), .B(n4536), .Z(n4537) );
  XNOR U8635 ( .A(b[3152]), .B(n4538), .Z(c[3152]) );
  XOR U8636 ( .A(n4539), .B(n4540), .Z(n4536) );
  ANDN U8637 ( .B(n4541), .A(n4542), .Z(n4539) );
  XNOR U8638 ( .A(b[3151]), .B(n4540), .Z(n4541) );
  XNOR U8639 ( .A(b[3151]), .B(n4542), .Z(c[3151]) );
  XOR U8640 ( .A(n4543), .B(n4544), .Z(n4540) );
  ANDN U8641 ( .B(n4545), .A(n4546), .Z(n4543) );
  XNOR U8642 ( .A(b[3150]), .B(n4544), .Z(n4545) );
  XNOR U8643 ( .A(b[3150]), .B(n4546), .Z(c[3150]) );
  XOR U8644 ( .A(n4547), .B(n4548), .Z(n4544) );
  ANDN U8645 ( .B(n4549), .A(n4550), .Z(n4547) );
  XNOR U8646 ( .A(b[3149]), .B(n4548), .Z(n4549) );
  XNOR U8647 ( .A(b[314]), .B(n4551), .Z(c[314]) );
  XNOR U8648 ( .A(b[3149]), .B(n4550), .Z(c[3149]) );
  XOR U8649 ( .A(n4552), .B(n4553), .Z(n4548) );
  ANDN U8650 ( .B(n4554), .A(n4555), .Z(n4552) );
  XNOR U8651 ( .A(b[3148]), .B(n4553), .Z(n4554) );
  XNOR U8652 ( .A(b[3148]), .B(n4555), .Z(c[3148]) );
  XOR U8653 ( .A(n4556), .B(n4557), .Z(n4553) );
  ANDN U8654 ( .B(n4558), .A(n4559), .Z(n4556) );
  XNOR U8655 ( .A(b[3147]), .B(n4557), .Z(n4558) );
  XNOR U8656 ( .A(b[3147]), .B(n4559), .Z(c[3147]) );
  XOR U8657 ( .A(n4560), .B(n4561), .Z(n4557) );
  ANDN U8658 ( .B(n4562), .A(n4563), .Z(n4560) );
  XNOR U8659 ( .A(b[3146]), .B(n4561), .Z(n4562) );
  XNOR U8660 ( .A(b[3146]), .B(n4563), .Z(c[3146]) );
  XOR U8661 ( .A(n4564), .B(n4565), .Z(n4561) );
  ANDN U8662 ( .B(n4566), .A(n4567), .Z(n4564) );
  XNOR U8663 ( .A(b[3145]), .B(n4565), .Z(n4566) );
  XNOR U8664 ( .A(b[3145]), .B(n4567), .Z(c[3145]) );
  XOR U8665 ( .A(n4568), .B(n4569), .Z(n4565) );
  ANDN U8666 ( .B(n4570), .A(n4571), .Z(n4568) );
  XNOR U8667 ( .A(b[3144]), .B(n4569), .Z(n4570) );
  XNOR U8668 ( .A(b[3144]), .B(n4571), .Z(c[3144]) );
  XOR U8669 ( .A(n4572), .B(n4573), .Z(n4569) );
  ANDN U8670 ( .B(n4574), .A(n4575), .Z(n4572) );
  XNOR U8671 ( .A(b[3143]), .B(n4573), .Z(n4574) );
  XNOR U8672 ( .A(b[3143]), .B(n4575), .Z(c[3143]) );
  XOR U8673 ( .A(n4576), .B(n4577), .Z(n4573) );
  ANDN U8674 ( .B(n4578), .A(n4579), .Z(n4576) );
  XNOR U8675 ( .A(b[3142]), .B(n4577), .Z(n4578) );
  XNOR U8676 ( .A(b[3142]), .B(n4579), .Z(c[3142]) );
  XOR U8677 ( .A(n4580), .B(n4581), .Z(n4577) );
  ANDN U8678 ( .B(n4582), .A(n4583), .Z(n4580) );
  XNOR U8679 ( .A(b[3141]), .B(n4581), .Z(n4582) );
  XNOR U8680 ( .A(b[3141]), .B(n4583), .Z(c[3141]) );
  XOR U8681 ( .A(n4584), .B(n4585), .Z(n4581) );
  ANDN U8682 ( .B(n4586), .A(n4587), .Z(n4584) );
  XNOR U8683 ( .A(b[3140]), .B(n4585), .Z(n4586) );
  XNOR U8684 ( .A(b[3140]), .B(n4587), .Z(c[3140]) );
  XOR U8685 ( .A(n4588), .B(n4589), .Z(n4585) );
  ANDN U8686 ( .B(n4590), .A(n4591), .Z(n4588) );
  XNOR U8687 ( .A(b[3139]), .B(n4589), .Z(n4590) );
  XNOR U8688 ( .A(b[313]), .B(n4592), .Z(c[313]) );
  XNOR U8689 ( .A(b[3139]), .B(n4591), .Z(c[3139]) );
  XOR U8690 ( .A(n4593), .B(n4594), .Z(n4589) );
  ANDN U8691 ( .B(n4595), .A(n4596), .Z(n4593) );
  XNOR U8692 ( .A(b[3138]), .B(n4594), .Z(n4595) );
  XNOR U8693 ( .A(b[3138]), .B(n4596), .Z(c[3138]) );
  XOR U8694 ( .A(n4597), .B(n4598), .Z(n4594) );
  ANDN U8695 ( .B(n4599), .A(n4600), .Z(n4597) );
  XNOR U8696 ( .A(b[3137]), .B(n4598), .Z(n4599) );
  XNOR U8697 ( .A(b[3137]), .B(n4600), .Z(c[3137]) );
  XOR U8698 ( .A(n4601), .B(n4602), .Z(n4598) );
  ANDN U8699 ( .B(n4603), .A(n4604), .Z(n4601) );
  XNOR U8700 ( .A(b[3136]), .B(n4602), .Z(n4603) );
  XNOR U8701 ( .A(b[3136]), .B(n4604), .Z(c[3136]) );
  XOR U8702 ( .A(n4605), .B(n4606), .Z(n4602) );
  ANDN U8703 ( .B(n4607), .A(n4608), .Z(n4605) );
  XNOR U8704 ( .A(b[3135]), .B(n4606), .Z(n4607) );
  XNOR U8705 ( .A(b[3135]), .B(n4608), .Z(c[3135]) );
  XOR U8706 ( .A(n4609), .B(n4610), .Z(n4606) );
  ANDN U8707 ( .B(n4611), .A(n4612), .Z(n4609) );
  XNOR U8708 ( .A(b[3134]), .B(n4610), .Z(n4611) );
  XNOR U8709 ( .A(b[3134]), .B(n4612), .Z(c[3134]) );
  XOR U8710 ( .A(n4613), .B(n4614), .Z(n4610) );
  ANDN U8711 ( .B(n4615), .A(n4616), .Z(n4613) );
  XNOR U8712 ( .A(b[3133]), .B(n4614), .Z(n4615) );
  XNOR U8713 ( .A(b[3133]), .B(n4616), .Z(c[3133]) );
  XOR U8714 ( .A(n4617), .B(n4618), .Z(n4614) );
  ANDN U8715 ( .B(n4619), .A(n4620), .Z(n4617) );
  XNOR U8716 ( .A(b[3132]), .B(n4618), .Z(n4619) );
  XNOR U8717 ( .A(b[3132]), .B(n4620), .Z(c[3132]) );
  XOR U8718 ( .A(n4621), .B(n4622), .Z(n4618) );
  ANDN U8719 ( .B(n4623), .A(n4624), .Z(n4621) );
  XNOR U8720 ( .A(b[3131]), .B(n4622), .Z(n4623) );
  XNOR U8721 ( .A(b[3131]), .B(n4624), .Z(c[3131]) );
  XOR U8722 ( .A(n4625), .B(n4626), .Z(n4622) );
  ANDN U8723 ( .B(n4627), .A(n4628), .Z(n4625) );
  XNOR U8724 ( .A(b[3130]), .B(n4626), .Z(n4627) );
  XNOR U8725 ( .A(b[3130]), .B(n4628), .Z(c[3130]) );
  XOR U8726 ( .A(n4629), .B(n4630), .Z(n4626) );
  ANDN U8727 ( .B(n4631), .A(n4632), .Z(n4629) );
  XNOR U8728 ( .A(b[3129]), .B(n4630), .Z(n4631) );
  XNOR U8729 ( .A(b[312]), .B(n4633), .Z(c[312]) );
  XNOR U8730 ( .A(b[3129]), .B(n4632), .Z(c[3129]) );
  XOR U8731 ( .A(n4634), .B(n4635), .Z(n4630) );
  ANDN U8732 ( .B(n4636), .A(n4637), .Z(n4634) );
  XNOR U8733 ( .A(b[3128]), .B(n4635), .Z(n4636) );
  XNOR U8734 ( .A(b[3128]), .B(n4637), .Z(c[3128]) );
  XOR U8735 ( .A(n4638), .B(n4639), .Z(n4635) );
  ANDN U8736 ( .B(n4640), .A(n4641), .Z(n4638) );
  XNOR U8737 ( .A(b[3127]), .B(n4639), .Z(n4640) );
  XNOR U8738 ( .A(b[3127]), .B(n4641), .Z(c[3127]) );
  XOR U8739 ( .A(n4642), .B(n4643), .Z(n4639) );
  ANDN U8740 ( .B(n4644), .A(n4645), .Z(n4642) );
  XNOR U8741 ( .A(b[3126]), .B(n4643), .Z(n4644) );
  XNOR U8742 ( .A(b[3126]), .B(n4645), .Z(c[3126]) );
  XOR U8743 ( .A(n4646), .B(n4647), .Z(n4643) );
  ANDN U8744 ( .B(n4648), .A(n4649), .Z(n4646) );
  XNOR U8745 ( .A(b[3125]), .B(n4647), .Z(n4648) );
  XNOR U8746 ( .A(b[3125]), .B(n4649), .Z(c[3125]) );
  XOR U8747 ( .A(n4650), .B(n4651), .Z(n4647) );
  ANDN U8748 ( .B(n4652), .A(n4653), .Z(n4650) );
  XNOR U8749 ( .A(b[3124]), .B(n4651), .Z(n4652) );
  XNOR U8750 ( .A(b[3124]), .B(n4653), .Z(c[3124]) );
  XOR U8751 ( .A(n4654), .B(n4655), .Z(n4651) );
  ANDN U8752 ( .B(n4656), .A(n4657), .Z(n4654) );
  XNOR U8753 ( .A(b[3123]), .B(n4655), .Z(n4656) );
  XNOR U8754 ( .A(b[3123]), .B(n4657), .Z(c[3123]) );
  XOR U8755 ( .A(n4658), .B(n4659), .Z(n4655) );
  ANDN U8756 ( .B(n4660), .A(n4661), .Z(n4658) );
  XNOR U8757 ( .A(b[3122]), .B(n4659), .Z(n4660) );
  XNOR U8758 ( .A(b[3122]), .B(n4661), .Z(c[3122]) );
  XOR U8759 ( .A(n4662), .B(n4663), .Z(n4659) );
  ANDN U8760 ( .B(n4664), .A(n4665), .Z(n4662) );
  XNOR U8761 ( .A(b[3121]), .B(n4663), .Z(n4664) );
  XNOR U8762 ( .A(b[3121]), .B(n4665), .Z(c[3121]) );
  XOR U8763 ( .A(n4666), .B(n4667), .Z(n4663) );
  ANDN U8764 ( .B(n4668), .A(n4669), .Z(n4666) );
  XNOR U8765 ( .A(b[3120]), .B(n4667), .Z(n4668) );
  XNOR U8766 ( .A(b[3120]), .B(n4669), .Z(c[3120]) );
  XOR U8767 ( .A(n4670), .B(n4671), .Z(n4667) );
  ANDN U8768 ( .B(n4672), .A(n4673), .Z(n4670) );
  XNOR U8769 ( .A(b[3119]), .B(n4671), .Z(n4672) );
  XNOR U8770 ( .A(b[311]), .B(n4674), .Z(c[311]) );
  XNOR U8771 ( .A(b[3119]), .B(n4673), .Z(c[3119]) );
  XOR U8772 ( .A(n4675), .B(n4676), .Z(n4671) );
  ANDN U8773 ( .B(n4677), .A(n4678), .Z(n4675) );
  XNOR U8774 ( .A(b[3118]), .B(n4676), .Z(n4677) );
  XNOR U8775 ( .A(b[3118]), .B(n4678), .Z(c[3118]) );
  XOR U8776 ( .A(n4679), .B(n4680), .Z(n4676) );
  ANDN U8777 ( .B(n4681), .A(n4682), .Z(n4679) );
  XNOR U8778 ( .A(b[3117]), .B(n4680), .Z(n4681) );
  XNOR U8779 ( .A(b[3117]), .B(n4682), .Z(c[3117]) );
  XOR U8780 ( .A(n4683), .B(n4684), .Z(n4680) );
  ANDN U8781 ( .B(n4685), .A(n4686), .Z(n4683) );
  XNOR U8782 ( .A(b[3116]), .B(n4684), .Z(n4685) );
  XNOR U8783 ( .A(b[3116]), .B(n4686), .Z(c[3116]) );
  XOR U8784 ( .A(n4687), .B(n4688), .Z(n4684) );
  ANDN U8785 ( .B(n4689), .A(n4690), .Z(n4687) );
  XNOR U8786 ( .A(b[3115]), .B(n4688), .Z(n4689) );
  XNOR U8787 ( .A(b[3115]), .B(n4690), .Z(c[3115]) );
  XOR U8788 ( .A(n4691), .B(n4692), .Z(n4688) );
  ANDN U8789 ( .B(n4693), .A(n4694), .Z(n4691) );
  XNOR U8790 ( .A(b[3114]), .B(n4692), .Z(n4693) );
  XNOR U8791 ( .A(b[3114]), .B(n4694), .Z(c[3114]) );
  XOR U8792 ( .A(n4695), .B(n4696), .Z(n4692) );
  ANDN U8793 ( .B(n4697), .A(n4698), .Z(n4695) );
  XNOR U8794 ( .A(b[3113]), .B(n4696), .Z(n4697) );
  XNOR U8795 ( .A(b[3113]), .B(n4698), .Z(c[3113]) );
  XOR U8796 ( .A(n4699), .B(n4700), .Z(n4696) );
  ANDN U8797 ( .B(n4701), .A(n4702), .Z(n4699) );
  XNOR U8798 ( .A(b[3112]), .B(n4700), .Z(n4701) );
  XNOR U8799 ( .A(b[3112]), .B(n4702), .Z(c[3112]) );
  XOR U8800 ( .A(n4703), .B(n4704), .Z(n4700) );
  ANDN U8801 ( .B(n4705), .A(n4706), .Z(n4703) );
  XNOR U8802 ( .A(b[3111]), .B(n4704), .Z(n4705) );
  XNOR U8803 ( .A(b[3111]), .B(n4706), .Z(c[3111]) );
  XOR U8804 ( .A(n4707), .B(n4708), .Z(n4704) );
  ANDN U8805 ( .B(n4709), .A(n4710), .Z(n4707) );
  XNOR U8806 ( .A(b[3110]), .B(n4708), .Z(n4709) );
  XNOR U8807 ( .A(b[3110]), .B(n4710), .Z(c[3110]) );
  XOR U8808 ( .A(n4711), .B(n4712), .Z(n4708) );
  ANDN U8809 ( .B(n4713), .A(n4714), .Z(n4711) );
  XNOR U8810 ( .A(b[3109]), .B(n4712), .Z(n4713) );
  XNOR U8811 ( .A(b[310]), .B(n4715), .Z(c[310]) );
  XNOR U8812 ( .A(b[3109]), .B(n4714), .Z(c[3109]) );
  XOR U8813 ( .A(n4716), .B(n4717), .Z(n4712) );
  ANDN U8814 ( .B(n4718), .A(n4719), .Z(n4716) );
  XNOR U8815 ( .A(b[3108]), .B(n4717), .Z(n4718) );
  XNOR U8816 ( .A(b[3108]), .B(n4719), .Z(c[3108]) );
  XOR U8817 ( .A(n4720), .B(n4721), .Z(n4717) );
  ANDN U8818 ( .B(n4722), .A(n4723), .Z(n4720) );
  XNOR U8819 ( .A(b[3107]), .B(n4721), .Z(n4722) );
  XNOR U8820 ( .A(b[3107]), .B(n4723), .Z(c[3107]) );
  XOR U8821 ( .A(n4724), .B(n4725), .Z(n4721) );
  ANDN U8822 ( .B(n4726), .A(n4727), .Z(n4724) );
  XNOR U8823 ( .A(b[3106]), .B(n4725), .Z(n4726) );
  XNOR U8824 ( .A(b[3106]), .B(n4727), .Z(c[3106]) );
  XOR U8825 ( .A(n4728), .B(n4729), .Z(n4725) );
  ANDN U8826 ( .B(n4730), .A(n4731), .Z(n4728) );
  XNOR U8827 ( .A(b[3105]), .B(n4729), .Z(n4730) );
  XNOR U8828 ( .A(b[3105]), .B(n4731), .Z(c[3105]) );
  XOR U8829 ( .A(n4732), .B(n4733), .Z(n4729) );
  ANDN U8830 ( .B(n4734), .A(n4735), .Z(n4732) );
  XNOR U8831 ( .A(b[3104]), .B(n4733), .Z(n4734) );
  XNOR U8832 ( .A(b[3104]), .B(n4735), .Z(c[3104]) );
  XOR U8833 ( .A(n4736), .B(n4737), .Z(n4733) );
  ANDN U8834 ( .B(n4738), .A(n4739), .Z(n4736) );
  XNOR U8835 ( .A(b[3103]), .B(n4737), .Z(n4738) );
  XNOR U8836 ( .A(b[3103]), .B(n4739), .Z(c[3103]) );
  XOR U8837 ( .A(n4740), .B(n4741), .Z(n4737) );
  ANDN U8838 ( .B(n4742), .A(n4743), .Z(n4740) );
  XNOR U8839 ( .A(b[3102]), .B(n4741), .Z(n4742) );
  XNOR U8840 ( .A(b[3102]), .B(n4743), .Z(c[3102]) );
  XOR U8841 ( .A(n4744), .B(n4745), .Z(n4741) );
  ANDN U8842 ( .B(n4746), .A(n4747), .Z(n4744) );
  XNOR U8843 ( .A(b[3101]), .B(n4745), .Z(n4746) );
  XNOR U8844 ( .A(b[3101]), .B(n4747), .Z(c[3101]) );
  XOR U8845 ( .A(n4748), .B(n4749), .Z(n4745) );
  ANDN U8846 ( .B(n4750), .A(n4751), .Z(n4748) );
  XNOR U8847 ( .A(b[3100]), .B(n4749), .Z(n4750) );
  XNOR U8848 ( .A(b[3100]), .B(n4751), .Z(c[3100]) );
  XOR U8849 ( .A(n4752), .B(n4753), .Z(n4749) );
  ANDN U8850 ( .B(n4754), .A(n4755), .Z(n4752) );
  XNOR U8851 ( .A(b[3099]), .B(n4753), .Z(n4754) );
  XNOR U8852 ( .A(b[30]), .B(n4756), .Z(c[30]) );
  XNOR U8853 ( .A(b[309]), .B(n4757), .Z(c[309]) );
  XNOR U8854 ( .A(b[3099]), .B(n4755), .Z(c[3099]) );
  XOR U8855 ( .A(n4758), .B(n4759), .Z(n4753) );
  ANDN U8856 ( .B(n4760), .A(n4761), .Z(n4758) );
  XNOR U8857 ( .A(b[3098]), .B(n4759), .Z(n4760) );
  XNOR U8858 ( .A(b[3098]), .B(n4761), .Z(c[3098]) );
  XOR U8859 ( .A(n4762), .B(n4763), .Z(n4759) );
  ANDN U8860 ( .B(n4764), .A(n4765), .Z(n4762) );
  XNOR U8861 ( .A(b[3097]), .B(n4763), .Z(n4764) );
  XNOR U8862 ( .A(b[3097]), .B(n4765), .Z(c[3097]) );
  XOR U8863 ( .A(n4766), .B(n4767), .Z(n4763) );
  ANDN U8864 ( .B(n4768), .A(n4769), .Z(n4766) );
  XNOR U8865 ( .A(b[3096]), .B(n4767), .Z(n4768) );
  XNOR U8866 ( .A(b[3096]), .B(n4769), .Z(c[3096]) );
  XOR U8867 ( .A(n4770), .B(n4771), .Z(n4767) );
  ANDN U8868 ( .B(n4772), .A(n4773), .Z(n4770) );
  XNOR U8869 ( .A(b[3095]), .B(n4771), .Z(n4772) );
  XNOR U8870 ( .A(b[3095]), .B(n4773), .Z(c[3095]) );
  XOR U8871 ( .A(n4774), .B(n4775), .Z(n4771) );
  ANDN U8872 ( .B(n4776), .A(n4777), .Z(n4774) );
  XNOR U8873 ( .A(b[3094]), .B(n4775), .Z(n4776) );
  XNOR U8874 ( .A(b[3094]), .B(n4777), .Z(c[3094]) );
  XOR U8875 ( .A(n4778), .B(n4779), .Z(n4775) );
  ANDN U8876 ( .B(n4780), .A(n4781), .Z(n4778) );
  XNOR U8877 ( .A(b[3093]), .B(n4779), .Z(n4780) );
  XNOR U8878 ( .A(b[3093]), .B(n4781), .Z(c[3093]) );
  XOR U8879 ( .A(n4782), .B(n4783), .Z(n4779) );
  ANDN U8880 ( .B(n4784), .A(n4785), .Z(n4782) );
  XNOR U8881 ( .A(b[3092]), .B(n4783), .Z(n4784) );
  XNOR U8882 ( .A(b[3092]), .B(n4785), .Z(c[3092]) );
  XOR U8883 ( .A(n4786), .B(n4787), .Z(n4783) );
  ANDN U8884 ( .B(n4788), .A(n4789), .Z(n4786) );
  XNOR U8885 ( .A(b[3091]), .B(n4787), .Z(n4788) );
  XNOR U8886 ( .A(b[3091]), .B(n4789), .Z(c[3091]) );
  XOR U8887 ( .A(n4790), .B(n4791), .Z(n4787) );
  ANDN U8888 ( .B(n4792), .A(n4793), .Z(n4790) );
  XNOR U8889 ( .A(b[3090]), .B(n4791), .Z(n4792) );
  XNOR U8890 ( .A(b[3090]), .B(n4793), .Z(c[3090]) );
  XOR U8891 ( .A(n4794), .B(n4795), .Z(n4791) );
  ANDN U8892 ( .B(n4796), .A(n4797), .Z(n4794) );
  XNOR U8893 ( .A(b[3089]), .B(n4795), .Z(n4796) );
  XNOR U8894 ( .A(b[308]), .B(n4798), .Z(c[308]) );
  XNOR U8895 ( .A(b[3089]), .B(n4797), .Z(c[3089]) );
  XOR U8896 ( .A(n4799), .B(n4800), .Z(n4795) );
  ANDN U8897 ( .B(n4801), .A(n4802), .Z(n4799) );
  XNOR U8898 ( .A(b[3088]), .B(n4800), .Z(n4801) );
  XNOR U8899 ( .A(b[3088]), .B(n4802), .Z(c[3088]) );
  XOR U8900 ( .A(n4803), .B(n4804), .Z(n4800) );
  ANDN U8901 ( .B(n4805), .A(n4806), .Z(n4803) );
  XNOR U8902 ( .A(b[3087]), .B(n4804), .Z(n4805) );
  XNOR U8903 ( .A(b[3087]), .B(n4806), .Z(c[3087]) );
  XOR U8904 ( .A(n4807), .B(n4808), .Z(n4804) );
  ANDN U8905 ( .B(n4809), .A(n4810), .Z(n4807) );
  XNOR U8906 ( .A(b[3086]), .B(n4808), .Z(n4809) );
  XNOR U8907 ( .A(b[3086]), .B(n4810), .Z(c[3086]) );
  XOR U8908 ( .A(n4811), .B(n4812), .Z(n4808) );
  ANDN U8909 ( .B(n4813), .A(n4814), .Z(n4811) );
  XNOR U8910 ( .A(b[3085]), .B(n4812), .Z(n4813) );
  XNOR U8911 ( .A(b[3085]), .B(n4814), .Z(c[3085]) );
  XOR U8912 ( .A(n4815), .B(n4816), .Z(n4812) );
  ANDN U8913 ( .B(n4817), .A(n4818), .Z(n4815) );
  XNOR U8914 ( .A(b[3084]), .B(n4816), .Z(n4817) );
  XNOR U8915 ( .A(b[3084]), .B(n4818), .Z(c[3084]) );
  XOR U8916 ( .A(n4819), .B(n4820), .Z(n4816) );
  ANDN U8917 ( .B(n4821), .A(n4822), .Z(n4819) );
  XNOR U8918 ( .A(b[3083]), .B(n4820), .Z(n4821) );
  XNOR U8919 ( .A(b[3083]), .B(n4822), .Z(c[3083]) );
  XOR U8920 ( .A(n4823), .B(n4824), .Z(n4820) );
  ANDN U8921 ( .B(n4825), .A(n4826), .Z(n4823) );
  XNOR U8922 ( .A(b[3082]), .B(n4824), .Z(n4825) );
  XNOR U8923 ( .A(b[3082]), .B(n4826), .Z(c[3082]) );
  XOR U8924 ( .A(n4827), .B(n4828), .Z(n4824) );
  ANDN U8925 ( .B(n4829), .A(n4830), .Z(n4827) );
  XNOR U8926 ( .A(b[3081]), .B(n4828), .Z(n4829) );
  XNOR U8927 ( .A(b[3081]), .B(n4830), .Z(c[3081]) );
  XOR U8928 ( .A(n4831), .B(n4832), .Z(n4828) );
  ANDN U8929 ( .B(n4833), .A(n4834), .Z(n4831) );
  XNOR U8930 ( .A(b[3080]), .B(n4832), .Z(n4833) );
  XNOR U8931 ( .A(b[3080]), .B(n4834), .Z(c[3080]) );
  XOR U8932 ( .A(n4835), .B(n4836), .Z(n4832) );
  ANDN U8933 ( .B(n4837), .A(n4838), .Z(n4835) );
  XNOR U8934 ( .A(b[3079]), .B(n4836), .Z(n4837) );
  XNOR U8935 ( .A(b[307]), .B(n4839), .Z(c[307]) );
  XNOR U8936 ( .A(b[3079]), .B(n4838), .Z(c[3079]) );
  XOR U8937 ( .A(n4840), .B(n4841), .Z(n4836) );
  ANDN U8938 ( .B(n4842), .A(n4843), .Z(n4840) );
  XNOR U8939 ( .A(b[3078]), .B(n4841), .Z(n4842) );
  XNOR U8940 ( .A(b[3078]), .B(n4843), .Z(c[3078]) );
  XOR U8941 ( .A(n4844), .B(n4845), .Z(n4841) );
  ANDN U8942 ( .B(n4846), .A(n4847), .Z(n4844) );
  XNOR U8943 ( .A(b[3077]), .B(n4845), .Z(n4846) );
  XNOR U8944 ( .A(b[3077]), .B(n4847), .Z(c[3077]) );
  XOR U8945 ( .A(n4848), .B(n4849), .Z(n4845) );
  ANDN U8946 ( .B(n4850), .A(n4851), .Z(n4848) );
  XNOR U8947 ( .A(b[3076]), .B(n4849), .Z(n4850) );
  XNOR U8948 ( .A(b[3076]), .B(n4851), .Z(c[3076]) );
  XOR U8949 ( .A(n4852), .B(n4853), .Z(n4849) );
  ANDN U8950 ( .B(n4854), .A(n4855), .Z(n4852) );
  XNOR U8951 ( .A(b[3075]), .B(n4853), .Z(n4854) );
  XNOR U8952 ( .A(b[3075]), .B(n4855), .Z(c[3075]) );
  XOR U8953 ( .A(n4856), .B(n4857), .Z(n4853) );
  ANDN U8954 ( .B(n4858), .A(n4859), .Z(n4856) );
  XNOR U8955 ( .A(b[3074]), .B(n4857), .Z(n4858) );
  XNOR U8956 ( .A(b[3074]), .B(n4859), .Z(c[3074]) );
  XOR U8957 ( .A(n4860), .B(n4861), .Z(n4857) );
  ANDN U8958 ( .B(n4862), .A(n4863), .Z(n4860) );
  XNOR U8959 ( .A(b[3073]), .B(n4861), .Z(n4862) );
  XNOR U8960 ( .A(b[3073]), .B(n4863), .Z(c[3073]) );
  XOR U8961 ( .A(n4864), .B(n4865), .Z(n4861) );
  ANDN U8962 ( .B(n4866), .A(n4867), .Z(n4864) );
  XNOR U8963 ( .A(b[3072]), .B(n4865), .Z(n4866) );
  XNOR U8964 ( .A(b[3072]), .B(n4867), .Z(c[3072]) );
  XOR U8965 ( .A(n4868), .B(n4869), .Z(n4865) );
  ANDN U8966 ( .B(n4870), .A(n4871), .Z(n4868) );
  XNOR U8967 ( .A(b[3071]), .B(n4869), .Z(n4870) );
  XNOR U8968 ( .A(b[3071]), .B(n4871), .Z(c[3071]) );
  XOR U8969 ( .A(n4872), .B(n4873), .Z(n4869) );
  ANDN U8970 ( .B(n4874), .A(n4875), .Z(n4872) );
  XNOR U8971 ( .A(b[3070]), .B(n4873), .Z(n4874) );
  XNOR U8972 ( .A(b[3070]), .B(n4875), .Z(c[3070]) );
  XOR U8973 ( .A(n4876), .B(n4877), .Z(n4873) );
  ANDN U8974 ( .B(n4878), .A(n4879), .Z(n4876) );
  XNOR U8975 ( .A(b[3069]), .B(n4877), .Z(n4878) );
  XNOR U8976 ( .A(b[306]), .B(n4880), .Z(c[306]) );
  XNOR U8977 ( .A(b[3069]), .B(n4879), .Z(c[3069]) );
  XOR U8978 ( .A(n4881), .B(n4882), .Z(n4877) );
  ANDN U8979 ( .B(n4883), .A(n4884), .Z(n4881) );
  XNOR U8980 ( .A(b[3068]), .B(n4882), .Z(n4883) );
  XNOR U8981 ( .A(b[3068]), .B(n4884), .Z(c[3068]) );
  XOR U8982 ( .A(n4885), .B(n4886), .Z(n4882) );
  ANDN U8983 ( .B(n4887), .A(n4888), .Z(n4885) );
  XNOR U8984 ( .A(b[3067]), .B(n4886), .Z(n4887) );
  XNOR U8985 ( .A(b[3067]), .B(n4888), .Z(c[3067]) );
  XOR U8986 ( .A(n4889), .B(n4890), .Z(n4886) );
  ANDN U8987 ( .B(n4891), .A(n4892), .Z(n4889) );
  XNOR U8988 ( .A(b[3066]), .B(n4890), .Z(n4891) );
  XNOR U8989 ( .A(b[3066]), .B(n4892), .Z(c[3066]) );
  XOR U8990 ( .A(n4893), .B(n4894), .Z(n4890) );
  ANDN U8991 ( .B(n4895), .A(n4896), .Z(n4893) );
  XNOR U8992 ( .A(b[3065]), .B(n4894), .Z(n4895) );
  XNOR U8993 ( .A(b[3065]), .B(n4896), .Z(c[3065]) );
  XOR U8994 ( .A(n4897), .B(n4898), .Z(n4894) );
  ANDN U8995 ( .B(n4899), .A(n4900), .Z(n4897) );
  XNOR U8996 ( .A(b[3064]), .B(n4898), .Z(n4899) );
  XNOR U8997 ( .A(b[3064]), .B(n4900), .Z(c[3064]) );
  XOR U8998 ( .A(n4901), .B(n4902), .Z(n4898) );
  ANDN U8999 ( .B(n4903), .A(n4904), .Z(n4901) );
  XNOR U9000 ( .A(b[3063]), .B(n4902), .Z(n4903) );
  XNOR U9001 ( .A(b[3063]), .B(n4904), .Z(c[3063]) );
  XOR U9002 ( .A(n4905), .B(n4906), .Z(n4902) );
  ANDN U9003 ( .B(n4907), .A(n4908), .Z(n4905) );
  XNOR U9004 ( .A(b[3062]), .B(n4906), .Z(n4907) );
  XNOR U9005 ( .A(b[3062]), .B(n4908), .Z(c[3062]) );
  XOR U9006 ( .A(n4909), .B(n4910), .Z(n4906) );
  ANDN U9007 ( .B(n4911), .A(n4912), .Z(n4909) );
  XNOR U9008 ( .A(b[3061]), .B(n4910), .Z(n4911) );
  XNOR U9009 ( .A(b[3061]), .B(n4912), .Z(c[3061]) );
  XOR U9010 ( .A(n4913), .B(n4914), .Z(n4910) );
  ANDN U9011 ( .B(n4915), .A(n4916), .Z(n4913) );
  XNOR U9012 ( .A(b[3060]), .B(n4914), .Z(n4915) );
  XNOR U9013 ( .A(b[3060]), .B(n4916), .Z(c[3060]) );
  XOR U9014 ( .A(n4917), .B(n4918), .Z(n4914) );
  ANDN U9015 ( .B(n4919), .A(n4920), .Z(n4917) );
  XNOR U9016 ( .A(b[3059]), .B(n4918), .Z(n4919) );
  XNOR U9017 ( .A(b[305]), .B(n4921), .Z(c[305]) );
  XNOR U9018 ( .A(b[3059]), .B(n4920), .Z(c[3059]) );
  XOR U9019 ( .A(n4922), .B(n4923), .Z(n4918) );
  ANDN U9020 ( .B(n4924), .A(n4925), .Z(n4922) );
  XNOR U9021 ( .A(b[3058]), .B(n4923), .Z(n4924) );
  XNOR U9022 ( .A(b[3058]), .B(n4925), .Z(c[3058]) );
  XOR U9023 ( .A(n4926), .B(n4927), .Z(n4923) );
  ANDN U9024 ( .B(n4928), .A(n4929), .Z(n4926) );
  XNOR U9025 ( .A(b[3057]), .B(n4927), .Z(n4928) );
  XNOR U9026 ( .A(b[3057]), .B(n4929), .Z(c[3057]) );
  XOR U9027 ( .A(n4930), .B(n4931), .Z(n4927) );
  ANDN U9028 ( .B(n4932), .A(n4933), .Z(n4930) );
  XNOR U9029 ( .A(b[3056]), .B(n4931), .Z(n4932) );
  XNOR U9030 ( .A(b[3056]), .B(n4933), .Z(c[3056]) );
  XOR U9031 ( .A(n4934), .B(n4935), .Z(n4931) );
  ANDN U9032 ( .B(n4936), .A(n4937), .Z(n4934) );
  XNOR U9033 ( .A(b[3055]), .B(n4935), .Z(n4936) );
  XNOR U9034 ( .A(b[3055]), .B(n4937), .Z(c[3055]) );
  XOR U9035 ( .A(n4938), .B(n4939), .Z(n4935) );
  ANDN U9036 ( .B(n4940), .A(n4941), .Z(n4938) );
  XNOR U9037 ( .A(b[3054]), .B(n4939), .Z(n4940) );
  XNOR U9038 ( .A(b[3054]), .B(n4941), .Z(c[3054]) );
  XOR U9039 ( .A(n4942), .B(n4943), .Z(n4939) );
  ANDN U9040 ( .B(n4944), .A(n4945), .Z(n4942) );
  XNOR U9041 ( .A(b[3053]), .B(n4943), .Z(n4944) );
  XNOR U9042 ( .A(b[3053]), .B(n4945), .Z(c[3053]) );
  XOR U9043 ( .A(n4946), .B(n4947), .Z(n4943) );
  ANDN U9044 ( .B(n4948), .A(n4949), .Z(n4946) );
  XNOR U9045 ( .A(b[3052]), .B(n4947), .Z(n4948) );
  XNOR U9046 ( .A(b[3052]), .B(n4949), .Z(c[3052]) );
  XOR U9047 ( .A(n4950), .B(n4951), .Z(n4947) );
  ANDN U9048 ( .B(n4952), .A(n4953), .Z(n4950) );
  XNOR U9049 ( .A(b[3051]), .B(n4951), .Z(n4952) );
  XNOR U9050 ( .A(b[3051]), .B(n4953), .Z(c[3051]) );
  XOR U9051 ( .A(n4954), .B(n4955), .Z(n4951) );
  ANDN U9052 ( .B(n4956), .A(n4957), .Z(n4954) );
  XNOR U9053 ( .A(b[3050]), .B(n4955), .Z(n4956) );
  XNOR U9054 ( .A(b[3050]), .B(n4957), .Z(c[3050]) );
  XOR U9055 ( .A(n4958), .B(n4959), .Z(n4955) );
  ANDN U9056 ( .B(n4960), .A(n4961), .Z(n4958) );
  XNOR U9057 ( .A(b[3049]), .B(n4959), .Z(n4960) );
  XNOR U9058 ( .A(b[304]), .B(n4962), .Z(c[304]) );
  XNOR U9059 ( .A(b[3049]), .B(n4961), .Z(c[3049]) );
  XOR U9060 ( .A(n4963), .B(n4964), .Z(n4959) );
  ANDN U9061 ( .B(n4965), .A(n4966), .Z(n4963) );
  XNOR U9062 ( .A(b[3048]), .B(n4964), .Z(n4965) );
  XNOR U9063 ( .A(b[3048]), .B(n4966), .Z(c[3048]) );
  XOR U9064 ( .A(n4967), .B(n4968), .Z(n4964) );
  ANDN U9065 ( .B(n4969), .A(n4970), .Z(n4967) );
  XNOR U9066 ( .A(b[3047]), .B(n4968), .Z(n4969) );
  XNOR U9067 ( .A(b[3047]), .B(n4970), .Z(c[3047]) );
  XOR U9068 ( .A(n4971), .B(n4972), .Z(n4968) );
  ANDN U9069 ( .B(n4973), .A(n4974), .Z(n4971) );
  XNOR U9070 ( .A(b[3046]), .B(n4972), .Z(n4973) );
  XNOR U9071 ( .A(b[3046]), .B(n4974), .Z(c[3046]) );
  XOR U9072 ( .A(n4975), .B(n4976), .Z(n4972) );
  ANDN U9073 ( .B(n4977), .A(n4978), .Z(n4975) );
  XNOR U9074 ( .A(b[3045]), .B(n4976), .Z(n4977) );
  XNOR U9075 ( .A(b[3045]), .B(n4978), .Z(c[3045]) );
  XOR U9076 ( .A(n4979), .B(n4980), .Z(n4976) );
  ANDN U9077 ( .B(n4981), .A(n4982), .Z(n4979) );
  XNOR U9078 ( .A(b[3044]), .B(n4980), .Z(n4981) );
  XNOR U9079 ( .A(b[3044]), .B(n4982), .Z(c[3044]) );
  XOR U9080 ( .A(n4983), .B(n4984), .Z(n4980) );
  ANDN U9081 ( .B(n4985), .A(n4986), .Z(n4983) );
  XNOR U9082 ( .A(b[3043]), .B(n4984), .Z(n4985) );
  XNOR U9083 ( .A(b[3043]), .B(n4986), .Z(c[3043]) );
  XOR U9084 ( .A(n4987), .B(n4988), .Z(n4984) );
  ANDN U9085 ( .B(n4989), .A(n4990), .Z(n4987) );
  XNOR U9086 ( .A(b[3042]), .B(n4988), .Z(n4989) );
  XNOR U9087 ( .A(b[3042]), .B(n4990), .Z(c[3042]) );
  XOR U9088 ( .A(n4991), .B(n4992), .Z(n4988) );
  ANDN U9089 ( .B(n4993), .A(n4994), .Z(n4991) );
  XNOR U9090 ( .A(b[3041]), .B(n4992), .Z(n4993) );
  XNOR U9091 ( .A(b[3041]), .B(n4994), .Z(c[3041]) );
  XOR U9092 ( .A(n4995), .B(n4996), .Z(n4992) );
  ANDN U9093 ( .B(n4997), .A(n4998), .Z(n4995) );
  XNOR U9094 ( .A(b[3040]), .B(n4996), .Z(n4997) );
  XNOR U9095 ( .A(b[3040]), .B(n4998), .Z(c[3040]) );
  XOR U9096 ( .A(n4999), .B(n5000), .Z(n4996) );
  ANDN U9097 ( .B(n5001), .A(n5002), .Z(n4999) );
  XNOR U9098 ( .A(b[3039]), .B(n5000), .Z(n5001) );
  XNOR U9099 ( .A(b[303]), .B(n5003), .Z(c[303]) );
  XNOR U9100 ( .A(b[3039]), .B(n5002), .Z(c[3039]) );
  XOR U9101 ( .A(n5004), .B(n5005), .Z(n5000) );
  ANDN U9102 ( .B(n5006), .A(n5007), .Z(n5004) );
  XNOR U9103 ( .A(b[3038]), .B(n5005), .Z(n5006) );
  XNOR U9104 ( .A(b[3038]), .B(n5007), .Z(c[3038]) );
  XOR U9105 ( .A(n5008), .B(n5009), .Z(n5005) );
  ANDN U9106 ( .B(n5010), .A(n5011), .Z(n5008) );
  XNOR U9107 ( .A(b[3037]), .B(n5009), .Z(n5010) );
  XNOR U9108 ( .A(b[3037]), .B(n5011), .Z(c[3037]) );
  XOR U9109 ( .A(n5012), .B(n5013), .Z(n5009) );
  ANDN U9110 ( .B(n5014), .A(n5015), .Z(n5012) );
  XNOR U9111 ( .A(b[3036]), .B(n5013), .Z(n5014) );
  XNOR U9112 ( .A(b[3036]), .B(n5015), .Z(c[3036]) );
  XOR U9113 ( .A(n5016), .B(n5017), .Z(n5013) );
  ANDN U9114 ( .B(n5018), .A(n5019), .Z(n5016) );
  XNOR U9115 ( .A(b[3035]), .B(n5017), .Z(n5018) );
  XNOR U9116 ( .A(b[3035]), .B(n5019), .Z(c[3035]) );
  XOR U9117 ( .A(n5020), .B(n5021), .Z(n5017) );
  ANDN U9118 ( .B(n5022), .A(n5023), .Z(n5020) );
  XNOR U9119 ( .A(b[3034]), .B(n5021), .Z(n5022) );
  XNOR U9120 ( .A(b[3034]), .B(n5023), .Z(c[3034]) );
  XOR U9121 ( .A(n5024), .B(n5025), .Z(n5021) );
  ANDN U9122 ( .B(n5026), .A(n5027), .Z(n5024) );
  XNOR U9123 ( .A(b[3033]), .B(n5025), .Z(n5026) );
  XNOR U9124 ( .A(b[3033]), .B(n5027), .Z(c[3033]) );
  XOR U9125 ( .A(n5028), .B(n5029), .Z(n5025) );
  ANDN U9126 ( .B(n5030), .A(n5031), .Z(n5028) );
  XNOR U9127 ( .A(b[3032]), .B(n5029), .Z(n5030) );
  XNOR U9128 ( .A(b[3032]), .B(n5031), .Z(c[3032]) );
  XOR U9129 ( .A(n5032), .B(n5033), .Z(n5029) );
  ANDN U9130 ( .B(n5034), .A(n5035), .Z(n5032) );
  XNOR U9131 ( .A(b[3031]), .B(n5033), .Z(n5034) );
  XNOR U9132 ( .A(b[3031]), .B(n5035), .Z(c[3031]) );
  XOR U9133 ( .A(n5036), .B(n5037), .Z(n5033) );
  ANDN U9134 ( .B(n5038), .A(n5039), .Z(n5036) );
  XNOR U9135 ( .A(b[3030]), .B(n5037), .Z(n5038) );
  XNOR U9136 ( .A(b[3030]), .B(n5039), .Z(c[3030]) );
  XOR U9137 ( .A(n5040), .B(n5041), .Z(n5037) );
  ANDN U9138 ( .B(n5042), .A(n5043), .Z(n5040) );
  XNOR U9139 ( .A(b[3029]), .B(n5041), .Z(n5042) );
  XNOR U9140 ( .A(b[302]), .B(n5044), .Z(c[302]) );
  XNOR U9141 ( .A(b[3029]), .B(n5043), .Z(c[3029]) );
  XOR U9142 ( .A(n5045), .B(n5046), .Z(n5041) );
  ANDN U9143 ( .B(n5047), .A(n5048), .Z(n5045) );
  XNOR U9144 ( .A(b[3028]), .B(n5046), .Z(n5047) );
  XNOR U9145 ( .A(b[3028]), .B(n5048), .Z(c[3028]) );
  XOR U9146 ( .A(n5049), .B(n5050), .Z(n5046) );
  ANDN U9147 ( .B(n5051), .A(n5052), .Z(n5049) );
  XNOR U9148 ( .A(b[3027]), .B(n5050), .Z(n5051) );
  XNOR U9149 ( .A(b[3027]), .B(n5052), .Z(c[3027]) );
  XOR U9150 ( .A(n5053), .B(n5054), .Z(n5050) );
  ANDN U9151 ( .B(n5055), .A(n5056), .Z(n5053) );
  XNOR U9152 ( .A(b[3026]), .B(n5054), .Z(n5055) );
  XNOR U9153 ( .A(b[3026]), .B(n5056), .Z(c[3026]) );
  XOR U9154 ( .A(n5057), .B(n5058), .Z(n5054) );
  ANDN U9155 ( .B(n5059), .A(n5060), .Z(n5057) );
  XNOR U9156 ( .A(b[3025]), .B(n5058), .Z(n5059) );
  XNOR U9157 ( .A(b[3025]), .B(n5060), .Z(c[3025]) );
  XOR U9158 ( .A(n5061), .B(n5062), .Z(n5058) );
  ANDN U9159 ( .B(n5063), .A(n5064), .Z(n5061) );
  XNOR U9160 ( .A(b[3024]), .B(n5062), .Z(n5063) );
  XNOR U9161 ( .A(b[3024]), .B(n5064), .Z(c[3024]) );
  XOR U9162 ( .A(n5065), .B(n5066), .Z(n5062) );
  ANDN U9163 ( .B(n5067), .A(n5068), .Z(n5065) );
  XNOR U9164 ( .A(b[3023]), .B(n5066), .Z(n5067) );
  XNOR U9165 ( .A(b[3023]), .B(n5068), .Z(c[3023]) );
  XOR U9166 ( .A(n5069), .B(n5070), .Z(n5066) );
  ANDN U9167 ( .B(n5071), .A(n5072), .Z(n5069) );
  XNOR U9168 ( .A(b[3022]), .B(n5070), .Z(n5071) );
  XNOR U9169 ( .A(b[3022]), .B(n5072), .Z(c[3022]) );
  XOR U9170 ( .A(n5073), .B(n5074), .Z(n5070) );
  ANDN U9171 ( .B(n5075), .A(n5076), .Z(n5073) );
  XNOR U9172 ( .A(b[3021]), .B(n5074), .Z(n5075) );
  XNOR U9173 ( .A(b[3021]), .B(n5076), .Z(c[3021]) );
  XOR U9174 ( .A(n5077), .B(n5078), .Z(n5074) );
  ANDN U9175 ( .B(n5079), .A(n5080), .Z(n5077) );
  XNOR U9176 ( .A(b[3020]), .B(n5078), .Z(n5079) );
  XNOR U9177 ( .A(b[3020]), .B(n5080), .Z(c[3020]) );
  XOR U9178 ( .A(n5081), .B(n5082), .Z(n5078) );
  ANDN U9179 ( .B(n5083), .A(n5084), .Z(n5081) );
  XNOR U9180 ( .A(b[3019]), .B(n5082), .Z(n5083) );
  XNOR U9181 ( .A(b[301]), .B(n5085), .Z(c[301]) );
  XNOR U9182 ( .A(b[3019]), .B(n5084), .Z(c[3019]) );
  XOR U9183 ( .A(n5086), .B(n5087), .Z(n5082) );
  ANDN U9184 ( .B(n5088), .A(n5089), .Z(n5086) );
  XNOR U9185 ( .A(b[3018]), .B(n5087), .Z(n5088) );
  XNOR U9186 ( .A(b[3018]), .B(n5089), .Z(c[3018]) );
  XOR U9187 ( .A(n5090), .B(n5091), .Z(n5087) );
  ANDN U9188 ( .B(n5092), .A(n5093), .Z(n5090) );
  XNOR U9189 ( .A(b[3017]), .B(n5091), .Z(n5092) );
  XNOR U9190 ( .A(b[3017]), .B(n5093), .Z(c[3017]) );
  XOR U9191 ( .A(n5094), .B(n5095), .Z(n5091) );
  ANDN U9192 ( .B(n5096), .A(n5097), .Z(n5094) );
  XNOR U9193 ( .A(b[3016]), .B(n5095), .Z(n5096) );
  XNOR U9194 ( .A(b[3016]), .B(n5097), .Z(c[3016]) );
  XOR U9195 ( .A(n5098), .B(n5099), .Z(n5095) );
  ANDN U9196 ( .B(n5100), .A(n5101), .Z(n5098) );
  XNOR U9197 ( .A(b[3015]), .B(n5099), .Z(n5100) );
  XNOR U9198 ( .A(b[3015]), .B(n5101), .Z(c[3015]) );
  XOR U9199 ( .A(n5102), .B(n5103), .Z(n5099) );
  ANDN U9200 ( .B(n5104), .A(n5105), .Z(n5102) );
  XNOR U9201 ( .A(b[3014]), .B(n5103), .Z(n5104) );
  XNOR U9202 ( .A(b[3014]), .B(n5105), .Z(c[3014]) );
  XOR U9203 ( .A(n5106), .B(n5107), .Z(n5103) );
  ANDN U9204 ( .B(n5108), .A(n5109), .Z(n5106) );
  XNOR U9205 ( .A(b[3013]), .B(n5107), .Z(n5108) );
  XNOR U9206 ( .A(b[3013]), .B(n5109), .Z(c[3013]) );
  XOR U9207 ( .A(n5110), .B(n5111), .Z(n5107) );
  ANDN U9208 ( .B(n5112), .A(n5113), .Z(n5110) );
  XNOR U9209 ( .A(b[3012]), .B(n5111), .Z(n5112) );
  XNOR U9210 ( .A(b[3012]), .B(n5113), .Z(c[3012]) );
  XOR U9211 ( .A(n5114), .B(n5115), .Z(n5111) );
  ANDN U9212 ( .B(n5116), .A(n5117), .Z(n5114) );
  XNOR U9213 ( .A(b[3011]), .B(n5115), .Z(n5116) );
  XNOR U9214 ( .A(b[3011]), .B(n5117), .Z(c[3011]) );
  XOR U9215 ( .A(n5118), .B(n5119), .Z(n5115) );
  ANDN U9216 ( .B(n5120), .A(n5121), .Z(n5118) );
  XNOR U9217 ( .A(b[3010]), .B(n5119), .Z(n5120) );
  XNOR U9218 ( .A(b[3010]), .B(n5121), .Z(c[3010]) );
  XOR U9219 ( .A(n5122), .B(n5123), .Z(n5119) );
  ANDN U9220 ( .B(n5124), .A(n5125), .Z(n5122) );
  XNOR U9221 ( .A(b[3009]), .B(n5123), .Z(n5124) );
  XNOR U9222 ( .A(b[300]), .B(n5126), .Z(c[300]) );
  XNOR U9223 ( .A(b[3009]), .B(n5125), .Z(c[3009]) );
  XOR U9224 ( .A(n5127), .B(n5128), .Z(n5123) );
  ANDN U9225 ( .B(n5129), .A(n5130), .Z(n5127) );
  XNOR U9226 ( .A(b[3008]), .B(n5128), .Z(n5129) );
  XNOR U9227 ( .A(b[3008]), .B(n5130), .Z(c[3008]) );
  XOR U9228 ( .A(n5131), .B(n5132), .Z(n5128) );
  ANDN U9229 ( .B(n5133), .A(n5134), .Z(n5131) );
  XNOR U9230 ( .A(b[3007]), .B(n5132), .Z(n5133) );
  XNOR U9231 ( .A(b[3007]), .B(n5134), .Z(c[3007]) );
  XOR U9232 ( .A(n5135), .B(n5136), .Z(n5132) );
  ANDN U9233 ( .B(n5137), .A(n5138), .Z(n5135) );
  XNOR U9234 ( .A(b[3006]), .B(n5136), .Z(n5137) );
  XNOR U9235 ( .A(b[3006]), .B(n5138), .Z(c[3006]) );
  XOR U9236 ( .A(n5139), .B(n5140), .Z(n5136) );
  ANDN U9237 ( .B(n5141), .A(n5142), .Z(n5139) );
  XNOR U9238 ( .A(b[3005]), .B(n5140), .Z(n5141) );
  XNOR U9239 ( .A(b[3005]), .B(n5142), .Z(c[3005]) );
  XOR U9240 ( .A(n5143), .B(n5144), .Z(n5140) );
  ANDN U9241 ( .B(n5145), .A(n5146), .Z(n5143) );
  XNOR U9242 ( .A(b[3004]), .B(n5144), .Z(n5145) );
  XNOR U9243 ( .A(b[3004]), .B(n5146), .Z(c[3004]) );
  XOR U9244 ( .A(n5147), .B(n5148), .Z(n5144) );
  ANDN U9245 ( .B(n5149), .A(n5150), .Z(n5147) );
  XNOR U9246 ( .A(b[3003]), .B(n5148), .Z(n5149) );
  XNOR U9247 ( .A(b[3003]), .B(n5150), .Z(c[3003]) );
  XOR U9248 ( .A(n5151), .B(n5152), .Z(n5148) );
  ANDN U9249 ( .B(n5153), .A(n5154), .Z(n5151) );
  XNOR U9250 ( .A(b[3002]), .B(n5152), .Z(n5153) );
  XNOR U9251 ( .A(b[3002]), .B(n5154), .Z(c[3002]) );
  XOR U9252 ( .A(n5155), .B(n5156), .Z(n5152) );
  ANDN U9253 ( .B(n5157), .A(n5158), .Z(n5155) );
  XNOR U9254 ( .A(b[3001]), .B(n5156), .Z(n5157) );
  XNOR U9255 ( .A(b[3001]), .B(n5158), .Z(c[3001]) );
  XOR U9256 ( .A(n5159), .B(n5160), .Z(n5156) );
  ANDN U9257 ( .B(n5161), .A(n5162), .Z(n5159) );
  XNOR U9258 ( .A(b[3000]), .B(n5160), .Z(n5161) );
  XNOR U9259 ( .A(b[3000]), .B(n5162), .Z(c[3000]) );
  XOR U9260 ( .A(n5163), .B(n5164), .Z(n5160) );
  ANDN U9261 ( .B(n5165), .A(n5166), .Z(n5163) );
  XNOR U9262 ( .A(b[2999]), .B(n5164), .Z(n5165) );
  XNOR U9263 ( .A(b[2]), .B(n5167), .Z(c[2]) );
  XNOR U9264 ( .A(b[29]), .B(n5168), .Z(c[29]) );
  XNOR U9265 ( .A(b[299]), .B(n5169), .Z(c[299]) );
  XNOR U9266 ( .A(b[2999]), .B(n5166), .Z(c[2999]) );
  XOR U9267 ( .A(n5170), .B(n5171), .Z(n5164) );
  ANDN U9268 ( .B(n5172), .A(n5173), .Z(n5170) );
  XNOR U9269 ( .A(b[2998]), .B(n5171), .Z(n5172) );
  XNOR U9270 ( .A(b[2998]), .B(n5173), .Z(c[2998]) );
  XOR U9271 ( .A(n5174), .B(n5175), .Z(n5171) );
  ANDN U9272 ( .B(n5176), .A(n5177), .Z(n5174) );
  XNOR U9273 ( .A(b[2997]), .B(n5175), .Z(n5176) );
  XNOR U9274 ( .A(b[2997]), .B(n5177), .Z(c[2997]) );
  XOR U9275 ( .A(n5178), .B(n5179), .Z(n5175) );
  ANDN U9276 ( .B(n5180), .A(n5181), .Z(n5178) );
  XNOR U9277 ( .A(b[2996]), .B(n5179), .Z(n5180) );
  XNOR U9278 ( .A(b[2996]), .B(n5181), .Z(c[2996]) );
  XOR U9279 ( .A(n5182), .B(n5183), .Z(n5179) );
  ANDN U9280 ( .B(n5184), .A(n5185), .Z(n5182) );
  XNOR U9281 ( .A(b[2995]), .B(n5183), .Z(n5184) );
  XNOR U9282 ( .A(b[2995]), .B(n5185), .Z(c[2995]) );
  XOR U9283 ( .A(n5186), .B(n5187), .Z(n5183) );
  ANDN U9284 ( .B(n5188), .A(n5189), .Z(n5186) );
  XNOR U9285 ( .A(b[2994]), .B(n5187), .Z(n5188) );
  XNOR U9286 ( .A(b[2994]), .B(n5189), .Z(c[2994]) );
  XOR U9287 ( .A(n5190), .B(n5191), .Z(n5187) );
  ANDN U9288 ( .B(n5192), .A(n5193), .Z(n5190) );
  XNOR U9289 ( .A(b[2993]), .B(n5191), .Z(n5192) );
  XNOR U9290 ( .A(b[2993]), .B(n5193), .Z(c[2993]) );
  XOR U9291 ( .A(n5194), .B(n5195), .Z(n5191) );
  ANDN U9292 ( .B(n5196), .A(n5197), .Z(n5194) );
  XNOR U9293 ( .A(b[2992]), .B(n5195), .Z(n5196) );
  XNOR U9294 ( .A(b[2992]), .B(n5197), .Z(c[2992]) );
  XOR U9295 ( .A(n5198), .B(n5199), .Z(n5195) );
  ANDN U9296 ( .B(n5200), .A(n5201), .Z(n5198) );
  XNOR U9297 ( .A(b[2991]), .B(n5199), .Z(n5200) );
  XNOR U9298 ( .A(b[2991]), .B(n5201), .Z(c[2991]) );
  XOR U9299 ( .A(n5202), .B(n5203), .Z(n5199) );
  ANDN U9300 ( .B(n5204), .A(n5205), .Z(n5202) );
  XNOR U9301 ( .A(b[2990]), .B(n5203), .Z(n5204) );
  XNOR U9302 ( .A(b[2990]), .B(n5205), .Z(c[2990]) );
  XOR U9303 ( .A(n5206), .B(n5207), .Z(n5203) );
  ANDN U9304 ( .B(n5208), .A(n5209), .Z(n5206) );
  XNOR U9305 ( .A(b[2989]), .B(n5207), .Z(n5208) );
  XNOR U9306 ( .A(b[298]), .B(n5210), .Z(c[298]) );
  XNOR U9307 ( .A(b[2989]), .B(n5209), .Z(c[2989]) );
  XOR U9308 ( .A(n5211), .B(n5212), .Z(n5207) );
  ANDN U9309 ( .B(n5213), .A(n5214), .Z(n5211) );
  XNOR U9310 ( .A(b[2988]), .B(n5212), .Z(n5213) );
  XNOR U9311 ( .A(b[2988]), .B(n5214), .Z(c[2988]) );
  XOR U9312 ( .A(n5215), .B(n5216), .Z(n5212) );
  ANDN U9313 ( .B(n5217), .A(n5218), .Z(n5215) );
  XNOR U9314 ( .A(b[2987]), .B(n5216), .Z(n5217) );
  XNOR U9315 ( .A(b[2987]), .B(n5218), .Z(c[2987]) );
  XOR U9316 ( .A(n5219), .B(n5220), .Z(n5216) );
  ANDN U9317 ( .B(n5221), .A(n5222), .Z(n5219) );
  XNOR U9318 ( .A(b[2986]), .B(n5220), .Z(n5221) );
  XNOR U9319 ( .A(b[2986]), .B(n5222), .Z(c[2986]) );
  XOR U9320 ( .A(n5223), .B(n5224), .Z(n5220) );
  ANDN U9321 ( .B(n5225), .A(n5226), .Z(n5223) );
  XNOR U9322 ( .A(b[2985]), .B(n5224), .Z(n5225) );
  XNOR U9323 ( .A(b[2985]), .B(n5226), .Z(c[2985]) );
  XOR U9324 ( .A(n5227), .B(n5228), .Z(n5224) );
  ANDN U9325 ( .B(n5229), .A(n5230), .Z(n5227) );
  XNOR U9326 ( .A(b[2984]), .B(n5228), .Z(n5229) );
  XNOR U9327 ( .A(b[2984]), .B(n5230), .Z(c[2984]) );
  XOR U9328 ( .A(n5231), .B(n5232), .Z(n5228) );
  ANDN U9329 ( .B(n5233), .A(n5234), .Z(n5231) );
  XNOR U9330 ( .A(b[2983]), .B(n5232), .Z(n5233) );
  XNOR U9331 ( .A(b[2983]), .B(n5234), .Z(c[2983]) );
  XOR U9332 ( .A(n5235), .B(n5236), .Z(n5232) );
  ANDN U9333 ( .B(n5237), .A(n5238), .Z(n5235) );
  XNOR U9334 ( .A(b[2982]), .B(n5236), .Z(n5237) );
  XNOR U9335 ( .A(b[2982]), .B(n5238), .Z(c[2982]) );
  XOR U9336 ( .A(n5239), .B(n5240), .Z(n5236) );
  ANDN U9337 ( .B(n5241), .A(n5242), .Z(n5239) );
  XNOR U9338 ( .A(b[2981]), .B(n5240), .Z(n5241) );
  XNOR U9339 ( .A(b[2981]), .B(n5242), .Z(c[2981]) );
  XOR U9340 ( .A(n5243), .B(n5244), .Z(n5240) );
  ANDN U9341 ( .B(n5245), .A(n5246), .Z(n5243) );
  XNOR U9342 ( .A(b[2980]), .B(n5244), .Z(n5245) );
  XNOR U9343 ( .A(b[2980]), .B(n5246), .Z(c[2980]) );
  XOR U9344 ( .A(n5247), .B(n5248), .Z(n5244) );
  ANDN U9345 ( .B(n5249), .A(n5250), .Z(n5247) );
  XNOR U9346 ( .A(b[2979]), .B(n5248), .Z(n5249) );
  XNOR U9347 ( .A(b[297]), .B(n5251), .Z(c[297]) );
  XNOR U9348 ( .A(b[2979]), .B(n5250), .Z(c[2979]) );
  XOR U9349 ( .A(n5252), .B(n5253), .Z(n5248) );
  ANDN U9350 ( .B(n5254), .A(n5255), .Z(n5252) );
  XNOR U9351 ( .A(b[2978]), .B(n5253), .Z(n5254) );
  XNOR U9352 ( .A(b[2978]), .B(n5255), .Z(c[2978]) );
  XOR U9353 ( .A(n5256), .B(n5257), .Z(n5253) );
  ANDN U9354 ( .B(n5258), .A(n5259), .Z(n5256) );
  XNOR U9355 ( .A(b[2977]), .B(n5257), .Z(n5258) );
  XNOR U9356 ( .A(b[2977]), .B(n5259), .Z(c[2977]) );
  XOR U9357 ( .A(n5260), .B(n5261), .Z(n5257) );
  ANDN U9358 ( .B(n5262), .A(n5263), .Z(n5260) );
  XNOR U9359 ( .A(b[2976]), .B(n5261), .Z(n5262) );
  XNOR U9360 ( .A(b[2976]), .B(n5263), .Z(c[2976]) );
  XOR U9361 ( .A(n5264), .B(n5265), .Z(n5261) );
  ANDN U9362 ( .B(n5266), .A(n5267), .Z(n5264) );
  XNOR U9363 ( .A(b[2975]), .B(n5265), .Z(n5266) );
  XNOR U9364 ( .A(b[2975]), .B(n5267), .Z(c[2975]) );
  XOR U9365 ( .A(n5268), .B(n5269), .Z(n5265) );
  ANDN U9366 ( .B(n5270), .A(n5271), .Z(n5268) );
  XNOR U9367 ( .A(b[2974]), .B(n5269), .Z(n5270) );
  XNOR U9368 ( .A(b[2974]), .B(n5271), .Z(c[2974]) );
  XOR U9369 ( .A(n5272), .B(n5273), .Z(n5269) );
  ANDN U9370 ( .B(n5274), .A(n5275), .Z(n5272) );
  XNOR U9371 ( .A(b[2973]), .B(n5273), .Z(n5274) );
  XNOR U9372 ( .A(b[2973]), .B(n5275), .Z(c[2973]) );
  XOR U9373 ( .A(n5276), .B(n5277), .Z(n5273) );
  ANDN U9374 ( .B(n5278), .A(n5279), .Z(n5276) );
  XNOR U9375 ( .A(b[2972]), .B(n5277), .Z(n5278) );
  XNOR U9376 ( .A(b[2972]), .B(n5279), .Z(c[2972]) );
  XOR U9377 ( .A(n5280), .B(n5281), .Z(n5277) );
  ANDN U9378 ( .B(n5282), .A(n5283), .Z(n5280) );
  XNOR U9379 ( .A(b[2971]), .B(n5281), .Z(n5282) );
  XNOR U9380 ( .A(b[2971]), .B(n5283), .Z(c[2971]) );
  XOR U9381 ( .A(n5284), .B(n5285), .Z(n5281) );
  ANDN U9382 ( .B(n5286), .A(n5287), .Z(n5284) );
  XNOR U9383 ( .A(b[2970]), .B(n5285), .Z(n5286) );
  XNOR U9384 ( .A(b[2970]), .B(n5287), .Z(c[2970]) );
  XOR U9385 ( .A(n5288), .B(n5289), .Z(n5285) );
  ANDN U9386 ( .B(n5290), .A(n5291), .Z(n5288) );
  XNOR U9387 ( .A(b[2969]), .B(n5289), .Z(n5290) );
  XNOR U9388 ( .A(b[296]), .B(n5292), .Z(c[296]) );
  XNOR U9389 ( .A(b[2969]), .B(n5291), .Z(c[2969]) );
  XOR U9390 ( .A(n5293), .B(n5294), .Z(n5289) );
  ANDN U9391 ( .B(n5295), .A(n5296), .Z(n5293) );
  XNOR U9392 ( .A(b[2968]), .B(n5294), .Z(n5295) );
  XNOR U9393 ( .A(b[2968]), .B(n5296), .Z(c[2968]) );
  XOR U9394 ( .A(n5297), .B(n5298), .Z(n5294) );
  ANDN U9395 ( .B(n5299), .A(n5300), .Z(n5297) );
  XNOR U9396 ( .A(b[2967]), .B(n5298), .Z(n5299) );
  XNOR U9397 ( .A(b[2967]), .B(n5300), .Z(c[2967]) );
  XOR U9398 ( .A(n5301), .B(n5302), .Z(n5298) );
  ANDN U9399 ( .B(n5303), .A(n5304), .Z(n5301) );
  XNOR U9400 ( .A(b[2966]), .B(n5302), .Z(n5303) );
  XNOR U9401 ( .A(b[2966]), .B(n5304), .Z(c[2966]) );
  XOR U9402 ( .A(n5305), .B(n5306), .Z(n5302) );
  ANDN U9403 ( .B(n5307), .A(n5308), .Z(n5305) );
  XNOR U9404 ( .A(b[2965]), .B(n5306), .Z(n5307) );
  XNOR U9405 ( .A(b[2965]), .B(n5308), .Z(c[2965]) );
  XOR U9406 ( .A(n5309), .B(n5310), .Z(n5306) );
  ANDN U9407 ( .B(n5311), .A(n5312), .Z(n5309) );
  XNOR U9408 ( .A(b[2964]), .B(n5310), .Z(n5311) );
  XNOR U9409 ( .A(b[2964]), .B(n5312), .Z(c[2964]) );
  XOR U9410 ( .A(n5313), .B(n5314), .Z(n5310) );
  ANDN U9411 ( .B(n5315), .A(n5316), .Z(n5313) );
  XNOR U9412 ( .A(b[2963]), .B(n5314), .Z(n5315) );
  XNOR U9413 ( .A(b[2963]), .B(n5316), .Z(c[2963]) );
  XOR U9414 ( .A(n5317), .B(n5318), .Z(n5314) );
  ANDN U9415 ( .B(n5319), .A(n5320), .Z(n5317) );
  XNOR U9416 ( .A(b[2962]), .B(n5318), .Z(n5319) );
  XNOR U9417 ( .A(b[2962]), .B(n5320), .Z(c[2962]) );
  XOR U9418 ( .A(n5321), .B(n5322), .Z(n5318) );
  ANDN U9419 ( .B(n5323), .A(n5324), .Z(n5321) );
  XNOR U9420 ( .A(b[2961]), .B(n5322), .Z(n5323) );
  XNOR U9421 ( .A(b[2961]), .B(n5324), .Z(c[2961]) );
  XOR U9422 ( .A(n5325), .B(n5326), .Z(n5322) );
  ANDN U9423 ( .B(n5327), .A(n5328), .Z(n5325) );
  XNOR U9424 ( .A(b[2960]), .B(n5326), .Z(n5327) );
  XNOR U9425 ( .A(b[2960]), .B(n5328), .Z(c[2960]) );
  XOR U9426 ( .A(n5329), .B(n5330), .Z(n5326) );
  ANDN U9427 ( .B(n5331), .A(n5332), .Z(n5329) );
  XNOR U9428 ( .A(b[2959]), .B(n5330), .Z(n5331) );
  XNOR U9429 ( .A(b[295]), .B(n5333), .Z(c[295]) );
  XNOR U9430 ( .A(b[2959]), .B(n5332), .Z(c[2959]) );
  XOR U9431 ( .A(n5334), .B(n5335), .Z(n5330) );
  ANDN U9432 ( .B(n5336), .A(n5337), .Z(n5334) );
  XNOR U9433 ( .A(b[2958]), .B(n5335), .Z(n5336) );
  XNOR U9434 ( .A(b[2958]), .B(n5337), .Z(c[2958]) );
  XOR U9435 ( .A(n5338), .B(n5339), .Z(n5335) );
  ANDN U9436 ( .B(n5340), .A(n5341), .Z(n5338) );
  XNOR U9437 ( .A(b[2957]), .B(n5339), .Z(n5340) );
  XNOR U9438 ( .A(b[2957]), .B(n5341), .Z(c[2957]) );
  XOR U9439 ( .A(n5342), .B(n5343), .Z(n5339) );
  ANDN U9440 ( .B(n5344), .A(n5345), .Z(n5342) );
  XNOR U9441 ( .A(b[2956]), .B(n5343), .Z(n5344) );
  XNOR U9442 ( .A(b[2956]), .B(n5345), .Z(c[2956]) );
  XOR U9443 ( .A(n5346), .B(n5347), .Z(n5343) );
  ANDN U9444 ( .B(n5348), .A(n5349), .Z(n5346) );
  XNOR U9445 ( .A(b[2955]), .B(n5347), .Z(n5348) );
  XNOR U9446 ( .A(b[2955]), .B(n5349), .Z(c[2955]) );
  XOR U9447 ( .A(n5350), .B(n5351), .Z(n5347) );
  ANDN U9448 ( .B(n5352), .A(n5353), .Z(n5350) );
  XNOR U9449 ( .A(b[2954]), .B(n5351), .Z(n5352) );
  XNOR U9450 ( .A(b[2954]), .B(n5353), .Z(c[2954]) );
  XOR U9451 ( .A(n5354), .B(n5355), .Z(n5351) );
  ANDN U9452 ( .B(n5356), .A(n5357), .Z(n5354) );
  XNOR U9453 ( .A(b[2953]), .B(n5355), .Z(n5356) );
  XNOR U9454 ( .A(b[2953]), .B(n5357), .Z(c[2953]) );
  XOR U9455 ( .A(n5358), .B(n5359), .Z(n5355) );
  ANDN U9456 ( .B(n5360), .A(n5361), .Z(n5358) );
  XNOR U9457 ( .A(b[2952]), .B(n5359), .Z(n5360) );
  XNOR U9458 ( .A(b[2952]), .B(n5361), .Z(c[2952]) );
  XOR U9459 ( .A(n5362), .B(n5363), .Z(n5359) );
  ANDN U9460 ( .B(n5364), .A(n5365), .Z(n5362) );
  XNOR U9461 ( .A(b[2951]), .B(n5363), .Z(n5364) );
  XNOR U9462 ( .A(b[2951]), .B(n5365), .Z(c[2951]) );
  XOR U9463 ( .A(n5366), .B(n5367), .Z(n5363) );
  ANDN U9464 ( .B(n5368), .A(n5369), .Z(n5366) );
  XNOR U9465 ( .A(b[2950]), .B(n5367), .Z(n5368) );
  XNOR U9466 ( .A(b[2950]), .B(n5369), .Z(c[2950]) );
  XOR U9467 ( .A(n5370), .B(n5371), .Z(n5367) );
  ANDN U9468 ( .B(n5372), .A(n5373), .Z(n5370) );
  XNOR U9469 ( .A(b[2949]), .B(n5371), .Z(n5372) );
  XNOR U9470 ( .A(b[294]), .B(n5374), .Z(c[294]) );
  XNOR U9471 ( .A(b[2949]), .B(n5373), .Z(c[2949]) );
  XOR U9472 ( .A(n5375), .B(n5376), .Z(n5371) );
  ANDN U9473 ( .B(n5377), .A(n5378), .Z(n5375) );
  XNOR U9474 ( .A(b[2948]), .B(n5376), .Z(n5377) );
  XNOR U9475 ( .A(b[2948]), .B(n5378), .Z(c[2948]) );
  XOR U9476 ( .A(n5379), .B(n5380), .Z(n5376) );
  ANDN U9477 ( .B(n5381), .A(n5382), .Z(n5379) );
  XNOR U9478 ( .A(b[2947]), .B(n5380), .Z(n5381) );
  XNOR U9479 ( .A(b[2947]), .B(n5382), .Z(c[2947]) );
  XOR U9480 ( .A(n5383), .B(n5384), .Z(n5380) );
  ANDN U9481 ( .B(n5385), .A(n5386), .Z(n5383) );
  XNOR U9482 ( .A(b[2946]), .B(n5384), .Z(n5385) );
  XNOR U9483 ( .A(b[2946]), .B(n5386), .Z(c[2946]) );
  XOR U9484 ( .A(n5387), .B(n5388), .Z(n5384) );
  ANDN U9485 ( .B(n5389), .A(n5390), .Z(n5387) );
  XNOR U9486 ( .A(b[2945]), .B(n5388), .Z(n5389) );
  XNOR U9487 ( .A(b[2945]), .B(n5390), .Z(c[2945]) );
  XOR U9488 ( .A(n5391), .B(n5392), .Z(n5388) );
  ANDN U9489 ( .B(n5393), .A(n5394), .Z(n5391) );
  XNOR U9490 ( .A(b[2944]), .B(n5392), .Z(n5393) );
  XNOR U9491 ( .A(b[2944]), .B(n5394), .Z(c[2944]) );
  XOR U9492 ( .A(n5395), .B(n5396), .Z(n5392) );
  ANDN U9493 ( .B(n5397), .A(n5398), .Z(n5395) );
  XNOR U9494 ( .A(b[2943]), .B(n5396), .Z(n5397) );
  XNOR U9495 ( .A(b[2943]), .B(n5398), .Z(c[2943]) );
  XOR U9496 ( .A(n5399), .B(n5400), .Z(n5396) );
  ANDN U9497 ( .B(n5401), .A(n5402), .Z(n5399) );
  XNOR U9498 ( .A(b[2942]), .B(n5400), .Z(n5401) );
  XNOR U9499 ( .A(b[2942]), .B(n5402), .Z(c[2942]) );
  XOR U9500 ( .A(n5403), .B(n5404), .Z(n5400) );
  ANDN U9501 ( .B(n5405), .A(n5406), .Z(n5403) );
  XNOR U9502 ( .A(b[2941]), .B(n5404), .Z(n5405) );
  XNOR U9503 ( .A(b[2941]), .B(n5406), .Z(c[2941]) );
  XOR U9504 ( .A(n5407), .B(n5408), .Z(n5404) );
  ANDN U9505 ( .B(n5409), .A(n5410), .Z(n5407) );
  XNOR U9506 ( .A(b[2940]), .B(n5408), .Z(n5409) );
  XNOR U9507 ( .A(b[2940]), .B(n5410), .Z(c[2940]) );
  XOR U9508 ( .A(n5411), .B(n5412), .Z(n5408) );
  ANDN U9509 ( .B(n5413), .A(n5414), .Z(n5411) );
  XNOR U9510 ( .A(b[2939]), .B(n5412), .Z(n5413) );
  XNOR U9511 ( .A(b[293]), .B(n5415), .Z(c[293]) );
  XNOR U9512 ( .A(b[2939]), .B(n5414), .Z(c[2939]) );
  XOR U9513 ( .A(n5416), .B(n5417), .Z(n5412) );
  ANDN U9514 ( .B(n5418), .A(n5419), .Z(n5416) );
  XNOR U9515 ( .A(b[2938]), .B(n5417), .Z(n5418) );
  XNOR U9516 ( .A(b[2938]), .B(n5419), .Z(c[2938]) );
  XOR U9517 ( .A(n5420), .B(n5421), .Z(n5417) );
  ANDN U9518 ( .B(n5422), .A(n5423), .Z(n5420) );
  XNOR U9519 ( .A(b[2937]), .B(n5421), .Z(n5422) );
  XNOR U9520 ( .A(b[2937]), .B(n5423), .Z(c[2937]) );
  XOR U9521 ( .A(n5424), .B(n5425), .Z(n5421) );
  ANDN U9522 ( .B(n5426), .A(n5427), .Z(n5424) );
  XNOR U9523 ( .A(b[2936]), .B(n5425), .Z(n5426) );
  XNOR U9524 ( .A(b[2936]), .B(n5427), .Z(c[2936]) );
  XOR U9525 ( .A(n5428), .B(n5429), .Z(n5425) );
  ANDN U9526 ( .B(n5430), .A(n5431), .Z(n5428) );
  XNOR U9527 ( .A(b[2935]), .B(n5429), .Z(n5430) );
  XNOR U9528 ( .A(b[2935]), .B(n5431), .Z(c[2935]) );
  XOR U9529 ( .A(n5432), .B(n5433), .Z(n5429) );
  ANDN U9530 ( .B(n5434), .A(n5435), .Z(n5432) );
  XNOR U9531 ( .A(b[2934]), .B(n5433), .Z(n5434) );
  XNOR U9532 ( .A(b[2934]), .B(n5435), .Z(c[2934]) );
  XOR U9533 ( .A(n5436), .B(n5437), .Z(n5433) );
  ANDN U9534 ( .B(n5438), .A(n5439), .Z(n5436) );
  XNOR U9535 ( .A(b[2933]), .B(n5437), .Z(n5438) );
  XNOR U9536 ( .A(b[2933]), .B(n5439), .Z(c[2933]) );
  XOR U9537 ( .A(n5440), .B(n5441), .Z(n5437) );
  ANDN U9538 ( .B(n5442), .A(n5443), .Z(n5440) );
  XNOR U9539 ( .A(b[2932]), .B(n5441), .Z(n5442) );
  XNOR U9540 ( .A(b[2932]), .B(n5443), .Z(c[2932]) );
  XOR U9541 ( .A(n5444), .B(n5445), .Z(n5441) );
  ANDN U9542 ( .B(n5446), .A(n5447), .Z(n5444) );
  XNOR U9543 ( .A(b[2931]), .B(n5445), .Z(n5446) );
  XNOR U9544 ( .A(b[2931]), .B(n5447), .Z(c[2931]) );
  XOR U9545 ( .A(n5448), .B(n5449), .Z(n5445) );
  ANDN U9546 ( .B(n5450), .A(n5451), .Z(n5448) );
  XNOR U9547 ( .A(b[2930]), .B(n5449), .Z(n5450) );
  XNOR U9548 ( .A(b[2930]), .B(n5451), .Z(c[2930]) );
  XOR U9549 ( .A(n5452), .B(n5453), .Z(n5449) );
  ANDN U9550 ( .B(n5454), .A(n5455), .Z(n5452) );
  XNOR U9551 ( .A(b[2929]), .B(n5453), .Z(n5454) );
  XNOR U9552 ( .A(b[292]), .B(n5456), .Z(c[292]) );
  XNOR U9553 ( .A(b[2929]), .B(n5455), .Z(c[2929]) );
  XOR U9554 ( .A(n5457), .B(n5458), .Z(n5453) );
  ANDN U9555 ( .B(n5459), .A(n5460), .Z(n5457) );
  XNOR U9556 ( .A(b[2928]), .B(n5458), .Z(n5459) );
  XNOR U9557 ( .A(b[2928]), .B(n5460), .Z(c[2928]) );
  XOR U9558 ( .A(n5461), .B(n5462), .Z(n5458) );
  ANDN U9559 ( .B(n5463), .A(n5464), .Z(n5461) );
  XNOR U9560 ( .A(b[2927]), .B(n5462), .Z(n5463) );
  XNOR U9561 ( .A(b[2927]), .B(n5464), .Z(c[2927]) );
  XOR U9562 ( .A(n5465), .B(n5466), .Z(n5462) );
  ANDN U9563 ( .B(n5467), .A(n5468), .Z(n5465) );
  XNOR U9564 ( .A(b[2926]), .B(n5466), .Z(n5467) );
  XNOR U9565 ( .A(b[2926]), .B(n5468), .Z(c[2926]) );
  XOR U9566 ( .A(n5469), .B(n5470), .Z(n5466) );
  ANDN U9567 ( .B(n5471), .A(n5472), .Z(n5469) );
  XNOR U9568 ( .A(b[2925]), .B(n5470), .Z(n5471) );
  XNOR U9569 ( .A(b[2925]), .B(n5472), .Z(c[2925]) );
  XOR U9570 ( .A(n5473), .B(n5474), .Z(n5470) );
  ANDN U9571 ( .B(n5475), .A(n5476), .Z(n5473) );
  XNOR U9572 ( .A(b[2924]), .B(n5474), .Z(n5475) );
  XNOR U9573 ( .A(b[2924]), .B(n5476), .Z(c[2924]) );
  XOR U9574 ( .A(n5477), .B(n5478), .Z(n5474) );
  ANDN U9575 ( .B(n5479), .A(n5480), .Z(n5477) );
  XNOR U9576 ( .A(b[2923]), .B(n5478), .Z(n5479) );
  XNOR U9577 ( .A(b[2923]), .B(n5480), .Z(c[2923]) );
  XOR U9578 ( .A(n5481), .B(n5482), .Z(n5478) );
  ANDN U9579 ( .B(n5483), .A(n5484), .Z(n5481) );
  XNOR U9580 ( .A(b[2922]), .B(n5482), .Z(n5483) );
  XNOR U9581 ( .A(b[2922]), .B(n5484), .Z(c[2922]) );
  XOR U9582 ( .A(n5485), .B(n5486), .Z(n5482) );
  ANDN U9583 ( .B(n5487), .A(n5488), .Z(n5485) );
  XNOR U9584 ( .A(b[2921]), .B(n5486), .Z(n5487) );
  XNOR U9585 ( .A(b[2921]), .B(n5488), .Z(c[2921]) );
  XOR U9586 ( .A(n5489), .B(n5490), .Z(n5486) );
  ANDN U9587 ( .B(n5491), .A(n5492), .Z(n5489) );
  XNOR U9588 ( .A(b[2920]), .B(n5490), .Z(n5491) );
  XNOR U9589 ( .A(b[2920]), .B(n5492), .Z(c[2920]) );
  XOR U9590 ( .A(n5493), .B(n5494), .Z(n5490) );
  ANDN U9591 ( .B(n5495), .A(n5496), .Z(n5493) );
  XNOR U9592 ( .A(b[2919]), .B(n5494), .Z(n5495) );
  XNOR U9593 ( .A(b[291]), .B(n5497), .Z(c[291]) );
  XNOR U9594 ( .A(b[2919]), .B(n5496), .Z(c[2919]) );
  XOR U9595 ( .A(n5498), .B(n5499), .Z(n5494) );
  ANDN U9596 ( .B(n5500), .A(n5501), .Z(n5498) );
  XNOR U9597 ( .A(b[2918]), .B(n5499), .Z(n5500) );
  XNOR U9598 ( .A(b[2918]), .B(n5501), .Z(c[2918]) );
  XOR U9599 ( .A(n5502), .B(n5503), .Z(n5499) );
  ANDN U9600 ( .B(n5504), .A(n5505), .Z(n5502) );
  XNOR U9601 ( .A(b[2917]), .B(n5503), .Z(n5504) );
  XNOR U9602 ( .A(b[2917]), .B(n5505), .Z(c[2917]) );
  XOR U9603 ( .A(n5506), .B(n5507), .Z(n5503) );
  ANDN U9604 ( .B(n5508), .A(n5509), .Z(n5506) );
  XNOR U9605 ( .A(b[2916]), .B(n5507), .Z(n5508) );
  XNOR U9606 ( .A(b[2916]), .B(n5509), .Z(c[2916]) );
  XOR U9607 ( .A(n5510), .B(n5511), .Z(n5507) );
  ANDN U9608 ( .B(n5512), .A(n5513), .Z(n5510) );
  XNOR U9609 ( .A(b[2915]), .B(n5511), .Z(n5512) );
  XNOR U9610 ( .A(b[2915]), .B(n5513), .Z(c[2915]) );
  XOR U9611 ( .A(n5514), .B(n5515), .Z(n5511) );
  ANDN U9612 ( .B(n5516), .A(n5517), .Z(n5514) );
  XNOR U9613 ( .A(b[2914]), .B(n5515), .Z(n5516) );
  XNOR U9614 ( .A(b[2914]), .B(n5517), .Z(c[2914]) );
  XOR U9615 ( .A(n5518), .B(n5519), .Z(n5515) );
  ANDN U9616 ( .B(n5520), .A(n5521), .Z(n5518) );
  XNOR U9617 ( .A(b[2913]), .B(n5519), .Z(n5520) );
  XNOR U9618 ( .A(b[2913]), .B(n5521), .Z(c[2913]) );
  XOR U9619 ( .A(n5522), .B(n5523), .Z(n5519) );
  ANDN U9620 ( .B(n5524), .A(n5525), .Z(n5522) );
  XNOR U9621 ( .A(b[2912]), .B(n5523), .Z(n5524) );
  XNOR U9622 ( .A(b[2912]), .B(n5525), .Z(c[2912]) );
  XOR U9623 ( .A(n5526), .B(n5527), .Z(n5523) );
  ANDN U9624 ( .B(n5528), .A(n5529), .Z(n5526) );
  XNOR U9625 ( .A(b[2911]), .B(n5527), .Z(n5528) );
  XNOR U9626 ( .A(b[2911]), .B(n5529), .Z(c[2911]) );
  XOR U9627 ( .A(n5530), .B(n5531), .Z(n5527) );
  ANDN U9628 ( .B(n5532), .A(n5533), .Z(n5530) );
  XNOR U9629 ( .A(b[2910]), .B(n5531), .Z(n5532) );
  XNOR U9630 ( .A(b[2910]), .B(n5533), .Z(c[2910]) );
  XOR U9631 ( .A(n5534), .B(n5535), .Z(n5531) );
  ANDN U9632 ( .B(n5536), .A(n5537), .Z(n5534) );
  XNOR U9633 ( .A(b[2909]), .B(n5535), .Z(n5536) );
  XNOR U9634 ( .A(b[290]), .B(n5538), .Z(c[290]) );
  XNOR U9635 ( .A(b[2909]), .B(n5537), .Z(c[2909]) );
  XOR U9636 ( .A(n5539), .B(n5540), .Z(n5535) );
  ANDN U9637 ( .B(n5541), .A(n5542), .Z(n5539) );
  XNOR U9638 ( .A(b[2908]), .B(n5540), .Z(n5541) );
  XNOR U9639 ( .A(b[2908]), .B(n5542), .Z(c[2908]) );
  XOR U9640 ( .A(n5543), .B(n5544), .Z(n5540) );
  ANDN U9641 ( .B(n5545), .A(n5546), .Z(n5543) );
  XNOR U9642 ( .A(b[2907]), .B(n5544), .Z(n5545) );
  XNOR U9643 ( .A(b[2907]), .B(n5546), .Z(c[2907]) );
  XOR U9644 ( .A(n5547), .B(n5548), .Z(n5544) );
  ANDN U9645 ( .B(n5549), .A(n5550), .Z(n5547) );
  XNOR U9646 ( .A(b[2906]), .B(n5548), .Z(n5549) );
  XNOR U9647 ( .A(b[2906]), .B(n5550), .Z(c[2906]) );
  XOR U9648 ( .A(n5551), .B(n5552), .Z(n5548) );
  ANDN U9649 ( .B(n5553), .A(n5554), .Z(n5551) );
  XNOR U9650 ( .A(b[2905]), .B(n5552), .Z(n5553) );
  XNOR U9651 ( .A(b[2905]), .B(n5554), .Z(c[2905]) );
  XOR U9652 ( .A(n5555), .B(n5556), .Z(n5552) );
  ANDN U9653 ( .B(n5557), .A(n5558), .Z(n5555) );
  XNOR U9654 ( .A(b[2904]), .B(n5556), .Z(n5557) );
  XNOR U9655 ( .A(b[2904]), .B(n5558), .Z(c[2904]) );
  XOR U9656 ( .A(n5559), .B(n5560), .Z(n5556) );
  ANDN U9657 ( .B(n5561), .A(n5562), .Z(n5559) );
  XNOR U9658 ( .A(b[2903]), .B(n5560), .Z(n5561) );
  XNOR U9659 ( .A(b[2903]), .B(n5562), .Z(c[2903]) );
  XOR U9660 ( .A(n5563), .B(n5564), .Z(n5560) );
  ANDN U9661 ( .B(n5565), .A(n5566), .Z(n5563) );
  XNOR U9662 ( .A(b[2902]), .B(n5564), .Z(n5565) );
  XNOR U9663 ( .A(b[2902]), .B(n5566), .Z(c[2902]) );
  XOR U9664 ( .A(n5567), .B(n5568), .Z(n5564) );
  ANDN U9665 ( .B(n5569), .A(n5570), .Z(n5567) );
  XNOR U9666 ( .A(b[2901]), .B(n5568), .Z(n5569) );
  XNOR U9667 ( .A(b[2901]), .B(n5570), .Z(c[2901]) );
  XOR U9668 ( .A(n5571), .B(n5572), .Z(n5568) );
  ANDN U9669 ( .B(n5573), .A(n5574), .Z(n5571) );
  XNOR U9670 ( .A(b[2900]), .B(n5572), .Z(n5573) );
  XNOR U9671 ( .A(b[2900]), .B(n5574), .Z(c[2900]) );
  XOR U9672 ( .A(n5575), .B(n5576), .Z(n5572) );
  ANDN U9673 ( .B(n5577), .A(n5578), .Z(n5575) );
  XNOR U9674 ( .A(b[2899]), .B(n5576), .Z(n5577) );
  XNOR U9675 ( .A(b[28]), .B(n5579), .Z(c[28]) );
  XNOR U9676 ( .A(b[289]), .B(n5580), .Z(c[289]) );
  XNOR U9677 ( .A(b[2899]), .B(n5578), .Z(c[2899]) );
  XOR U9678 ( .A(n5581), .B(n5582), .Z(n5576) );
  ANDN U9679 ( .B(n5583), .A(n5584), .Z(n5581) );
  XNOR U9680 ( .A(b[2898]), .B(n5582), .Z(n5583) );
  XNOR U9681 ( .A(b[2898]), .B(n5584), .Z(c[2898]) );
  XOR U9682 ( .A(n5585), .B(n5586), .Z(n5582) );
  ANDN U9683 ( .B(n5587), .A(n5588), .Z(n5585) );
  XNOR U9684 ( .A(b[2897]), .B(n5586), .Z(n5587) );
  XNOR U9685 ( .A(b[2897]), .B(n5588), .Z(c[2897]) );
  XOR U9686 ( .A(n5589), .B(n5590), .Z(n5586) );
  ANDN U9687 ( .B(n5591), .A(n5592), .Z(n5589) );
  XNOR U9688 ( .A(b[2896]), .B(n5590), .Z(n5591) );
  XNOR U9689 ( .A(b[2896]), .B(n5592), .Z(c[2896]) );
  XOR U9690 ( .A(n5593), .B(n5594), .Z(n5590) );
  ANDN U9691 ( .B(n5595), .A(n5596), .Z(n5593) );
  XNOR U9692 ( .A(b[2895]), .B(n5594), .Z(n5595) );
  XNOR U9693 ( .A(b[2895]), .B(n5596), .Z(c[2895]) );
  XOR U9694 ( .A(n5597), .B(n5598), .Z(n5594) );
  ANDN U9695 ( .B(n5599), .A(n5600), .Z(n5597) );
  XNOR U9696 ( .A(b[2894]), .B(n5598), .Z(n5599) );
  XNOR U9697 ( .A(b[2894]), .B(n5600), .Z(c[2894]) );
  XOR U9698 ( .A(n5601), .B(n5602), .Z(n5598) );
  ANDN U9699 ( .B(n5603), .A(n5604), .Z(n5601) );
  XNOR U9700 ( .A(b[2893]), .B(n5602), .Z(n5603) );
  XNOR U9701 ( .A(b[2893]), .B(n5604), .Z(c[2893]) );
  XOR U9702 ( .A(n5605), .B(n5606), .Z(n5602) );
  ANDN U9703 ( .B(n5607), .A(n5608), .Z(n5605) );
  XNOR U9704 ( .A(b[2892]), .B(n5606), .Z(n5607) );
  XNOR U9705 ( .A(b[2892]), .B(n5608), .Z(c[2892]) );
  XOR U9706 ( .A(n5609), .B(n5610), .Z(n5606) );
  ANDN U9707 ( .B(n5611), .A(n5612), .Z(n5609) );
  XNOR U9708 ( .A(b[2891]), .B(n5610), .Z(n5611) );
  XNOR U9709 ( .A(b[2891]), .B(n5612), .Z(c[2891]) );
  XOR U9710 ( .A(n5613), .B(n5614), .Z(n5610) );
  ANDN U9711 ( .B(n5615), .A(n5616), .Z(n5613) );
  XNOR U9712 ( .A(b[2890]), .B(n5614), .Z(n5615) );
  XNOR U9713 ( .A(b[2890]), .B(n5616), .Z(c[2890]) );
  XOR U9714 ( .A(n5617), .B(n5618), .Z(n5614) );
  ANDN U9715 ( .B(n5619), .A(n5620), .Z(n5617) );
  XNOR U9716 ( .A(b[2889]), .B(n5618), .Z(n5619) );
  XNOR U9717 ( .A(b[288]), .B(n5621), .Z(c[288]) );
  XNOR U9718 ( .A(b[2889]), .B(n5620), .Z(c[2889]) );
  XOR U9719 ( .A(n5622), .B(n5623), .Z(n5618) );
  ANDN U9720 ( .B(n5624), .A(n5625), .Z(n5622) );
  XNOR U9721 ( .A(b[2888]), .B(n5623), .Z(n5624) );
  XNOR U9722 ( .A(b[2888]), .B(n5625), .Z(c[2888]) );
  XOR U9723 ( .A(n5626), .B(n5627), .Z(n5623) );
  ANDN U9724 ( .B(n5628), .A(n5629), .Z(n5626) );
  XNOR U9725 ( .A(b[2887]), .B(n5627), .Z(n5628) );
  XNOR U9726 ( .A(b[2887]), .B(n5629), .Z(c[2887]) );
  XOR U9727 ( .A(n5630), .B(n5631), .Z(n5627) );
  ANDN U9728 ( .B(n5632), .A(n5633), .Z(n5630) );
  XNOR U9729 ( .A(b[2886]), .B(n5631), .Z(n5632) );
  XNOR U9730 ( .A(b[2886]), .B(n5633), .Z(c[2886]) );
  XOR U9731 ( .A(n5634), .B(n5635), .Z(n5631) );
  ANDN U9732 ( .B(n5636), .A(n5637), .Z(n5634) );
  XNOR U9733 ( .A(b[2885]), .B(n5635), .Z(n5636) );
  XNOR U9734 ( .A(b[2885]), .B(n5637), .Z(c[2885]) );
  XOR U9735 ( .A(n5638), .B(n5639), .Z(n5635) );
  ANDN U9736 ( .B(n5640), .A(n5641), .Z(n5638) );
  XNOR U9737 ( .A(b[2884]), .B(n5639), .Z(n5640) );
  XNOR U9738 ( .A(b[2884]), .B(n5641), .Z(c[2884]) );
  XOR U9739 ( .A(n5642), .B(n5643), .Z(n5639) );
  ANDN U9740 ( .B(n5644), .A(n5645), .Z(n5642) );
  XNOR U9741 ( .A(b[2883]), .B(n5643), .Z(n5644) );
  XNOR U9742 ( .A(b[2883]), .B(n5645), .Z(c[2883]) );
  XOR U9743 ( .A(n5646), .B(n5647), .Z(n5643) );
  ANDN U9744 ( .B(n5648), .A(n5649), .Z(n5646) );
  XNOR U9745 ( .A(b[2882]), .B(n5647), .Z(n5648) );
  XNOR U9746 ( .A(b[2882]), .B(n5649), .Z(c[2882]) );
  XOR U9747 ( .A(n5650), .B(n5651), .Z(n5647) );
  ANDN U9748 ( .B(n5652), .A(n5653), .Z(n5650) );
  XNOR U9749 ( .A(b[2881]), .B(n5651), .Z(n5652) );
  XNOR U9750 ( .A(b[2881]), .B(n5653), .Z(c[2881]) );
  XOR U9751 ( .A(n5654), .B(n5655), .Z(n5651) );
  ANDN U9752 ( .B(n5656), .A(n5657), .Z(n5654) );
  XNOR U9753 ( .A(b[2880]), .B(n5655), .Z(n5656) );
  XNOR U9754 ( .A(b[2880]), .B(n5657), .Z(c[2880]) );
  XOR U9755 ( .A(n5658), .B(n5659), .Z(n5655) );
  ANDN U9756 ( .B(n5660), .A(n5661), .Z(n5658) );
  XNOR U9757 ( .A(b[2879]), .B(n5659), .Z(n5660) );
  XNOR U9758 ( .A(b[287]), .B(n5662), .Z(c[287]) );
  XNOR U9759 ( .A(b[2879]), .B(n5661), .Z(c[2879]) );
  XOR U9760 ( .A(n5663), .B(n5664), .Z(n5659) );
  ANDN U9761 ( .B(n5665), .A(n5666), .Z(n5663) );
  XNOR U9762 ( .A(b[2878]), .B(n5664), .Z(n5665) );
  XNOR U9763 ( .A(b[2878]), .B(n5666), .Z(c[2878]) );
  XOR U9764 ( .A(n5667), .B(n5668), .Z(n5664) );
  ANDN U9765 ( .B(n5669), .A(n5670), .Z(n5667) );
  XNOR U9766 ( .A(b[2877]), .B(n5668), .Z(n5669) );
  XNOR U9767 ( .A(b[2877]), .B(n5670), .Z(c[2877]) );
  XOR U9768 ( .A(n5671), .B(n5672), .Z(n5668) );
  ANDN U9769 ( .B(n5673), .A(n5674), .Z(n5671) );
  XNOR U9770 ( .A(b[2876]), .B(n5672), .Z(n5673) );
  XNOR U9771 ( .A(b[2876]), .B(n5674), .Z(c[2876]) );
  XOR U9772 ( .A(n5675), .B(n5676), .Z(n5672) );
  ANDN U9773 ( .B(n5677), .A(n5678), .Z(n5675) );
  XNOR U9774 ( .A(b[2875]), .B(n5676), .Z(n5677) );
  XNOR U9775 ( .A(b[2875]), .B(n5678), .Z(c[2875]) );
  XOR U9776 ( .A(n5679), .B(n5680), .Z(n5676) );
  ANDN U9777 ( .B(n5681), .A(n5682), .Z(n5679) );
  XNOR U9778 ( .A(b[2874]), .B(n5680), .Z(n5681) );
  XNOR U9779 ( .A(b[2874]), .B(n5682), .Z(c[2874]) );
  XOR U9780 ( .A(n5683), .B(n5684), .Z(n5680) );
  ANDN U9781 ( .B(n5685), .A(n5686), .Z(n5683) );
  XNOR U9782 ( .A(b[2873]), .B(n5684), .Z(n5685) );
  XNOR U9783 ( .A(b[2873]), .B(n5686), .Z(c[2873]) );
  XOR U9784 ( .A(n5687), .B(n5688), .Z(n5684) );
  ANDN U9785 ( .B(n5689), .A(n5690), .Z(n5687) );
  XNOR U9786 ( .A(b[2872]), .B(n5688), .Z(n5689) );
  XNOR U9787 ( .A(b[2872]), .B(n5690), .Z(c[2872]) );
  XOR U9788 ( .A(n5691), .B(n5692), .Z(n5688) );
  ANDN U9789 ( .B(n5693), .A(n5694), .Z(n5691) );
  XNOR U9790 ( .A(b[2871]), .B(n5692), .Z(n5693) );
  XNOR U9791 ( .A(b[2871]), .B(n5694), .Z(c[2871]) );
  XOR U9792 ( .A(n5695), .B(n5696), .Z(n5692) );
  ANDN U9793 ( .B(n5697), .A(n5698), .Z(n5695) );
  XNOR U9794 ( .A(b[2870]), .B(n5696), .Z(n5697) );
  XNOR U9795 ( .A(b[2870]), .B(n5698), .Z(c[2870]) );
  XOR U9796 ( .A(n5699), .B(n5700), .Z(n5696) );
  ANDN U9797 ( .B(n5701), .A(n5702), .Z(n5699) );
  XNOR U9798 ( .A(b[2869]), .B(n5700), .Z(n5701) );
  XNOR U9799 ( .A(b[286]), .B(n5703), .Z(c[286]) );
  XNOR U9800 ( .A(b[2869]), .B(n5702), .Z(c[2869]) );
  XOR U9801 ( .A(n5704), .B(n5705), .Z(n5700) );
  ANDN U9802 ( .B(n5706), .A(n5707), .Z(n5704) );
  XNOR U9803 ( .A(b[2868]), .B(n5705), .Z(n5706) );
  XNOR U9804 ( .A(b[2868]), .B(n5707), .Z(c[2868]) );
  XOR U9805 ( .A(n5708), .B(n5709), .Z(n5705) );
  ANDN U9806 ( .B(n5710), .A(n5711), .Z(n5708) );
  XNOR U9807 ( .A(b[2867]), .B(n5709), .Z(n5710) );
  XNOR U9808 ( .A(b[2867]), .B(n5711), .Z(c[2867]) );
  XOR U9809 ( .A(n5712), .B(n5713), .Z(n5709) );
  ANDN U9810 ( .B(n5714), .A(n5715), .Z(n5712) );
  XNOR U9811 ( .A(b[2866]), .B(n5713), .Z(n5714) );
  XNOR U9812 ( .A(b[2866]), .B(n5715), .Z(c[2866]) );
  XOR U9813 ( .A(n5716), .B(n5717), .Z(n5713) );
  ANDN U9814 ( .B(n5718), .A(n5719), .Z(n5716) );
  XNOR U9815 ( .A(b[2865]), .B(n5717), .Z(n5718) );
  XNOR U9816 ( .A(b[2865]), .B(n5719), .Z(c[2865]) );
  XOR U9817 ( .A(n5720), .B(n5721), .Z(n5717) );
  ANDN U9818 ( .B(n5722), .A(n5723), .Z(n5720) );
  XNOR U9819 ( .A(b[2864]), .B(n5721), .Z(n5722) );
  XNOR U9820 ( .A(b[2864]), .B(n5723), .Z(c[2864]) );
  XOR U9821 ( .A(n5724), .B(n5725), .Z(n5721) );
  ANDN U9822 ( .B(n5726), .A(n5727), .Z(n5724) );
  XNOR U9823 ( .A(b[2863]), .B(n5725), .Z(n5726) );
  XNOR U9824 ( .A(b[2863]), .B(n5727), .Z(c[2863]) );
  XOR U9825 ( .A(n5728), .B(n5729), .Z(n5725) );
  ANDN U9826 ( .B(n5730), .A(n5731), .Z(n5728) );
  XNOR U9827 ( .A(b[2862]), .B(n5729), .Z(n5730) );
  XNOR U9828 ( .A(b[2862]), .B(n5731), .Z(c[2862]) );
  XOR U9829 ( .A(n5732), .B(n5733), .Z(n5729) );
  ANDN U9830 ( .B(n5734), .A(n5735), .Z(n5732) );
  XNOR U9831 ( .A(b[2861]), .B(n5733), .Z(n5734) );
  XNOR U9832 ( .A(b[2861]), .B(n5735), .Z(c[2861]) );
  XOR U9833 ( .A(n5736), .B(n5737), .Z(n5733) );
  ANDN U9834 ( .B(n5738), .A(n5739), .Z(n5736) );
  XNOR U9835 ( .A(b[2860]), .B(n5737), .Z(n5738) );
  XNOR U9836 ( .A(b[2860]), .B(n5739), .Z(c[2860]) );
  XOR U9837 ( .A(n5740), .B(n5741), .Z(n5737) );
  ANDN U9838 ( .B(n5742), .A(n5743), .Z(n5740) );
  XNOR U9839 ( .A(b[2859]), .B(n5741), .Z(n5742) );
  XNOR U9840 ( .A(b[285]), .B(n5744), .Z(c[285]) );
  XNOR U9841 ( .A(b[2859]), .B(n5743), .Z(c[2859]) );
  XOR U9842 ( .A(n5745), .B(n5746), .Z(n5741) );
  ANDN U9843 ( .B(n5747), .A(n5748), .Z(n5745) );
  XNOR U9844 ( .A(b[2858]), .B(n5746), .Z(n5747) );
  XNOR U9845 ( .A(b[2858]), .B(n5748), .Z(c[2858]) );
  XOR U9846 ( .A(n5749), .B(n5750), .Z(n5746) );
  ANDN U9847 ( .B(n5751), .A(n5752), .Z(n5749) );
  XNOR U9848 ( .A(b[2857]), .B(n5750), .Z(n5751) );
  XNOR U9849 ( .A(b[2857]), .B(n5752), .Z(c[2857]) );
  XOR U9850 ( .A(n5753), .B(n5754), .Z(n5750) );
  ANDN U9851 ( .B(n5755), .A(n5756), .Z(n5753) );
  XNOR U9852 ( .A(b[2856]), .B(n5754), .Z(n5755) );
  XNOR U9853 ( .A(b[2856]), .B(n5756), .Z(c[2856]) );
  XOR U9854 ( .A(n5757), .B(n5758), .Z(n5754) );
  ANDN U9855 ( .B(n5759), .A(n5760), .Z(n5757) );
  XNOR U9856 ( .A(b[2855]), .B(n5758), .Z(n5759) );
  XNOR U9857 ( .A(b[2855]), .B(n5760), .Z(c[2855]) );
  XOR U9858 ( .A(n5761), .B(n5762), .Z(n5758) );
  ANDN U9859 ( .B(n5763), .A(n5764), .Z(n5761) );
  XNOR U9860 ( .A(b[2854]), .B(n5762), .Z(n5763) );
  XNOR U9861 ( .A(b[2854]), .B(n5764), .Z(c[2854]) );
  XOR U9862 ( .A(n5765), .B(n5766), .Z(n5762) );
  ANDN U9863 ( .B(n5767), .A(n5768), .Z(n5765) );
  XNOR U9864 ( .A(b[2853]), .B(n5766), .Z(n5767) );
  XNOR U9865 ( .A(b[2853]), .B(n5768), .Z(c[2853]) );
  XOR U9866 ( .A(n5769), .B(n5770), .Z(n5766) );
  ANDN U9867 ( .B(n5771), .A(n5772), .Z(n5769) );
  XNOR U9868 ( .A(b[2852]), .B(n5770), .Z(n5771) );
  XNOR U9869 ( .A(b[2852]), .B(n5772), .Z(c[2852]) );
  XOR U9870 ( .A(n5773), .B(n5774), .Z(n5770) );
  ANDN U9871 ( .B(n5775), .A(n5776), .Z(n5773) );
  XNOR U9872 ( .A(b[2851]), .B(n5774), .Z(n5775) );
  XNOR U9873 ( .A(b[2851]), .B(n5776), .Z(c[2851]) );
  XOR U9874 ( .A(n5777), .B(n5778), .Z(n5774) );
  ANDN U9875 ( .B(n5779), .A(n5780), .Z(n5777) );
  XNOR U9876 ( .A(b[2850]), .B(n5778), .Z(n5779) );
  XNOR U9877 ( .A(b[2850]), .B(n5780), .Z(c[2850]) );
  XOR U9878 ( .A(n5781), .B(n5782), .Z(n5778) );
  ANDN U9879 ( .B(n5783), .A(n5784), .Z(n5781) );
  XNOR U9880 ( .A(b[2849]), .B(n5782), .Z(n5783) );
  XNOR U9881 ( .A(b[284]), .B(n5785), .Z(c[284]) );
  XNOR U9882 ( .A(b[2849]), .B(n5784), .Z(c[2849]) );
  XOR U9883 ( .A(n5786), .B(n5787), .Z(n5782) );
  ANDN U9884 ( .B(n5788), .A(n5789), .Z(n5786) );
  XNOR U9885 ( .A(b[2848]), .B(n5787), .Z(n5788) );
  XNOR U9886 ( .A(b[2848]), .B(n5789), .Z(c[2848]) );
  XOR U9887 ( .A(n5790), .B(n5791), .Z(n5787) );
  ANDN U9888 ( .B(n5792), .A(n5793), .Z(n5790) );
  XNOR U9889 ( .A(b[2847]), .B(n5791), .Z(n5792) );
  XNOR U9890 ( .A(b[2847]), .B(n5793), .Z(c[2847]) );
  XOR U9891 ( .A(n5794), .B(n5795), .Z(n5791) );
  ANDN U9892 ( .B(n5796), .A(n5797), .Z(n5794) );
  XNOR U9893 ( .A(b[2846]), .B(n5795), .Z(n5796) );
  XNOR U9894 ( .A(b[2846]), .B(n5797), .Z(c[2846]) );
  XOR U9895 ( .A(n5798), .B(n5799), .Z(n5795) );
  ANDN U9896 ( .B(n5800), .A(n5801), .Z(n5798) );
  XNOR U9897 ( .A(b[2845]), .B(n5799), .Z(n5800) );
  XNOR U9898 ( .A(b[2845]), .B(n5801), .Z(c[2845]) );
  XOR U9899 ( .A(n5802), .B(n5803), .Z(n5799) );
  ANDN U9900 ( .B(n5804), .A(n5805), .Z(n5802) );
  XNOR U9901 ( .A(b[2844]), .B(n5803), .Z(n5804) );
  XNOR U9902 ( .A(b[2844]), .B(n5805), .Z(c[2844]) );
  XOR U9903 ( .A(n5806), .B(n5807), .Z(n5803) );
  ANDN U9904 ( .B(n5808), .A(n5809), .Z(n5806) );
  XNOR U9905 ( .A(b[2843]), .B(n5807), .Z(n5808) );
  XNOR U9906 ( .A(b[2843]), .B(n5809), .Z(c[2843]) );
  XOR U9907 ( .A(n5810), .B(n5811), .Z(n5807) );
  ANDN U9908 ( .B(n5812), .A(n5813), .Z(n5810) );
  XNOR U9909 ( .A(b[2842]), .B(n5811), .Z(n5812) );
  XNOR U9910 ( .A(b[2842]), .B(n5813), .Z(c[2842]) );
  XOR U9911 ( .A(n5814), .B(n5815), .Z(n5811) );
  ANDN U9912 ( .B(n5816), .A(n5817), .Z(n5814) );
  XNOR U9913 ( .A(b[2841]), .B(n5815), .Z(n5816) );
  XNOR U9914 ( .A(b[2841]), .B(n5817), .Z(c[2841]) );
  XOR U9915 ( .A(n5818), .B(n5819), .Z(n5815) );
  ANDN U9916 ( .B(n5820), .A(n5821), .Z(n5818) );
  XNOR U9917 ( .A(b[2840]), .B(n5819), .Z(n5820) );
  XNOR U9918 ( .A(b[2840]), .B(n5821), .Z(c[2840]) );
  XOR U9919 ( .A(n5822), .B(n5823), .Z(n5819) );
  ANDN U9920 ( .B(n5824), .A(n5825), .Z(n5822) );
  XNOR U9921 ( .A(b[2839]), .B(n5823), .Z(n5824) );
  XNOR U9922 ( .A(b[283]), .B(n5826), .Z(c[283]) );
  XNOR U9923 ( .A(b[2839]), .B(n5825), .Z(c[2839]) );
  XOR U9924 ( .A(n5827), .B(n5828), .Z(n5823) );
  ANDN U9925 ( .B(n5829), .A(n5830), .Z(n5827) );
  XNOR U9926 ( .A(b[2838]), .B(n5828), .Z(n5829) );
  XNOR U9927 ( .A(b[2838]), .B(n5830), .Z(c[2838]) );
  XOR U9928 ( .A(n5831), .B(n5832), .Z(n5828) );
  ANDN U9929 ( .B(n5833), .A(n5834), .Z(n5831) );
  XNOR U9930 ( .A(b[2837]), .B(n5832), .Z(n5833) );
  XNOR U9931 ( .A(b[2837]), .B(n5834), .Z(c[2837]) );
  XOR U9932 ( .A(n5835), .B(n5836), .Z(n5832) );
  ANDN U9933 ( .B(n5837), .A(n5838), .Z(n5835) );
  XNOR U9934 ( .A(b[2836]), .B(n5836), .Z(n5837) );
  XNOR U9935 ( .A(b[2836]), .B(n5838), .Z(c[2836]) );
  XOR U9936 ( .A(n5839), .B(n5840), .Z(n5836) );
  ANDN U9937 ( .B(n5841), .A(n5842), .Z(n5839) );
  XNOR U9938 ( .A(b[2835]), .B(n5840), .Z(n5841) );
  XNOR U9939 ( .A(b[2835]), .B(n5842), .Z(c[2835]) );
  XOR U9940 ( .A(n5843), .B(n5844), .Z(n5840) );
  ANDN U9941 ( .B(n5845), .A(n5846), .Z(n5843) );
  XNOR U9942 ( .A(b[2834]), .B(n5844), .Z(n5845) );
  XNOR U9943 ( .A(b[2834]), .B(n5846), .Z(c[2834]) );
  XOR U9944 ( .A(n5847), .B(n5848), .Z(n5844) );
  ANDN U9945 ( .B(n5849), .A(n5850), .Z(n5847) );
  XNOR U9946 ( .A(b[2833]), .B(n5848), .Z(n5849) );
  XNOR U9947 ( .A(b[2833]), .B(n5850), .Z(c[2833]) );
  XOR U9948 ( .A(n5851), .B(n5852), .Z(n5848) );
  ANDN U9949 ( .B(n5853), .A(n5854), .Z(n5851) );
  XNOR U9950 ( .A(b[2832]), .B(n5852), .Z(n5853) );
  XNOR U9951 ( .A(b[2832]), .B(n5854), .Z(c[2832]) );
  XOR U9952 ( .A(n5855), .B(n5856), .Z(n5852) );
  ANDN U9953 ( .B(n5857), .A(n5858), .Z(n5855) );
  XNOR U9954 ( .A(b[2831]), .B(n5856), .Z(n5857) );
  XNOR U9955 ( .A(b[2831]), .B(n5858), .Z(c[2831]) );
  XOR U9956 ( .A(n5859), .B(n5860), .Z(n5856) );
  ANDN U9957 ( .B(n5861), .A(n5862), .Z(n5859) );
  XNOR U9958 ( .A(b[2830]), .B(n5860), .Z(n5861) );
  XNOR U9959 ( .A(b[2830]), .B(n5862), .Z(c[2830]) );
  XOR U9960 ( .A(n5863), .B(n5864), .Z(n5860) );
  ANDN U9961 ( .B(n5865), .A(n5866), .Z(n5863) );
  XNOR U9962 ( .A(b[2829]), .B(n5864), .Z(n5865) );
  XNOR U9963 ( .A(b[282]), .B(n5867), .Z(c[282]) );
  XNOR U9964 ( .A(b[2829]), .B(n5866), .Z(c[2829]) );
  XOR U9965 ( .A(n5868), .B(n5869), .Z(n5864) );
  ANDN U9966 ( .B(n5870), .A(n5871), .Z(n5868) );
  XNOR U9967 ( .A(b[2828]), .B(n5869), .Z(n5870) );
  XNOR U9968 ( .A(b[2828]), .B(n5871), .Z(c[2828]) );
  XOR U9969 ( .A(n5872), .B(n5873), .Z(n5869) );
  ANDN U9970 ( .B(n5874), .A(n5875), .Z(n5872) );
  XNOR U9971 ( .A(b[2827]), .B(n5873), .Z(n5874) );
  XNOR U9972 ( .A(b[2827]), .B(n5875), .Z(c[2827]) );
  XOR U9973 ( .A(n5876), .B(n5877), .Z(n5873) );
  ANDN U9974 ( .B(n5878), .A(n5879), .Z(n5876) );
  XNOR U9975 ( .A(b[2826]), .B(n5877), .Z(n5878) );
  XNOR U9976 ( .A(b[2826]), .B(n5879), .Z(c[2826]) );
  XOR U9977 ( .A(n5880), .B(n5881), .Z(n5877) );
  ANDN U9978 ( .B(n5882), .A(n5883), .Z(n5880) );
  XNOR U9979 ( .A(b[2825]), .B(n5881), .Z(n5882) );
  XNOR U9980 ( .A(b[2825]), .B(n5883), .Z(c[2825]) );
  XOR U9981 ( .A(n5884), .B(n5885), .Z(n5881) );
  ANDN U9982 ( .B(n5886), .A(n5887), .Z(n5884) );
  XNOR U9983 ( .A(b[2824]), .B(n5885), .Z(n5886) );
  XNOR U9984 ( .A(b[2824]), .B(n5887), .Z(c[2824]) );
  XOR U9985 ( .A(n5888), .B(n5889), .Z(n5885) );
  ANDN U9986 ( .B(n5890), .A(n5891), .Z(n5888) );
  XNOR U9987 ( .A(b[2823]), .B(n5889), .Z(n5890) );
  XNOR U9988 ( .A(b[2823]), .B(n5891), .Z(c[2823]) );
  XOR U9989 ( .A(n5892), .B(n5893), .Z(n5889) );
  ANDN U9990 ( .B(n5894), .A(n5895), .Z(n5892) );
  XNOR U9991 ( .A(b[2822]), .B(n5893), .Z(n5894) );
  XNOR U9992 ( .A(b[2822]), .B(n5895), .Z(c[2822]) );
  XOR U9993 ( .A(n5896), .B(n5897), .Z(n5893) );
  ANDN U9994 ( .B(n5898), .A(n5899), .Z(n5896) );
  XNOR U9995 ( .A(b[2821]), .B(n5897), .Z(n5898) );
  XNOR U9996 ( .A(b[2821]), .B(n5899), .Z(c[2821]) );
  XOR U9997 ( .A(n5900), .B(n5901), .Z(n5897) );
  ANDN U9998 ( .B(n5902), .A(n5903), .Z(n5900) );
  XNOR U9999 ( .A(b[2820]), .B(n5901), .Z(n5902) );
  XNOR U10000 ( .A(b[2820]), .B(n5903), .Z(c[2820]) );
  XOR U10001 ( .A(n5904), .B(n5905), .Z(n5901) );
  ANDN U10002 ( .B(n5906), .A(n5907), .Z(n5904) );
  XNOR U10003 ( .A(b[2819]), .B(n5905), .Z(n5906) );
  XNOR U10004 ( .A(b[281]), .B(n5908), .Z(c[281]) );
  XNOR U10005 ( .A(b[2819]), .B(n5907), .Z(c[2819]) );
  XOR U10006 ( .A(n5909), .B(n5910), .Z(n5905) );
  ANDN U10007 ( .B(n5911), .A(n5912), .Z(n5909) );
  XNOR U10008 ( .A(b[2818]), .B(n5910), .Z(n5911) );
  XNOR U10009 ( .A(b[2818]), .B(n5912), .Z(c[2818]) );
  XOR U10010 ( .A(n5913), .B(n5914), .Z(n5910) );
  ANDN U10011 ( .B(n5915), .A(n5916), .Z(n5913) );
  XNOR U10012 ( .A(b[2817]), .B(n5914), .Z(n5915) );
  XNOR U10013 ( .A(b[2817]), .B(n5916), .Z(c[2817]) );
  XOR U10014 ( .A(n5917), .B(n5918), .Z(n5914) );
  ANDN U10015 ( .B(n5919), .A(n5920), .Z(n5917) );
  XNOR U10016 ( .A(b[2816]), .B(n5918), .Z(n5919) );
  XNOR U10017 ( .A(b[2816]), .B(n5920), .Z(c[2816]) );
  XOR U10018 ( .A(n5921), .B(n5922), .Z(n5918) );
  ANDN U10019 ( .B(n5923), .A(n5924), .Z(n5921) );
  XNOR U10020 ( .A(b[2815]), .B(n5922), .Z(n5923) );
  XNOR U10021 ( .A(b[2815]), .B(n5924), .Z(c[2815]) );
  XOR U10022 ( .A(n5925), .B(n5926), .Z(n5922) );
  ANDN U10023 ( .B(n5927), .A(n5928), .Z(n5925) );
  XNOR U10024 ( .A(b[2814]), .B(n5926), .Z(n5927) );
  XNOR U10025 ( .A(b[2814]), .B(n5928), .Z(c[2814]) );
  XOR U10026 ( .A(n5929), .B(n5930), .Z(n5926) );
  ANDN U10027 ( .B(n5931), .A(n5932), .Z(n5929) );
  XNOR U10028 ( .A(b[2813]), .B(n5930), .Z(n5931) );
  XNOR U10029 ( .A(b[2813]), .B(n5932), .Z(c[2813]) );
  XOR U10030 ( .A(n5933), .B(n5934), .Z(n5930) );
  ANDN U10031 ( .B(n5935), .A(n5936), .Z(n5933) );
  XNOR U10032 ( .A(b[2812]), .B(n5934), .Z(n5935) );
  XNOR U10033 ( .A(b[2812]), .B(n5936), .Z(c[2812]) );
  XOR U10034 ( .A(n5937), .B(n5938), .Z(n5934) );
  ANDN U10035 ( .B(n5939), .A(n5940), .Z(n5937) );
  XNOR U10036 ( .A(b[2811]), .B(n5938), .Z(n5939) );
  XNOR U10037 ( .A(b[2811]), .B(n5940), .Z(c[2811]) );
  XOR U10038 ( .A(n5941), .B(n5942), .Z(n5938) );
  ANDN U10039 ( .B(n5943), .A(n5944), .Z(n5941) );
  XNOR U10040 ( .A(b[2810]), .B(n5942), .Z(n5943) );
  XNOR U10041 ( .A(b[2810]), .B(n5944), .Z(c[2810]) );
  XOR U10042 ( .A(n5945), .B(n5946), .Z(n5942) );
  ANDN U10043 ( .B(n5947), .A(n5948), .Z(n5945) );
  XNOR U10044 ( .A(b[2809]), .B(n5946), .Z(n5947) );
  XNOR U10045 ( .A(b[280]), .B(n5949), .Z(c[280]) );
  XNOR U10046 ( .A(b[2809]), .B(n5948), .Z(c[2809]) );
  XOR U10047 ( .A(n5950), .B(n5951), .Z(n5946) );
  ANDN U10048 ( .B(n5952), .A(n5953), .Z(n5950) );
  XNOR U10049 ( .A(b[2808]), .B(n5951), .Z(n5952) );
  XNOR U10050 ( .A(b[2808]), .B(n5953), .Z(c[2808]) );
  XOR U10051 ( .A(n5954), .B(n5955), .Z(n5951) );
  ANDN U10052 ( .B(n5956), .A(n5957), .Z(n5954) );
  XNOR U10053 ( .A(b[2807]), .B(n5955), .Z(n5956) );
  XNOR U10054 ( .A(b[2807]), .B(n5957), .Z(c[2807]) );
  XOR U10055 ( .A(n5958), .B(n5959), .Z(n5955) );
  ANDN U10056 ( .B(n5960), .A(n5961), .Z(n5958) );
  XNOR U10057 ( .A(b[2806]), .B(n5959), .Z(n5960) );
  XNOR U10058 ( .A(b[2806]), .B(n5961), .Z(c[2806]) );
  XOR U10059 ( .A(n5962), .B(n5963), .Z(n5959) );
  ANDN U10060 ( .B(n5964), .A(n5965), .Z(n5962) );
  XNOR U10061 ( .A(b[2805]), .B(n5963), .Z(n5964) );
  XNOR U10062 ( .A(b[2805]), .B(n5965), .Z(c[2805]) );
  XOR U10063 ( .A(n5966), .B(n5967), .Z(n5963) );
  ANDN U10064 ( .B(n5968), .A(n5969), .Z(n5966) );
  XNOR U10065 ( .A(b[2804]), .B(n5967), .Z(n5968) );
  XNOR U10066 ( .A(b[2804]), .B(n5969), .Z(c[2804]) );
  XOR U10067 ( .A(n5970), .B(n5971), .Z(n5967) );
  ANDN U10068 ( .B(n5972), .A(n5973), .Z(n5970) );
  XNOR U10069 ( .A(b[2803]), .B(n5971), .Z(n5972) );
  XNOR U10070 ( .A(b[2803]), .B(n5973), .Z(c[2803]) );
  XOR U10071 ( .A(n5974), .B(n5975), .Z(n5971) );
  ANDN U10072 ( .B(n5976), .A(n5977), .Z(n5974) );
  XNOR U10073 ( .A(b[2802]), .B(n5975), .Z(n5976) );
  XNOR U10074 ( .A(b[2802]), .B(n5977), .Z(c[2802]) );
  XOR U10075 ( .A(n5978), .B(n5979), .Z(n5975) );
  ANDN U10076 ( .B(n5980), .A(n5981), .Z(n5978) );
  XNOR U10077 ( .A(b[2801]), .B(n5979), .Z(n5980) );
  XNOR U10078 ( .A(b[2801]), .B(n5981), .Z(c[2801]) );
  XOR U10079 ( .A(n5982), .B(n5983), .Z(n5979) );
  ANDN U10080 ( .B(n5984), .A(n5985), .Z(n5982) );
  XNOR U10081 ( .A(b[2800]), .B(n5983), .Z(n5984) );
  XNOR U10082 ( .A(b[2800]), .B(n5985), .Z(c[2800]) );
  XOR U10083 ( .A(n5986), .B(n5987), .Z(n5983) );
  ANDN U10084 ( .B(n5988), .A(n5989), .Z(n5986) );
  XNOR U10085 ( .A(b[2799]), .B(n5987), .Z(n5988) );
  XNOR U10086 ( .A(b[27]), .B(n5990), .Z(c[27]) );
  XNOR U10087 ( .A(b[279]), .B(n5991), .Z(c[279]) );
  XNOR U10088 ( .A(b[2799]), .B(n5989), .Z(c[2799]) );
  XOR U10089 ( .A(n5992), .B(n5993), .Z(n5987) );
  ANDN U10090 ( .B(n5994), .A(n5995), .Z(n5992) );
  XNOR U10091 ( .A(b[2798]), .B(n5993), .Z(n5994) );
  XNOR U10092 ( .A(b[2798]), .B(n5995), .Z(c[2798]) );
  XOR U10093 ( .A(n5996), .B(n5997), .Z(n5993) );
  ANDN U10094 ( .B(n5998), .A(n5999), .Z(n5996) );
  XNOR U10095 ( .A(b[2797]), .B(n5997), .Z(n5998) );
  XNOR U10096 ( .A(b[2797]), .B(n5999), .Z(c[2797]) );
  XOR U10097 ( .A(n6000), .B(n6001), .Z(n5997) );
  ANDN U10098 ( .B(n6002), .A(n6003), .Z(n6000) );
  XNOR U10099 ( .A(b[2796]), .B(n6001), .Z(n6002) );
  XNOR U10100 ( .A(b[2796]), .B(n6003), .Z(c[2796]) );
  XOR U10101 ( .A(n6004), .B(n6005), .Z(n6001) );
  ANDN U10102 ( .B(n6006), .A(n6007), .Z(n6004) );
  XNOR U10103 ( .A(b[2795]), .B(n6005), .Z(n6006) );
  XNOR U10104 ( .A(b[2795]), .B(n6007), .Z(c[2795]) );
  XOR U10105 ( .A(n6008), .B(n6009), .Z(n6005) );
  ANDN U10106 ( .B(n6010), .A(n6011), .Z(n6008) );
  XNOR U10107 ( .A(b[2794]), .B(n6009), .Z(n6010) );
  XNOR U10108 ( .A(b[2794]), .B(n6011), .Z(c[2794]) );
  XOR U10109 ( .A(n6012), .B(n6013), .Z(n6009) );
  ANDN U10110 ( .B(n6014), .A(n6015), .Z(n6012) );
  XNOR U10111 ( .A(b[2793]), .B(n6013), .Z(n6014) );
  XNOR U10112 ( .A(b[2793]), .B(n6015), .Z(c[2793]) );
  XOR U10113 ( .A(n6016), .B(n6017), .Z(n6013) );
  ANDN U10114 ( .B(n6018), .A(n6019), .Z(n6016) );
  XNOR U10115 ( .A(b[2792]), .B(n6017), .Z(n6018) );
  XNOR U10116 ( .A(b[2792]), .B(n6019), .Z(c[2792]) );
  XOR U10117 ( .A(n6020), .B(n6021), .Z(n6017) );
  ANDN U10118 ( .B(n6022), .A(n6023), .Z(n6020) );
  XNOR U10119 ( .A(b[2791]), .B(n6021), .Z(n6022) );
  XNOR U10120 ( .A(b[2791]), .B(n6023), .Z(c[2791]) );
  XOR U10121 ( .A(n6024), .B(n6025), .Z(n6021) );
  ANDN U10122 ( .B(n6026), .A(n6027), .Z(n6024) );
  XNOR U10123 ( .A(b[2790]), .B(n6025), .Z(n6026) );
  XNOR U10124 ( .A(b[2790]), .B(n6027), .Z(c[2790]) );
  XOR U10125 ( .A(n6028), .B(n6029), .Z(n6025) );
  ANDN U10126 ( .B(n6030), .A(n6031), .Z(n6028) );
  XNOR U10127 ( .A(b[2789]), .B(n6029), .Z(n6030) );
  XNOR U10128 ( .A(b[278]), .B(n6032), .Z(c[278]) );
  XNOR U10129 ( .A(b[2789]), .B(n6031), .Z(c[2789]) );
  XOR U10130 ( .A(n6033), .B(n6034), .Z(n6029) );
  ANDN U10131 ( .B(n6035), .A(n6036), .Z(n6033) );
  XNOR U10132 ( .A(b[2788]), .B(n6034), .Z(n6035) );
  XNOR U10133 ( .A(b[2788]), .B(n6036), .Z(c[2788]) );
  XOR U10134 ( .A(n6037), .B(n6038), .Z(n6034) );
  ANDN U10135 ( .B(n6039), .A(n6040), .Z(n6037) );
  XNOR U10136 ( .A(b[2787]), .B(n6038), .Z(n6039) );
  XNOR U10137 ( .A(b[2787]), .B(n6040), .Z(c[2787]) );
  XOR U10138 ( .A(n6041), .B(n6042), .Z(n6038) );
  ANDN U10139 ( .B(n6043), .A(n6044), .Z(n6041) );
  XNOR U10140 ( .A(b[2786]), .B(n6042), .Z(n6043) );
  XNOR U10141 ( .A(b[2786]), .B(n6044), .Z(c[2786]) );
  XOR U10142 ( .A(n6045), .B(n6046), .Z(n6042) );
  ANDN U10143 ( .B(n6047), .A(n6048), .Z(n6045) );
  XNOR U10144 ( .A(b[2785]), .B(n6046), .Z(n6047) );
  XNOR U10145 ( .A(b[2785]), .B(n6048), .Z(c[2785]) );
  XOR U10146 ( .A(n6049), .B(n6050), .Z(n6046) );
  ANDN U10147 ( .B(n6051), .A(n6052), .Z(n6049) );
  XNOR U10148 ( .A(b[2784]), .B(n6050), .Z(n6051) );
  XNOR U10149 ( .A(b[2784]), .B(n6052), .Z(c[2784]) );
  XOR U10150 ( .A(n6053), .B(n6054), .Z(n6050) );
  ANDN U10151 ( .B(n6055), .A(n6056), .Z(n6053) );
  XNOR U10152 ( .A(b[2783]), .B(n6054), .Z(n6055) );
  XNOR U10153 ( .A(b[2783]), .B(n6056), .Z(c[2783]) );
  XOR U10154 ( .A(n6057), .B(n6058), .Z(n6054) );
  ANDN U10155 ( .B(n6059), .A(n6060), .Z(n6057) );
  XNOR U10156 ( .A(b[2782]), .B(n6058), .Z(n6059) );
  XNOR U10157 ( .A(b[2782]), .B(n6060), .Z(c[2782]) );
  XOR U10158 ( .A(n6061), .B(n6062), .Z(n6058) );
  ANDN U10159 ( .B(n6063), .A(n6064), .Z(n6061) );
  XNOR U10160 ( .A(b[2781]), .B(n6062), .Z(n6063) );
  XNOR U10161 ( .A(b[2781]), .B(n6064), .Z(c[2781]) );
  XOR U10162 ( .A(n6065), .B(n6066), .Z(n6062) );
  ANDN U10163 ( .B(n6067), .A(n6068), .Z(n6065) );
  XNOR U10164 ( .A(b[2780]), .B(n6066), .Z(n6067) );
  XNOR U10165 ( .A(b[2780]), .B(n6068), .Z(c[2780]) );
  XOR U10166 ( .A(n6069), .B(n6070), .Z(n6066) );
  ANDN U10167 ( .B(n6071), .A(n6072), .Z(n6069) );
  XNOR U10168 ( .A(b[2779]), .B(n6070), .Z(n6071) );
  XNOR U10169 ( .A(b[277]), .B(n6073), .Z(c[277]) );
  XNOR U10170 ( .A(b[2779]), .B(n6072), .Z(c[2779]) );
  XOR U10171 ( .A(n6074), .B(n6075), .Z(n6070) );
  ANDN U10172 ( .B(n6076), .A(n6077), .Z(n6074) );
  XNOR U10173 ( .A(b[2778]), .B(n6075), .Z(n6076) );
  XNOR U10174 ( .A(b[2778]), .B(n6077), .Z(c[2778]) );
  XOR U10175 ( .A(n6078), .B(n6079), .Z(n6075) );
  ANDN U10176 ( .B(n6080), .A(n6081), .Z(n6078) );
  XNOR U10177 ( .A(b[2777]), .B(n6079), .Z(n6080) );
  XNOR U10178 ( .A(b[2777]), .B(n6081), .Z(c[2777]) );
  XOR U10179 ( .A(n6082), .B(n6083), .Z(n6079) );
  ANDN U10180 ( .B(n6084), .A(n6085), .Z(n6082) );
  XNOR U10181 ( .A(b[2776]), .B(n6083), .Z(n6084) );
  XNOR U10182 ( .A(b[2776]), .B(n6085), .Z(c[2776]) );
  XOR U10183 ( .A(n6086), .B(n6087), .Z(n6083) );
  ANDN U10184 ( .B(n6088), .A(n6089), .Z(n6086) );
  XNOR U10185 ( .A(b[2775]), .B(n6087), .Z(n6088) );
  XNOR U10186 ( .A(b[2775]), .B(n6089), .Z(c[2775]) );
  XOR U10187 ( .A(n6090), .B(n6091), .Z(n6087) );
  ANDN U10188 ( .B(n6092), .A(n6093), .Z(n6090) );
  XNOR U10189 ( .A(b[2774]), .B(n6091), .Z(n6092) );
  XNOR U10190 ( .A(b[2774]), .B(n6093), .Z(c[2774]) );
  XOR U10191 ( .A(n6094), .B(n6095), .Z(n6091) );
  ANDN U10192 ( .B(n6096), .A(n6097), .Z(n6094) );
  XNOR U10193 ( .A(b[2773]), .B(n6095), .Z(n6096) );
  XNOR U10194 ( .A(b[2773]), .B(n6097), .Z(c[2773]) );
  XOR U10195 ( .A(n6098), .B(n6099), .Z(n6095) );
  ANDN U10196 ( .B(n6100), .A(n6101), .Z(n6098) );
  XNOR U10197 ( .A(b[2772]), .B(n6099), .Z(n6100) );
  XNOR U10198 ( .A(b[2772]), .B(n6101), .Z(c[2772]) );
  XOR U10199 ( .A(n6102), .B(n6103), .Z(n6099) );
  ANDN U10200 ( .B(n6104), .A(n6105), .Z(n6102) );
  XNOR U10201 ( .A(b[2771]), .B(n6103), .Z(n6104) );
  XNOR U10202 ( .A(b[2771]), .B(n6105), .Z(c[2771]) );
  XOR U10203 ( .A(n6106), .B(n6107), .Z(n6103) );
  ANDN U10204 ( .B(n6108), .A(n6109), .Z(n6106) );
  XNOR U10205 ( .A(b[2770]), .B(n6107), .Z(n6108) );
  XNOR U10206 ( .A(b[2770]), .B(n6109), .Z(c[2770]) );
  XOR U10207 ( .A(n6110), .B(n6111), .Z(n6107) );
  ANDN U10208 ( .B(n6112), .A(n6113), .Z(n6110) );
  XNOR U10209 ( .A(b[2769]), .B(n6111), .Z(n6112) );
  XNOR U10210 ( .A(b[276]), .B(n6114), .Z(c[276]) );
  XNOR U10211 ( .A(b[2769]), .B(n6113), .Z(c[2769]) );
  XOR U10212 ( .A(n6115), .B(n6116), .Z(n6111) );
  ANDN U10213 ( .B(n6117), .A(n6118), .Z(n6115) );
  XNOR U10214 ( .A(b[2768]), .B(n6116), .Z(n6117) );
  XNOR U10215 ( .A(b[2768]), .B(n6118), .Z(c[2768]) );
  XOR U10216 ( .A(n6119), .B(n6120), .Z(n6116) );
  ANDN U10217 ( .B(n6121), .A(n6122), .Z(n6119) );
  XNOR U10218 ( .A(b[2767]), .B(n6120), .Z(n6121) );
  XNOR U10219 ( .A(b[2767]), .B(n6122), .Z(c[2767]) );
  XOR U10220 ( .A(n6123), .B(n6124), .Z(n6120) );
  ANDN U10221 ( .B(n6125), .A(n6126), .Z(n6123) );
  XNOR U10222 ( .A(b[2766]), .B(n6124), .Z(n6125) );
  XNOR U10223 ( .A(b[2766]), .B(n6126), .Z(c[2766]) );
  XOR U10224 ( .A(n6127), .B(n6128), .Z(n6124) );
  ANDN U10225 ( .B(n6129), .A(n6130), .Z(n6127) );
  XNOR U10226 ( .A(b[2765]), .B(n6128), .Z(n6129) );
  XNOR U10227 ( .A(b[2765]), .B(n6130), .Z(c[2765]) );
  XOR U10228 ( .A(n6131), .B(n6132), .Z(n6128) );
  ANDN U10229 ( .B(n6133), .A(n6134), .Z(n6131) );
  XNOR U10230 ( .A(b[2764]), .B(n6132), .Z(n6133) );
  XNOR U10231 ( .A(b[2764]), .B(n6134), .Z(c[2764]) );
  XOR U10232 ( .A(n6135), .B(n6136), .Z(n6132) );
  ANDN U10233 ( .B(n6137), .A(n6138), .Z(n6135) );
  XNOR U10234 ( .A(b[2763]), .B(n6136), .Z(n6137) );
  XNOR U10235 ( .A(b[2763]), .B(n6138), .Z(c[2763]) );
  XOR U10236 ( .A(n6139), .B(n6140), .Z(n6136) );
  ANDN U10237 ( .B(n6141), .A(n6142), .Z(n6139) );
  XNOR U10238 ( .A(b[2762]), .B(n6140), .Z(n6141) );
  XNOR U10239 ( .A(b[2762]), .B(n6142), .Z(c[2762]) );
  XOR U10240 ( .A(n6143), .B(n6144), .Z(n6140) );
  ANDN U10241 ( .B(n6145), .A(n6146), .Z(n6143) );
  XNOR U10242 ( .A(b[2761]), .B(n6144), .Z(n6145) );
  XNOR U10243 ( .A(b[2761]), .B(n6146), .Z(c[2761]) );
  XOR U10244 ( .A(n6147), .B(n6148), .Z(n6144) );
  ANDN U10245 ( .B(n6149), .A(n6150), .Z(n6147) );
  XNOR U10246 ( .A(b[2760]), .B(n6148), .Z(n6149) );
  XNOR U10247 ( .A(b[2760]), .B(n6150), .Z(c[2760]) );
  XOR U10248 ( .A(n6151), .B(n6152), .Z(n6148) );
  ANDN U10249 ( .B(n6153), .A(n6154), .Z(n6151) );
  XNOR U10250 ( .A(b[2759]), .B(n6152), .Z(n6153) );
  XNOR U10251 ( .A(b[275]), .B(n6155), .Z(c[275]) );
  XNOR U10252 ( .A(b[2759]), .B(n6154), .Z(c[2759]) );
  XOR U10253 ( .A(n6156), .B(n6157), .Z(n6152) );
  ANDN U10254 ( .B(n6158), .A(n6159), .Z(n6156) );
  XNOR U10255 ( .A(b[2758]), .B(n6157), .Z(n6158) );
  XNOR U10256 ( .A(b[2758]), .B(n6159), .Z(c[2758]) );
  XOR U10257 ( .A(n6160), .B(n6161), .Z(n6157) );
  ANDN U10258 ( .B(n6162), .A(n6163), .Z(n6160) );
  XNOR U10259 ( .A(b[2757]), .B(n6161), .Z(n6162) );
  XNOR U10260 ( .A(b[2757]), .B(n6163), .Z(c[2757]) );
  XOR U10261 ( .A(n6164), .B(n6165), .Z(n6161) );
  ANDN U10262 ( .B(n6166), .A(n6167), .Z(n6164) );
  XNOR U10263 ( .A(b[2756]), .B(n6165), .Z(n6166) );
  XNOR U10264 ( .A(b[2756]), .B(n6167), .Z(c[2756]) );
  XOR U10265 ( .A(n6168), .B(n6169), .Z(n6165) );
  ANDN U10266 ( .B(n6170), .A(n6171), .Z(n6168) );
  XNOR U10267 ( .A(b[2755]), .B(n6169), .Z(n6170) );
  XNOR U10268 ( .A(b[2755]), .B(n6171), .Z(c[2755]) );
  XOR U10269 ( .A(n6172), .B(n6173), .Z(n6169) );
  ANDN U10270 ( .B(n6174), .A(n6175), .Z(n6172) );
  XNOR U10271 ( .A(b[2754]), .B(n6173), .Z(n6174) );
  XNOR U10272 ( .A(b[2754]), .B(n6175), .Z(c[2754]) );
  XOR U10273 ( .A(n6176), .B(n6177), .Z(n6173) );
  ANDN U10274 ( .B(n6178), .A(n6179), .Z(n6176) );
  XNOR U10275 ( .A(b[2753]), .B(n6177), .Z(n6178) );
  XNOR U10276 ( .A(b[2753]), .B(n6179), .Z(c[2753]) );
  XOR U10277 ( .A(n6180), .B(n6181), .Z(n6177) );
  ANDN U10278 ( .B(n6182), .A(n6183), .Z(n6180) );
  XNOR U10279 ( .A(b[2752]), .B(n6181), .Z(n6182) );
  XNOR U10280 ( .A(b[2752]), .B(n6183), .Z(c[2752]) );
  XOR U10281 ( .A(n6184), .B(n6185), .Z(n6181) );
  ANDN U10282 ( .B(n6186), .A(n6187), .Z(n6184) );
  XNOR U10283 ( .A(b[2751]), .B(n6185), .Z(n6186) );
  XNOR U10284 ( .A(b[2751]), .B(n6187), .Z(c[2751]) );
  XOR U10285 ( .A(n6188), .B(n6189), .Z(n6185) );
  ANDN U10286 ( .B(n6190), .A(n6191), .Z(n6188) );
  XNOR U10287 ( .A(b[2750]), .B(n6189), .Z(n6190) );
  XNOR U10288 ( .A(b[2750]), .B(n6191), .Z(c[2750]) );
  XOR U10289 ( .A(n6192), .B(n6193), .Z(n6189) );
  ANDN U10290 ( .B(n6194), .A(n6195), .Z(n6192) );
  XNOR U10291 ( .A(b[2749]), .B(n6193), .Z(n6194) );
  XNOR U10292 ( .A(b[274]), .B(n6196), .Z(c[274]) );
  XNOR U10293 ( .A(b[2749]), .B(n6195), .Z(c[2749]) );
  XOR U10294 ( .A(n6197), .B(n6198), .Z(n6193) );
  ANDN U10295 ( .B(n6199), .A(n6200), .Z(n6197) );
  XNOR U10296 ( .A(b[2748]), .B(n6198), .Z(n6199) );
  XNOR U10297 ( .A(b[2748]), .B(n6200), .Z(c[2748]) );
  XOR U10298 ( .A(n6201), .B(n6202), .Z(n6198) );
  ANDN U10299 ( .B(n6203), .A(n6204), .Z(n6201) );
  XNOR U10300 ( .A(b[2747]), .B(n6202), .Z(n6203) );
  XNOR U10301 ( .A(b[2747]), .B(n6204), .Z(c[2747]) );
  XOR U10302 ( .A(n6205), .B(n6206), .Z(n6202) );
  ANDN U10303 ( .B(n6207), .A(n6208), .Z(n6205) );
  XNOR U10304 ( .A(b[2746]), .B(n6206), .Z(n6207) );
  XNOR U10305 ( .A(b[2746]), .B(n6208), .Z(c[2746]) );
  XOR U10306 ( .A(n6209), .B(n6210), .Z(n6206) );
  ANDN U10307 ( .B(n6211), .A(n6212), .Z(n6209) );
  XNOR U10308 ( .A(b[2745]), .B(n6210), .Z(n6211) );
  XNOR U10309 ( .A(b[2745]), .B(n6212), .Z(c[2745]) );
  XOR U10310 ( .A(n6213), .B(n6214), .Z(n6210) );
  ANDN U10311 ( .B(n6215), .A(n6216), .Z(n6213) );
  XNOR U10312 ( .A(b[2744]), .B(n6214), .Z(n6215) );
  XNOR U10313 ( .A(b[2744]), .B(n6216), .Z(c[2744]) );
  XOR U10314 ( .A(n6217), .B(n6218), .Z(n6214) );
  ANDN U10315 ( .B(n6219), .A(n6220), .Z(n6217) );
  XNOR U10316 ( .A(b[2743]), .B(n6218), .Z(n6219) );
  XNOR U10317 ( .A(b[2743]), .B(n6220), .Z(c[2743]) );
  XOR U10318 ( .A(n6221), .B(n6222), .Z(n6218) );
  ANDN U10319 ( .B(n6223), .A(n6224), .Z(n6221) );
  XNOR U10320 ( .A(b[2742]), .B(n6222), .Z(n6223) );
  XNOR U10321 ( .A(b[2742]), .B(n6224), .Z(c[2742]) );
  XOR U10322 ( .A(n6225), .B(n6226), .Z(n6222) );
  ANDN U10323 ( .B(n6227), .A(n6228), .Z(n6225) );
  XNOR U10324 ( .A(b[2741]), .B(n6226), .Z(n6227) );
  XNOR U10325 ( .A(b[2741]), .B(n6228), .Z(c[2741]) );
  XOR U10326 ( .A(n6229), .B(n6230), .Z(n6226) );
  ANDN U10327 ( .B(n6231), .A(n6232), .Z(n6229) );
  XNOR U10328 ( .A(b[2740]), .B(n6230), .Z(n6231) );
  XNOR U10329 ( .A(b[2740]), .B(n6232), .Z(c[2740]) );
  XOR U10330 ( .A(n6233), .B(n6234), .Z(n6230) );
  ANDN U10331 ( .B(n6235), .A(n6236), .Z(n6233) );
  XNOR U10332 ( .A(b[2739]), .B(n6234), .Z(n6235) );
  XNOR U10333 ( .A(b[273]), .B(n6237), .Z(c[273]) );
  XNOR U10334 ( .A(b[2739]), .B(n6236), .Z(c[2739]) );
  XOR U10335 ( .A(n6238), .B(n6239), .Z(n6234) );
  ANDN U10336 ( .B(n6240), .A(n6241), .Z(n6238) );
  XNOR U10337 ( .A(b[2738]), .B(n6239), .Z(n6240) );
  XNOR U10338 ( .A(b[2738]), .B(n6241), .Z(c[2738]) );
  XOR U10339 ( .A(n6242), .B(n6243), .Z(n6239) );
  ANDN U10340 ( .B(n6244), .A(n6245), .Z(n6242) );
  XNOR U10341 ( .A(b[2737]), .B(n6243), .Z(n6244) );
  XNOR U10342 ( .A(b[2737]), .B(n6245), .Z(c[2737]) );
  XOR U10343 ( .A(n6246), .B(n6247), .Z(n6243) );
  ANDN U10344 ( .B(n6248), .A(n6249), .Z(n6246) );
  XNOR U10345 ( .A(b[2736]), .B(n6247), .Z(n6248) );
  XNOR U10346 ( .A(b[2736]), .B(n6249), .Z(c[2736]) );
  XOR U10347 ( .A(n6250), .B(n6251), .Z(n6247) );
  ANDN U10348 ( .B(n6252), .A(n6253), .Z(n6250) );
  XNOR U10349 ( .A(b[2735]), .B(n6251), .Z(n6252) );
  XNOR U10350 ( .A(b[2735]), .B(n6253), .Z(c[2735]) );
  XOR U10351 ( .A(n6254), .B(n6255), .Z(n6251) );
  ANDN U10352 ( .B(n6256), .A(n6257), .Z(n6254) );
  XNOR U10353 ( .A(b[2734]), .B(n6255), .Z(n6256) );
  XNOR U10354 ( .A(b[2734]), .B(n6257), .Z(c[2734]) );
  XOR U10355 ( .A(n6258), .B(n6259), .Z(n6255) );
  ANDN U10356 ( .B(n6260), .A(n6261), .Z(n6258) );
  XNOR U10357 ( .A(b[2733]), .B(n6259), .Z(n6260) );
  XNOR U10358 ( .A(b[2733]), .B(n6261), .Z(c[2733]) );
  XOR U10359 ( .A(n6262), .B(n6263), .Z(n6259) );
  ANDN U10360 ( .B(n6264), .A(n6265), .Z(n6262) );
  XNOR U10361 ( .A(b[2732]), .B(n6263), .Z(n6264) );
  XNOR U10362 ( .A(b[2732]), .B(n6265), .Z(c[2732]) );
  XOR U10363 ( .A(n6266), .B(n6267), .Z(n6263) );
  ANDN U10364 ( .B(n6268), .A(n6269), .Z(n6266) );
  XNOR U10365 ( .A(b[2731]), .B(n6267), .Z(n6268) );
  XNOR U10366 ( .A(b[2731]), .B(n6269), .Z(c[2731]) );
  XOR U10367 ( .A(n6270), .B(n6271), .Z(n6267) );
  ANDN U10368 ( .B(n6272), .A(n6273), .Z(n6270) );
  XNOR U10369 ( .A(b[2730]), .B(n6271), .Z(n6272) );
  XNOR U10370 ( .A(b[2730]), .B(n6273), .Z(c[2730]) );
  XOR U10371 ( .A(n6274), .B(n6275), .Z(n6271) );
  ANDN U10372 ( .B(n6276), .A(n6277), .Z(n6274) );
  XNOR U10373 ( .A(b[2729]), .B(n6275), .Z(n6276) );
  XNOR U10374 ( .A(b[272]), .B(n6278), .Z(c[272]) );
  XNOR U10375 ( .A(b[2729]), .B(n6277), .Z(c[2729]) );
  XOR U10376 ( .A(n6279), .B(n6280), .Z(n6275) );
  ANDN U10377 ( .B(n6281), .A(n6282), .Z(n6279) );
  XNOR U10378 ( .A(b[2728]), .B(n6280), .Z(n6281) );
  XNOR U10379 ( .A(b[2728]), .B(n6282), .Z(c[2728]) );
  XOR U10380 ( .A(n6283), .B(n6284), .Z(n6280) );
  ANDN U10381 ( .B(n6285), .A(n6286), .Z(n6283) );
  XNOR U10382 ( .A(b[2727]), .B(n6284), .Z(n6285) );
  XNOR U10383 ( .A(b[2727]), .B(n6286), .Z(c[2727]) );
  XOR U10384 ( .A(n6287), .B(n6288), .Z(n6284) );
  ANDN U10385 ( .B(n6289), .A(n6290), .Z(n6287) );
  XNOR U10386 ( .A(b[2726]), .B(n6288), .Z(n6289) );
  XNOR U10387 ( .A(b[2726]), .B(n6290), .Z(c[2726]) );
  XOR U10388 ( .A(n6291), .B(n6292), .Z(n6288) );
  ANDN U10389 ( .B(n6293), .A(n6294), .Z(n6291) );
  XNOR U10390 ( .A(b[2725]), .B(n6292), .Z(n6293) );
  XNOR U10391 ( .A(b[2725]), .B(n6294), .Z(c[2725]) );
  XOR U10392 ( .A(n6295), .B(n6296), .Z(n6292) );
  ANDN U10393 ( .B(n6297), .A(n6298), .Z(n6295) );
  XNOR U10394 ( .A(b[2724]), .B(n6296), .Z(n6297) );
  XNOR U10395 ( .A(b[2724]), .B(n6298), .Z(c[2724]) );
  XOR U10396 ( .A(n6299), .B(n6300), .Z(n6296) );
  ANDN U10397 ( .B(n6301), .A(n6302), .Z(n6299) );
  XNOR U10398 ( .A(b[2723]), .B(n6300), .Z(n6301) );
  XNOR U10399 ( .A(b[2723]), .B(n6302), .Z(c[2723]) );
  XOR U10400 ( .A(n6303), .B(n6304), .Z(n6300) );
  ANDN U10401 ( .B(n6305), .A(n6306), .Z(n6303) );
  XNOR U10402 ( .A(b[2722]), .B(n6304), .Z(n6305) );
  XNOR U10403 ( .A(b[2722]), .B(n6306), .Z(c[2722]) );
  XOR U10404 ( .A(n6307), .B(n6308), .Z(n6304) );
  ANDN U10405 ( .B(n6309), .A(n6310), .Z(n6307) );
  XNOR U10406 ( .A(b[2721]), .B(n6308), .Z(n6309) );
  XNOR U10407 ( .A(b[2721]), .B(n6310), .Z(c[2721]) );
  XOR U10408 ( .A(n6311), .B(n6312), .Z(n6308) );
  ANDN U10409 ( .B(n6313), .A(n6314), .Z(n6311) );
  XNOR U10410 ( .A(b[2720]), .B(n6312), .Z(n6313) );
  XNOR U10411 ( .A(b[2720]), .B(n6314), .Z(c[2720]) );
  XOR U10412 ( .A(n6315), .B(n6316), .Z(n6312) );
  ANDN U10413 ( .B(n6317), .A(n6318), .Z(n6315) );
  XNOR U10414 ( .A(b[2719]), .B(n6316), .Z(n6317) );
  XNOR U10415 ( .A(b[271]), .B(n6319), .Z(c[271]) );
  XNOR U10416 ( .A(b[2719]), .B(n6318), .Z(c[2719]) );
  XOR U10417 ( .A(n6320), .B(n6321), .Z(n6316) );
  ANDN U10418 ( .B(n6322), .A(n6323), .Z(n6320) );
  XNOR U10419 ( .A(b[2718]), .B(n6321), .Z(n6322) );
  XNOR U10420 ( .A(b[2718]), .B(n6323), .Z(c[2718]) );
  XOR U10421 ( .A(n6324), .B(n6325), .Z(n6321) );
  ANDN U10422 ( .B(n6326), .A(n6327), .Z(n6324) );
  XNOR U10423 ( .A(b[2717]), .B(n6325), .Z(n6326) );
  XNOR U10424 ( .A(b[2717]), .B(n6327), .Z(c[2717]) );
  XOR U10425 ( .A(n6328), .B(n6329), .Z(n6325) );
  ANDN U10426 ( .B(n6330), .A(n6331), .Z(n6328) );
  XNOR U10427 ( .A(b[2716]), .B(n6329), .Z(n6330) );
  XNOR U10428 ( .A(b[2716]), .B(n6331), .Z(c[2716]) );
  XOR U10429 ( .A(n6332), .B(n6333), .Z(n6329) );
  ANDN U10430 ( .B(n6334), .A(n6335), .Z(n6332) );
  XNOR U10431 ( .A(b[2715]), .B(n6333), .Z(n6334) );
  XNOR U10432 ( .A(b[2715]), .B(n6335), .Z(c[2715]) );
  XOR U10433 ( .A(n6336), .B(n6337), .Z(n6333) );
  ANDN U10434 ( .B(n6338), .A(n6339), .Z(n6336) );
  XNOR U10435 ( .A(b[2714]), .B(n6337), .Z(n6338) );
  XNOR U10436 ( .A(b[2714]), .B(n6339), .Z(c[2714]) );
  XOR U10437 ( .A(n6340), .B(n6341), .Z(n6337) );
  ANDN U10438 ( .B(n6342), .A(n6343), .Z(n6340) );
  XNOR U10439 ( .A(b[2713]), .B(n6341), .Z(n6342) );
  XNOR U10440 ( .A(b[2713]), .B(n6343), .Z(c[2713]) );
  XOR U10441 ( .A(n6344), .B(n6345), .Z(n6341) );
  ANDN U10442 ( .B(n6346), .A(n6347), .Z(n6344) );
  XNOR U10443 ( .A(b[2712]), .B(n6345), .Z(n6346) );
  XNOR U10444 ( .A(b[2712]), .B(n6347), .Z(c[2712]) );
  XOR U10445 ( .A(n6348), .B(n6349), .Z(n6345) );
  ANDN U10446 ( .B(n6350), .A(n6351), .Z(n6348) );
  XNOR U10447 ( .A(b[2711]), .B(n6349), .Z(n6350) );
  XNOR U10448 ( .A(b[2711]), .B(n6351), .Z(c[2711]) );
  XOR U10449 ( .A(n6352), .B(n6353), .Z(n6349) );
  ANDN U10450 ( .B(n6354), .A(n6355), .Z(n6352) );
  XNOR U10451 ( .A(b[2710]), .B(n6353), .Z(n6354) );
  XNOR U10452 ( .A(b[2710]), .B(n6355), .Z(c[2710]) );
  XOR U10453 ( .A(n6356), .B(n6357), .Z(n6353) );
  ANDN U10454 ( .B(n6358), .A(n6359), .Z(n6356) );
  XNOR U10455 ( .A(b[2709]), .B(n6357), .Z(n6358) );
  XNOR U10456 ( .A(b[270]), .B(n6360), .Z(c[270]) );
  XNOR U10457 ( .A(b[2709]), .B(n6359), .Z(c[2709]) );
  XOR U10458 ( .A(n6361), .B(n6362), .Z(n6357) );
  ANDN U10459 ( .B(n6363), .A(n6364), .Z(n6361) );
  XNOR U10460 ( .A(b[2708]), .B(n6362), .Z(n6363) );
  XNOR U10461 ( .A(b[2708]), .B(n6364), .Z(c[2708]) );
  XOR U10462 ( .A(n6365), .B(n6366), .Z(n6362) );
  ANDN U10463 ( .B(n6367), .A(n6368), .Z(n6365) );
  XNOR U10464 ( .A(b[2707]), .B(n6366), .Z(n6367) );
  XNOR U10465 ( .A(b[2707]), .B(n6368), .Z(c[2707]) );
  XOR U10466 ( .A(n6369), .B(n6370), .Z(n6366) );
  ANDN U10467 ( .B(n6371), .A(n6372), .Z(n6369) );
  XNOR U10468 ( .A(b[2706]), .B(n6370), .Z(n6371) );
  XNOR U10469 ( .A(b[2706]), .B(n6372), .Z(c[2706]) );
  XOR U10470 ( .A(n6373), .B(n6374), .Z(n6370) );
  ANDN U10471 ( .B(n6375), .A(n6376), .Z(n6373) );
  XNOR U10472 ( .A(b[2705]), .B(n6374), .Z(n6375) );
  XNOR U10473 ( .A(b[2705]), .B(n6376), .Z(c[2705]) );
  XOR U10474 ( .A(n6377), .B(n6378), .Z(n6374) );
  ANDN U10475 ( .B(n6379), .A(n6380), .Z(n6377) );
  XNOR U10476 ( .A(b[2704]), .B(n6378), .Z(n6379) );
  XNOR U10477 ( .A(b[2704]), .B(n6380), .Z(c[2704]) );
  XOR U10478 ( .A(n6381), .B(n6382), .Z(n6378) );
  ANDN U10479 ( .B(n6383), .A(n6384), .Z(n6381) );
  XNOR U10480 ( .A(b[2703]), .B(n6382), .Z(n6383) );
  XNOR U10481 ( .A(b[2703]), .B(n6384), .Z(c[2703]) );
  XOR U10482 ( .A(n6385), .B(n6386), .Z(n6382) );
  ANDN U10483 ( .B(n6387), .A(n6388), .Z(n6385) );
  XNOR U10484 ( .A(b[2702]), .B(n6386), .Z(n6387) );
  XNOR U10485 ( .A(b[2702]), .B(n6388), .Z(c[2702]) );
  XOR U10486 ( .A(n6389), .B(n6390), .Z(n6386) );
  ANDN U10487 ( .B(n6391), .A(n6392), .Z(n6389) );
  XNOR U10488 ( .A(b[2701]), .B(n6390), .Z(n6391) );
  XNOR U10489 ( .A(b[2701]), .B(n6392), .Z(c[2701]) );
  XOR U10490 ( .A(n6393), .B(n6394), .Z(n6390) );
  ANDN U10491 ( .B(n6395), .A(n6396), .Z(n6393) );
  XNOR U10492 ( .A(b[2700]), .B(n6394), .Z(n6395) );
  XNOR U10493 ( .A(b[2700]), .B(n6396), .Z(c[2700]) );
  XOR U10494 ( .A(n6397), .B(n6398), .Z(n6394) );
  ANDN U10495 ( .B(n6399), .A(n6400), .Z(n6397) );
  XNOR U10496 ( .A(b[2699]), .B(n6398), .Z(n6399) );
  XNOR U10497 ( .A(b[26]), .B(n6401), .Z(c[26]) );
  XNOR U10498 ( .A(b[269]), .B(n6402), .Z(c[269]) );
  XNOR U10499 ( .A(b[2699]), .B(n6400), .Z(c[2699]) );
  XOR U10500 ( .A(n6403), .B(n6404), .Z(n6398) );
  ANDN U10501 ( .B(n6405), .A(n6406), .Z(n6403) );
  XNOR U10502 ( .A(b[2698]), .B(n6404), .Z(n6405) );
  XNOR U10503 ( .A(b[2698]), .B(n6406), .Z(c[2698]) );
  XOR U10504 ( .A(n6407), .B(n6408), .Z(n6404) );
  ANDN U10505 ( .B(n6409), .A(n6410), .Z(n6407) );
  XNOR U10506 ( .A(b[2697]), .B(n6408), .Z(n6409) );
  XNOR U10507 ( .A(b[2697]), .B(n6410), .Z(c[2697]) );
  XOR U10508 ( .A(n6411), .B(n6412), .Z(n6408) );
  ANDN U10509 ( .B(n6413), .A(n6414), .Z(n6411) );
  XNOR U10510 ( .A(b[2696]), .B(n6412), .Z(n6413) );
  XNOR U10511 ( .A(b[2696]), .B(n6414), .Z(c[2696]) );
  XOR U10512 ( .A(n6415), .B(n6416), .Z(n6412) );
  ANDN U10513 ( .B(n6417), .A(n6418), .Z(n6415) );
  XNOR U10514 ( .A(b[2695]), .B(n6416), .Z(n6417) );
  XNOR U10515 ( .A(b[2695]), .B(n6418), .Z(c[2695]) );
  XOR U10516 ( .A(n6419), .B(n6420), .Z(n6416) );
  ANDN U10517 ( .B(n6421), .A(n6422), .Z(n6419) );
  XNOR U10518 ( .A(b[2694]), .B(n6420), .Z(n6421) );
  XNOR U10519 ( .A(b[2694]), .B(n6422), .Z(c[2694]) );
  XOR U10520 ( .A(n6423), .B(n6424), .Z(n6420) );
  ANDN U10521 ( .B(n6425), .A(n6426), .Z(n6423) );
  XNOR U10522 ( .A(b[2693]), .B(n6424), .Z(n6425) );
  XNOR U10523 ( .A(b[2693]), .B(n6426), .Z(c[2693]) );
  XOR U10524 ( .A(n6427), .B(n6428), .Z(n6424) );
  ANDN U10525 ( .B(n6429), .A(n6430), .Z(n6427) );
  XNOR U10526 ( .A(b[2692]), .B(n6428), .Z(n6429) );
  XNOR U10527 ( .A(b[2692]), .B(n6430), .Z(c[2692]) );
  XOR U10528 ( .A(n6431), .B(n6432), .Z(n6428) );
  ANDN U10529 ( .B(n6433), .A(n6434), .Z(n6431) );
  XNOR U10530 ( .A(b[2691]), .B(n6432), .Z(n6433) );
  XNOR U10531 ( .A(b[2691]), .B(n6434), .Z(c[2691]) );
  XOR U10532 ( .A(n6435), .B(n6436), .Z(n6432) );
  ANDN U10533 ( .B(n6437), .A(n6438), .Z(n6435) );
  XNOR U10534 ( .A(b[2690]), .B(n6436), .Z(n6437) );
  XNOR U10535 ( .A(b[2690]), .B(n6438), .Z(c[2690]) );
  XOR U10536 ( .A(n6439), .B(n6440), .Z(n6436) );
  ANDN U10537 ( .B(n6441), .A(n6442), .Z(n6439) );
  XNOR U10538 ( .A(b[2689]), .B(n6440), .Z(n6441) );
  XNOR U10539 ( .A(b[268]), .B(n6443), .Z(c[268]) );
  XNOR U10540 ( .A(b[2689]), .B(n6442), .Z(c[2689]) );
  XOR U10541 ( .A(n6444), .B(n6445), .Z(n6440) );
  ANDN U10542 ( .B(n6446), .A(n6447), .Z(n6444) );
  XNOR U10543 ( .A(b[2688]), .B(n6445), .Z(n6446) );
  XNOR U10544 ( .A(b[2688]), .B(n6447), .Z(c[2688]) );
  XOR U10545 ( .A(n6448), .B(n6449), .Z(n6445) );
  ANDN U10546 ( .B(n6450), .A(n6451), .Z(n6448) );
  XNOR U10547 ( .A(b[2687]), .B(n6449), .Z(n6450) );
  XNOR U10548 ( .A(b[2687]), .B(n6451), .Z(c[2687]) );
  XOR U10549 ( .A(n6452), .B(n6453), .Z(n6449) );
  ANDN U10550 ( .B(n6454), .A(n6455), .Z(n6452) );
  XNOR U10551 ( .A(b[2686]), .B(n6453), .Z(n6454) );
  XNOR U10552 ( .A(b[2686]), .B(n6455), .Z(c[2686]) );
  XOR U10553 ( .A(n6456), .B(n6457), .Z(n6453) );
  ANDN U10554 ( .B(n6458), .A(n6459), .Z(n6456) );
  XNOR U10555 ( .A(b[2685]), .B(n6457), .Z(n6458) );
  XNOR U10556 ( .A(b[2685]), .B(n6459), .Z(c[2685]) );
  XOR U10557 ( .A(n6460), .B(n6461), .Z(n6457) );
  ANDN U10558 ( .B(n6462), .A(n6463), .Z(n6460) );
  XNOR U10559 ( .A(b[2684]), .B(n6461), .Z(n6462) );
  XNOR U10560 ( .A(b[2684]), .B(n6463), .Z(c[2684]) );
  XOR U10561 ( .A(n6464), .B(n6465), .Z(n6461) );
  ANDN U10562 ( .B(n6466), .A(n6467), .Z(n6464) );
  XNOR U10563 ( .A(b[2683]), .B(n6465), .Z(n6466) );
  XNOR U10564 ( .A(b[2683]), .B(n6467), .Z(c[2683]) );
  XOR U10565 ( .A(n6468), .B(n6469), .Z(n6465) );
  ANDN U10566 ( .B(n6470), .A(n6471), .Z(n6468) );
  XNOR U10567 ( .A(b[2682]), .B(n6469), .Z(n6470) );
  XNOR U10568 ( .A(b[2682]), .B(n6471), .Z(c[2682]) );
  XOR U10569 ( .A(n6472), .B(n6473), .Z(n6469) );
  ANDN U10570 ( .B(n6474), .A(n6475), .Z(n6472) );
  XNOR U10571 ( .A(b[2681]), .B(n6473), .Z(n6474) );
  XNOR U10572 ( .A(b[2681]), .B(n6475), .Z(c[2681]) );
  XOR U10573 ( .A(n6476), .B(n6477), .Z(n6473) );
  ANDN U10574 ( .B(n6478), .A(n6479), .Z(n6476) );
  XNOR U10575 ( .A(b[2680]), .B(n6477), .Z(n6478) );
  XNOR U10576 ( .A(b[2680]), .B(n6479), .Z(c[2680]) );
  XOR U10577 ( .A(n6480), .B(n6481), .Z(n6477) );
  ANDN U10578 ( .B(n6482), .A(n6483), .Z(n6480) );
  XNOR U10579 ( .A(b[2679]), .B(n6481), .Z(n6482) );
  XNOR U10580 ( .A(b[267]), .B(n6484), .Z(c[267]) );
  XNOR U10581 ( .A(b[2679]), .B(n6483), .Z(c[2679]) );
  XOR U10582 ( .A(n6485), .B(n6486), .Z(n6481) );
  ANDN U10583 ( .B(n6487), .A(n6488), .Z(n6485) );
  XNOR U10584 ( .A(b[2678]), .B(n6486), .Z(n6487) );
  XNOR U10585 ( .A(b[2678]), .B(n6488), .Z(c[2678]) );
  XOR U10586 ( .A(n6489), .B(n6490), .Z(n6486) );
  ANDN U10587 ( .B(n6491), .A(n6492), .Z(n6489) );
  XNOR U10588 ( .A(b[2677]), .B(n6490), .Z(n6491) );
  XNOR U10589 ( .A(b[2677]), .B(n6492), .Z(c[2677]) );
  XOR U10590 ( .A(n6493), .B(n6494), .Z(n6490) );
  ANDN U10591 ( .B(n6495), .A(n6496), .Z(n6493) );
  XNOR U10592 ( .A(b[2676]), .B(n6494), .Z(n6495) );
  XNOR U10593 ( .A(b[2676]), .B(n6496), .Z(c[2676]) );
  XOR U10594 ( .A(n6497), .B(n6498), .Z(n6494) );
  ANDN U10595 ( .B(n6499), .A(n6500), .Z(n6497) );
  XNOR U10596 ( .A(b[2675]), .B(n6498), .Z(n6499) );
  XNOR U10597 ( .A(b[2675]), .B(n6500), .Z(c[2675]) );
  XOR U10598 ( .A(n6501), .B(n6502), .Z(n6498) );
  ANDN U10599 ( .B(n6503), .A(n6504), .Z(n6501) );
  XNOR U10600 ( .A(b[2674]), .B(n6502), .Z(n6503) );
  XNOR U10601 ( .A(b[2674]), .B(n6504), .Z(c[2674]) );
  XOR U10602 ( .A(n6505), .B(n6506), .Z(n6502) );
  ANDN U10603 ( .B(n6507), .A(n6508), .Z(n6505) );
  XNOR U10604 ( .A(b[2673]), .B(n6506), .Z(n6507) );
  XNOR U10605 ( .A(b[2673]), .B(n6508), .Z(c[2673]) );
  XOR U10606 ( .A(n6509), .B(n6510), .Z(n6506) );
  ANDN U10607 ( .B(n6511), .A(n6512), .Z(n6509) );
  XNOR U10608 ( .A(b[2672]), .B(n6510), .Z(n6511) );
  XNOR U10609 ( .A(b[2672]), .B(n6512), .Z(c[2672]) );
  XOR U10610 ( .A(n6513), .B(n6514), .Z(n6510) );
  ANDN U10611 ( .B(n6515), .A(n6516), .Z(n6513) );
  XNOR U10612 ( .A(b[2671]), .B(n6514), .Z(n6515) );
  XNOR U10613 ( .A(b[2671]), .B(n6516), .Z(c[2671]) );
  XOR U10614 ( .A(n6517), .B(n6518), .Z(n6514) );
  ANDN U10615 ( .B(n6519), .A(n6520), .Z(n6517) );
  XNOR U10616 ( .A(b[2670]), .B(n6518), .Z(n6519) );
  XNOR U10617 ( .A(b[2670]), .B(n6520), .Z(c[2670]) );
  XOR U10618 ( .A(n6521), .B(n6522), .Z(n6518) );
  ANDN U10619 ( .B(n6523), .A(n6524), .Z(n6521) );
  XNOR U10620 ( .A(b[2669]), .B(n6522), .Z(n6523) );
  XNOR U10621 ( .A(b[266]), .B(n6525), .Z(c[266]) );
  XNOR U10622 ( .A(b[2669]), .B(n6524), .Z(c[2669]) );
  XOR U10623 ( .A(n6526), .B(n6527), .Z(n6522) );
  ANDN U10624 ( .B(n6528), .A(n6529), .Z(n6526) );
  XNOR U10625 ( .A(b[2668]), .B(n6527), .Z(n6528) );
  XNOR U10626 ( .A(b[2668]), .B(n6529), .Z(c[2668]) );
  XOR U10627 ( .A(n6530), .B(n6531), .Z(n6527) );
  ANDN U10628 ( .B(n6532), .A(n6533), .Z(n6530) );
  XNOR U10629 ( .A(b[2667]), .B(n6531), .Z(n6532) );
  XNOR U10630 ( .A(b[2667]), .B(n6533), .Z(c[2667]) );
  XOR U10631 ( .A(n6534), .B(n6535), .Z(n6531) );
  ANDN U10632 ( .B(n6536), .A(n6537), .Z(n6534) );
  XNOR U10633 ( .A(b[2666]), .B(n6535), .Z(n6536) );
  XNOR U10634 ( .A(b[2666]), .B(n6537), .Z(c[2666]) );
  XOR U10635 ( .A(n6538), .B(n6539), .Z(n6535) );
  ANDN U10636 ( .B(n6540), .A(n6541), .Z(n6538) );
  XNOR U10637 ( .A(b[2665]), .B(n6539), .Z(n6540) );
  XNOR U10638 ( .A(b[2665]), .B(n6541), .Z(c[2665]) );
  XOR U10639 ( .A(n6542), .B(n6543), .Z(n6539) );
  ANDN U10640 ( .B(n6544), .A(n6545), .Z(n6542) );
  XNOR U10641 ( .A(b[2664]), .B(n6543), .Z(n6544) );
  XNOR U10642 ( .A(b[2664]), .B(n6545), .Z(c[2664]) );
  XOR U10643 ( .A(n6546), .B(n6547), .Z(n6543) );
  ANDN U10644 ( .B(n6548), .A(n6549), .Z(n6546) );
  XNOR U10645 ( .A(b[2663]), .B(n6547), .Z(n6548) );
  XNOR U10646 ( .A(b[2663]), .B(n6549), .Z(c[2663]) );
  XOR U10647 ( .A(n6550), .B(n6551), .Z(n6547) );
  ANDN U10648 ( .B(n6552), .A(n6553), .Z(n6550) );
  XNOR U10649 ( .A(b[2662]), .B(n6551), .Z(n6552) );
  XNOR U10650 ( .A(b[2662]), .B(n6553), .Z(c[2662]) );
  XOR U10651 ( .A(n6554), .B(n6555), .Z(n6551) );
  ANDN U10652 ( .B(n6556), .A(n6557), .Z(n6554) );
  XNOR U10653 ( .A(b[2661]), .B(n6555), .Z(n6556) );
  XNOR U10654 ( .A(b[2661]), .B(n6557), .Z(c[2661]) );
  XOR U10655 ( .A(n6558), .B(n6559), .Z(n6555) );
  ANDN U10656 ( .B(n6560), .A(n6561), .Z(n6558) );
  XNOR U10657 ( .A(b[2660]), .B(n6559), .Z(n6560) );
  XNOR U10658 ( .A(b[2660]), .B(n6561), .Z(c[2660]) );
  XOR U10659 ( .A(n6562), .B(n6563), .Z(n6559) );
  ANDN U10660 ( .B(n6564), .A(n6565), .Z(n6562) );
  XNOR U10661 ( .A(b[2659]), .B(n6563), .Z(n6564) );
  XNOR U10662 ( .A(b[265]), .B(n6566), .Z(c[265]) );
  XNOR U10663 ( .A(b[2659]), .B(n6565), .Z(c[2659]) );
  XOR U10664 ( .A(n6567), .B(n6568), .Z(n6563) );
  ANDN U10665 ( .B(n6569), .A(n6570), .Z(n6567) );
  XNOR U10666 ( .A(b[2658]), .B(n6568), .Z(n6569) );
  XNOR U10667 ( .A(b[2658]), .B(n6570), .Z(c[2658]) );
  XOR U10668 ( .A(n6571), .B(n6572), .Z(n6568) );
  ANDN U10669 ( .B(n6573), .A(n6574), .Z(n6571) );
  XNOR U10670 ( .A(b[2657]), .B(n6572), .Z(n6573) );
  XNOR U10671 ( .A(b[2657]), .B(n6574), .Z(c[2657]) );
  XOR U10672 ( .A(n6575), .B(n6576), .Z(n6572) );
  ANDN U10673 ( .B(n6577), .A(n6578), .Z(n6575) );
  XNOR U10674 ( .A(b[2656]), .B(n6576), .Z(n6577) );
  XNOR U10675 ( .A(b[2656]), .B(n6578), .Z(c[2656]) );
  XOR U10676 ( .A(n6579), .B(n6580), .Z(n6576) );
  ANDN U10677 ( .B(n6581), .A(n6582), .Z(n6579) );
  XNOR U10678 ( .A(b[2655]), .B(n6580), .Z(n6581) );
  XNOR U10679 ( .A(b[2655]), .B(n6582), .Z(c[2655]) );
  XOR U10680 ( .A(n6583), .B(n6584), .Z(n6580) );
  ANDN U10681 ( .B(n6585), .A(n6586), .Z(n6583) );
  XNOR U10682 ( .A(b[2654]), .B(n6584), .Z(n6585) );
  XNOR U10683 ( .A(b[2654]), .B(n6586), .Z(c[2654]) );
  XOR U10684 ( .A(n6587), .B(n6588), .Z(n6584) );
  ANDN U10685 ( .B(n6589), .A(n6590), .Z(n6587) );
  XNOR U10686 ( .A(b[2653]), .B(n6588), .Z(n6589) );
  XNOR U10687 ( .A(b[2653]), .B(n6590), .Z(c[2653]) );
  XOR U10688 ( .A(n6591), .B(n6592), .Z(n6588) );
  ANDN U10689 ( .B(n6593), .A(n6594), .Z(n6591) );
  XNOR U10690 ( .A(b[2652]), .B(n6592), .Z(n6593) );
  XNOR U10691 ( .A(b[2652]), .B(n6594), .Z(c[2652]) );
  XOR U10692 ( .A(n6595), .B(n6596), .Z(n6592) );
  ANDN U10693 ( .B(n6597), .A(n6598), .Z(n6595) );
  XNOR U10694 ( .A(b[2651]), .B(n6596), .Z(n6597) );
  XNOR U10695 ( .A(b[2651]), .B(n6598), .Z(c[2651]) );
  XOR U10696 ( .A(n6599), .B(n6600), .Z(n6596) );
  ANDN U10697 ( .B(n6601), .A(n6602), .Z(n6599) );
  XNOR U10698 ( .A(b[2650]), .B(n6600), .Z(n6601) );
  XNOR U10699 ( .A(b[2650]), .B(n6602), .Z(c[2650]) );
  XOR U10700 ( .A(n6603), .B(n6604), .Z(n6600) );
  ANDN U10701 ( .B(n6605), .A(n6606), .Z(n6603) );
  XNOR U10702 ( .A(b[2649]), .B(n6604), .Z(n6605) );
  XNOR U10703 ( .A(b[264]), .B(n6607), .Z(c[264]) );
  XNOR U10704 ( .A(b[2649]), .B(n6606), .Z(c[2649]) );
  XOR U10705 ( .A(n6608), .B(n6609), .Z(n6604) );
  ANDN U10706 ( .B(n6610), .A(n6611), .Z(n6608) );
  XNOR U10707 ( .A(b[2648]), .B(n6609), .Z(n6610) );
  XNOR U10708 ( .A(b[2648]), .B(n6611), .Z(c[2648]) );
  XOR U10709 ( .A(n6612), .B(n6613), .Z(n6609) );
  ANDN U10710 ( .B(n6614), .A(n6615), .Z(n6612) );
  XNOR U10711 ( .A(b[2647]), .B(n6613), .Z(n6614) );
  XNOR U10712 ( .A(b[2647]), .B(n6615), .Z(c[2647]) );
  XOR U10713 ( .A(n6616), .B(n6617), .Z(n6613) );
  ANDN U10714 ( .B(n6618), .A(n6619), .Z(n6616) );
  XNOR U10715 ( .A(b[2646]), .B(n6617), .Z(n6618) );
  XNOR U10716 ( .A(b[2646]), .B(n6619), .Z(c[2646]) );
  XOR U10717 ( .A(n6620), .B(n6621), .Z(n6617) );
  ANDN U10718 ( .B(n6622), .A(n6623), .Z(n6620) );
  XNOR U10719 ( .A(b[2645]), .B(n6621), .Z(n6622) );
  XNOR U10720 ( .A(b[2645]), .B(n6623), .Z(c[2645]) );
  XOR U10721 ( .A(n6624), .B(n6625), .Z(n6621) );
  ANDN U10722 ( .B(n6626), .A(n6627), .Z(n6624) );
  XNOR U10723 ( .A(b[2644]), .B(n6625), .Z(n6626) );
  XNOR U10724 ( .A(b[2644]), .B(n6627), .Z(c[2644]) );
  XOR U10725 ( .A(n6628), .B(n6629), .Z(n6625) );
  ANDN U10726 ( .B(n6630), .A(n6631), .Z(n6628) );
  XNOR U10727 ( .A(b[2643]), .B(n6629), .Z(n6630) );
  XNOR U10728 ( .A(b[2643]), .B(n6631), .Z(c[2643]) );
  XOR U10729 ( .A(n6632), .B(n6633), .Z(n6629) );
  ANDN U10730 ( .B(n6634), .A(n6635), .Z(n6632) );
  XNOR U10731 ( .A(b[2642]), .B(n6633), .Z(n6634) );
  XNOR U10732 ( .A(b[2642]), .B(n6635), .Z(c[2642]) );
  XOR U10733 ( .A(n6636), .B(n6637), .Z(n6633) );
  ANDN U10734 ( .B(n6638), .A(n6639), .Z(n6636) );
  XNOR U10735 ( .A(b[2641]), .B(n6637), .Z(n6638) );
  XNOR U10736 ( .A(b[2641]), .B(n6639), .Z(c[2641]) );
  XOR U10737 ( .A(n6640), .B(n6641), .Z(n6637) );
  ANDN U10738 ( .B(n6642), .A(n6643), .Z(n6640) );
  XNOR U10739 ( .A(b[2640]), .B(n6641), .Z(n6642) );
  XNOR U10740 ( .A(b[2640]), .B(n6643), .Z(c[2640]) );
  XOR U10741 ( .A(n6644), .B(n6645), .Z(n6641) );
  ANDN U10742 ( .B(n6646), .A(n6647), .Z(n6644) );
  XNOR U10743 ( .A(b[2639]), .B(n6645), .Z(n6646) );
  XNOR U10744 ( .A(b[263]), .B(n6648), .Z(c[263]) );
  XNOR U10745 ( .A(b[2639]), .B(n6647), .Z(c[2639]) );
  XOR U10746 ( .A(n6649), .B(n6650), .Z(n6645) );
  ANDN U10747 ( .B(n6651), .A(n6652), .Z(n6649) );
  XNOR U10748 ( .A(b[2638]), .B(n6650), .Z(n6651) );
  XNOR U10749 ( .A(b[2638]), .B(n6652), .Z(c[2638]) );
  XOR U10750 ( .A(n6653), .B(n6654), .Z(n6650) );
  ANDN U10751 ( .B(n6655), .A(n6656), .Z(n6653) );
  XNOR U10752 ( .A(b[2637]), .B(n6654), .Z(n6655) );
  XNOR U10753 ( .A(b[2637]), .B(n6656), .Z(c[2637]) );
  XOR U10754 ( .A(n6657), .B(n6658), .Z(n6654) );
  ANDN U10755 ( .B(n6659), .A(n6660), .Z(n6657) );
  XNOR U10756 ( .A(b[2636]), .B(n6658), .Z(n6659) );
  XNOR U10757 ( .A(b[2636]), .B(n6660), .Z(c[2636]) );
  XOR U10758 ( .A(n6661), .B(n6662), .Z(n6658) );
  ANDN U10759 ( .B(n6663), .A(n6664), .Z(n6661) );
  XNOR U10760 ( .A(b[2635]), .B(n6662), .Z(n6663) );
  XNOR U10761 ( .A(b[2635]), .B(n6664), .Z(c[2635]) );
  XOR U10762 ( .A(n6665), .B(n6666), .Z(n6662) );
  ANDN U10763 ( .B(n6667), .A(n6668), .Z(n6665) );
  XNOR U10764 ( .A(b[2634]), .B(n6666), .Z(n6667) );
  XNOR U10765 ( .A(b[2634]), .B(n6668), .Z(c[2634]) );
  XOR U10766 ( .A(n6669), .B(n6670), .Z(n6666) );
  ANDN U10767 ( .B(n6671), .A(n6672), .Z(n6669) );
  XNOR U10768 ( .A(b[2633]), .B(n6670), .Z(n6671) );
  XNOR U10769 ( .A(b[2633]), .B(n6672), .Z(c[2633]) );
  XOR U10770 ( .A(n6673), .B(n6674), .Z(n6670) );
  ANDN U10771 ( .B(n6675), .A(n6676), .Z(n6673) );
  XNOR U10772 ( .A(b[2632]), .B(n6674), .Z(n6675) );
  XNOR U10773 ( .A(b[2632]), .B(n6676), .Z(c[2632]) );
  XOR U10774 ( .A(n6677), .B(n6678), .Z(n6674) );
  ANDN U10775 ( .B(n6679), .A(n6680), .Z(n6677) );
  XNOR U10776 ( .A(b[2631]), .B(n6678), .Z(n6679) );
  XNOR U10777 ( .A(b[2631]), .B(n6680), .Z(c[2631]) );
  XOR U10778 ( .A(n6681), .B(n6682), .Z(n6678) );
  ANDN U10779 ( .B(n6683), .A(n6684), .Z(n6681) );
  XNOR U10780 ( .A(b[2630]), .B(n6682), .Z(n6683) );
  XNOR U10781 ( .A(b[2630]), .B(n6684), .Z(c[2630]) );
  XOR U10782 ( .A(n6685), .B(n6686), .Z(n6682) );
  ANDN U10783 ( .B(n6687), .A(n6688), .Z(n6685) );
  XNOR U10784 ( .A(b[2629]), .B(n6686), .Z(n6687) );
  XNOR U10785 ( .A(b[262]), .B(n6689), .Z(c[262]) );
  XNOR U10786 ( .A(b[2629]), .B(n6688), .Z(c[2629]) );
  XOR U10787 ( .A(n6690), .B(n6691), .Z(n6686) );
  ANDN U10788 ( .B(n6692), .A(n6693), .Z(n6690) );
  XNOR U10789 ( .A(b[2628]), .B(n6691), .Z(n6692) );
  XNOR U10790 ( .A(b[2628]), .B(n6693), .Z(c[2628]) );
  XOR U10791 ( .A(n6694), .B(n6695), .Z(n6691) );
  ANDN U10792 ( .B(n6696), .A(n6697), .Z(n6694) );
  XNOR U10793 ( .A(b[2627]), .B(n6695), .Z(n6696) );
  XNOR U10794 ( .A(b[2627]), .B(n6697), .Z(c[2627]) );
  XOR U10795 ( .A(n6698), .B(n6699), .Z(n6695) );
  ANDN U10796 ( .B(n6700), .A(n6701), .Z(n6698) );
  XNOR U10797 ( .A(b[2626]), .B(n6699), .Z(n6700) );
  XNOR U10798 ( .A(b[2626]), .B(n6701), .Z(c[2626]) );
  XOR U10799 ( .A(n6702), .B(n6703), .Z(n6699) );
  ANDN U10800 ( .B(n6704), .A(n6705), .Z(n6702) );
  XNOR U10801 ( .A(b[2625]), .B(n6703), .Z(n6704) );
  XNOR U10802 ( .A(b[2625]), .B(n6705), .Z(c[2625]) );
  XOR U10803 ( .A(n6706), .B(n6707), .Z(n6703) );
  ANDN U10804 ( .B(n6708), .A(n6709), .Z(n6706) );
  XNOR U10805 ( .A(b[2624]), .B(n6707), .Z(n6708) );
  XNOR U10806 ( .A(b[2624]), .B(n6709), .Z(c[2624]) );
  XOR U10807 ( .A(n6710), .B(n6711), .Z(n6707) );
  ANDN U10808 ( .B(n6712), .A(n6713), .Z(n6710) );
  XNOR U10809 ( .A(b[2623]), .B(n6711), .Z(n6712) );
  XNOR U10810 ( .A(b[2623]), .B(n6713), .Z(c[2623]) );
  XOR U10811 ( .A(n6714), .B(n6715), .Z(n6711) );
  ANDN U10812 ( .B(n6716), .A(n6717), .Z(n6714) );
  XNOR U10813 ( .A(b[2622]), .B(n6715), .Z(n6716) );
  XNOR U10814 ( .A(b[2622]), .B(n6717), .Z(c[2622]) );
  XOR U10815 ( .A(n6718), .B(n6719), .Z(n6715) );
  ANDN U10816 ( .B(n6720), .A(n6721), .Z(n6718) );
  XNOR U10817 ( .A(b[2621]), .B(n6719), .Z(n6720) );
  XNOR U10818 ( .A(b[2621]), .B(n6721), .Z(c[2621]) );
  XOR U10819 ( .A(n6722), .B(n6723), .Z(n6719) );
  ANDN U10820 ( .B(n6724), .A(n6725), .Z(n6722) );
  XNOR U10821 ( .A(b[2620]), .B(n6723), .Z(n6724) );
  XNOR U10822 ( .A(b[2620]), .B(n6725), .Z(c[2620]) );
  XOR U10823 ( .A(n6726), .B(n6727), .Z(n6723) );
  ANDN U10824 ( .B(n6728), .A(n6729), .Z(n6726) );
  XNOR U10825 ( .A(b[2619]), .B(n6727), .Z(n6728) );
  XNOR U10826 ( .A(b[261]), .B(n6730), .Z(c[261]) );
  XNOR U10827 ( .A(b[2619]), .B(n6729), .Z(c[2619]) );
  XOR U10828 ( .A(n6731), .B(n6732), .Z(n6727) );
  ANDN U10829 ( .B(n6733), .A(n6734), .Z(n6731) );
  XNOR U10830 ( .A(b[2618]), .B(n6732), .Z(n6733) );
  XNOR U10831 ( .A(b[2618]), .B(n6734), .Z(c[2618]) );
  XOR U10832 ( .A(n6735), .B(n6736), .Z(n6732) );
  ANDN U10833 ( .B(n6737), .A(n6738), .Z(n6735) );
  XNOR U10834 ( .A(b[2617]), .B(n6736), .Z(n6737) );
  XNOR U10835 ( .A(b[2617]), .B(n6738), .Z(c[2617]) );
  XOR U10836 ( .A(n6739), .B(n6740), .Z(n6736) );
  ANDN U10837 ( .B(n6741), .A(n6742), .Z(n6739) );
  XNOR U10838 ( .A(b[2616]), .B(n6740), .Z(n6741) );
  XNOR U10839 ( .A(b[2616]), .B(n6742), .Z(c[2616]) );
  XOR U10840 ( .A(n6743), .B(n6744), .Z(n6740) );
  ANDN U10841 ( .B(n6745), .A(n6746), .Z(n6743) );
  XNOR U10842 ( .A(b[2615]), .B(n6744), .Z(n6745) );
  XNOR U10843 ( .A(b[2615]), .B(n6746), .Z(c[2615]) );
  XOR U10844 ( .A(n6747), .B(n6748), .Z(n6744) );
  ANDN U10845 ( .B(n6749), .A(n6750), .Z(n6747) );
  XNOR U10846 ( .A(b[2614]), .B(n6748), .Z(n6749) );
  XNOR U10847 ( .A(b[2614]), .B(n6750), .Z(c[2614]) );
  XOR U10848 ( .A(n6751), .B(n6752), .Z(n6748) );
  ANDN U10849 ( .B(n6753), .A(n6754), .Z(n6751) );
  XNOR U10850 ( .A(b[2613]), .B(n6752), .Z(n6753) );
  XNOR U10851 ( .A(b[2613]), .B(n6754), .Z(c[2613]) );
  XOR U10852 ( .A(n6755), .B(n6756), .Z(n6752) );
  ANDN U10853 ( .B(n6757), .A(n6758), .Z(n6755) );
  XNOR U10854 ( .A(b[2612]), .B(n6756), .Z(n6757) );
  XNOR U10855 ( .A(b[2612]), .B(n6758), .Z(c[2612]) );
  XOR U10856 ( .A(n6759), .B(n6760), .Z(n6756) );
  ANDN U10857 ( .B(n6761), .A(n6762), .Z(n6759) );
  XNOR U10858 ( .A(b[2611]), .B(n6760), .Z(n6761) );
  XNOR U10859 ( .A(b[2611]), .B(n6762), .Z(c[2611]) );
  XOR U10860 ( .A(n6763), .B(n6764), .Z(n6760) );
  ANDN U10861 ( .B(n6765), .A(n6766), .Z(n6763) );
  XNOR U10862 ( .A(b[2610]), .B(n6764), .Z(n6765) );
  XNOR U10863 ( .A(b[2610]), .B(n6766), .Z(c[2610]) );
  XOR U10864 ( .A(n6767), .B(n6768), .Z(n6764) );
  ANDN U10865 ( .B(n6769), .A(n6770), .Z(n6767) );
  XNOR U10866 ( .A(b[2609]), .B(n6768), .Z(n6769) );
  XNOR U10867 ( .A(b[260]), .B(n6771), .Z(c[260]) );
  XNOR U10868 ( .A(b[2609]), .B(n6770), .Z(c[2609]) );
  XOR U10869 ( .A(n6772), .B(n6773), .Z(n6768) );
  ANDN U10870 ( .B(n6774), .A(n6775), .Z(n6772) );
  XNOR U10871 ( .A(b[2608]), .B(n6773), .Z(n6774) );
  XNOR U10872 ( .A(b[2608]), .B(n6775), .Z(c[2608]) );
  XOR U10873 ( .A(n6776), .B(n6777), .Z(n6773) );
  ANDN U10874 ( .B(n6778), .A(n6779), .Z(n6776) );
  XNOR U10875 ( .A(b[2607]), .B(n6777), .Z(n6778) );
  XNOR U10876 ( .A(b[2607]), .B(n6779), .Z(c[2607]) );
  XOR U10877 ( .A(n6780), .B(n6781), .Z(n6777) );
  ANDN U10878 ( .B(n6782), .A(n6783), .Z(n6780) );
  XNOR U10879 ( .A(b[2606]), .B(n6781), .Z(n6782) );
  XNOR U10880 ( .A(b[2606]), .B(n6783), .Z(c[2606]) );
  XOR U10881 ( .A(n6784), .B(n6785), .Z(n6781) );
  ANDN U10882 ( .B(n6786), .A(n6787), .Z(n6784) );
  XNOR U10883 ( .A(b[2605]), .B(n6785), .Z(n6786) );
  XNOR U10884 ( .A(b[2605]), .B(n6787), .Z(c[2605]) );
  XOR U10885 ( .A(n6788), .B(n6789), .Z(n6785) );
  ANDN U10886 ( .B(n6790), .A(n6791), .Z(n6788) );
  XNOR U10887 ( .A(b[2604]), .B(n6789), .Z(n6790) );
  XNOR U10888 ( .A(b[2604]), .B(n6791), .Z(c[2604]) );
  XOR U10889 ( .A(n6792), .B(n6793), .Z(n6789) );
  ANDN U10890 ( .B(n6794), .A(n6795), .Z(n6792) );
  XNOR U10891 ( .A(b[2603]), .B(n6793), .Z(n6794) );
  XNOR U10892 ( .A(b[2603]), .B(n6795), .Z(c[2603]) );
  XOR U10893 ( .A(n6796), .B(n6797), .Z(n6793) );
  ANDN U10894 ( .B(n6798), .A(n6799), .Z(n6796) );
  XNOR U10895 ( .A(b[2602]), .B(n6797), .Z(n6798) );
  XNOR U10896 ( .A(b[2602]), .B(n6799), .Z(c[2602]) );
  XOR U10897 ( .A(n6800), .B(n6801), .Z(n6797) );
  ANDN U10898 ( .B(n6802), .A(n6803), .Z(n6800) );
  XNOR U10899 ( .A(b[2601]), .B(n6801), .Z(n6802) );
  XNOR U10900 ( .A(b[2601]), .B(n6803), .Z(c[2601]) );
  XOR U10901 ( .A(n6804), .B(n6805), .Z(n6801) );
  ANDN U10902 ( .B(n6806), .A(n6807), .Z(n6804) );
  XNOR U10903 ( .A(b[2600]), .B(n6805), .Z(n6806) );
  XNOR U10904 ( .A(b[2600]), .B(n6807), .Z(c[2600]) );
  XOR U10905 ( .A(n6808), .B(n6809), .Z(n6805) );
  ANDN U10906 ( .B(n6810), .A(n6811), .Z(n6808) );
  XNOR U10907 ( .A(b[2599]), .B(n6809), .Z(n6810) );
  XNOR U10908 ( .A(b[25]), .B(n6812), .Z(c[25]) );
  XNOR U10909 ( .A(b[259]), .B(n6813), .Z(c[259]) );
  XNOR U10910 ( .A(b[2599]), .B(n6811), .Z(c[2599]) );
  XOR U10911 ( .A(n6814), .B(n6815), .Z(n6809) );
  ANDN U10912 ( .B(n6816), .A(n6817), .Z(n6814) );
  XNOR U10913 ( .A(b[2598]), .B(n6815), .Z(n6816) );
  XNOR U10914 ( .A(b[2598]), .B(n6817), .Z(c[2598]) );
  XOR U10915 ( .A(n6818), .B(n6819), .Z(n6815) );
  ANDN U10916 ( .B(n6820), .A(n6821), .Z(n6818) );
  XNOR U10917 ( .A(b[2597]), .B(n6819), .Z(n6820) );
  XNOR U10918 ( .A(b[2597]), .B(n6821), .Z(c[2597]) );
  XOR U10919 ( .A(n6822), .B(n6823), .Z(n6819) );
  ANDN U10920 ( .B(n6824), .A(n6825), .Z(n6822) );
  XNOR U10921 ( .A(b[2596]), .B(n6823), .Z(n6824) );
  XNOR U10922 ( .A(b[2596]), .B(n6825), .Z(c[2596]) );
  XOR U10923 ( .A(n6826), .B(n6827), .Z(n6823) );
  ANDN U10924 ( .B(n6828), .A(n6829), .Z(n6826) );
  XNOR U10925 ( .A(b[2595]), .B(n6827), .Z(n6828) );
  XNOR U10926 ( .A(b[2595]), .B(n6829), .Z(c[2595]) );
  XOR U10927 ( .A(n6830), .B(n6831), .Z(n6827) );
  ANDN U10928 ( .B(n6832), .A(n6833), .Z(n6830) );
  XNOR U10929 ( .A(b[2594]), .B(n6831), .Z(n6832) );
  XNOR U10930 ( .A(b[2594]), .B(n6833), .Z(c[2594]) );
  XOR U10931 ( .A(n6834), .B(n6835), .Z(n6831) );
  ANDN U10932 ( .B(n6836), .A(n6837), .Z(n6834) );
  XNOR U10933 ( .A(b[2593]), .B(n6835), .Z(n6836) );
  XNOR U10934 ( .A(b[2593]), .B(n6837), .Z(c[2593]) );
  XOR U10935 ( .A(n6838), .B(n6839), .Z(n6835) );
  ANDN U10936 ( .B(n6840), .A(n6841), .Z(n6838) );
  XNOR U10937 ( .A(b[2592]), .B(n6839), .Z(n6840) );
  XNOR U10938 ( .A(b[2592]), .B(n6841), .Z(c[2592]) );
  XOR U10939 ( .A(n6842), .B(n6843), .Z(n6839) );
  ANDN U10940 ( .B(n6844), .A(n6845), .Z(n6842) );
  XNOR U10941 ( .A(b[2591]), .B(n6843), .Z(n6844) );
  XNOR U10942 ( .A(b[2591]), .B(n6845), .Z(c[2591]) );
  XOR U10943 ( .A(n6846), .B(n6847), .Z(n6843) );
  ANDN U10944 ( .B(n6848), .A(n6849), .Z(n6846) );
  XNOR U10945 ( .A(b[2590]), .B(n6847), .Z(n6848) );
  XNOR U10946 ( .A(b[2590]), .B(n6849), .Z(c[2590]) );
  XOR U10947 ( .A(n6850), .B(n6851), .Z(n6847) );
  ANDN U10948 ( .B(n6852), .A(n6853), .Z(n6850) );
  XNOR U10949 ( .A(b[2589]), .B(n6851), .Z(n6852) );
  XNOR U10950 ( .A(b[258]), .B(n6854), .Z(c[258]) );
  XNOR U10951 ( .A(b[2589]), .B(n6853), .Z(c[2589]) );
  XOR U10952 ( .A(n6855), .B(n6856), .Z(n6851) );
  ANDN U10953 ( .B(n6857), .A(n6858), .Z(n6855) );
  XNOR U10954 ( .A(b[2588]), .B(n6856), .Z(n6857) );
  XNOR U10955 ( .A(b[2588]), .B(n6858), .Z(c[2588]) );
  XOR U10956 ( .A(n6859), .B(n6860), .Z(n6856) );
  ANDN U10957 ( .B(n6861), .A(n6862), .Z(n6859) );
  XNOR U10958 ( .A(b[2587]), .B(n6860), .Z(n6861) );
  XNOR U10959 ( .A(b[2587]), .B(n6862), .Z(c[2587]) );
  XOR U10960 ( .A(n6863), .B(n6864), .Z(n6860) );
  ANDN U10961 ( .B(n6865), .A(n6866), .Z(n6863) );
  XNOR U10962 ( .A(b[2586]), .B(n6864), .Z(n6865) );
  XNOR U10963 ( .A(b[2586]), .B(n6866), .Z(c[2586]) );
  XOR U10964 ( .A(n6867), .B(n6868), .Z(n6864) );
  ANDN U10965 ( .B(n6869), .A(n6870), .Z(n6867) );
  XNOR U10966 ( .A(b[2585]), .B(n6868), .Z(n6869) );
  XNOR U10967 ( .A(b[2585]), .B(n6870), .Z(c[2585]) );
  XOR U10968 ( .A(n6871), .B(n6872), .Z(n6868) );
  ANDN U10969 ( .B(n6873), .A(n6874), .Z(n6871) );
  XNOR U10970 ( .A(b[2584]), .B(n6872), .Z(n6873) );
  XNOR U10971 ( .A(b[2584]), .B(n6874), .Z(c[2584]) );
  XOR U10972 ( .A(n6875), .B(n6876), .Z(n6872) );
  ANDN U10973 ( .B(n6877), .A(n6878), .Z(n6875) );
  XNOR U10974 ( .A(b[2583]), .B(n6876), .Z(n6877) );
  XNOR U10975 ( .A(b[2583]), .B(n6878), .Z(c[2583]) );
  XOR U10976 ( .A(n6879), .B(n6880), .Z(n6876) );
  ANDN U10977 ( .B(n6881), .A(n6882), .Z(n6879) );
  XNOR U10978 ( .A(b[2582]), .B(n6880), .Z(n6881) );
  XNOR U10979 ( .A(b[2582]), .B(n6882), .Z(c[2582]) );
  XOR U10980 ( .A(n6883), .B(n6884), .Z(n6880) );
  ANDN U10981 ( .B(n6885), .A(n6886), .Z(n6883) );
  XNOR U10982 ( .A(b[2581]), .B(n6884), .Z(n6885) );
  XNOR U10983 ( .A(b[2581]), .B(n6886), .Z(c[2581]) );
  XOR U10984 ( .A(n6887), .B(n6888), .Z(n6884) );
  ANDN U10985 ( .B(n6889), .A(n6890), .Z(n6887) );
  XNOR U10986 ( .A(b[2580]), .B(n6888), .Z(n6889) );
  XNOR U10987 ( .A(b[2580]), .B(n6890), .Z(c[2580]) );
  XOR U10988 ( .A(n6891), .B(n6892), .Z(n6888) );
  ANDN U10989 ( .B(n6893), .A(n6894), .Z(n6891) );
  XNOR U10990 ( .A(b[2579]), .B(n6892), .Z(n6893) );
  XNOR U10991 ( .A(b[257]), .B(n6895), .Z(c[257]) );
  XNOR U10992 ( .A(b[2579]), .B(n6894), .Z(c[2579]) );
  XOR U10993 ( .A(n6896), .B(n6897), .Z(n6892) );
  ANDN U10994 ( .B(n6898), .A(n6899), .Z(n6896) );
  XNOR U10995 ( .A(b[2578]), .B(n6897), .Z(n6898) );
  XNOR U10996 ( .A(b[2578]), .B(n6899), .Z(c[2578]) );
  XOR U10997 ( .A(n6900), .B(n6901), .Z(n6897) );
  ANDN U10998 ( .B(n6902), .A(n6903), .Z(n6900) );
  XNOR U10999 ( .A(b[2577]), .B(n6901), .Z(n6902) );
  XNOR U11000 ( .A(b[2577]), .B(n6903), .Z(c[2577]) );
  XOR U11001 ( .A(n6904), .B(n6905), .Z(n6901) );
  ANDN U11002 ( .B(n6906), .A(n6907), .Z(n6904) );
  XNOR U11003 ( .A(b[2576]), .B(n6905), .Z(n6906) );
  XNOR U11004 ( .A(b[2576]), .B(n6907), .Z(c[2576]) );
  XOR U11005 ( .A(n6908), .B(n6909), .Z(n6905) );
  ANDN U11006 ( .B(n6910), .A(n6911), .Z(n6908) );
  XNOR U11007 ( .A(b[2575]), .B(n6909), .Z(n6910) );
  XNOR U11008 ( .A(b[2575]), .B(n6911), .Z(c[2575]) );
  XOR U11009 ( .A(n6912), .B(n6913), .Z(n6909) );
  ANDN U11010 ( .B(n6914), .A(n6915), .Z(n6912) );
  XNOR U11011 ( .A(b[2574]), .B(n6913), .Z(n6914) );
  XNOR U11012 ( .A(b[2574]), .B(n6915), .Z(c[2574]) );
  XOR U11013 ( .A(n6916), .B(n6917), .Z(n6913) );
  ANDN U11014 ( .B(n6918), .A(n6919), .Z(n6916) );
  XNOR U11015 ( .A(b[2573]), .B(n6917), .Z(n6918) );
  XNOR U11016 ( .A(b[2573]), .B(n6919), .Z(c[2573]) );
  XOR U11017 ( .A(n6920), .B(n6921), .Z(n6917) );
  ANDN U11018 ( .B(n6922), .A(n6923), .Z(n6920) );
  XNOR U11019 ( .A(b[2572]), .B(n6921), .Z(n6922) );
  XNOR U11020 ( .A(b[2572]), .B(n6923), .Z(c[2572]) );
  XOR U11021 ( .A(n6924), .B(n6925), .Z(n6921) );
  ANDN U11022 ( .B(n6926), .A(n6927), .Z(n6924) );
  XNOR U11023 ( .A(b[2571]), .B(n6925), .Z(n6926) );
  XNOR U11024 ( .A(b[2571]), .B(n6927), .Z(c[2571]) );
  XOR U11025 ( .A(n6928), .B(n6929), .Z(n6925) );
  ANDN U11026 ( .B(n6930), .A(n6931), .Z(n6928) );
  XNOR U11027 ( .A(b[2570]), .B(n6929), .Z(n6930) );
  XNOR U11028 ( .A(b[2570]), .B(n6931), .Z(c[2570]) );
  XOR U11029 ( .A(n6932), .B(n6933), .Z(n6929) );
  ANDN U11030 ( .B(n6934), .A(n6935), .Z(n6932) );
  XNOR U11031 ( .A(b[2569]), .B(n6933), .Z(n6934) );
  XNOR U11032 ( .A(b[256]), .B(n6936), .Z(c[256]) );
  XNOR U11033 ( .A(b[2569]), .B(n6935), .Z(c[2569]) );
  XOR U11034 ( .A(n6937), .B(n6938), .Z(n6933) );
  ANDN U11035 ( .B(n6939), .A(n6940), .Z(n6937) );
  XNOR U11036 ( .A(b[2568]), .B(n6938), .Z(n6939) );
  XNOR U11037 ( .A(b[2568]), .B(n6940), .Z(c[2568]) );
  XOR U11038 ( .A(n6941), .B(n6942), .Z(n6938) );
  ANDN U11039 ( .B(n6943), .A(n6944), .Z(n6941) );
  XNOR U11040 ( .A(b[2567]), .B(n6942), .Z(n6943) );
  XNOR U11041 ( .A(b[2567]), .B(n6944), .Z(c[2567]) );
  XOR U11042 ( .A(n6945), .B(n6946), .Z(n6942) );
  ANDN U11043 ( .B(n6947), .A(n6948), .Z(n6945) );
  XNOR U11044 ( .A(b[2566]), .B(n6946), .Z(n6947) );
  XNOR U11045 ( .A(b[2566]), .B(n6948), .Z(c[2566]) );
  XOR U11046 ( .A(n6949), .B(n6950), .Z(n6946) );
  ANDN U11047 ( .B(n6951), .A(n6952), .Z(n6949) );
  XNOR U11048 ( .A(b[2565]), .B(n6950), .Z(n6951) );
  XNOR U11049 ( .A(b[2565]), .B(n6952), .Z(c[2565]) );
  XOR U11050 ( .A(n6953), .B(n6954), .Z(n6950) );
  ANDN U11051 ( .B(n6955), .A(n6956), .Z(n6953) );
  XNOR U11052 ( .A(b[2564]), .B(n6954), .Z(n6955) );
  XNOR U11053 ( .A(b[2564]), .B(n6956), .Z(c[2564]) );
  XOR U11054 ( .A(n6957), .B(n6958), .Z(n6954) );
  ANDN U11055 ( .B(n6959), .A(n6960), .Z(n6957) );
  XNOR U11056 ( .A(b[2563]), .B(n6958), .Z(n6959) );
  XNOR U11057 ( .A(b[2563]), .B(n6960), .Z(c[2563]) );
  XOR U11058 ( .A(n6961), .B(n6962), .Z(n6958) );
  ANDN U11059 ( .B(n6963), .A(n6964), .Z(n6961) );
  XNOR U11060 ( .A(b[2562]), .B(n6962), .Z(n6963) );
  XNOR U11061 ( .A(b[2562]), .B(n6964), .Z(c[2562]) );
  XOR U11062 ( .A(n6965), .B(n6966), .Z(n6962) );
  ANDN U11063 ( .B(n6967), .A(n6968), .Z(n6965) );
  XNOR U11064 ( .A(b[2561]), .B(n6966), .Z(n6967) );
  XNOR U11065 ( .A(b[2561]), .B(n6968), .Z(c[2561]) );
  XOR U11066 ( .A(n6969), .B(n6970), .Z(n6966) );
  ANDN U11067 ( .B(n6971), .A(n6972), .Z(n6969) );
  XNOR U11068 ( .A(b[2560]), .B(n6970), .Z(n6971) );
  XNOR U11069 ( .A(b[2560]), .B(n6972), .Z(c[2560]) );
  XOR U11070 ( .A(n6973), .B(n6974), .Z(n6970) );
  ANDN U11071 ( .B(n6975), .A(n6976), .Z(n6973) );
  XNOR U11072 ( .A(b[2559]), .B(n6974), .Z(n6975) );
  XNOR U11073 ( .A(b[255]), .B(n6977), .Z(c[255]) );
  XNOR U11074 ( .A(b[2559]), .B(n6976), .Z(c[2559]) );
  XOR U11075 ( .A(n6978), .B(n6979), .Z(n6974) );
  ANDN U11076 ( .B(n6980), .A(n6981), .Z(n6978) );
  XNOR U11077 ( .A(b[2558]), .B(n6979), .Z(n6980) );
  XNOR U11078 ( .A(b[2558]), .B(n6981), .Z(c[2558]) );
  XOR U11079 ( .A(n6982), .B(n6983), .Z(n6979) );
  ANDN U11080 ( .B(n6984), .A(n6985), .Z(n6982) );
  XNOR U11081 ( .A(b[2557]), .B(n6983), .Z(n6984) );
  XNOR U11082 ( .A(b[2557]), .B(n6985), .Z(c[2557]) );
  XOR U11083 ( .A(n6986), .B(n6987), .Z(n6983) );
  ANDN U11084 ( .B(n6988), .A(n6989), .Z(n6986) );
  XNOR U11085 ( .A(b[2556]), .B(n6987), .Z(n6988) );
  XNOR U11086 ( .A(b[2556]), .B(n6989), .Z(c[2556]) );
  XOR U11087 ( .A(n6990), .B(n6991), .Z(n6987) );
  ANDN U11088 ( .B(n6992), .A(n6993), .Z(n6990) );
  XNOR U11089 ( .A(b[2555]), .B(n6991), .Z(n6992) );
  XNOR U11090 ( .A(b[2555]), .B(n6993), .Z(c[2555]) );
  XOR U11091 ( .A(n6994), .B(n6995), .Z(n6991) );
  ANDN U11092 ( .B(n6996), .A(n6997), .Z(n6994) );
  XNOR U11093 ( .A(b[2554]), .B(n6995), .Z(n6996) );
  XNOR U11094 ( .A(b[2554]), .B(n6997), .Z(c[2554]) );
  XOR U11095 ( .A(n6998), .B(n6999), .Z(n6995) );
  ANDN U11096 ( .B(n7000), .A(n7001), .Z(n6998) );
  XNOR U11097 ( .A(b[2553]), .B(n6999), .Z(n7000) );
  XNOR U11098 ( .A(b[2553]), .B(n7001), .Z(c[2553]) );
  XOR U11099 ( .A(n7002), .B(n7003), .Z(n6999) );
  ANDN U11100 ( .B(n7004), .A(n7005), .Z(n7002) );
  XNOR U11101 ( .A(b[2552]), .B(n7003), .Z(n7004) );
  XNOR U11102 ( .A(b[2552]), .B(n7005), .Z(c[2552]) );
  XOR U11103 ( .A(n7006), .B(n7007), .Z(n7003) );
  ANDN U11104 ( .B(n7008), .A(n7009), .Z(n7006) );
  XNOR U11105 ( .A(b[2551]), .B(n7007), .Z(n7008) );
  XNOR U11106 ( .A(b[2551]), .B(n7009), .Z(c[2551]) );
  XOR U11107 ( .A(n7010), .B(n7011), .Z(n7007) );
  ANDN U11108 ( .B(n7012), .A(n7013), .Z(n7010) );
  XNOR U11109 ( .A(b[2550]), .B(n7011), .Z(n7012) );
  XNOR U11110 ( .A(b[2550]), .B(n7013), .Z(c[2550]) );
  XOR U11111 ( .A(n7014), .B(n7015), .Z(n7011) );
  ANDN U11112 ( .B(n7016), .A(n7017), .Z(n7014) );
  XNOR U11113 ( .A(b[2549]), .B(n7015), .Z(n7016) );
  XNOR U11114 ( .A(b[254]), .B(n7018), .Z(c[254]) );
  XNOR U11115 ( .A(b[2549]), .B(n7017), .Z(c[2549]) );
  XOR U11116 ( .A(n7019), .B(n7020), .Z(n7015) );
  ANDN U11117 ( .B(n7021), .A(n7022), .Z(n7019) );
  XNOR U11118 ( .A(b[2548]), .B(n7020), .Z(n7021) );
  XNOR U11119 ( .A(b[2548]), .B(n7022), .Z(c[2548]) );
  XOR U11120 ( .A(n7023), .B(n7024), .Z(n7020) );
  ANDN U11121 ( .B(n7025), .A(n7026), .Z(n7023) );
  XNOR U11122 ( .A(b[2547]), .B(n7024), .Z(n7025) );
  XNOR U11123 ( .A(b[2547]), .B(n7026), .Z(c[2547]) );
  XOR U11124 ( .A(n7027), .B(n7028), .Z(n7024) );
  ANDN U11125 ( .B(n7029), .A(n7030), .Z(n7027) );
  XNOR U11126 ( .A(b[2546]), .B(n7028), .Z(n7029) );
  XNOR U11127 ( .A(b[2546]), .B(n7030), .Z(c[2546]) );
  XOR U11128 ( .A(n7031), .B(n7032), .Z(n7028) );
  ANDN U11129 ( .B(n7033), .A(n7034), .Z(n7031) );
  XNOR U11130 ( .A(b[2545]), .B(n7032), .Z(n7033) );
  XNOR U11131 ( .A(b[2545]), .B(n7034), .Z(c[2545]) );
  XOR U11132 ( .A(n7035), .B(n7036), .Z(n7032) );
  ANDN U11133 ( .B(n7037), .A(n7038), .Z(n7035) );
  XNOR U11134 ( .A(b[2544]), .B(n7036), .Z(n7037) );
  XNOR U11135 ( .A(b[2544]), .B(n7038), .Z(c[2544]) );
  XOR U11136 ( .A(n7039), .B(n7040), .Z(n7036) );
  ANDN U11137 ( .B(n7041), .A(n7042), .Z(n7039) );
  XNOR U11138 ( .A(b[2543]), .B(n7040), .Z(n7041) );
  XNOR U11139 ( .A(b[2543]), .B(n7042), .Z(c[2543]) );
  XOR U11140 ( .A(n7043), .B(n7044), .Z(n7040) );
  ANDN U11141 ( .B(n7045), .A(n7046), .Z(n7043) );
  XNOR U11142 ( .A(b[2542]), .B(n7044), .Z(n7045) );
  XNOR U11143 ( .A(b[2542]), .B(n7046), .Z(c[2542]) );
  XOR U11144 ( .A(n7047), .B(n7048), .Z(n7044) );
  ANDN U11145 ( .B(n7049), .A(n7050), .Z(n7047) );
  XNOR U11146 ( .A(b[2541]), .B(n7048), .Z(n7049) );
  XNOR U11147 ( .A(b[2541]), .B(n7050), .Z(c[2541]) );
  XOR U11148 ( .A(n7051), .B(n7052), .Z(n7048) );
  ANDN U11149 ( .B(n7053), .A(n7054), .Z(n7051) );
  XNOR U11150 ( .A(b[2540]), .B(n7052), .Z(n7053) );
  XNOR U11151 ( .A(b[2540]), .B(n7054), .Z(c[2540]) );
  XOR U11152 ( .A(n7055), .B(n7056), .Z(n7052) );
  ANDN U11153 ( .B(n7057), .A(n7058), .Z(n7055) );
  XNOR U11154 ( .A(b[2539]), .B(n7056), .Z(n7057) );
  XNOR U11155 ( .A(b[253]), .B(n7059), .Z(c[253]) );
  XNOR U11156 ( .A(b[2539]), .B(n7058), .Z(c[2539]) );
  XOR U11157 ( .A(n7060), .B(n7061), .Z(n7056) );
  ANDN U11158 ( .B(n7062), .A(n7063), .Z(n7060) );
  XNOR U11159 ( .A(b[2538]), .B(n7061), .Z(n7062) );
  XNOR U11160 ( .A(b[2538]), .B(n7063), .Z(c[2538]) );
  XOR U11161 ( .A(n7064), .B(n7065), .Z(n7061) );
  ANDN U11162 ( .B(n7066), .A(n7067), .Z(n7064) );
  XNOR U11163 ( .A(b[2537]), .B(n7065), .Z(n7066) );
  XNOR U11164 ( .A(b[2537]), .B(n7067), .Z(c[2537]) );
  XOR U11165 ( .A(n7068), .B(n7069), .Z(n7065) );
  ANDN U11166 ( .B(n7070), .A(n7071), .Z(n7068) );
  XNOR U11167 ( .A(b[2536]), .B(n7069), .Z(n7070) );
  XNOR U11168 ( .A(b[2536]), .B(n7071), .Z(c[2536]) );
  XOR U11169 ( .A(n7072), .B(n7073), .Z(n7069) );
  ANDN U11170 ( .B(n7074), .A(n7075), .Z(n7072) );
  XNOR U11171 ( .A(b[2535]), .B(n7073), .Z(n7074) );
  XNOR U11172 ( .A(b[2535]), .B(n7075), .Z(c[2535]) );
  XOR U11173 ( .A(n7076), .B(n7077), .Z(n7073) );
  ANDN U11174 ( .B(n7078), .A(n7079), .Z(n7076) );
  XNOR U11175 ( .A(b[2534]), .B(n7077), .Z(n7078) );
  XNOR U11176 ( .A(b[2534]), .B(n7079), .Z(c[2534]) );
  XOR U11177 ( .A(n7080), .B(n7081), .Z(n7077) );
  ANDN U11178 ( .B(n7082), .A(n7083), .Z(n7080) );
  XNOR U11179 ( .A(b[2533]), .B(n7081), .Z(n7082) );
  XNOR U11180 ( .A(b[2533]), .B(n7083), .Z(c[2533]) );
  XOR U11181 ( .A(n7084), .B(n7085), .Z(n7081) );
  ANDN U11182 ( .B(n7086), .A(n7087), .Z(n7084) );
  XNOR U11183 ( .A(b[2532]), .B(n7085), .Z(n7086) );
  XNOR U11184 ( .A(b[2532]), .B(n7087), .Z(c[2532]) );
  XOR U11185 ( .A(n7088), .B(n7089), .Z(n7085) );
  ANDN U11186 ( .B(n7090), .A(n7091), .Z(n7088) );
  XNOR U11187 ( .A(b[2531]), .B(n7089), .Z(n7090) );
  XNOR U11188 ( .A(b[2531]), .B(n7091), .Z(c[2531]) );
  XOR U11189 ( .A(n7092), .B(n7093), .Z(n7089) );
  ANDN U11190 ( .B(n7094), .A(n7095), .Z(n7092) );
  XNOR U11191 ( .A(b[2530]), .B(n7093), .Z(n7094) );
  XNOR U11192 ( .A(b[2530]), .B(n7095), .Z(c[2530]) );
  XOR U11193 ( .A(n7096), .B(n7097), .Z(n7093) );
  ANDN U11194 ( .B(n7098), .A(n7099), .Z(n7096) );
  XNOR U11195 ( .A(b[2529]), .B(n7097), .Z(n7098) );
  XNOR U11196 ( .A(b[252]), .B(n7100), .Z(c[252]) );
  XNOR U11197 ( .A(b[2529]), .B(n7099), .Z(c[2529]) );
  XOR U11198 ( .A(n7101), .B(n7102), .Z(n7097) );
  ANDN U11199 ( .B(n7103), .A(n7104), .Z(n7101) );
  XNOR U11200 ( .A(b[2528]), .B(n7102), .Z(n7103) );
  XNOR U11201 ( .A(b[2528]), .B(n7104), .Z(c[2528]) );
  XOR U11202 ( .A(n7105), .B(n7106), .Z(n7102) );
  ANDN U11203 ( .B(n7107), .A(n7108), .Z(n7105) );
  XNOR U11204 ( .A(b[2527]), .B(n7106), .Z(n7107) );
  XNOR U11205 ( .A(b[2527]), .B(n7108), .Z(c[2527]) );
  XOR U11206 ( .A(n7109), .B(n7110), .Z(n7106) );
  ANDN U11207 ( .B(n7111), .A(n7112), .Z(n7109) );
  XNOR U11208 ( .A(b[2526]), .B(n7110), .Z(n7111) );
  XNOR U11209 ( .A(b[2526]), .B(n7112), .Z(c[2526]) );
  XOR U11210 ( .A(n7113), .B(n7114), .Z(n7110) );
  ANDN U11211 ( .B(n7115), .A(n7116), .Z(n7113) );
  XNOR U11212 ( .A(b[2525]), .B(n7114), .Z(n7115) );
  XNOR U11213 ( .A(b[2525]), .B(n7116), .Z(c[2525]) );
  XOR U11214 ( .A(n7117), .B(n7118), .Z(n7114) );
  ANDN U11215 ( .B(n7119), .A(n7120), .Z(n7117) );
  XNOR U11216 ( .A(b[2524]), .B(n7118), .Z(n7119) );
  XNOR U11217 ( .A(b[2524]), .B(n7120), .Z(c[2524]) );
  XOR U11218 ( .A(n7121), .B(n7122), .Z(n7118) );
  ANDN U11219 ( .B(n7123), .A(n7124), .Z(n7121) );
  XNOR U11220 ( .A(b[2523]), .B(n7122), .Z(n7123) );
  XNOR U11221 ( .A(b[2523]), .B(n7124), .Z(c[2523]) );
  XOR U11222 ( .A(n7125), .B(n7126), .Z(n7122) );
  ANDN U11223 ( .B(n7127), .A(n7128), .Z(n7125) );
  XNOR U11224 ( .A(b[2522]), .B(n7126), .Z(n7127) );
  XNOR U11225 ( .A(b[2522]), .B(n7128), .Z(c[2522]) );
  XOR U11226 ( .A(n7129), .B(n7130), .Z(n7126) );
  ANDN U11227 ( .B(n7131), .A(n7132), .Z(n7129) );
  XNOR U11228 ( .A(b[2521]), .B(n7130), .Z(n7131) );
  XNOR U11229 ( .A(b[2521]), .B(n7132), .Z(c[2521]) );
  XOR U11230 ( .A(n7133), .B(n7134), .Z(n7130) );
  ANDN U11231 ( .B(n7135), .A(n7136), .Z(n7133) );
  XNOR U11232 ( .A(b[2520]), .B(n7134), .Z(n7135) );
  XNOR U11233 ( .A(b[2520]), .B(n7136), .Z(c[2520]) );
  XOR U11234 ( .A(n7137), .B(n7138), .Z(n7134) );
  ANDN U11235 ( .B(n7139), .A(n7140), .Z(n7137) );
  XNOR U11236 ( .A(b[2519]), .B(n7138), .Z(n7139) );
  XNOR U11237 ( .A(b[251]), .B(n7141), .Z(c[251]) );
  XNOR U11238 ( .A(b[2519]), .B(n7140), .Z(c[2519]) );
  XOR U11239 ( .A(n7142), .B(n7143), .Z(n7138) );
  ANDN U11240 ( .B(n7144), .A(n7145), .Z(n7142) );
  XNOR U11241 ( .A(b[2518]), .B(n7143), .Z(n7144) );
  XNOR U11242 ( .A(b[2518]), .B(n7145), .Z(c[2518]) );
  XOR U11243 ( .A(n7146), .B(n7147), .Z(n7143) );
  ANDN U11244 ( .B(n7148), .A(n7149), .Z(n7146) );
  XNOR U11245 ( .A(b[2517]), .B(n7147), .Z(n7148) );
  XNOR U11246 ( .A(b[2517]), .B(n7149), .Z(c[2517]) );
  XOR U11247 ( .A(n7150), .B(n7151), .Z(n7147) );
  ANDN U11248 ( .B(n7152), .A(n7153), .Z(n7150) );
  XNOR U11249 ( .A(b[2516]), .B(n7151), .Z(n7152) );
  XNOR U11250 ( .A(b[2516]), .B(n7153), .Z(c[2516]) );
  XOR U11251 ( .A(n7154), .B(n7155), .Z(n7151) );
  ANDN U11252 ( .B(n7156), .A(n7157), .Z(n7154) );
  XNOR U11253 ( .A(b[2515]), .B(n7155), .Z(n7156) );
  XNOR U11254 ( .A(b[2515]), .B(n7157), .Z(c[2515]) );
  XOR U11255 ( .A(n7158), .B(n7159), .Z(n7155) );
  ANDN U11256 ( .B(n7160), .A(n7161), .Z(n7158) );
  XNOR U11257 ( .A(b[2514]), .B(n7159), .Z(n7160) );
  XNOR U11258 ( .A(b[2514]), .B(n7161), .Z(c[2514]) );
  XOR U11259 ( .A(n7162), .B(n7163), .Z(n7159) );
  ANDN U11260 ( .B(n7164), .A(n7165), .Z(n7162) );
  XNOR U11261 ( .A(b[2513]), .B(n7163), .Z(n7164) );
  XNOR U11262 ( .A(b[2513]), .B(n7165), .Z(c[2513]) );
  XOR U11263 ( .A(n7166), .B(n7167), .Z(n7163) );
  ANDN U11264 ( .B(n7168), .A(n7169), .Z(n7166) );
  XNOR U11265 ( .A(b[2512]), .B(n7167), .Z(n7168) );
  XNOR U11266 ( .A(b[2512]), .B(n7169), .Z(c[2512]) );
  XOR U11267 ( .A(n7170), .B(n7171), .Z(n7167) );
  ANDN U11268 ( .B(n7172), .A(n7173), .Z(n7170) );
  XNOR U11269 ( .A(b[2511]), .B(n7171), .Z(n7172) );
  XNOR U11270 ( .A(b[2511]), .B(n7173), .Z(c[2511]) );
  XOR U11271 ( .A(n7174), .B(n7175), .Z(n7171) );
  ANDN U11272 ( .B(n7176), .A(n7177), .Z(n7174) );
  XNOR U11273 ( .A(b[2510]), .B(n7175), .Z(n7176) );
  XNOR U11274 ( .A(b[2510]), .B(n7177), .Z(c[2510]) );
  XOR U11275 ( .A(n7178), .B(n7179), .Z(n7175) );
  ANDN U11276 ( .B(n7180), .A(n7181), .Z(n7178) );
  XNOR U11277 ( .A(b[2509]), .B(n7179), .Z(n7180) );
  XNOR U11278 ( .A(b[250]), .B(n7182), .Z(c[250]) );
  XNOR U11279 ( .A(b[2509]), .B(n7181), .Z(c[2509]) );
  XOR U11280 ( .A(n7183), .B(n7184), .Z(n7179) );
  ANDN U11281 ( .B(n7185), .A(n7186), .Z(n7183) );
  XNOR U11282 ( .A(b[2508]), .B(n7184), .Z(n7185) );
  XNOR U11283 ( .A(b[2508]), .B(n7186), .Z(c[2508]) );
  XOR U11284 ( .A(n7187), .B(n7188), .Z(n7184) );
  ANDN U11285 ( .B(n7189), .A(n7190), .Z(n7187) );
  XNOR U11286 ( .A(b[2507]), .B(n7188), .Z(n7189) );
  XNOR U11287 ( .A(b[2507]), .B(n7190), .Z(c[2507]) );
  XOR U11288 ( .A(n7191), .B(n7192), .Z(n7188) );
  ANDN U11289 ( .B(n7193), .A(n7194), .Z(n7191) );
  XNOR U11290 ( .A(b[2506]), .B(n7192), .Z(n7193) );
  XNOR U11291 ( .A(b[2506]), .B(n7194), .Z(c[2506]) );
  XOR U11292 ( .A(n7195), .B(n7196), .Z(n7192) );
  ANDN U11293 ( .B(n7197), .A(n7198), .Z(n7195) );
  XNOR U11294 ( .A(b[2505]), .B(n7196), .Z(n7197) );
  XNOR U11295 ( .A(b[2505]), .B(n7198), .Z(c[2505]) );
  XOR U11296 ( .A(n7199), .B(n7200), .Z(n7196) );
  ANDN U11297 ( .B(n7201), .A(n7202), .Z(n7199) );
  XNOR U11298 ( .A(b[2504]), .B(n7200), .Z(n7201) );
  XNOR U11299 ( .A(b[2504]), .B(n7202), .Z(c[2504]) );
  XOR U11300 ( .A(n7203), .B(n7204), .Z(n7200) );
  ANDN U11301 ( .B(n7205), .A(n7206), .Z(n7203) );
  XNOR U11302 ( .A(b[2503]), .B(n7204), .Z(n7205) );
  XNOR U11303 ( .A(b[2503]), .B(n7206), .Z(c[2503]) );
  XOR U11304 ( .A(n7207), .B(n7208), .Z(n7204) );
  ANDN U11305 ( .B(n7209), .A(n7210), .Z(n7207) );
  XNOR U11306 ( .A(b[2502]), .B(n7208), .Z(n7209) );
  XNOR U11307 ( .A(b[2502]), .B(n7210), .Z(c[2502]) );
  XOR U11308 ( .A(n7211), .B(n7212), .Z(n7208) );
  ANDN U11309 ( .B(n7213), .A(n7214), .Z(n7211) );
  XNOR U11310 ( .A(b[2501]), .B(n7212), .Z(n7213) );
  XNOR U11311 ( .A(b[2501]), .B(n7214), .Z(c[2501]) );
  XOR U11312 ( .A(n7215), .B(n7216), .Z(n7212) );
  ANDN U11313 ( .B(n7217), .A(n7218), .Z(n7215) );
  XNOR U11314 ( .A(b[2500]), .B(n7216), .Z(n7217) );
  XNOR U11315 ( .A(b[2500]), .B(n7218), .Z(c[2500]) );
  XOR U11316 ( .A(n7219), .B(n7220), .Z(n7216) );
  ANDN U11317 ( .B(n7221), .A(n7222), .Z(n7219) );
  XNOR U11318 ( .A(b[2499]), .B(n7220), .Z(n7221) );
  XNOR U11319 ( .A(b[24]), .B(n7223), .Z(c[24]) );
  XNOR U11320 ( .A(b[249]), .B(n7224), .Z(c[249]) );
  XNOR U11321 ( .A(b[2499]), .B(n7222), .Z(c[2499]) );
  XOR U11322 ( .A(n7225), .B(n7226), .Z(n7220) );
  ANDN U11323 ( .B(n7227), .A(n7228), .Z(n7225) );
  XNOR U11324 ( .A(b[2498]), .B(n7226), .Z(n7227) );
  XNOR U11325 ( .A(b[2498]), .B(n7228), .Z(c[2498]) );
  XOR U11326 ( .A(n7229), .B(n7230), .Z(n7226) );
  ANDN U11327 ( .B(n7231), .A(n7232), .Z(n7229) );
  XNOR U11328 ( .A(b[2497]), .B(n7230), .Z(n7231) );
  XNOR U11329 ( .A(b[2497]), .B(n7232), .Z(c[2497]) );
  XOR U11330 ( .A(n7233), .B(n7234), .Z(n7230) );
  ANDN U11331 ( .B(n7235), .A(n7236), .Z(n7233) );
  XNOR U11332 ( .A(b[2496]), .B(n7234), .Z(n7235) );
  XNOR U11333 ( .A(b[2496]), .B(n7236), .Z(c[2496]) );
  XOR U11334 ( .A(n7237), .B(n7238), .Z(n7234) );
  ANDN U11335 ( .B(n7239), .A(n7240), .Z(n7237) );
  XNOR U11336 ( .A(b[2495]), .B(n7238), .Z(n7239) );
  XNOR U11337 ( .A(b[2495]), .B(n7240), .Z(c[2495]) );
  XOR U11338 ( .A(n7241), .B(n7242), .Z(n7238) );
  ANDN U11339 ( .B(n7243), .A(n7244), .Z(n7241) );
  XNOR U11340 ( .A(b[2494]), .B(n7242), .Z(n7243) );
  XNOR U11341 ( .A(b[2494]), .B(n7244), .Z(c[2494]) );
  XOR U11342 ( .A(n7245), .B(n7246), .Z(n7242) );
  ANDN U11343 ( .B(n7247), .A(n7248), .Z(n7245) );
  XNOR U11344 ( .A(b[2493]), .B(n7246), .Z(n7247) );
  XNOR U11345 ( .A(b[2493]), .B(n7248), .Z(c[2493]) );
  XOR U11346 ( .A(n7249), .B(n7250), .Z(n7246) );
  ANDN U11347 ( .B(n7251), .A(n7252), .Z(n7249) );
  XNOR U11348 ( .A(b[2492]), .B(n7250), .Z(n7251) );
  XNOR U11349 ( .A(b[2492]), .B(n7252), .Z(c[2492]) );
  XOR U11350 ( .A(n7253), .B(n7254), .Z(n7250) );
  ANDN U11351 ( .B(n7255), .A(n7256), .Z(n7253) );
  XNOR U11352 ( .A(b[2491]), .B(n7254), .Z(n7255) );
  XNOR U11353 ( .A(b[2491]), .B(n7256), .Z(c[2491]) );
  XOR U11354 ( .A(n7257), .B(n7258), .Z(n7254) );
  ANDN U11355 ( .B(n7259), .A(n7260), .Z(n7257) );
  XNOR U11356 ( .A(b[2490]), .B(n7258), .Z(n7259) );
  XNOR U11357 ( .A(b[2490]), .B(n7260), .Z(c[2490]) );
  XOR U11358 ( .A(n7261), .B(n7262), .Z(n7258) );
  ANDN U11359 ( .B(n7263), .A(n7264), .Z(n7261) );
  XNOR U11360 ( .A(b[2489]), .B(n7262), .Z(n7263) );
  XNOR U11361 ( .A(b[248]), .B(n7265), .Z(c[248]) );
  XNOR U11362 ( .A(b[2489]), .B(n7264), .Z(c[2489]) );
  XOR U11363 ( .A(n7266), .B(n7267), .Z(n7262) );
  ANDN U11364 ( .B(n7268), .A(n7269), .Z(n7266) );
  XNOR U11365 ( .A(b[2488]), .B(n7267), .Z(n7268) );
  XNOR U11366 ( .A(b[2488]), .B(n7269), .Z(c[2488]) );
  XOR U11367 ( .A(n7270), .B(n7271), .Z(n7267) );
  ANDN U11368 ( .B(n7272), .A(n7273), .Z(n7270) );
  XNOR U11369 ( .A(b[2487]), .B(n7271), .Z(n7272) );
  XNOR U11370 ( .A(b[2487]), .B(n7273), .Z(c[2487]) );
  XOR U11371 ( .A(n7274), .B(n7275), .Z(n7271) );
  ANDN U11372 ( .B(n7276), .A(n7277), .Z(n7274) );
  XNOR U11373 ( .A(b[2486]), .B(n7275), .Z(n7276) );
  XNOR U11374 ( .A(b[2486]), .B(n7277), .Z(c[2486]) );
  XOR U11375 ( .A(n7278), .B(n7279), .Z(n7275) );
  ANDN U11376 ( .B(n7280), .A(n7281), .Z(n7278) );
  XNOR U11377 ( .A(b[2485]), .B(n7279), .Z(n7280) );
  XNOR U11378 ( .A(b[2485]), .B(n7281), .Z(c[2485]) );
  XOR U11379 ( .A(n7282), .B(n7283), .Z(n7279) );
  ANDN U11380 ( .B(n7284), .A(n7285), .Z(n7282) );
  XNOR U11381 ( .A(b[2484]), .B(n7283), .Z(n7284) );
  XNOR U11382 ( .A(b[2484]), .B(n7285), .Z(c[2484]) );
  XOR U11383 ( .A(n7286), .B(n7287), .Z(n7283) );
  ANDN U11384 ( .B(n7288), .A(n7289), .Z(n7286) );
  XNOR U11385 ( .A(b[2483]), .B(n7287), .Z(n7288) );
  XNOR U11386 ( .A(b[2483]), .B(n7289), .Z(c[2483]) );
  XOR U11387 ( .A(n7290), .B(n7291), .Z(n7287) );
  ANDN U11388 ( .B(n7292), .A(n7293), .Z(n7290) );
  XNOR U11389 ( .A(b[2482]), .B(n7291), .Z(n7292) );
  XNOR U11390 ( .A(b[2482]), .B(n7293), .Z(c[2482]) );
  XOR U11391 ( .A(n7294), .B(n7295), .Z(n7291) );
  ANDN U11392 ( .B(n7296), .A(n7297), .Z(n7294) );
  XNOR U11393 ( .A(b[2481]), .B(n7295), .Z(n7296) );
  XNOR U11394 ( .A(b[2481]), .B(n7297), .Z(c[2481]) );
  XOR U11395 ( .A(n7298), .B(n7299), .Z(n7295) );
  ANDN U11396 ( .B(n7300), .A(n7301), .Z(n7298) );
  XNOR U11397 ( .A(b[2480]), .B(n7299), .Z(n7300) );
  XNOR U11398 ( .A(b[2480]), .B(n7301), .Z(c[2480]) );
  XOR U11399 ( .A(n7302), .B(n7303), .Z(n7299) );
  ANDN U11400 ( .B(n7304), .A(n7305), .Z(n7302) );
  XNOR U11401 ( .A(b[2479]), .B(n7303), .Z(n7304) );
  XNOR U11402 ( .A(b[247]), .B(n7306), .Z(c[247]) );
  XNOR U11403 ( .A(b[2479]), .B(n7305), .Z(c[2479]) );
  XOR U11404 ( .A(n7307), .B(n7308), .Z(n7303) );
  ANDN U11405 ( .B(n7309), .A(n7310), .Z(n7307) );
  XNOR U11406 ( .A(b[2478]), .B(n7308), .Z(n7309) );
  XNOR U11407 ( .A(b[2478]), .B(n7310), .Z(c[2478]) );
  XOR U11408 ( .A(n7311), .B(n7312), .Z(n7308) );
  ANDN U11409 ( .B(n7313), .A(n7314), .Z(n7311) );
  XNOR U11410 ( .A(b[2477]), .B(n7312), .Z(n7313) );
  XNOR U11411 ( .A(b[2477]), .B(n7314), .Z(c[2477]) );
  XOR U11412 ( .A(n7315), .B(n7316), .Z(n7312) );
  ANDN U11413 ( .B(n7317), .A(n7318), .Z(n7315) );
  XNOR U11414 ( .A(b[2476]), .B(n7316), .Z(n7317) );
  XNOR U11415 ( .A(b[2476]), .B(n7318), .Z(c[2476]) );
  XOR U11416 ( .A(n7319), .B(n7320), .Z(n7316) );
  ANDN U11417 ( .B(n7321), .A(n7322), .Z(n7319) );
  XNOR U11418 ( .A(b[2475]), .B(n7320), .Z(n7321) );
  XNOR U11419 ( .A(b[2475]), .B(n7322), .Z(c[2475]) );
  XOR U11420 ( .A(n7323), .B(n7324), .Z(n7320) );
  ANDN U11421 ( .B(n7325), .A(n7326), .Z(n7323) );
  XNOR U11422 ( .A(b[2474]), .B(n7324), .Z(n7325) );
  XNOR U11423 ( .A(b[2474]), .B(n7326), .Z(c[2474]) );
  XOR U11424 ( .A(n7327), .B(n7328), .Z(n7324) );
  ANDN U11425 ( .B(n7329), .A(n7330), .Z(n7327) );
  XNOR U11426 ( .A(b[2473]), .B(n7328), .Z(n7329) );
  XNOR U11427 ( .A(b[2473]), .B(n7330), .Z(c[2473]) );
  XOR U11428 ( .A(n7331), .B(n7332), .Z(n7328) );
  ANDN U11429 ( .B(n7333), .A(n7334), .Z(n7331) );
  XNOR U11430 ( .A(b[2472]), .B(n7332), .Z(n7333) );
  XNOR U11431 ( .A(b[2472]), .B(n7334), .Z(c[2472]) );
  XOR U11432 ( .A(n7335), .B(n7336), .Z(n7332) );
  ANDN U11433 ( .B(n7337), .A(n7338), .Z(n7335) );
  XNOR U11434 ( .A(b[2471]), .B(n7336), .Z(n7337) );
  XNOR U11435 ( .A(b[2471]), .B(n7338), .Z(c[2471]) );
  XOR U11436 ( .A(n7339), .B(n7340), .Z(n7336) );
  ANDN U11437 ( .B(n7341), .A(n7342), .Z(n7339) );
  XNOR U11438 ( .A(b[2470]), .B(n7340), .Z(n7341) );
  XNOR U11439 ( .A(b[2470]), .B(n7342), .Z(c[2470]) );
  XOR U11440 ( .A(n7343), .B(n7344), .Z(n7340) );
  ANDN U11441 ( .B(n7345), .A(n7346), .Z(n7343) );
  XNOR U11442 ( .A(b[2469]), .B(n7344), .Z(n7345) );
  XNOR U11443 ( .A(b[246]), .B(n7347), .Z(c[246]) );
  XNOR U11444 ( .A(b[2469]), .B(n7346), .Z(c[2469]) );
  XOR U11445 ( .A(n7348), .B(n7349), .Z(n7344) );
  ANDN U11446 ( .B(n7350), .A(n7351), .Z(n7348) );
  XNOR U11447 ( .A(b[2468]), .B(n7349), .Z(n7350) );
  XNOR U11448 ( .A(b[2468]), .B(n7351), .Z(c[2468]) );
  XOR U11449 ( .A(n7352), .B(n7353), .Z(n7349) );
  ANDN U11450 ( .B(n7354), .A(n7355), .Z(n7352) );
  XNOR U11451 ( .A(b[2467]), .B(n7353), .Z(n7354) );
  XNOR U11452 ( .A(b[2467]), .B(n7355), .Z(c[2467]) );
  XOR U11453 ( .A(n7356), .B(n7357), .Z(n7353) );
  ANDN U11454 ( .B(n7358), .A(n7359), .Z(n7356) );
  XNOR U11455 ( .A(b[2466]), .B(n7357), .Z(n7358) );
  XNOR U11456 ( .A(b[2466]), .B(n7359), .Z(c[2466]) );
  XOR U11457 ( .A(n7360), .B(n7361), .Z(n7357) );
  ANDN U11458 ( .B(n7362), .A(n7363), .Z(n7360) );
  XNOR U11459 ( .A(b[2465]), .B(n7361), .Z(n7362) );
  XNOR U11460 ( .A(b[2465]), .B(n7363), .Z(c[2465]) );
  XOR U11461 ( .A(n7364), .B(n7365), .Z(n7361) );
  ANDN U11462 ( .B(n7366), .A(n7367), .Z(n7364) );
  XNOR U11463 ( .A(b[2464]), .B(n7365), .Z(n7366) );
  XNOR U11464 ( .A(b[2464]), .B(n7367), .Z(c[2464]) );
  XOR U11465 ( .A(n7368), .B(n7369), .Z(n7365) );
  ANDN U11466 ( .B(n7370), .A(n7371), .Z(n7368) );
  XNOR U11467 ( .A(b[2463]), .B(n7369), .Z(n7370) );
  XNOR U11468 ( .A(b[2463]), .B(n7371), .Z(c[2463]) );
  XOR U11469 ( .A(n7372), .B(n7373), .Z(n7369) );
  ANDN U11470 ( .B(n7374), .A(n7375), .Z(n7372) );
  XNOR U11471 ( .A(b[2462]), .B(n7373), .Z(n7374) );
  XNOR U11472 ( .A(b[2462]), .B(n7375), .Z(c[2462]) );
  XOR U11473 ( .A(n7376), .B(n7377), .Z(n7373) );
  ANDN U11474 ( .B(n7378), .A(n7379), .Z(n7376) );
  XNOR U11475 ( .A(b[2461]), .B(n7377), .Z(n7378) );
  XNOR U11476 ( .A(b[2461]), .B(n7379), .Z(c[2461]) );
  XOR U11477 ( .A(n7380), .B(n7381), .Z(n7377) );
  ANDN U11478 ( .B(n7382), .A(n7383), .Z(n7380) );
  XNOR U11479 ( .A(b[2460]), .B(n7381), .Z(n7382) );
  XNOR U11480 ( .A(b[2460]), .B(n7383), .Z(c[2460]) );
  XOR U11481 ( .A(n7384), .B(n7385), .Z(n7381) );
  ANDN U11482 ( .B(n7386), .A(n7387), .Z(n7384) );
  XNOR U11483 ( .A(b[2459]), .B(n7385), .Z(n7386) );
  XNOR U11484 ( .A(b[245]), .B(n7388), .Z(c[245]) );
  XNOR U11485 ( .A(b[2459]), .B(n7387), .Z(c[2459]) );
  XOR U11486 ( .A(n7389), .B(n7390), .Z(n7385) );
  ANDN U11487 ( .B(n7391), .A(n7392), .Z(n7389) );
  XNOR U11488 ( .A(b[2458]), .B(n7390), .Z(n7391) );
  XNOR U11489 ( .A(b[2458]), .B(n7392), .Z(c[2458]) );
  XOR U11490 ( .A(n7393), .B(n7394), .Z(n7390) );
  ANDN U11491 ( .B(n7395), .A(n7396), .Z(n7393) );
  XNOR U11492 ( .A(b[2457]), .B(n7394), .Z(n7395) );
  XNOR U11493 ( .A(b[2457]), .B(n7396), .Z(c[2457]) );
  XOR U11494 ( .A(n7397), .B(n7398), .Z(n7394) );
  ANDN U11495 ( .B(n7399), .A(n7400), .Z(n7397) );
  XNOR U11496 ( .A(b[2456]), .B(n7398), .Z(n7399) );
  XNOR U11497 ( .A(b[2456]), .B(n7400), .Z(c[2456]) );
  XOR U11498 ( .A(n7401), .B(n7402), .Z(n7398) );
  ANDN U11499 ( .B(n7403), .A(n7404), .Z(n7401) );
  XNOR U11500 ( .A(b[2455]), .B(n7402), .Z(n7403) );
  XNOR U11501 ( .A(b[2455]), .B(n7404), .Z(c[2455]) );
  XOR U11502 ( .A(n7405), .B(n7406), .Z(n7402) );
  ANDN U11503 ( .B(n7407), .A(n7408), .Z(n7405) );
  XNOR U11504 ( .A(b[2454]), .B(n7406), .Z(n7407) );
  XNOR U11505 ( .A(b[2454]), .B(n7408), .Z(c[2454]) );
  XOR U11506 ( .A(n7409), .B(n7410), .Z(n7406) );
  ANDN U11507 ( .B(n7411), .A(n7412), .Z(n7409) );
  XNOR U11508 ( .A(b[2453]), .B(n7410), .Z(n7411) );
  XNOR U11509 ( .A(b[2453]), .B(n7412), .Z(c[2453]) );
  XOR U11510 ( .A(n7413), .B(n7414), .Z(n7410) );
  ANDN U11511 ( .B(n7415), .A(n7416), .Z(n7413) );
  XNOR U11512 ( .A(b[2452]), .B(n7414), .Z(n7415) );
  XNOR U11513 ( .A(b[2452]), .B(n7416), .Z(c[2452]) );
  XOR U11514 ( .A(n7417), .B(n7418), .Z(n7414) );
  ANDN U11515 ( .B(n7419), .A(n7420), .Z(n7417) );
  XNOR U11516 ( .A(b[2451]), .B(n7418), .Z(n7419) );
  XNOR U11517 ( .A(b[2451]), .B(n7420), .Z(c[2451]) );
  XOR U11518 ( .A(n7421), .B(n7422), .Z(n7418) );
  ANDN U11519 ( .B(n7423), .A(n7424), .Z(n7421) );
  XNOR U11520 ( .A(b[2450]), .B(n7422), .Z(n7423) );
  XNOR U11521 ( .A(b[2450]), .B(n7424), .Z(c[2450]) );
  XOR U11522 ( .A(n7425), .B(n7426), .Z(n7422) );
  ANDN U11523 ( .B(n7427), .A(n7428), .Z(n7425) );
  XNOR U11524 ( .A(b[2449]), .B(n7426), .Z(n7427) );
  XNOR U11525 ( .A(b[244]), .B(n7429), .Z(c[244]) );
  XNOR U11526 ( .A(b[2449]), .B(n7428), .Z(c[2449]) );
  XOR U11527 ( .A(n7430), .B(n7431), .Z(n7426) );
  ANDN U11528 ( .B(n7432), .A(n7433), .Z(n7430) );
  XNOR U11529 ( .A(b[2448]), .B(n7431), .Z(n7432) );
  XNOR U11530 ( .A(b[2448]), .B(n7433), .Z(c[2448]) );
  XOR U11531 ( .A(n7434), .B(n7435), .Z(n7431) );
  ANDN U11532 ( .B(n7436), .A(n7437), .Z(n7434) );
  XNOR U11533 ( .A(b[2447]), .B(n7435), .Z(n7436) );
  XNOR U11534 ( .A(b[2447]), .B(n7437), .Z(c[2447]) );
  XOR U11535 ( .A(n7438), .B(n7439), .Z(n7435) );
  ANDN U11536 ( .B(n7440), .A(n7441), .Z(n7438) );
  XNOR U11537 ( .A(b[2446]), .B(n7439), .Z(n7440) );
  XNOR U11538 ( .A(b[2446]), .B(n7441), .Z(c[2446]) );
  XOR U11539 ( .A(n7442), .B(n7443), .Z(n7439) );
  ANDN U11540 ( .B(n7444), .A(n7445), .Z(n7442) );
  XNOR U11541 ( .A(b[2445]), .B(n7443), .Z(n7444) );
  XNOR U11542 ( .A(b[2445]), .B(n7445), .Z(c[2445]) );
  XOR U11543 ( .A(n7446), .B(n7447), .Z(n7443) );
  ANDN U11544 ( .B(n7448), .A(n7449), .Z(n7446) );
  XNOR U11545 ( .A(b[2444]), .B(n7447), .Z(n7448) );
  XNOR U11546 ( .A(b[2444]), .B(n7449), .Z(c[2444]) );
  XOR U11547 ( .A(n7450), .B(n7451), .Z(n7447) );
  ANDN U11548 ( .B(n7452), .A(n7453), .Z(n7450) );
  XNOR U11549 ( .A(b[2443]), .B(n7451), .Z(n7452) );
  XNOR U11550 ( .A(b[2443]), .B(n7453), .Z(c[2443]) );
  XOR U11551 ( .A(n7454), .B(n7455), .Z(n7451) );
  ANDN U11552 ( .B(n7456), .A(n7457), .Z(n7454) );
  XNOR U11553 ( .A(b[2442]), .B(n7455), .Z(n7456) );
  XNOR U11554 ( .A(b[2442]), .B(n7457), .Z(c[2442]) );
  XOR U11555 ( .A(n7458), .B(n7459), .Z(n7455) );
  ANDN U11556 ( .B(n7460), .A(n7461), .Z(n7458) );
  XNOR U11557 ( .A(b[2441]), .B(n7459), .Z(n7460) );
  XNOR U11558 ( .A(b[2441]), .B(n7461), .Z(c[2441]) );
  XOR U11559 ( .A(n7462), .B(n7463), .Z(n7459) );
  ANDN U11560 ( .B(n7464), .A(n7465), .Z(n7462) );
  XNOR U11561 ( .A(b[2440]), .B(n7463), .Z(n7464) );
  XNOR U11562 ( .A(b[2440]), .B(n7465), .Z(c[2440]) );
  XOR U11563 ( .A(n7466), .B(n7467), .Z(n7463) );
  ANDN U11564 ( .B(n7468), .A(n7469), .Z(n7466) );
  XNOR U11565 ( .A(b[2439]), .B(n7467), .Z(n7468) );
  XNOR U11566 ( .A(b[243]), .B(n7470), .Z(c[243]) );
  XNOR U11567 ( .A(b[2439]), .B(n7469), .Z(c[2439]) );
  XOR U11568 ( .A(n7471), .B(n7472), .Z(n7467) );
  ANDN U11569 ( .B(n7473), .A(n7474), .Z(n7471) );
  XNOR U11570 ( .A(b[2438]), .B(n7472), .Z(n7473) );
  XNOR U11571 ( .A(b[2438]), .B(n7474), .Z(c[2438]) );
  XOR U11572 ( .A(n7475), .B(n7476), .Z(n7472) );
  ANDN U11573 ( .B(n7477), .A(n7478), .Z(n7475) );
  XNOR U11574 ( .A(b[2437]), .B(n7476), .Z(n7477) );
  XNOR U11575 ( .A(b[2437]), .B(n7478), .Z(c[2437]) );
  XOR U11576 ( .A(n7479), .B(n7480), .Z(n7476) );
  ANDN U11577 ( .B(n7481), .A(n7482), .Z(n7479) );
  XNOR U11578 ( .A(b[2436]), .B(n7480), .Z(n7481) );
  XNOR U11579 ( .A(b[2436]), .B(n7482), .Z(c[2436]) );
  XOR U11580 ( .A(n7483), .B(n7484), .Z(n7480) );
  ANDN U11581 ( .B(n7485), .A(n7486), .Z(n7483) );
  XNOR U11582 ( .A(b[2435]), .B(n7484), .Z(n7485) );
  XNOR U11583 ( .A(b[2435]), .B(n7486), .Z(c[2435]) );
  XOR U11584 ( .A(n7487), .B(n7488), .Z(n7484) );
  ANDN U11585 ( .B(n7489), .A(n7490), .Z(n7487) );
  XNOR U11586 ( .A(b[2434]), .B(n7488), .Z(n7489) );
  XNOR U11587 ( .A(b[2434]), .B(n7490), .Z(c[2434]) );
  XOR U11588 ( .A(n7491), .B(n7492), .Z(n7488) );
  ANDN U11589 ( .B(n7493), .A(n7494), .Z(n7491) );
  XNOR U11590 ( .A(b[2433]), .B(n7492), .Z(n7493) );
  XNOR U11591 ( .A(b[2433]), .B(n7494), .Z(c[2433]) );
  XOR U11592 ( .A(n7495), .B(n7496), .Z(n7492) );
  ANDN U11593 ( .B(n7497), .A(n7498), .Z(n7495) );
  XNOR U11594 ( .A(b[2432]), .B(n7496), .Z(n7497) );
  XNOR U11595 ( .A(b[2432]), .B(n7498), .Z(c[2432]) );
  XOR U11596 ( .A(n7499), .B(n7500), .Z(n7496) );
  ANDN U11597 ( .B(n7501), .A(n7502), .Z(n7499) );
  XNOR U11598 ( .A(b[2431]), .B(n7500), .Z(n7501) );
  XNOR U11599 ( .A(b[2431]), .B(n7502), .Z(c[2431]) );
  XOR U11600 ( .A(n7503), .B(n7504), .Z(n7500) );
  ANDN U11601 ( .B(n7505), .A(n7506), .Z(n7503) );
  XNOR U11602 ( .A(b[2430]), .B(n7504), .Z(n7505) );
  XNOR U11603 ( .A(b[2430]), .B(n7506), .Z(c[2430]) );
  XOR U11604 ( .A(n7507), .B(n7508), .Z(n7504) );
  ANDN U11605 ( .B(n7509), .A(n7510), .Z(n7507) );
  XNOR U11606 ( .A(b[2429]), .B(n7508), .Z(n7509) );
  XNOR U11607 ( .A(b[242]), .B(n7511), .Z(c[242]) );
  XNOR U11608 ( .A(b[2429]), .B(n7510), .Z(c[2429]) );
  XOR U11609 ( .A(n7512), .B(n7513), .Z(n7508) );
  ANDN U11610 ( .B(n7514), .A(n7515), .Z(n7512) );
  XNOR U11611 ( .A(b[2428]), .B(n7513), .Z(n7514) );
  XNOR U11612 ( .A(b[2428]), .B(n7515), .Z(c[2428]) );
  XOR U11613 ( .A(n7516), .B(n7517), .Z(n7513) );
  ANDN U11614 ( .B(n7518), .A(n7519), .Z(n7516) );
  XNOR U11615 ( .A(b[2427]), .B(n7517), .Z(n7518) );
  XNOR U11616 ( .A(b[2427]), .B(n7519), .Z(c[2427]) );
  XOR U11617 ( .A(n7520), .B(n7521), .Z(n7517) );
  ANDN U11618 ( .B(n7522), .A(n7523), .Z(n7520) );
  XNOR U11619 ( .A(b[2426]), .B(n7521), .Z(n7522) );
  XNOR U11620 ( .A(b[2426]), .B(n7523), .Z(c[2426]) );
  XOR U11621 ( .A(n7524), .B(n7525), .Z(n7521) );
  ANDN U11622 ( .B(n7526), .A(n7527), .Z(n7524) );
  XNOR U11623 ( .A(b[2425]), .B(n7525), .Z(n7526) );
  XNOR U11624 ( .A(b[2425]), .B(n7527), .Z(c[2425]) );
  XOR U11625 ( .A(n7528), .B(n7529), .Z(n7525) );
  ANDN U11626 ( .B(n7530), .A(n7531), .Z(n7528) );
  XNOR U11627 ( .A(b[2424]), .B(n7529), .Z(n7530) );
  XNOR U11628 ( .A(b[2424]), .B(n7531), .Z(c[2424]) );
  XOR U11629 ( .A(n7532), .B(n7533), .Z(n7529) );
  ANDN U11630 ( .B(n7534), .A(n7535), .Z(n7532) );
  XNOR U11631 ( .A(b[2423]), .B(n7533), .Z(n7534) );
  XNOR U11632 ( .A(b[2423]), .B(n7535), .Z(c[2423]) );
  XOR U11633 ( .A(n7536), .B(n7537), .Z(n7533) );
  ANDN U11634 ( .B(n7538), .A(n7539), .Z(n7536) );
  XNOR U11635 ( .A(b[2422]), .B(n7537), .Z(n7538) );
  XNOR U11636 ( .A(b[2422]), .B(n7539), .Z(c[2422]) );
  XOR U11637 ( .A(n7540), .B(n7541), .Z(n7537) );
  ANDN U11638 ( .B(n7542), .A(n7543), .Z(n7540) );
  XNOR U11639 ( .A(b[2421]), .B(n7541), .Z(n7542) );
  XNOR U11640 ( .A(b[2421]), .B(n7543), .Z(c[2421]) );
  XOR U11641 ( .A(n7544), .B(n7545), .Z(n7541) );
  ANDN U11642 ( .B(n7546), .A(n7547), .Z(n7544) );
  XNOR U11643 ( .A(b[2420]), .B(n7545), .Z(n7546) );
  XNOR U11644 ( .A(b[2420]), .B(n7547), .Z(c[2420]) );
  XOR U11645 ( .A(n7548), .B(n7549), .Z(n7545) );
  ANDN U11646 ( .B(n7550), .A(n7551), .Z(n7548) );
  XNOR U11647 ( .A(b[2419]), .B(n7549), .Z(n7550) );
  XNOR U11648 ( .A(b[241]), .B(n7552), .Z(c[241]) );
  XNOR U11649 ( .A(b[2419]), .B(n7551), .Z(c[2419]) );
  XOR U11650 ( .A(n7553), .B(n7554), .Z(n7549) );
  ANDN U11651 ( .B(n7555), .A(n7556), .Z(n7553) );
  XNOR U11652 ( .A(b[2418]), .B(n7554), .Z(n7555) );
  XNOR U11653 ( .A(b[2418]), .B(n7556), .Z(c[2418]) );
  XOR U11654 ( .A(n7557), .B(n7558), .Z(n7554) );
  ANDN U11655 ( .B(n7559), .A(n7560), .Z(n7557) );
  XNOR U11656 ( .A(b[2417]), .B(n7558), .Z(n7559) );
  XNOR U11657 ( .A(b[2417]), .B(n7560), .Z(c[2417]) );
  XOR U11658 ( .A(n7561), .B(n7562), .Z(n7558) );
  ANDN U11659 ( .B(n7563), .A(n7564), .Z(n7561) );
  XNOR U11660 ( .A(b[2416]), .B(n7562), .Z(n7563) );
  XNOR U11661 ( .A(b[2416]), .B(n7564), .Z(c[2416]) );
  XOR U11662 ( .A(n7565), .B(n7566), .Z(n7562) );
  ANDN U11663 ( .B(n7567), .A(n7568), .Z(n7565) );
  XNOR U11664 ( .A(b[2415]), .B(n7566), .Z(n7567) );
  XNOR U11665 ( .A(b[2415]), .B(n7568), .Z(c[2415]) );
  XOR U11666 ( .A(n7569), .B(n7570), .Z(n7566) );
  ANDN U11667 ( .B(n7571), .A(n7572), .Z(n7569) );
  XNOR U11668 ( .A(b[2414]), .B(n7570), .Z(n7571) );
  XNOR U11669 ( .A(b[2414]), .B(n7572), .Z(c[2414]) );
  XOR U11670 ( .A(n7573), .B(n7574), .Z(n7570) );
  ANDN U11671 ( .B(n7575), .A(n7576), .Z(n7573) );
  XNOR U11672 ( .A(b[2413]), .B(n7574), .Z(n7575) );
  XNOR U11673 ( .A(b[2413]), .B(n7576), .Z(c[2413]) );
  XOR U11674 ( .A(n7577), .B(n7578), .Z(n7574) );
  ANDN U11675 ( .B(n7579), .A(n7580), .Z(n7577) );
  XNOR U11676 ( .A(b[2412]), .B(n7578), .Z(n7579) );
  XNOR U11677 ( .A(b[2412]), .B(n7580), .Z(c[2412]) );
  XOR U11678 ( .A(n7581), .B(n7582), .Z(n7578) );
  ANDN U11679 ( .B(n7583), .A(n7584), .Z(n7581) );
  XNOR U11680 ( .A(b[2411]), .B(n7582), .Z(n7583) );
  XNOR U11681 ( .A(b[2411]), .B(n7584), .Z(c[2411]) );
  XOR U11682 ( .A(n7585), .B(n7586), .Z(n7582) );
  ANDN U11683 ( .B(n7587), .A(n7588), .Z(n7585) );
  XNOR U11684 ( .A(b[2410]), .B(n7586), .Z(n7587) );
  XNOR U11685 ( .A(b[2410]), .B(n7588), .Z(c[2410]) );
  XOR U11686 ( .A(n7589), .B(n7590), .Z(n7586) );
  ANDN U11687 ( .B(n7591), .A(n7592), .Z(n7589) );
  XNOR U11688 ( .A(b[2409]), .B(n7590), .Z(n7591) );
  XNOR U11689 ( .A(b[240]), .B(n7593), .Z(c[240]) );
  XNOR U11690 ( .A(b[2409]), .B(n7592), .Z(c[2409]) );
  XOR U11691 ( .A(n7594), .B(n7595), .Z(n7590) );
  ANDN U11692 ( .B(n7596), .A(n7597), .Z(n7594) );
  XNOR U11693 ( .A(b[2408]), .B(n7595), .Z(n7596) );
  XNOR U11694 ( .A(b[2408]), .B(n7597), .Z(c[2408]) );
  XOR U11695 ( .A(n7598), .B(n7599), .Z(n7595) );
  ANDN U11696 ( .B(n7600), .A(n7601), .Z(n7598) );
  XNOR U11697 ( .A(b[2407]), .B(n7599), .Z(n7600) );
  XNOR U11698 ( .A(b[2407]), .B(n7601), .Z(c[2407]) );
  XOR U11699 ( .A(n7602), .B(n7603), .Z(n7599) );
  ANDN U11700 ( .B(n7604), .A(n7605), .Z(n7602) );
  XNOR U11701 ( .A(b[2406]), .B(n7603), .Z(n7604) );
  XNOR U11702 ( .A(b[2406]), .B(n7605), .Z(c[2406]) );
  XOR U11703 ( .A(n7606), .B(n7607), .Z(n7603) );
  ANDN U11704 ( .B(n7608), .A(n7609), .Z(n7606) );
  XNOR U11705 ( .A(b[2405]), .B(n7607), .Z(n7608) );
  XNOR U11706 ( .A(b[2405]), .B(n7609), .Z(c[2405]) );
  XOR U11707 ( .A(n7610), .B(n7611), .Z(n7607) );
  ANDN U11708 ( .B(n7612), .A(n7613), .Z(n7610) );
  XNOR U11709 ( .A(b[2404]), .B(n7611), .Z(n7612) );
  XNOR U11710 ( .A(b[2404]), .B(n7613), .Z(c[2404]) );
  XOR U11711 ( .A(n7614), .B(n7615), .Z(n7611) );
  ANDN U11712 ( .B(n7616), .A(n7617), .Z(n7614) );
  XNOR U11713 ( .A(b[2403]), .B(n7615), .Z(n7616) );
  XNOR U11714 ( .A(b[2403]), .B(n7617), .Z(c[2403]) );
  XOR U11715 ( .A(n7618), .B(n7619), .Z(n7615) );
  ANDN U11716 ( .B(n7620), .A(n7621), .Z(n7618) );
  XNOR U11717 ( .A(b[2402]), .B(n7619), .Z(n7620) );
  XNOR U11718 ( .A(b[2402]), .B(n7621), .Z(c[2402]) );
  XOR U11719 ( .A(n7622), .B(n7623), .Z(n7619) );
  ANDN U11720 ( .B(n7624), .A(n7625), .Z(n7622) );
  XNOR U11721 ( .A(b[2401]), .B(n7623), .Z(n7624) );
  XNOR U11722 ( .A(b[2401]), .B(n7625), .Z(c[2401]) );
  XOR U11723 ( .A(n7626), .B(n7627), .Z(n7623) );
  ANDN U11724 ( .B(n7628), .A(n7629), .Z(n7626) );
  XNOR U11725 ( .A(b[2400]), .B(n7627), .Z(n7628) );
  XNOR U11726 ( .A(b[2400]), .B(n7629), .Z(c[2400]) );
  XOR U11727 ( .A(n7630), .B(n7631), .Z(n7627) );
  ANDN U11728 ( .B(n7632), .A(n7633), .Z(n7630) );
  XNOR U11729 ( .A(b[2399]), .B(n7631), .Z(n7632) );
  XNOR U11730 ( .A(b[23]), .B(n7634), .Z(c[23]) );
  XNOR U11731 ( .A(b[239]), .B(n7635), .Z(c[239]) );
  XNOR U11732 ( .A(b[2399]), .B(n7633), .Z(c[2399]) );
  XOR U11733 ( .A(n7636), .B(n7637), .Z(n7631) );
  ANDN U11734 ( .B(n7638), .A(n7639), .Z(n7636) );
  XNOR U11735 ( .A(b[2398]), .B(n7637), .Z(n7638) );
  XNOR U11736 ( .A(b[2398]), .B(n7639), .Z(c[2398]) );
  XOR U11737 ( .A(n7640), .B(n7641), .Z(n7637) );
  ANDN U11738 ( .B(n7642), .A(n7643), .Z(n7640) );
  XNOR U11739 ( .A(b[2397]), .B(n7641), .Z(n7642) );
  XNOR U11740 ( .A(b[2397]), .B(n7643), .Z(c[2397]) );
  XOR U11741 ( .A(n7644), .B(n7645), .Z(n7641) );
  ANDN U11742 ( .B(n7646), .A(n7647), .Z(n7644) );
  XNOR U11743 ( .A(b[2396]), .B(n7645), .Z(n7646) );
  XNOR U11744 ( .A(b[2396]), .B(n7647), .Z(c[2396]) );
  XOR U11745 ( .A(n7648), .B(n7649), .Z(n7645) );
  ANDN U11746 ( .B(n7650), .A(n7651), .Z(n7648) );
  XNOR U11747 ( .A(b[2395]), .B(n7649), .Z(n7650) );
  XNOR U11748 ( .A(b[2395]), .B(n7651), .Z(c[2395]) );
  XOR U11749 ( .A(n7652), .B(n7653), .Z(n7649) );
  ANDN U11750 ( .B(n7654), .A(n7655), .Z(n7652) );
  XNOR U11751 ( .A(b[2394]), .B(n7653), .Z(n7654) );
  XNOR U11752 ( .A(b[2394]), .B(n7655), .Z(c[2394]) );
  XOR U11753 ( .A(n7656), .B(n7657), .Z(n7653) );
  ANDN U11754 ( .B(n7658), .A(n7659), .Z(n7656) );
  XNOR U11755 ( .A(b[2393]), .B(n7657), .Z(n7658) );
  XNOR U11756 ( .A(b[2393]), .B(n7659), .Z(c[2393]) );
  XOR U11757 ( .A(n7660), .B(n7661), .Z(n7657) );
  ANDN U11758 ( .B(n7662), .A(n7663), .Z(n7660) );
  XNOR U11759 ( .A(b[2392]), .B(n7661), .Z(n7662) );
  XNOR U11760 ( .A(b[2392]), .B(n7663), .Z(c[2392]) );
  XOR U11761 ( .A(n7664), .B(n7665), .Z(n7661) );
  ANDN U11762 ( .B(n7666), .A(n7667), .Z(n7664) );
  XNOR U11763 ( .A(b[2391]), .B(n7665), .Z(n7666) );
  XNOR U11764 ( .A(b[2391]), .B(n7667), .Z(c[2391]) );
  XOR U11765 ( .A(n7668), .B(n7669), .Z(n7665) );
  ANDN U11766 ( .B(n7670), .A(n7671), .Z(n7668) );
  XNOR U11767 ( .A(b[2390]), .B(n7669), .Z(n7670) );
  XNOR U11768 ( .A(b[2390]), .B(n7671), .Z(c[2390]) );
  XOR U11769 ( .A(n7672), .B(n7673), .Z(n7669) );
  ANDN U11770 ( .B(n7674), .A(n7675), .Z(n7672) );
  XNOR U11771 ( .A(b[2389]), .B(n7673), .Z(n7674) );
  XNOR U11772 ( .A(b[238]), .B(n7676), .Z(c[238]) );
  XNOR U11773 ( .A(b[2389]), .B(n7675), .Z(c[2389]) );
  XOR U11774 ( .A(n7677), .B(n7678), .Z(n7673) );
  ANDN U11775 ( .B(n7679), .A(n7680), .Z(n7677) );
  XNOR U11776 ( .A(b[2388]), .B(n7678), .Z(n7679) );
  XNOR U11777 ( .A(b[2388]), .B(n7680), .Z(c[2388]) );
  XOR U11778 ( .A(n7681), .B(n7682), .Z(n7678) );
  ANDN U11779 ( .B(n7683), .A(n7684), .Z(n7681) );
  XNOR U11780 ( .A(b[2387]), .B(n7682), .Z(n7683) );
  XNOR U11781 ( .A(b[2387]), .B(n7684), .Z(c[2387]) );
  XOR U11782 ( .A(n7685), .B(n7686), .Z(n7682) );
  ANDN U11783 ( .B(n7687), .A(n7688), .Z(n7685) );
  XNOR U11784 ( .A(b[2386]), .B(n7686), .Z(n7687) );
  XNOR U11785 ( .A(b[2386]), .B(n7688), .Z(c[2386]) );
  XOR U11786 ( .A(n7689), .B(n7690), .Z(n7686) );
  ANDN U11787 ( .B(n7691), .A(n7692), .Z(n7689) );
  XNOR U11788 ( .A(b[2385]), .B(n7690), .Z(n7691) );
  XNOR U11789 ( .A(b[2385]), .B(n7692), .Z(c[2385]) );
  XOR U11790 ( .A(n7693), .B(n7694), .Z(n7690) );
  ANDN U11791 ( .B(n7695), .A(n7696), .Z(n7693) );
  XNOR U11792 ( .A(b[2384]), .B(n7694), .Z(n7695) );
  XNOR U11793 ( .A(b[2384]), .B(n7696), .Z(c[2384]) );
  XOR U11794 ( .A(n7697), .B(n7698), .Z(n7694) );
  ANDN U11795 ( .B(n7699), .A(n7700), .Z(n7697) );
  XNOR U11796 ( .A(b[2383]), .B(n7698), .Z(n7699) );
  XNOR U11797 ( .A(b[2383]), .B(n7700), .Z(c[2383]) );
  XOR U11798 ( .A(n7701), .B(n7702), .Z(n7698) );
  ANDN U11799 ( .B(n7703), .A(n7704), .Z(n7701) );
  XNOR U11800 ( .A(b[2382]), .B(n7702), .Z(n7703) );
  XNOR U11801 ( .A(b[2382]), .B(n7704), .Z(c[2382]) );
  XOR U11802 ( .A(n7705), .B(n7706), .Z(n7702) );
  ANDN U11803 ( .B(n7707), .A(n7708), .Z(n7705) );
  XNOR U11804 ( .A(b[2381]), .B(n7706), .Z(n7707) );
  XNOR U11805 ( .A(b[2381]), .B(n7708), .Z(c[2381]) );
  XOR U11806 ( .A(n7709), .B(n7710), .Z(n7706) );
  ANDN U11807 ( .B(n7711), .A(n7712), .Z(n7709) );
  XNOR U11808 ( .A(b[2380]), .B(n7710), .Z(n7711) );
  XNOR U11809 ( .A(b[2380]), .B(n7712), .Z(c[2380]) );
  XOR U11810 ( .A(n7713), .B(n7714), .Z(n7710) );
  ANDN U11811 ( .B(n7715), .A(n7716), .Z(n7713) );
  XNOR U11812 ( .A(b[2379]), .B(n7714), .Z(n7715) );
  XNOR U11813 ( .A(b[237]), .B(n7717), .Z(c[237]) );
  XNOR U11814 ( .A(b[2379]), .B(n7716), .Z(c[2379]) );
  XOR U11815 ( .A(n7718), .B(n7719), .Z(n7714) );
  ANDN U11816 ( .B(n7720), .A(n7721), .Z(n7718) );
  XNOR U11817 ( .A(b[2378]), .B(n7719), .Z(n7720) );
  XNOR U11818 ( .A(b[2378]), .B(n7721), .Z(c[2378]) );
  XOR U11819 ( .A(n7722), .B(n7723), .Z(n7719) );
  ANDN U11820 ( .B(n7724), .A(n7725), .Z(n7722) );
  XNOR U11821 ( .A(b[2377]), .B(n7723), .Z(n7724) );
  XNOR U11822 ( .A(b[2377]), .B(n7725), .Z(c[2377]) );
  XOR U11823 ( .A(n7726), .B(n7727), .Z(n7723) );
  ANDN U11824 ( .B(n7728), .A(n7729), .Z(n7726) );
  XNOR U11825 ( .A(b[2376]), .B(n7727), .Z(n7728) );
  XNOR U11826 ( .A(b[2376]), .B(n7729), .Z(c[2376]) );
  XOR U11827 ( .A(n7730), .B(n7731), .Z(n7727) );
  ANDN U11828 ( .B(n7732), .A(n7733), .Z(n7730) );
  XNOR U11829 ( .A(b[2375]), .B(n7731), .Z(n7732) );
  XNOR U11830 ( .A(b[2375]), .B(n7733), .Z(c[2375]) );
  XOR U11831 ( .A(n7734), .B(n7735), .Z(n7731) );
  ANDN U11832 ( .B(n7736), .A(n7737), .Z(n7734) );
  XNOR U11833 ( .A(b[2374]), .B(n7735), .Z(n7736) );
  XNOR U11834 ( .A(b[2374]), .B(n7737), .Z(c[2374]) );
  XOR U11835 ( .A(n7738), .B(n7739), .Z(n7735) );
  ANDN U11836 ( .B(n7740), .A(n7741), .Z(n7738) );
  XNOR U11837 ( .A(b[2373]), .B(n7739), .Z(n7740) );
  XNOR U11838 ( .A(b[2373]), .B(n7741), .Z(c[2373]) );
  XOR U11839 ( .A(n7742), .B(n7743), .Z(n7739) );
  ANDN U11840 ( .B(n7744), .A(n7745), .Z(n7742) );
  XNOR U11841 ( .A(b[2372]), .B(n7743), .Z(n7744) );
  XNOR U11842 ( .A(b[2372]), .B(n7745), .Z(c[2372]) );
  XOR U11843 ( .A(n7746), .B(n7747), .Z(n7743) );
  ANDN U11844 ( .B(n7748), .A(n7749), .Z(n7746) );
  XNOR U11845 ( .A(b[2371]), .B(n7747), .Z(n7748) );
  XNOR U11846 ( .A(b[2371]), .B(n7749), .Z(c[2371]) );
  XOR U11847 ( .A(n7750), .B(n7751), .Z(n7747) );
  ANDN U11848 ( .B(n7752), .A(n7753), .Z(n7750) );
  XNOR U11849 ( .A(b[2370]), .B(n7751), .Z(n7752) );
  XNOR U11850 ( .A(b[2370]), .B(n7753), .Z(c[2370]) );
  XOR U11851 ( .A(n7754), .B(n7755), .Z(n7751) );
  ANDN U11852 ( .B(n7756), .A(n7757), .Z(n7754) );
  XNOR U11853 ( .A(b[2369]), .B(n7755), .Z(n7756) );
  XNOR U11854 ( .A(b[236]), .B(n7758), .Z(c[236]) );
  XNOR U11855 ( .A(b[2369]), .B(n7757), .Z(c[2369]) );
  XOR U11856 ( .A(n7759), .B(n7760), .Z(n7755) );
  ANDN U11857 ( .B(n7761), .A(n7762), .Z(n7759) );
  XNOR U11858 ( .A(b[2368]), .B(n7760), .Z(n7761) );
  XNOR U11859 ( .A(b[2368]), .B(n7762), .Z(c[2368]) );
  XOR U11860 ( .A(n7763), .B(n7764), .Z(n7760) );
  ANDN U11861 ( .B(n7765), .A(n7766), .Z(n7763) );
  XNOR U11862 ( .A(b[2367]), .B(n7764), .Z(n7765) );
  XNOR U11863 ( .A(b[2367]), .B(n7766), .Z(c[2367]) );
  XOR U11864 ( .A(n7767), .B(n7768), .Z(n7764) );
  ANDN U11865 ( .B(n7769), .A(n7770), .Z(n7767) );
  XNOR U11866 ( .A(b[2366]), .B(n7768), .Z(n7769) );
  XNOR U11867 ( .A(b[2366]), .B(n7770), .Z(c[2366]) );
  XOR U11868 ( .A(n7771), .B(n7772), .Z(n7768) );
  ANDN U11869 ( .B(n7773), .A(n7774), .Z(n7771) );
  XNOR U11870 ( .A(b[2365]), .B(n7772), .Z(n7773) );
  XNOR U11871 ( .A(b[2365]), .B(n7774), .Z(c[2365]) );
  XOR U11872 ( .A(n7775), .B(n7776), .Z(n7772) );
  ANDN U11873 ( .B(n7777), .A(n7778), .Z(n7775) );
  XNOR U11874 ( .A(b[2364]), .B(n7776), .Z(n7777) );
  XNOR U11875 ( .A(b[2364]), .B(n7778), .Z(c[2364]) );
  XOR U11876 ( .A(n7779), .B(n7780), .Z(n7776) );
  ANDN U11877 ( .B(n7781), .A(n7782), .Z(n7779) );
  XNOR U11878 ( .A(b[2363]), .B(n7780), .Z(n7781) );
  XNOR U11879 ( .A(b[2363]), .B(n7782), .Z(c[2363]) );
  XOR U11880 ( .A(n7783), .B(n7784), .Z(n7780) );
  ANDN U11881 ( .B(n7785), .A(n7786), .Z(n7783) );
  XNOR U11882 ( .A(b[2362]), .B(n7784), .Z(n7785) );
  XNOR U11883 ( .A(b[2362]), .B(n7786), .Z(c[2362]) );
  XOR U11884 ( .A(n7787), .B(n7788), .Z(n7784) );
  ANDN U11885 ( .B(n7789), .A(n7790), .Z(n7787) );
  XNOR U11886 ( .A(b[2361]), .B(n7788), .Z(n7789) );
  XNOR U11887 ( .A(b[2361]), .B(n7790), .Z(c[2361]) );
  XOR U11888 ( .A(n7791), .B(n7792), .Z(n7788) );
  ANDN U11889 ( .B(n7793), .A(n7794), .Z(n7791) );
  XNOR U11890 ( .A(b[2360]), .B(n7792), .Z(n7793) );
  XNOR U11891 ( .A(b[2360]), .B(n7794), .Z(c[2360]) );
  XOR U11892 ( .A(n7795), .B(n7796), .Z(n7792) );
  ANDN U11893 ( .B(n7797), .A(n7798), .Z(n7795) );
  XNOR U11894 ( .A(b[2359]), .B(n7796), .Z(n7797) );
  XNOR U11895 ( .A(b[235]), .B(n7799), .Z(c[235]) );
  XNOR U11896 ( .A(b[2359]), .B(n7798), .Z(c[2359]) );
  XOR U11897 ( .A(n7800), .B(n7801), .Z(n7796) );
  ANDN U11898 ( .B(n7802), .A(n7803), .Z(n7800) );
  XNOR U11899 ( .A(b[2358]), .B(n7801), .Z(n7802) );
  XNOR U11900 ( .A(b[2358]), .B(n7803), .Z(c[2358]) );
  XOR U11901 ( .A(n7804), .B(n7805), .Z(n7801) );
  ANDN U11902 ( .B(n7806), .A(n7807), .Z(n7804) );
  XNOR U11903 ( .A(b[2357]), .B(n7805), .Z(n7806) );
  XNOR U11904 ( .A(b[2357]), .B(n7807), .Z(c[2357]) );
  XOR U11905 ( .A(n7808), .B(n7809), .Z(n7805) );
  ANDN U11906 ( .B(n7810), .A(n7811), .Z(n7808) );
  XNOR U11907 ( .A(b[2356]), .B(n7809), .Z(n7810) );
  XNOR U11908 ( .A(b[2356]), .B(n7811), .Z(c[2356]) );
  XOR U11909 ( .A(n7812), .B(n7813), .Z(n7809) );
  ANDN U11910 ( .B(n7814), .A(n7815), .Z(n7812) );
  XNOR U11911 ( .A(b[2355]), .B(n7813), .Z(n7814) );
  XNOR U11912 ( .A(b[2355]), .B(n7815), .Z(c[2355]) );
  XOR U11913 ( .A(n7816), .B(n7817), .Z(n7813) );
  ANDN U11914 ( .B(n7818), .A(n7819), .Z(n7816) );
  XNOR U11915 ( .A(b[2354]), .B(n7817), .Z(n7818) );
  XNOR U11916 ( .A(b[2354]), .B(n7819), .Z(c[2354]) );
  XOR U11917 ( .A(n7820), .B(n7821), .Z(n7817) );
  ANDN U11918 ( .B(n7822), .A(n7823), .Z(n7820) );
  XNOR U11919 ( .A(b[2353]), .B(n7821), .Z(n7822) );
  XNOR U11920 ( .A(b[2353]), .B(n7823), .Z(c[2353]) );
  XOR U11921 ( .A(n7824), .B(n7825), .Z(n7821) );
  ANDN U11922 ( .B(n7826), .A(n7827), .Z(n7824) );
  XNOR U11923 ( .A(b[2352]), .B(n7825), .Z(n7826) );
  XNOR U11924 ( .A(b[2352]), .B(n7827), .Z(c[2352]) );
  XOR U11925 ( .A(n7828), .B(n7829), .Z(n7825) );
  ANDN U11926 ( .B(n7830), .A(n7831), .Z(n7828) );
  XNOR U11927 ( .A(b[2351]), .B(n7829), .Z(n7830) );
  XNOR U11928 ( .A(b[2351]), .B(n7831), .Z(c[2351]) );
  XOR U11929 ( .A(n7832), .B(n7833), .Z(n7829) );
  ANDN U11930 ( .B(n7834), .A(n7835), .Z(n7832) );
  XNOR U11931 ( .A(b[2350]), .B(n7833), .Z(n7834) );
  XNOR U11932 ( .A(b[2350]), .B(n7835), .Z(c[2350]) );
  XOR U11933 ( .A(n7836), .B(n7837), .Z(n7833) );
  ANDN U11934 ( .B(n7838), .A(n7839), .Z(n7836) );
  XNOR U11935 ( .A(b[2349]), .B(n7837), .Z(n7838) );
  XNOR U11936 ( .A(b[234]), .B(n7840), .Z(c[234]) );
  XNOR U11937 ( .A(b[2349]), .B(n7839), .Z(c[2349]) );
  XOR U11938 ( .A(n7841), .B(n7842), .Z(n7837) );
  ANDN U11939 ( .B(n7843), .A(n7844), .Z(n7841) );
  XNOR U11940 ( .A(b[2348]), .B(n7842), .Z(n7843) );
  XNOR U11941 ( .A(b[2348]), .B(n7844), .Z(c[2348]) );
  XOR U11942 ( .A(n7845), .B(n7846), .Z(n7842) );
  ANDN U11943 ( .B(n7847), .A(n7848), .Z(n7845) );
  XNOR U11944 ( .A(b[2347]), .B(n7846), .Z(n7847) );
  XNOR U11945 ( .A(b[2347]), .B(n7848), .Z(c[2347]) );
  XOR U11946 ( .A(n7849), .B(n7850), .Z(n7846) );
  ANDN U11947 ( .B(n7851), .A(n7852), .Z(n7849) );
  XNOR U11948 ( .A(b[2346]), .B(n7850), .Z(n7851) );
  XNOR U11949 ( .A(b[2346]), .B(n7852), .Z(c[2346]) );
  XOR U11950 ( .A(n7853), .B(n7854), .Z(n7850) );
  ANDN U11951 ( .B(n7855), .A(n7856), .Z(n7853) );
  XNOR U11952 ( .A(b[2345]), .B(n7854), .Z(n7855) );
  XNOR U11953 ( .A(b[2345]), .B(n7856), .Z(c[2345]) );
  XOR U11954 ( .A(n7857), .B(n7858), .Z(n7854) );
  ANDN U11955 ( .B(n7859), .A(n7860), .Z(n7857) );
  XNOR U11956 ( .A(b[2344]), .B(n7858), .Z(n7859) );
  XNOR U11957 ( .A(b[2344]), .B(n7860), .Z(c[2344]) );
  XOR U11958 ( .A(n7861), .B(n7862), .Z(n7858) );
  ANDN U11959 ( .B(n7863), .A(n7864), .Z(n7861) );
  XNOR U11960 ( .A(b[2343]), .B(n7862), .Z(n7863) );
  XNOR U11961 ( .A(b[2343]), .B(n7864), .Z(c[2343]) );
  XOR U11962 ( .A(n7865), .B(n7866), .Z(n7862) );
  ANDN U11963 ( .B(n7867), .A(n7868), .Z(n7865) );
  XNOR U11964 ( .A(b[2342]), .B(n7866), .Z(n7867) );
  XNOR U11965 ( .A(b[2342]), .B(n7868), .Z(c[2342]) );
  XOR U11966 ( .A(n7869), .B(n7870), .Z(n7866) );
  ANDN U11967 ( .B(n7871), .A(n7872), .Z(n7869) );
  XNOR U11968 ( .A(b[2341]), .B(n7870), .Z(n7871) );
  XNOR U11969 ( .A(b[2341]), .B(n7872), .Z(c[2341]) );
  XOR U11970 ( .A(n7873), .B(n7874), .Z(n7870) );
  ANDN U11971 ( .B(n7875), .A(n7876), .Z(n7873) );
  XNOR U11972 ( .A(b[2340]), .B(n7874), .Z(n7875) );
  XNOR U11973 ( .A(b[2340]), .B(n7876), .Z(c[2340]) );
  XOR U11974 ( .A(n7877), .B(n7878), .Z(n7874) );
  ANDN U11975 ( .B(n7879), .A(n7880), .Z(n7877) );
  XNOR U11976 ( .A(b[2339]), .B(n7878), .Z(n7879) );
  XNOR U11977 ( .A(b[233]), .B(n7881), .Z(c[233]) );
  XNOR U11978 ( .A(b[2339]), .B(n7880), .Z(c[2339]) );
  XOR U11979 ( .A(n7882), .B(n7883), .Z(n7878) );
  ANDN U11980 ( .B(n7884), .A(n7885), .Z(n7882) );
  XNOR U11981 ( .A(b[2338]), .B(n7883), .Z(n7884) );
  XNOR U11982 ( .A(b[2338]), .B(n7885), .Z(c[2338]) );
  XOR U11983 ( .A(n7886), .B(n7887), .Z(n7883) );
  ANDN U11984 ( .B(n7888), .A(n7889), .Z(n7886) );
  XNOR U11985 ( .A(b[2337]), .B(n7887), .Z(n7888) );
  XNOR U11986 ( .A(b[2337]), .B(n7889), .Z(c[2337]) );
  XOR U11987 ( .A(n7890), .B(n7891), .Z(n7887) );
  ANDN U11988 ( .B(n7892), .A(n7893), .Z(n7890) );
  XNOR U11989 ( .A(b[2336]), .B(n7891), .Z(n7892) );
  XNOR U11990 ( .A(b[2336]), .B(n7893), .Z(c[2336]) );
  XOR U11991 ( .A(n7894), .B(n7895), .Z(n7891) );
  ANDN U11992 ( .B(n7896), .A(n7897), .Z(n7894) );
  XNOR U11993 ( .A(b[2335]), .B(n7895), .Z(n7896) );
  XNOR U11994 ( .A(b[2335]), .B(n7897), .Z(c[2335]) );
  XOR U11995 ( .A(n7898), .B(n7899), .Z(n7895) );
  ANDN U11996 ( .B(n7900), .A(n7901), .Z(n7898) );
  XNOR U11997 ( .A(b[2334]), .B(n7899), .Z(n7900) );
  XNOR U11998 ( .A(b[2334]), .B(n7901), .Z(c[2334]) );
  XOR U11999 ( .A(n7902), .B(n7903), .Z(n7899) );
  ANDN U12000 ( .B(n7904), .A(n7905), .Z(n7902) );
  XNOR U12001 ( .A(b[2333]), .B(n7903), .Z(n7904) );
  XNOR U12002 ( .A(b[2333]), .B(n7905), .Z(c[2333]) );
  XOR U12003 ( .A(n7906), .B(n7907), .Z(n7903) );
  ANDN U12004 ( .B(n7908), .A(n7909), .Z(n7906) );
  XNOR U12005 ( .A(b[2332]), .B(n7907), .Z(n7908) );
  XNOR U12006 ( .A(b[2332]), .B(n7909), .Z(c[2332]) );
  XOR U12007 ( .A(n7910), .B(n7911), .Z(n7907) );
  ANDN U12008 ( .B(n7912), .A(n7913), .Z(n7910) );
  XNOR U12009 ( .A(b[2331]), .B(n7911), .Z(n7912) );
  XNOR U12010 ( .A(b[2331]), .B(n7913), .Z(c[2331]) );
  XOR U12011 ( .A(n7914), .B(n7915), .Z(n7911) );
  ANDN U12012 ( .B(n7916), .A(n7917), .Z(n7914) );
  XNOR U12013 ( .A(b[2330]), .B(n7915), .Z(n7916) );
  XNOR U12014 ( .A(b[2330]), .B(n7917), .Z(c[2330]) );
  XOR U12015 ( .A(n7918), .B(n7919), .Z(n7915) );
  ANDN U12016 ( .B(n7920), .A(n7921), .Z(n7918) );
  XNOR U12017 ( .A(b[2329]), .B(n7919), .Z(n7920) );
  XNOR U12018 ( .A(b[232]), .B(n7922), .Z(c[232]) );
  XNOR U12019 ( .A(b[2329]), .B(n7921), .Z(c[2329]) );
  XOR U12020 ( .A(n7923), .B(n7924), .Z(n7919) );
  ANDN U12021 ( .B(n7925), .A(n7926), .Z(n7923) );
  XNOR U12022 ( .A(b[2328]), .B(n7924), .Z(n7925) );
  XNOR U12023 ( .A(b[2328]), .B(n7926), .Z(c[2328]) );
  XOR U12024 ( .A(n7927), .B(n7928), .Z(n7924) );
  ANDN U12025 ( .B(n7929), .A(n7930), .Z(n7927) );
  XNOR U12026 ( .A(b[2327]), .B(n7928), .Z(n7929) );
  XNOR U12027 ( .A(b[2327]), .B(n7930), .Z(c[2327]) );
  XOR U12028 ( .A(n7931), .B(n7932), .Z(n7928) );
  ANDN U12029 ( .B(n7933), .A(n7934), .Z(n7931) );
  XNOR U12030 ( .A(b[2326]), .B(n7932), .Z(n7933) );
  XNOR U12031 ( .A(b[2326]), .B(n7934), .Z(c[2326]) );
  XOR U12032 ( .A(n7935), .B(n7936), .Z(n7932) );
  ANDN U12033 ( .B(n7937), .A(n7938), .Z(n7935) );
  XNOR U12034 ( .A(b[2325]), .B(n7936), .Z(n7937) );
  XNOR U12035 ( .A(b[2325]), .B(n7938), .Z(c[2325]) );
  XOR U12036 ( .A(n7939), .B(n7940), .Z(n7936) );
  ANDN U12037 ( .B(n7941), .A(n7942), .Z(n7939) );
  XNOR U12038 ( .A(b[2324]), .B(n7940), .Z(n7941) );
  XNOR U12039 ( .A(b[2324]), .B(n7942), .Z(c[2324]) );
  XOR U12040 ( .A(n7943), .B(n7944), .Z(n7940) );
  ANDN U12041 ( .B(n7945), .A(n7946), .Z(n7943) );
  XNOR U12042 ( .A(b[2323]), .B(n7944), .Z(n7945) );
  XNOR U12043 ( .A(b[2323]), .B(n7946), .Z(c[2323]) );
  XOR U12044 ( .A(n7947), .B(n7948), .Z(n7944) );
  ANDN U12045 ( .B(n7949), .A(n7950), .Z(n7947) );
  XNOR U12046 ( .A(b[2322]), .B(n7948), .Z(n7949) );
  XNOR U12047 ( .A(b[2322]), .B(n7950), .Z(c[2322]) );
  XOR U12048 ( .A(n7951), .B(n7952), .Z(n7948) );
  ANDN U12049 ( .B(n7953), .A(n7954), .Z(n7951) );
  XNOR U12050 ( .A(b[2321]), .B(n7952), .Z(n7953) );
  XNOR U12051 ( .A(b[2321]), .B(n7954), .Z(c[2321]) );
  XOR U12052 ( .A(n7955), .B(n7956), .Z(n7952) );
  ANDN U12053 ( .B(n7957), .A(n7958), .Z(n7955) );
  XNOR U12054 ( .A(b[2320]), .B(n7956), .Z(n7957) );
  XNOR U12055 ( .A(b[2320]), .B(n7958), .Z(c[2320]) );
  XOR U12056 ( .A(n7959), .B(n7960), .Z(n7956) );
  ANDN U12057 ( .B(n7961), .A(n7962), .Z(n7959) );
  XNOR U12058 ( .A(b[2319]), .B(n7960), .Z(n7961) );
  XNOR U12059 ( .A(b[231]), .B(n7963), .Z(c[231]) );
  XNOR U12060 ( .A(b[2319]), .B(n7962), .Z(c[2319]) );
  XOR U12061 ( .A(n7964), .B(n7965), .Z(n7960) );
  ANDN U12062 ( .B(n7966), .A(n7967), .Z(n7964) );
  XNOR U12063 ( .A(b[2318]), .B(n7965), .Z(n7966) );
  XNOR U12064 ( .A(b[2318]), .B(n7967), .Z(c[2318]) );
  XOR U12065 ( .A(n7968), .B(n7969), .Z(n7965) );
  ANDN U12066 ( .B(n7970), .A(n7971), .Z(n7968) );
  XNOR U12067 ( .A(b[2317]), .B(n7969), .Z(n7970) );
  XNOR U12068 ( .A(b[2317]), .B(n7971), .Z(c[2317]) );
  XOR U12069 ( .A(n7972), .B(n7973), .Z(n7969) );
  ANDN U12070 ( .B(n7974), .A(n7975), .Z(n7972) );
  XNOR U12071 ( .A(b[2316]), .B(n7973), .Z(n7974) );
  XNOR U12072 ( .A(b[2316]), .B(n7975), .Z(c[2316]) );
  XOR U12073 ( .A(n7976), .B(n7977), .Z(n7973) );
  ANDN U12074 ( .B(n7978), .A(n7979), .Z(n7976) );
  XNOR U12075 ( .A(b[2315]), .B(n7977), .Z(n7978) );
  XNOR U12076 ( .A(b[2315]), .B(n7979), .Z(c[2315]) );
  XOR U12077 ( .A(n7980), .B(n7981), .Z(n7977) );
  ANDN U12078 ( .B(n7982), .A(n7983), .Z(n7980) );
  XNOR U12079 ( .A(b[2314]), .B(n7981), .Z(n7982) );
  XNOR U12080 ( .A(b[2314]), .B(n7983), .Z(c[2314]) );
  XOR U12081 ( .A(n7984), .B(n7985), .Z(n7981) );
  ANDN U12082 ( .B(n7986), .A(n7987), .Z(n7984) );
  XNOR U12083 ( .A(b[2313]), .B(n7985), .Z(n7986) );
  XNOR U12084 ( .A(b[2313]), .B(n7987), .Z(c[2313]) );
  XOR U12085 ( .A(n7988), .B(n7989), .Z(n7985) );
  ANDN U12086 ( .B(n7990), .A(n7991), .Z(n7988) );
  XNOR U12087 ( .A(b[2312]), .B(n7989), .Z(n7990) );
  XNOR U12088 ( .A(b[2312]), .B(n7991), .Z(c[2312]) );
  XOR U12089 ( .A(n7992), .B(n7993), .Z(n7989) );
  ANDN U12090 ( .B(n7994), .A(n7995), .Z(n7992) );
  XNOR U12091 ( .A(b[2311]), .B(n7993), .Z(n7994) );
  XNOR U12092 ( .A(b[2311]), .B(n7995), .Z(c[2311]) );
  XOR U12093 ( .A(n7996), .B(n7997), .Z(n7993) );
  ANDN U12094 ( .B(n7998), .A(n7999), .Z(n7996) );
  XNOR U12095 ( .A(b[2310]), .B(n7997), .Z(n7998) );
  XNOR U12096 ( .A(b[2310]), .B(n7999), .Z(c[2310]) );
  XOR U12097 ( .A(n8000), .B(n8001), .Z(n7997) );
  ANDN U12098 ( .B(n8002), .A(n8003), .Z(n8000) );
  XNOR U12099 ( .A(b[2309]), .B(n8001), .Z(n8002) );
  XNOR U12100 ( .A(b[230]), .B(n8004), .Z(c[230]) );
  XNOR U12101 ( .A(b[2309]), .B(n8003), .Z(c[2309]) );
  XOR U12102 ( .A(n8005), .B(n8006), .Z(n8001) );
  ANDN U12103 ( .B(n8007), .A(n8008), .Z(n8005) );
  XNOR U12104 ( .A(b[2308]), .B(n8006), .Z(n8007) );
  XNOR U12105 ( .A(b[2308]), .B(n8008), .Z(c[2308]) );
  XOR U12106 ( .A(n8009), .B(n8010), .Z(n8006) );
  ANDN U12107 ( .B(n8011), .A(n8012), .Z(n8009) );
  XNOR U12108 ( .A(b[2307]), .B(n8010), .Z(n8011) );
  XNOR U12109 ( .A(b[2307]), .B(n8012), .Z(c[2307]) );
  XOR U12110 ( .A(n8013), .B(n8014), .Z(n8010) );
  ANDN U12111 ( .B(n8015), .A(n8016), .Z(n8013) );
  XNOR U12112 ( .A(b[2306]), .B(n8014), .Z(n8015) );
  XNOR U12113 ( .A(b[2306]), .B(n8016), .Z(c[2306]) );
  XOR U12114 ( .A(n8017), .B(n8018), .Z(n8014) );
  ANDN U12115 ( .B(n8019), .A(n8020), .Z(n8017) );
  XNOR U12116 ( .A(b[2305]), .B(n8018), .Z(n8019) );
  XNOR U12117 ( .A(b[2305]), .B(n8020), .Z(c[2305]) );
  XOR U12118 ( .A(n8021), .B(n8022), .Z(n8018) );
  ANDN U12119 ( .B(n8023), .A(n8024), .Z(n8021) );
  XNOR U12120 ( .A(b[2304]), .B(n8022), .Z(n8023) );
  XNOR U12121 ( .A(b[2304]), .B(n8024), .Z(c[2304]) );
  XOR U12122 ( .A(n8025), .B(n8026), .Z(n8022) );
  ANDN U12123 ( .B(n8027), .A(n8028), .Z(n8025) );
  XNOR U12124 ( .A(b[2303]), .B(n8026), .Z(n8027) );
  XNOR U12125 ( .A(b[2303]), .B(n8028), .Z(c[2303]) );
  XOR U12126 ( .A(n8029), .B(n8030), .Z(n8026) );
  ANDN U12127 ( .B(n8031), .A(n8032), .Z(n8029) );
  XNOR U12128 ( .A(b[2302]), .B(n8030), .Z(n8031) );
  XNOR U12129 ( .A(b[2302]), .B(n8032), .Z(c[2302]) );
  XOR U12130 ( .A(n8033), .B(n8034), .Z(n8030) );
  ANDN U12131 ( .B(n8035), .A(n8036), .Z(n8033) );
  XNOR U12132 ( .A(b[2301]), .B(n8034), .Z(n8035) );
  XNOR U12133 ( .A(b[2301]), .B(n8036), .Z(c[2301]) );
  XOR U12134 ( .A(n8037), .B(n8038), .Z(n8034) );
  ANDN U12135 ( .B(n8039), .A(n8040), .Z(n8037) );
  XNOR U12136 ( .A(b[2300]), .B(n8038), .Z(n8039) );
  XNOR U12137 ( .A(b[2300]), .B(n8040), .Z(c[2300]) );
  XOR U12138 ( .A(n8041), .B(n8042), .Z(n8038) );
  ANDN U12139 ( .B(n8043), .A(n8044), .Z(n8041) );
  XNOR U12140 ( .A(b[2299]), .B(n8042), .Z(n8043) );
  XNOR U12141 ( .A(b[22]), .B(n8045), .Z(c[22]) );
  XNOR U12142 ( .A(b[229]), .B(n8046), .Z(c[229]) );
  XNOR U12143 ( .A(b[2299]), .B(n8044), .Z(c[2299]) );
  XOR U12144 ( .A(n8047), .B(n8048), .Z(n8042) );
  ANDN U12145 ( .B(n8049), .A(n8050), .Z(n8047) );
  XNOR U12146 ( .A(b[2298]), .B(n8048), .Z(n8049) );
  XNOR U12147 ( .A(b[2298]), .B(n8050), .Z(c[2298]) );
  XOR U12148 ( .A(n8051), .B(n8052), .Z(n8048) );
  ANDN U12149 ( .B(n8053), .A(n8054), .Z(n8051) );
  XNOR U12150 ( .A(b[2297]), .B(n8052), .Z(n8053) );
  XNOR U12151 ( .A(b[2297]), .B(n8054), .Z(c[2297]) );
  XOR U12152 ( .A(n8055), .B(n8056), .Z(n8052) );
  ANDN U12153 ( .B(n8057), .A(n8058), .Z(n8055) );
  XNOR U12154 ( .A(b[2296]), .B(n8056), .Z(n8057) );
  XNOR U12155 ( .A(b[2296]), .B(n8058), .Z(c[2296]) );
  XOR U12156 ( .A(n8059), .B(n8060), .Z(n8056) );
  ANDN U12157 ( .B(n8061), .A(n8062), .Z(n8059) );
  XNOR U12158 ( .A(b[2295]), .B(n8060), .Z(n8061) );
  XNOR U12159 ( .A(b[2295]), .B(n8062), .Z(c[2295]) );
  XOR U12160 ( .A(n8063), .B(n8064), .Z(n8060) );
  ANDN U12161 ( .B(n8065), .A(n8066), .Z(n8063) );
  XNOR U12162 ( .A(b[2294]), .B(n8064), .Z(n8065) );
  XNOR U12163 ( .A(b[2294]), .B(n8066), .Z(c[2294]) );
  XOR U12164 ( .A(n8067), .B(n8068), .Z(n8064) );
  ANDN U12165 ( .B(n8069), .A(n8070), .Z(n8067) );
  XNOR U12166 ( .A(b[2293]), .B(n8068), .Z(n8069) );
  XNOR U12167 ( .A(b[2293]), .B(n8070), .Z(c[2293]) );
  XOR U12168 ( .A(n8071), .B(n8072), .Z(n8068) );
  ANDN U12169 ( .B(n8073), .A(n8074), .Z(n8071) );
  XNOR U12170 ( .A(b[2292]), .B(n8072), .Z(n8073) );
  XNOR U12171 ( .A(b[2292]), .B(n8074), .Z(c[2292]) );
  XOR U12172 ( .A(n8075), .B(n8076), .Z(n8072) );
  ANDN U12173 ( .B(n8077), .A(n8078), .Z(n8075) );
  XNOR U12174 ( .A(b[2291]), .B(n8076), .Z(n8077) );
  XNOR U12175 ( .A(b[2291]), .B(n8078), .Z(c[2291]) );
  XOR U12176 ( .A(n8079), .B(n8080), .Z(n8076) );
  ANDN U12177 ( .B(n8081), .A(n8082), .Z(n8079) );
  XNOR U12178 ( .A(b[2290]), .B(n8080), .Z(n8081) );
  XNOR U12179 ( .A(b[2290]), .B(n8082), .Z(c[2290]) );
  XOR U12180 ( .A(n8083), .B(n8084), .Z(n8080) );
  ANDN U12181 ( .B(n8085), .A(n8086), .Z(n8083) );
  XNOR U12182 ( .A(b[2289]), .B(n8084), .Z(n8085) );
  XNOR U12183 ( .A(b[228]), .B(n8087), .Z(c[228]) );
  XNOR U12184 ( .A(b[2289]), .B(n8086), .Z(c[2289]) );
  XOR U12185 ( .A(n8088), .B(n8089), .Z(n8084) );
  ANDN U12186 ( .B(n8090), .A(n8091), .Z(n8088) );
  XNOR U12187 ( .A(b[2288]), .B(n8089), .Z(n8090) );
  XNOR U12188 ( .A(b[2288]), .B(n8091), .Z(c[2288]) );
  XOR U12189 ( .A(n8092), .B(n8093), .Z(n8089) );
  ANDN U12190 ( .B(n8094), .A(n8095), .Z(n8092) );
  XNOR U12191 ( .A(b[2287]), .B(n8093), .Z(n8094) );
  XNOR U12192 ( .A(b[2287]), .B(n8095), .Z(c[2287]) );
  XOR U12193 ( .A(n8096), .B(n8097), .Z(n8093) );
  ANDN U12194 ( .B(n8098), .A(n8099), .Z(n8096) );
  XNOR U12195 ( .A(b[2286]), .B(n8097), .Z(n8098) );
  XNOR U12196 ( .A(b[2286]), .B(n8099), .Z(c[2286]) );
  XOR U12197 ( .A(n8100), .B(n8101), .Z(n8097) );
  ANDN U12198 ( .B(n8102), .A(n8103), .Z(n8100) );
  XNOR U12199 ( .A(b[2285]), .B(n8101), .Z(n8102) );
  XNOR U12200 ( .A(b[2285]), .B(n8103), .Z(c[2285]) );
  XOR U12201 ( .A(n8104), .B(n8105), .Z(n8101) );
  ANDN U12202 ( .B(n8106), .A(n8107), .Z(n8104) );
  XNOR U12203 ( .A(b[2284]), .B(n8105), .Z(n8106) );
  XNOR U12204 ( .A(b[2284]), .B(n8107), .Z(c[2284]) );
  XOR U12205 ( .A(n8108), .B(n8109), .Z(n8105) );
  ANDN U12206 ( .B(n8110), .A(n8111), .Z(n8108) );
  XNOR U12207 ( .A(b[2283]), .B(n8109), .Z(n8110) );
  XNOR U12208 ( .A(b[2283]), .B(n8111), .Z(c[2283]) );
  XOR U12209 ( .A(n8112), .B(n8113), .Z(n8109) );
  ANDN U12210 ( .B(n8114), .A(n8115), .Z(n8112) );
  XNOR U12211 ( .A(b[2282]), .B(n8113), .Z(n8114) );
  XNOR U12212 ( .A(b[2282]), .B(n8115), .Z(c[2282]) );
  XOR U12213 ( .A(n8116), .B(n8117), .Z(n8113) );
  ANDN U12214 ( .B(n8118), .A(n8119), .Z(n8116) );
  XNOR U12215 ( .A(b[2281]), .B(n8117), .Z(n8118) );
  XNOR U12216 ( .A(b[2281]), .B(n8119), .Z(c[2281]) );
  XOR U12217 ( .A(n8120), .B(n8121), .Z(n8117) );
  ANDN U12218 ( .B(n8122), .A(n8123), .Z(n8120) );
  XNOR U12219 ( .A(b[2280]), .B(n8121), .Z(n8122) );
  XNOR U12220 ( .A(b[2280]), .B(n8123), .Z(c[2280]) );
  XOR U12221 ( .A(n8124), .B(n8125), .Z(n8121) );
  ANDN U12222 ( .B(n8126), .A(n8127), .Z(n8124) );
  XNOR U12223 ( .A(b[2279]), .B(n8125), .Z(n8126) );
  XNOR U12224 ( .A(b[227]), .B(n8128), .Z(c[227]) );
  XNOR U12225 ( .A(b[2279]), .B(n8127), .Z(c[2279]) );
  XOR U12226 ( .A(n8129), .B(n8130), .Z(n8125) );
  ANDN U12227 ( .B(n8131), .A(n8132), .Z(n8129) );
  XNOR U12228 ( .A(b[2278]), .B(n8130), .Z(n8131) );
  XNOR U12229 ( .A(b[2278]), .B(n8132), .Z(c[2278]) );
  XOR U12230 ( .A(n8133), .B(n8134), .Z(n8130) );
  ANDN U12231 ( .B(n8135), .A(n8136), .Z(n8133) );
  XNOR U12232 ( .A(b[2277]), .B(n8134), .Z(n8135) );
  XNOR U12233 ( .A(b[2277]), .B(n8136), .Z(c[2277]) );
  XOR U12234 ( .A(n8137), .B(n8138), .Z(n8134) );
  ANDN U12235 ( .B(n8139), .A(n8140), .Z(n8137) );
  XNOR U12236 ( .A(b[2276]), .B(n8138), .Z(n8139) );
  XNOR U12237 ( .A(b[2276]), .B(n8140), .Z(c[2276]) );
  XOR U12238 ( .A(n8141), .B(n8142), .Z(n8138) );
  ANDN U12239 ( .B(n8143), .A(n8144), .Z(n8141) );
  XNOR U12240 ( .A(b[2275]), .B(n8142), .Z(n8143) );
  XNOR U12241 ( .A(b[2275]), .B(n8144), .Z(c[2275]) );
  XOR U12242 ( .A(n8145), .B(n8146), .Z(n8142) );
  ANDN U12243 ( .B(n8147), .A(n8148), .Z(n8145) );
  XNOR U12244 ( .A(b[2274]), .B(n8146), .Z(n8147) );
  XNOR U12245 ( .A(b[2274]), .B(n8148), .Z(c[2274]) );
  XOR U12246 ( .A(n8149), .B(n8150), .Z(n8146) );
  ANDN U12247 ( .B(n8151), .A(n8152), .Z(n8149) );
  XNOR U12248 ( .A(b[2273]), .B(n8150), .Z(n8151) );
  XNOR U12249 ( .A(b[2273]), .B(n8152), .Z(c[2273]) );
  XOR U12250 ( .A(n8153), .B(n8154), .Z(n8150) );
  ANDN U12251 ( .B(n8155), .A(n8156), .Z(n8153) );
  XNOR U12252 ( .A(b[2272]), .B(n8154), .Z(n8155) );
  XNOR U12253 ( .A(b[2272]), .B(n8156), .Z(c[2272]) );
  XOR U12254 ( .A(n8157), .B(n8158), .Z(n8154) );
  ANDN U12255 ( .B(n8159), .A(n8160), .Z(n8157) );
  XNOR U12256 ( .A(b[2271]), .B(n8158), .Z(n8159) );
  XNOR U12257 ( .A(b[2271]), .B(n8160), .Z(c[2271]) );
  XOR U12258 ( .A(n8161), .B(n8162), .Z(n8158) );
  ANDN U12259 ( .B(n8163), .A(n8164), .Z(n8161) );
  XNOR U12260 ( .A(b[2270]), .B(n8162), .Z(n8163) );
  XNOR U12261 ( .A(b[2270]), .B(n8164), .Z(c[2270]) );
  XOR U12262 ( .A(n8165), .B(n8166), .Z(n8162) );
  ANDN U12263 ( .B(n8167), .A(n8168), .Z(n8165) );
  XNOR U12264 ( .A(b[2269]), .B(n8166), .Z(n8167) );
  XNOR U12265 ( .A(b[226]), .B(n8169), .Z(c[226]) );
  XNOR U12266 ( .A(b[2269]), .B(n8168), .Z(c[2269]) );
  XOR U12267 ( .A(n8170), .B(n8171), .Z(n8166) );
  ANDN U12268 ( .B(n8172), .A(n8173), .Z(n8170) );
  XNOR U12269 ( .A(b[2268]), .B(n8171), .Z(n8172) );
  XNOR U12270 ( .A(b[2268]), .B(n8173), .Z(c[2268]) );
  XOR U12271 ( .A(n8174), .B(n8175), .Z(n8171) );
  ANDN U12272 ( .B(n8176), .A(n8177), .Z(n8174) );
  XNOR U12273 ( .A(b[2267]), .B(n8175), .Z(n8176) );
  XNOR U12274 ( .A(b[2267]), .B(n8177), .Z(c[2267]) );
  XOR U12275 ( .A(n8178), .B(n8179), .Z(n8175) );
  ANDN U12276 ( .B(n8180), .A(n8181), .Z(n8178) );
  XNOR U12277 ( .A(b[2266]), .B(n8179), .Z(n8180) );
  XNOR U12278 ( .A(b[2266]), .B(n8181), .Z(c[2266]) );
  XOR U12279 ( .A(n8182), .B(n8183), .Z(n8179) );
  ANDN U12280 ( .B(n8184), .A(n8185), .Z(n8182) );
  XNOR U12281 ( .A(b[2265]), .B(n8183), .Z(n8184) );
  XNOR U12282 ( .A(b[2265]), .B(n8185), .Z(c[2265]) );
  XOR U12283 ( .A(n8186), .B(n8187), .Z(n8183) );
  ANDN U12284 ( .B(n8188), .A(n8189), .Z(n8186) );
  XNOR U12285 ( .A(b[2264]), .B(n8187), .Z(n8188) );
  XNOR U12286 ( .A(b[2264]), .B(n8189), .Z(c[2264]) );
  XOR U12287 ( .A(n8190), .B(n8191), .Z(n8187) );
  ANDN U12288 ( .B(n8192), .A(n8193), .Z(n8190) );
  XNOR U12289 ( .A(b[2263]), .B(n8191), .Z(n8192) );
  XNOR U12290 ( .A(b[2263]), .B(n8193), .Z(c[2263]) );
  XOR U12291 ( .A(n8194), .B(n8195), .Z(n8191) );
  ANDN U12292 ( .B(n8196), .A(n8197), .Z(n8194) );
  XNOR U12293 ( .A(b[2262]), .B(n8195), .Z(n8196) );
  XNOR U12294 ( .A(b[2262]), .B(n8197), .Z(c[2262]) );
  XOR U12295 ( .A(n8198), .B(n8199), .Z(n8195) );
  ANDN U12296 ( .B(n8200), .A(n8201), .Z(n8198) );
  XNOR U12297 ( .A(b[2261]), .B(n8199), .Z(n8200) );
  XNOR U12298 ( .A(b[2261]), .B(n8201), .Z(c[2261]) );
  XOR U12299 ( .A(n8202), .B(n8203), .Z(n8199) );
  ANDN U12300 ( .B(n8204), .A(n8205), .Z(n8202) );
  XNOR U12301 ( .A(b[2260]), .B(n8203), .Z(n8204) );
  XNOR U12302 ( .A(b[2260]), .B(n8205), .Z(c[2260]) );
  XOR U12303 ( .A(n8206), .B(n8207), .Z(n8203) );
  ANDN U12304 ( .B(n8208), .A(n8209), .Z(n8206) );
  XNOR U12305 ( .A(b[2259]), .B(n8207), .Z(n8208) );
  XNOR U12306 ( .A(b[225]), .B(n8210), .Z(c[225]) );
  XNOR U12307 ( .A(b[2259]), .B(n8209), .Z(c[2259]) );
  XOR U12308 ( .A(n8211), .B(n8212), .Z(n8207) );
  ANDN U12309 ( .B(n8213), .A(n8214), .Z(n8211) );
  XNOR U12310 ( .A(b[2258]), .B(n8212), .Z(n8213) );
  XNOR U12311 ( .A(b[2258]), .B(n8214), .Z(c[2258]) );
  XOR U12312 ( .A(n8215), .B(n8216), .Z(n8212) );
  ANDN U12313 ( .B(n8217), .A(n8218), .Z(n8215) );
  XNOR U12314 ( .A(b[2257]), .B(n8216), .Z(n8217) );
  XNOR U12315 ( .A(b[2257]), .B(n8218), .Z(c[2257]) );
  XOR U12316 ( .A(n8219), .B(n8220), .Z(n8216) );
  ANDN U12317 ( .B(n8221), .A(n8222), .Z(n8219) );
  XNOR U12318 ( .A(b[2256]), .B(n8220), .Z(n8221) );
  XNOR U12319 ( .A(b[2256]), .B(n8222), .Z(c[2256]) );
  XOR U12320 ( .A(n8223), .B(n8224), .Z(n8220) );
  ANDN U12321 ( .B(n8225), .A(n8226), .Z(n8223) );
  XNOR U12322 ( .A(b[2255]), .B(n8224), .Z(n8225) );
  XNOR U12323 ( .A(b[2255]), .B(n8226), .Z(c[2255]) );
  XOR U12324 ( .A(n8227), .B(n8228), .Z(n8224) );
  ANDN U12325 ( .B(n8229), .A(n8230), .Z(n8227) );
  XNOR U12326 ( .A(b[2254]), .B(n8228), .Z(n8229) );
  XNOR U12327 ( .A(b[2254]), .B(n8230), .Z(c[2254]) );
  XOR U12328 ( .A(n8231), .B(n8232), .Z(n8228) );
  ANDN U12329 ( .B(n8233), .A(n8234), .Z(n8231) );
  XNOR U12330 ( .A(b[2253]), .B(n8232), .Z(n8233) );
  XNOR U12331 ( .A(b[2253]), .B(n8234), .Z(c[2253]) );
  XOR U12332 ( .A(n8235), .B(n8236), .Z(n8232) );
  ANDN U12333 ( .B(n8237), .A(n8238), .Z(n8235) );
  XNOR U12334 ( .A(b[2252]), .B(n8236), .Z(n8237) );
  XNOR U12335 ( .A(b[2252]), .B(n8238), .Z(c[2252]) );
  XOR U12336 ( .A(n8239), .B(n8240), .Z(n8236) );
  ANDN U12337 ( .B(n8241), .A(n8242), .Z(n8239) );
  XNOR U12338 ( .A(b[2251]), .B(n8240), .Z(n8241) );
  XNOR U12339 ( .A(b[2251]), .B(n8242), .Z(c[2251]) );
  XOR U12340 ( .A(n8243), .B(n8244), .Z(n8240) );
  ANDN U12341 ( .B(n8245), .A(n8246), .Z(n8243) );
  XNOR U12342 ( .A(b[2250]), .B(n8244), .Z(n8245) );
  XNOR U12343 ( .A(b[2250]), .B(n8246), .Z(c[2250]) );
  XOR U12344 ( .A(n8247), .B(n8248), .Z(n8244) );
  ANDN U12345 ( .B(n8249), .A(n8250), .Z(n8247) );
  XNOR U12346 ( .A(b[2249]), .B(n8248), .Z(n8249) );
  XNOR U12347 ( .A(b[224]), .B(n8251), .Z(c[224]) );
  XNOR U12348 ( .A(b[2249]), .B(n8250), .Z(c[2249]) );
  XOR U12349 ( .A(n8252), .B(n8253), .Z(n8248) );
  ANDN U12350 ( .B(n8254), .A(n8255), .Z(n8252) );
  XNOR U12351 ( .A(b[2248]), .B(n8253), .Z(n8254) );
  XNOR U12352 ( .A(b[2248]), .B(n8255), .Z(c[2248]) );
  XOR U12353 ( .A(n8256), .B(n8257), .Z(n8253) );
  ANDN U12354 ( .B(n8258), .A(n8259), .Z(n8256) );
  XNOR U12355 ( .A(b[2247]), .B(n8257), .Z(n8258) );
  XNOR U12356 ( .A(b[2247]), .B(n8259), .Z(c[2247]) );
  XOR U12357 ( .A(n8260), .B(n8261), .Z(n8257) );
  ANDN U12358 ( .B(n8262), .A(n8263), .Z(n8260) );
  XNOR U12359 ( .A(b[2246]), .B(n8261), .Z(n8262) );
  XNOR U12360 ( .A(b[2246]), .B(n8263), .Z(c[2246]) );
  XOR U12361 ( .A(n8264), .B(n8265), .Z(n8261) );
  ANDN U12362 ( .B(n8266), .A(n8267), .Z(n8264) );
  XNOR U12363 ( .A(b[2245]), .B(n8265), .Z(n8266) );
  XNOR U12364 ( .A(b[2245]), .B(n8267), .Z(c[2245]) );
  XOR U12365 ( .A(n8268), .B(n8269), .Z(n8265) );
  ANDN U12366 ( .B(n8270), .A(n8271), .Z(n8268) );
  XNOR U12367 ( .A(b[2244]), .B(n8269), .Z(n8270) );
  XNOR U12368 ( .A(b[2244]), .B(n8271), .Z(c[2244]) );
  XOR U12369 ( .A(n8272), .B(n8273), .Z(n8269) );
  ANDN U12370 ( .B(n8274), .A(n8275), .Z(n8272) );
  XNOR U12371 ( .A(b[2243]), .B(n8273), .Z(n8274) );
  XNOR U12372 ( .A(b[2243]), .B(n8275), .Z(c[2243]) );
  XOR U12373 ( .A(n8276), .B(n8277), .Z(n8273) );
  ANDN U12374 ( .B(n8278), .A(n8279), .Z(n8276) );
  XNOR U12375 ( .A(b[2242]), .B(n8277), .Z(n8278) );
  XNOR U12376 ( .A(b[2242]), .B(n8279), .Z(c[2242]) );
  XOR U12377 ( .A(n8280), .B(n8281), .Z(n8277) );
  ANDN U12378 ( .B(n8282), .A(n8283), .Z(n8280) );
  XNOR U12379 ( .A(b[2241]), .B(n8281), .Z(n8282) );
  XNOR U12380 ( .A(b[2241]), .B(n8283), .Z(c[2241]) );
  XOR U12381 ( .A(n8284), .B(n8285), .Z(n8281) );
  ANDN U12382 ( .B(n8286), .A(n8287), .Z(n8284) );
  XNOR U12383 ( .A(b[2240]), .B(n8285), .Z(n8286) );
  XNOR U12384 ( .A(b[2240]), .B(n8287), .Z(c[2240]) );
  XOR U12385 ( .A(n8288), .B(n8289), .Z(n8285) );
  ANDN U12386 ( .B(n8290), .A(n8291), .Z(n8288) );
  XNOR U12387 ( .A(b[2239]), .B(n8289), .Z(n8290) );
  XNOR U12388 ( .A(b[223]), .B(n8292), .Z(c[223]) );
  XNOR U12389 ( .A(b[2239]), .B(n8291), .Z(c[2239]) );
  XOR U12390 ( .A(n8293), .B(n8294), .Z(n8289) );
  ANDN U12391 ( .B(n8295), .A(n8296), .Z(n8293) );
  XNOR U12392 ( .A(b[2238]), .B(n8294), .Z(n8295) );
  XNOR U12393 ( .A(b[2238]), .B(n8296), .Z(c[2238]) );
  XOR U12394 ( .A(n8297), .B(n8298), .Z(n8294) );
  ANDN U12395 ( .B(n8299), .A(n8300), .Z(n8297) );
  XNOR U12396 ( .A(b[2237]), .B(n8298), .Z(n8299) );
  XNOR U12397 ( .A(b[2237]), .B(n8300), .Z(c[2237]) );
  XOR U12398 ( .A(n8301), .B(n8302), .Z(n8298) );
  ANDN U12399 ( .B(n8303), .A(n8304), .Z(n8301) );
  XNOR U12400 ( .A(b[2236]), .B(n8302), .Z(n8303) );
  XNOR U12401 ( .A(b[2236]), .B(n8304), .Z(c[2236]) );
  XOR U12402 ( .A(n8305), .B(n8306), .Z(n8302) );
  ANDN U12403 ( .B(n8307), .A(n8308), .Z(n8305) );
  XNOR U12404 ( .A(b[2235]), .B(n8306), .Z(n8307) );
  XNOR U12405 ( .A(b[2235]), .B(n8308), .Z(c[2235]) );
  XOR U12406 ( .A(n8309), .B(n8310), .Z(n8306) );
  ANDN U12407 ( .B(n8311), .A(n8312), .Z(n8309) );
  XNOR U12408 ( .A(b[2234]), .B(n8310), .Z(n8311) );
  XNOR U12409 ( .A(b[2234]), .B(n8312), .Z(c[2234]) );
  XOR U12410 ( .A(n8313), .B(n8314), .Z(n8310) );
  ANDN U12411 ( .B(n8315), .A(n8316), .Z(n8313) );
  XNOR U12412 ( .A(b[2233]), .B(n8314), .Z(n8315) );
  XNOR U12413 ( .A(b[2233]), .B(n8316), .Z(c[2233]) );
  XOR U12414 ( .A(n8317), .B(n8318), .Z(n8314) );
  ANDN U12415 ( .B(n8319), .A(n8320), .Z(n8317) );
  XNOR U12416 ( .A(b[2232]), .B(n8318), .Z(n8319) );
  XNOR U12417 ( .A(b[2232]), .B(n8320), .Z(c[2232]) );
  XOR U12418 ( .A(n8321), .B(n8322), .Z(n8318) );
  ANDN U12419 ( .B(n8323), .A(n8324), .Z(n8321) );
  XNOR U12420 ( .A(b[2231]), .B(n8322), .Z(n8323) );
  XNOR U12421 ( .A(b[2231]), .B(n8324), .Z(c[2231]) );
  XOR U12422 ( .A(n8325), .B(n8326), .Z(n8322) );
  ANDN U12423 ( .B(n8327), .A(n8328), .Z(n8325) );
  XNOR U12424 ( .A(b[2230]), .B(n8326), .Z(n8327) );
  XNOR U12425 ( .A(b[2230]), .B(n8328), .Z(c[2230]) );
  XOR U12426 ( .A(n8329), .B(n8330), .Z(n8326) );
  ANDN U12427 ( .B(n8331), .A(n8332), .Z(n8329) );
  XNOR U12428 ( .A(b[2229]), .B(n8330), .Z(n8331) );
  XNOR U12429 ( .A(b[222]), .B(n8333), .Z(c[222]) );
  XNOR U12430 ( .A(b[2229]), .B(n8332), .Z(c[2229]) );
  XOR U12431 ( .A(n8334), .B(n8335), .Z(n8330) );
  ANDN U12432 ( .B(n8336), .A(n8337), .Z(n8334) );
  XNOR U12433 ( .A(b[2228]), .B(n8335), .Z(n8336) );
  XNOR U12434 ( .A(b[2228]), .B(n8337), .Z(c[2228]) );
  XOR U12435 ( .A(n8338), .B(n8339), .Z(n8335) );
  ANDN U12436 ( .B(n8340), .A(n8341), .Z(n8338) );
  XNOR U12437 ( .A(b[2227]), .B(n8339), .Z(n8340) );
  XNOR U12438 ( .A(b[2227]), .B(n8341), .Z(c[2227]) );
  XOR U12439 ( .A(n8342), .B(n8343), .Z(n8339) );
  ANDN U12440 ( .B(n8344), .A(n8345), .Z(n8342) );
  XNOR U12441 ( .A(b[2226]), .B(n8343), .Z(n8344) );
  XNOR U12442 ( .A(b[2226]), .B(n8345), .Z(c[2226]) );
  XOR U12443 ( .A(n8346), .B(n8347), .Z(n8343) );
  ANDN U12444 ( .B(n8348), .A(n8349), .Z(n8346) );
  XNOR U12445 ( .A(b[2225]), .B(n8347), .Z(n8348) );
  XNOR U12446 ( .A(b[2225]), .B(n8349), .Z(c[2225]) );
  XOR U12447 ( .A(n8350), .B(n8351), .Z(n8347) );
  ANDN U12448 ( .B(n8352), .A(n8353), .Z(n8350) );
  XNOR U12449 ( .A(b[2224]), .B(n8351), .Z(n8352) );
  XNOR U12450 ( .A(b[2224]), .B(n8353), .Z(c[2224]) );
  XOR U12451 ( .A(n8354), .B(n8355), .Z(n8351) );
  ANDN U12452 ( .B(n8356), .A(n8357), .Z(n8354) );
  XNOR U12453 ( .A(b[2223]), .B(n8355), .Z(n8356) );
  XNOR U12454 ( .A(b[2223]), .B(n8357), .Z(c[2223]) );
  XOR U12455 ( .A(n8358), .B(n8359), .Z(n8355) );
  ANDN U12456 ( .B(n8360), .A(n8361), .Z(n8358) );
  XNOR U12457 ( .A(b[2222]), .B(n8359), .Z(n8360) );
  XNOR U12458 ( .A(b[2222]), .B(n8361), .Z(c[2222]) );
  XOR U12459 ( .A(n8362), .B(n8363), .Z(n8359) );
  ANDN U12460 ( .B(n8364), .A(n8365), .Z(n8362) );
  XNOR U12461 ( .A(b[2221]), .B(n8363), .Z(n8364) );
  XNOR U12462 ( .A(b[2221]), .B(n8365), .Z(c[2221]) );
  XOR U12463 ( .A(n8366), .B(n8367), .Z(n8363) );
  ANDN U12464 ( .B(n8368), .A(n8369), .Z(n8366) );
  XNOR U12465 ( .A(b[2220]), .B(n8367), .Z(n8368) );
  XNOR U12466 ( .A(b[2220]), .B(n8369), .Z(c[2220]) );
  XOR U12467 ( .A(n8370), .B(n8371), .Z(n8367) );
  ANDN U12468 ( .B(n8372), .A(n8373), .Z(n8370) );
  XNOR U12469 ( .A(b[2219]), .B(n8371), .Z(n8372) );
  XNOR U12470 ( .A(b[221]), .B(n8374), .Z(c[221]) );
  XNOR U12471 ( .A(b[2219]), .B(n8373), .Z(c[2219]) );
  XOR U12472 ( .A(n8375), .B(n8376), .Z(n8371) );
  ANDN U12473 ( .B(n8377), .A(n8378), .Z(n8375) );
  XNOR U12474 ( .A(b[2218]), .B(n8376), .Z(n8377) );
  XNOR U12475 ( .A(b[2218]), .B(n8378), .Z(c[2218]) );
  XOR U12476 ( .A(n8379), .B(n8380), .Z(n8376) );
  ANDN U12477 ( .B(n8381), .A(n8382), .Z(n8379) );
  XNOR U12478 ( .A(b[2217]), .B(n8380), .Z(n8381) );
  XNOR U12479 ( .A(b[2217]), .B(n8382), .Z(c[2217]) );
  XOR U12480 ( .A(n8383), .B(n8384), .Z(n8380) );
  ANDN U12481 ( .B(n8385), .A(n8386), .Z(n8383) );
  XNOR U12482 ( .A(b[2216]), .B(n8384), .Z(n8385) );
  XNOR U12483 ( .A(b[2216]), .B(n8386), .Z(c[2216]) );
  XOR U12484 ( .A(n8387), .B(n8388), .Z(n8384) );
  ANDN U12485 ( .B(n8389), .A(n8390), .Z(n8387) );
  XNOR U12486 ( .A(b[2215]), .B(n8388), .Z(n8389) );
  XNOR U12487 ( .A(b[2215]), .B(n8390), .Z(c[2215]) );
  XOR U12488 ( .A(n8391), .B(n8392), .Z(n8388) );
  ANDN U12489 ( .B(n8393), .A(n8394), .Z(n8391) );
  XNOR U12490 ( .A(b[2214]), .B(n8392), .Z(n8393) );
  XNOR U12491 ( .A(b[2214]), .B(n8394), .Z(c[2214]) );
  XOR U12492 ( .A(n8395), .B(n8396), .Z(n8392) );
  ANDN U12493 ( .B(n8397), .A(n8398), .Z(n8395) );
  XNOR U12494 ( .A(b[2213]), .B(n8396), .Z(n8397) );
  XNOR U12495 ( .A(b[2213]), .B(n8398), .Z(c[2213]) );
  XOR U12496 ( .A(n8399), .B(n8400), .Z(n8396) );
  ANDN U12497 ( .B(n8401), .A(n8402), .Z(n8399) );
  XNOR U12498 ( .A(b[2212]), .B(n8400), .Z(n8401) );
  XNOR U12499 ( .A(b[2212]), .B(n8402), .Z(c[2212]) );
  XOR U12500 ( .A(n8403), .B(n8404), .Z(n8400) );
  ANDN U12501 ( .B(n8405), .A(n8406), .Z(n8403) );
  XNOR U12502 ( .A(b[2211]), .B(n8404), .Z(n8405) );
  XNOR U12503 ( .A(b[2211]), .B(n8406), .Z(c[2211]) );
  XOR U12504 ( .A(n8407), .B(n8408), .Z(n8404) );
  ANDN U12505 ( .B(n8409), .A(n8410), .Z(n8407) );
  XNOR U12506 ( .A(b[2210]), .B(n8408), .Z(n8409) );
  XNOR U12507 ( .A(b[2210]), .B(n8410), .Z(c[2210]) );
  XOR U12508 ( .A(n8411), .B(n8412), .Z(n8408) );
  ANDN U12509 ( .B(n8413), .A(n8414), .Z(n8411) );
  XNOR U12510 ( .A(b[2209]), .B(n8412), .Z(n8413) );
  XNOR U12511 ( .A(b[220]), .B(n8415), .Z(c[220]) );
  XNOR U12512 ( .A(b[2209]), .B(n8414), .Z(c[2209]) );
  XOR U12513 ( .A(n8416), .B(n8417), .Z(n8412) );
  ANDN U12514 ( .B(n8418), .A(n8419), .Z(n8416) );
  XNOR U12515 ( .A(b[2208]), .B(n8417), .Z(n8418) );
  XNOR U12516 ( .A(b[2208]), .B(n8419), .Z(c[2208]) );
  XOR U12517 ( .A(n8420), .B(n8421), .Z(n8417) );
  ANDN U12518 ( .B(n8422), .A(n8423), .Z(n8420) );
  XNOR U12519 ( .A(b[2207]), .B(n8421), .Z(n8422) );
  XNOR U12520 ( .A(b[2207]), .B(n8423), .Z(c[2207]) );
  XOR U12521 ( .A(n8424), .B(n8425), .Z(n8421) );
  ANDN U12522 ( .B(n8426), .A(n8427), .Z(n8424) );
  XNOR U12523 ( .A(b[2206]), .B(n8425), .Z(n8426) );
  XNOR U12524 ( .A(b[2206]), .B(n8427), .Z(c[2206]) );
  XOR U12525 ( .A(n8428), .B(n8429), .Z(n8425) );
  ANDN U12526 ( .B(n8430), .A(n8431), .Z(n8428) );
  XNOR U12527 ( .A(b[2205]), .B(n8429), .Z(n8430) );
  XNOR U12528 ( .A(b[2205]), .B(n8431), .Z(c[2205]) );
  XOR U12529 ( .A(n8432), .B(n8433), .Z(n8429) );
  ANDN U12530 ( .B(n8434), .A(n8435), .Z(n8432) );
  XNOR U12531 ( .A(b[2204]), .B(n8433), .Z(n8434) );
  XNOR U12532 ( .A(b[2204]), .B(n8435), .Z(c[2204]) );
  XOR U12533 ( .A(n8436), .B(n8437), .Z(n8433) );
  ANDN U12534 ( .B(n8438), .A(n8439), .Z(n8436) );
  XNOR U12535 ( .A(b[2203]), .B(n8437), .Z(n8438) );
  XNOR U12536 ( .A(b[2203]), .B(n8439), .Z(c[2203]) );
  XOR U12537 ( .A(n8440), .B(n8441), .Z(n8437) );
  ANDN U12538 ( .B(n8442), .A(n8443), .Z(n8440) );
  XNOR U12539 ( .A(b[2202]), .B(n8441), .Z(n8442) );
  XNOR U12540 ( .A(b[2202]), .B(n8443), .Z(c[2202]) );
  XOR U12541 ( .A(n8444), .B(n8445), .Z(n8441) );
  ANDN U12542 ( .B(n8446), .A(n8447), .Z(n8444) );
  XNOR U12543 ( .A(b[2201]), .B(n8445), .Z(n8446) );
  XNOR U12544 ( .A(b[2201]), .B(n8447), .Z(c[2201]) );
  XOR U12545 ( .A(n8448), .B(n8449), .Z(n8445) );
  ANDN U12546 ( .B(n8450), .A(n8451), .Z(n8448) );
  XNOR U12547 ( .A(b[2200]), .B(n8449), .Z(n8450) );
  XNOR U12548 ( .A(b[2200]), .B(n8451), .Z(c[2200]) );
  XOR U12549 ( .A(n8452), .B(n8453), .Z(n8449) );
  ANDN U12550 ( .B(n8454), .A(n8455), .Z(n8452) );
  XNOR U12551 ( .A(b[2199]), .B(n8453), .Z(n8454) );
  XNOR U12552 ( .A(b[21]), .B(n8456), .Z(c[21]) );
  XNOR U12553 ( .A(b[219]), .B(n8457), .Z(c[219]) );
  XNOR U12554 ( .A(b[2199]), .B(n8455), .Z(c[2199]) );
  XOR U12555 ( .A(n8458), .B(n8459), .Z(n8453) );
  ANDN U12556 ( .B(n8460), .A(n8461), .Z(n8458) );
  XNOR U12557 ( .A(b[2198]), .B(n8459), .Z(n8460) );
  XNOR U12558 ( .A(b[2198]), .B(n8461), .Z(c[2198]) );
  XOR U12559 ( .A(n8462), .B(n8463), .Z(n8459) );
  ANDN U12560 ( .B(n8464), .A(n8465), .Z(n8462) );
  XNOR U12561 ( .A(b[2197]), .B(n8463), .Z(n8464) );
  XNOR U12562 ( .A(b[2197]), .B(n8465), .Z(c[2197]) );
  XOR U12563 ( .A(n8466), .B(n8467), .Z(n8463) );
  ANDN U12564 ( .B(n8468), .A(n8469), .Z(n8466) );
  XNOR U12565 ( .A(b[2196]), .B(n8467), .Z(n8468) );
  XNOR U12566 ( .A(b[2196]), .B(n8469), .Z(c[2196]) );
  XOR U12567 ( .A(n8470), .B(n8471), .Z(n8467) );
  ANDN U12568 ( .B(n8472), .A(n8473), .Z(n8470) );
  XNOR U12569 ( .A(b[2195]), .B(n8471), .Z(n8472) );
  XNOR U12570 ( .A(b[2195]), .B(n8473), .Z(c[2195]) );
  XOR U12571 ( .A(n8474), .B(n8475), .Z(n8471) );
  ANDN U12572 ( .B(n8476), .A(n8477), .Z(n8474) );
  XNOR U12573 ( .A(b[2194]), .B(n8475), .Z(n8476) );
  XNOR U12574 ( .A(b[2194]), .B(n8477), .Z(c[2194]) );
  XOR U12575 ( .A(n8478), .B(n8479), .Z(n8475) );
  ANDN U12576 ( .B(n8480), .A(n8481), .Z(n8478) );
  XNOR U12577 ( .A(b[2193]), .B(n8479), .Z(n8480) );
  XNOR U12578 ( .A(b[2193]), .B(n8481), .Z(c[2193]) );
  XOR U12579 ( .A(n8482), .B(n8483), .Z(n8479) );
  ANDN U12580 ( .B(n8484), .A(n8485), .Z(n8482) );
  XNOR U12581 ( .A(b[2192]), .B(n8483), .Z(n8484) );
  XNOR U12582 ( .A(b[2192]), .B(n8485), .Z(c[2192]) );
  XOR U12583 ( .A(n8486), .B(n8487), .Z(n8483) );
  ANDN U12584 ( .B(n8488), .A(n8489), .Z(n8486) );
  XNOR U12585 ( .A(b[2191]), .B(n8487), .Z(n8488) );
  XNOR U12586 ( .A(b[2191]), .B(n8489), .Z(c[2191]) );
  XOR U12587 ( .A(n8490), .B(n8491), .Z(n8487) );
  ANDN U12588 ( .B(n8492), .A(n8493), .Z(n8490) );
  XNOR U12589 ( .A(b[2190]), .B(n8491), .Z(n8492) );
  XNOR U12590 ( .A(b[2190]), .B(n8493), .Z(c[2190]) );
  XOR U12591 ( .A(n8494), .B(n8495), .Z(n8491) );
  ANDN U12592 ( .B(n8496), .A(n8497), .Z(n8494) );
  XNOR U12593 ( .A(b[2189]), .B(n8495), .Z(n8496) );
  XNOR U12594 ( .A(b[218]), .B(n8498), .Z(c[218]) );
  XNOR U12595 ( .A(b[2189]), .B(n8497), .Z(c[2189]) );
  XOR U12596 ( .A(n8499), .B(n8500), .Z(n8495) );
  ANDN U12597 ( .B(n8501), .A(n8502), .Z(n8499) );
  XNOR U12598 ( .A(b[2188]), .B(n8500), .Z(n8501) );
  XNOR U12599 ( .A(b[2188]), .B(n8502), .Z(c[2188]) );
  XOR U12600 ( .A(n8503), .B(n8504), .Z(n8500) );
  ANDN U12601 ( .B(n8505), .A(n8506), .Z(n8503) );
  XNOR U12602 ( .A(b[2187]), .B(n8504), .Z(n8505) );
  XNOR U12603 ( .A(b[2187]), .B(n8506), .Z(c[2187]) );
  XOR U12604 ( .A(n8507), .B(n8508), .Z(n8504) );
  ANDN U12605 ( .B(n8509), .A(n8510), .Z(n8507) );
  XNOR U12606 ( .A(b[2186]), .B(n8508), .Z(n8509) );
  XNOR U12607 ( .A(b[2186]), .B(n8510), .Z(c[2186]) );
  XOR U12608 ( .A(n8511), .B(n8512), .Z(n8508) );
  ANDN U12609 ( .B(n8513), .A(n8514), .Z(n8511) );
  XNOR U12610 ( .A(b[2185]), .B(n8512), .Z(n8513) );
  XNOR U12611 ( .A(b[2185]), .B(n8514), .Z(c[2185]) );
  XOR U12612 ( .A(n8515), .B(n8516), .Z(n8512) );
  ANDN U12613 ( .B(n8517), .A(n8518), .Z(n8515) );
  XNOR U12614 ( .A(b[2184]), .B(n8516), .Z(n8517) );
  XNOR U12615 ( .A(b[2184]), .B(n8518), .Z(c[2184]) );
  XOR U12616 ( .A(n8519), .B(n8520), .Z(n8516) );
  ANDN U12617 ( .B(n8521), .A(n8522), .Z(n8519) );
  XNOR U12618 ( .A(b[2183]), .B(n8520), .Z(n8521) );
  XNOR U12619 ( .A(b[2183]), .B(n8522), .Z(c[2183]) );
  XOR U12620 ( .A(n8523), .B(n8524), .Z(n8520) );
  ANDN U12621 ( .B(n8525), .A(n8526), .Z(n8523) );
  XNOR U12622 ( .A(b[2182]), .B(n8524), .Z(n8525) );
  XNOR U12623 ( .A(b[2182]), .B(n8526), .Z(c[2182]) );
  XOR U12624 ( .A(n8527), .B(n8528), .Z(n8524) );
  ANDN U12625 ( .B(n8529), .A(n8530), .Z(n8527) );
  XNOR U12626 ( .A(b[2181]), .B(n8528), .Z(n8529) );
  XNOR U12627 ( .A(b[2181]), .B(n8530), .Z(c[2181]) );
  XOR U12628 ( .A(n8531), .B(n8532), .Z(n8528) );
  ANDN U12629 ( .B(n8533), .A(n8534), .Z(n8531) );
  XNOR U12630 ( .A(b[2180]), .B(n8532), .Z(n8533) );
  XNOR U12631 ( .A(b[2180]), .B(n8534), .Z(c[2180]) );
  XOR U12632 ( .A(n8535), .B(n8536), .Z(n8532) );
  ANDN U12633 ( .B(n8537), .A(n8538), .Z(n8535) );
  XNOR U12634 ( .A(b[2179]), .B(n8536), .Z(n8537) );
  XNOR U12635 ( .A(b[217]), .B(n8539), .Z(c[217]) );
  XNOR U12636 ( .A(b[2179]), .B(n8538), .Z(c[2179]) );
  XOR U12637 ( .A(n8540), .B(n8541), .Z(n8536) );
  ANDN U12638 ( .B(n8542), .A(n8543), .Z(n8540) );
  XNOR U12639 ( .A(b[2178]), .B(n8541), .Z(n8542) );
  XNOR U12640 ( .A(b[2178]), .B(n8543), .Z(c[2178]) );
  XOR U12641 ( .A(n8544), .B(n8545), .Z(n8541) );
  ANDN U12642 ( .B(n8546), .A(n8547), .Z(n8544) );
  XNOR U12643 ( .A(b[2177]), .B(n8545), .Z(n8546) );
  XNOR U12644 ( .A(b[2177]), .B(n8547), .Z(c[2177]) );
  XOR U12645 ( .A(n8548), .B(n8549), .Z(n8545) );
  ANDN U12646 ( .B(n8550), .A(n8551), .Z(n8548) );
  XNOR U12647 ( .A(b[2176]), .B(n8549), .Z(n8550) );
  XNOR U12648 ( .A(b[2176]), .B(n8551), .Z(c[2176]) );
  XOR U12649 ( .A(n8552), .B(n8553), .Z(n8549) );
  ANDN U12650 ( .B(n8554), .A(n8555), .Z(n8552) );
  XNOR U12651 ( .A(b[2175]), .B(n8553), .Z(n8554) );
  XNOR U12652 ( .A(b[2175]), .B(n8555), .Z(c[2175]) );
  XOR U12653 ( .A(n8556), .B(n8557), .Z(n8553) );
  ANDN U12654 ( .B(n8558), .A(n8559), .Z(n8556) );
  XNOR U12655 ( .A(b[2174]), .B(n8557), .Z(n8558) );
  XNOR U12656 ( .A(b[2174]), .B(n8559), .Z(c[2174]) );
  XOR U12657 ( .A(n8560), .B(n8561), .Z(n8557) );
  ANDN U12658 ( .B(n8562), .A(n8563), .Z(n8560) );
  XNOR U12659 ( .A(b[2173]), .B(n8561), .Z(n8562) );
  XNOR U12660 ( .A(b[2173]), .B(n8563), .Z(c[2173]) );
  XOR U12661 ( .A(n8564), .B(n8565), .Z(n8561) );
  ANDN U12662 ( .B(n8566), .A(n8567), .Z(n8564) );
  XNOR U12663 ( .A(b[2172]), .B(n8565), .Z(n8566) );
  XNOR U12664 ( .A(b[2172]), .B(n8567), .Z(c[2172]) );
  XOR U12665 ( .A(n8568), .B(n8569), .Z(n8565) );
  ANDN U12666 ( .B(n8570), .A(n8571), .Z(n8568) );
  XNOR U12667 ( .A(b[2171]), .B(n8569), .Z(n8570) );
  XNOR U12668 ( .A(b[2171]), .B(n8571), .Z(c[2171]) );
  XOR U12669 ( .A(n8572), .B(n8573), .Z(n8569) );
  ANDN U12670 ( .B(n8574), .A(n8575), .Z(n8572) );
  XNOR U12671 ( .A(b[2170]), .B(n8573), .Z(n8574) );
  XNOR U12672 ( .A(b[2170]), .B(n8575), .Z(c[2170]) );
  XOR U12673 ( .A(n8576), .B(n8577), .Z(n8573) );
  ANDN U12674 ( .B(n8578), .A(n8579), .Z(n8576) );
  XNOR U12675 ( .A(b[2169]), .B(n8577), .Z(n8578) );
  XNOR U12676 ( .A(b[216]), .B(n8580), .Z(c[216]) );
  XNOR U12677 ( .A(b[2169]), .B(n8579), .Z(c[2169]) );
  XOR U12678 ( .A(n8581), .B(n8582), .Z(n8577) );
  ANDN U12679 ( .B(n8583), .A(n8584), .Z(n8581) );
  XNOR U12680 ( .A(b[2168]), .B(n8582), .Z(n8583) );
  XNOR U12681 ( .A(b[2168]), .B(n8584), .Z(c[2168]) );
  XOR U12682 ( .A(n8585), .B(n8586), .Z(n8582) );
  ANDN U12683 ( .B(n8587), .A(n8588), .Z(n8585) );
  XNOR U12684 ( .A(b[2167]), .B(n8586), .Z(n8587) );
  XNOR U12685 ( .A(b[2167]), .B(n8588), .Z(c[2167]) );
  XOR U12686 ( .A(n8589), .B(n8590), .Z(n8586) );
  ANDN U12687 ( .B(n8591), .A(n8592), .Z(n8589) );
  XNOR U12688 ( .A(b[2166]), .B(n8590), .Z(n8591) );
  XNOR U12689 ( .A(b[2166]), .B(n8592), .Z(c[2166]) );
  XOR U12690 ( .A(n8593), .B(n8594), .Z(n8590) );
  ANDN U12691 ( .B(n8595), .A(n8596), .Z(n8593) );
  XNOR U12692 ( .A(b[2165]), .B(n8594), .Z(n8595) );
  XNOR U12693 ( .A(b[2165]), .B(n8596), .Z(c[2165]) );
  XOR U12694 ( .A(n8597), .B(n8598), .Z(n8594) );
  ANDN U12695 ( .B(n8599), .A(n8600), .Z(n8597) );
  XNOR U12696 ( .A(b[2164]), .B(n8598), .Z(n8599) );
  XNOR U12697 ( .A(b[2164]), .B(n8600), .Z(c[2164]) );
  XOR U12698 ( .A(n8601), .B(n8602), .Z(n8598) );
  ANDN U12699 ( .B(n8603), .A(n8604), .Z(n8601) );
  XNOR U12700 ( .A(b[2163]), .B(n8602), .Z(n8603) );
  XNOR U12701 ( .A(b[2163]), .B(n8604), .Z(c[2163]) );
  XOR U12702 ( .A(n8605), .B(n8606), .Z(n8602) );
  ANDN U12703 ( .B(n8607), .A(n8608), .Z(n8605) );
  XNOR U12704 ( .A(b[2162]), .B(n8606), .Z(n8607) );
  XNOR U12705 ( .A(b[2162]), .B(n8608), .Z(c[2162]) );
  XOR U12706 ( .A(n8609), .B(n8610), .Z(n8606) );
  ANDN U12707 ( .B(n8611), .A(n8612), .Z(n8609) );
  XNOR U12708 ( .A(b[2161]), .B(n8610), .Z(n8611) );
  XNOR U12709 ( .A(b[2161]), .B(n8612), .Z(c[2161]) );
  XOR U12710 ( .A(n8613), .B(n8614), .Z(n8610) );
  ANDN U12711 ( .B(n8615), .A(n8616), .Z(n8613) );
  XNOR U12712 ( .A(b[2160]), .B(n8614), .Z(n8615) );
  XNOR U12713 ( .A(b[2160]), .B(n8616), .Z(c[2160]) );
  XOR U12714 ( .A(n8617), .B(n8618), .Z(n8614) );
  ANDN U12715 ( .B(n8619), .A(n8620), .Z(n8617) );
  XNOR U12716 ( .A(b[2159]), .B(n8618), .Z(n8619) );
  XNOR U12717 ( .A(b[215]), .B(n8621), .Z(c[215]) );
  XNOR U12718 ( .A(b[2159]), .B(n8620), .Z(c[2159]) );
  XOR U12719 ( .A(n8622), .B(n8623), .Z(n8618) );
  ANDN U12720 ( .B(n8624), .A(n8625), .Z(n8622) );
  XNOR U12721 ( .A(b[2158]), .B(n8623), .Z(n8624) );
  XNOR U12722 ( .A(b[2158]), .B(n8625), .Z(c[2158]) );
  XOR U12723 ( .A(n8626), .B(n8627), .Z(n8623) );
  ANDN U12724 ( .B(n8628), .A(n8629), .Z(n8626) );
  XNOR U12725 ( .A(b[2157]), .B(n8627), .Z(n8628) );
  XNOR U12726 ( .A(b[2157]), .B(n8629), .Z(c[2157]) );
  XOR U12727 ( .A(n8630), .B(n8631), .Z(n8627) );
  ANDN U12728 ( .B(n8632), .A(n8633), .Z(n8630) );
  XNOR U12729 ( .A(b[2156]), .B(n8631), .Z(n8632) );
  XNOR U12730 ( .A(b[2156]), .B(n8633), .Z(c[2156]) );
  XOR U12731 ( .A(n8634), .B(n8635), .Z(n8631) );
  ANDN U12732 ( .B(n8636), .A(n8637), .Z(n8634) );
  XNOR U12733 ( .A(b[2155]), .B(n8635), .Z(n8636) );
  XNOR U12734 ( .A(b[2155]), .B(n8637), .Z(c[2155]) );
  XOR U12735 ( .A(n8638), .B(n8639), .Z(n8635) );
  ANDN U12736 ( .B(n8640), .A(n8641), .Z(n8638) );
  XNOR U12737 ( .A(b[2154]), .B(n8639), .Z(n8640) );
  XNOR U12738 ( .A(b[2154]), .B(n8641), .Z(c[2154]) );
  XOR U12739 ( .A(n8642), .B(n8643), .Z(n8639) );
  ANDN U12740 ( .B(n8644), .A(n8645), .Z(n8642) );
  XNOR U12741 ( .A(b[2153]), .B(n8643), .Z(n8644) );
  XNOR U12742 ( .A(b[2153]), .B(n8645), .Z(c[2153]) );
  XOR U12743 ( .A(n8646), .B(n8647), .Z(n8643) );
  ANDN U12744 ( .B(n8648), .A(n8649), .Z(n8646) );
  XNOR U12745 ( .A(b[2152]), .B(n8647), .Z(n8648) );
  XNOR U12746 ( .A(b[2152]), .B(n8649), .Z(c[2152]) );
  XOR U12747 ( .A(n8650), .B(n8651), .Z(n8647) );
  ANDN U12748 ( .B(n8652), .A(n8653), .Z(n8650) );
  XNOR U12749 ( .A(b[2151]), .B(n8651), .Z(n8652) );
  XNOR U12750 ( .A(b[2151]), .B(n8653), .Z(c[2151]) );
  XOR U12751 ( .A(n8654), .B(n8655), .Z(n8651) );
  ANDN U12752 ( .B(n8656), .A(n8657), .Z(n8654) );
  XNOR U12753 ( .A(b[2150]), .B(n8655), .Z(n8656) );
  XNOR U12754 ( .A(b[2150]), .B(n8657), .Z(c[2150]) );
  XOR U12755 ( .A(n8658), .B(n8659), .Z(n8655) );
  ANDN U12756 ( .B(n8660), .A(n8661), .Z(n8658) );
  XNOR U12757 ( .A(b[2149]), .B(n8659), .Z(n8660) );
  XNOR U12758 ( .A(b[214]), .B(n8662), .Z(c[214]) );
  XNOR U12759 ( .A(b[2149]), .B(n8661), .Z(c[2149]) );
  XOR U12760 ( .A(n8663), .B(n8664), .Z(n8659) );
  ANDN U12761 ( .B(n8665), .A(n8666), .Z(n8663) );
  XNOR U12762 ( .A(b[2148]), .B(n8664), .Z(n8665) );
  XNOR U12763 ( .A(b[2148]), .B(n8666), .Z(c[2148]) );
  XOR U12764 ( .A(n8667), .B(n8668), .Z(n8664) );
  ANDN U12765 ( .B(n8669), .A(n8670), .Z(n8667) );
  XNOR U12766 ( .A(b[2147]), .B(n8668), .Z(n8669) );
  XNOR U12767 ( .A(b[2147]), .B(n8670), .Z(c[2147]) );
  XOR U12768 ( .A(n8671), .B(n8672), .Z(n8668) );
  ANDN U12769 ( .B(n8673), .A(n8674), .Z(n8671) );
  XNOR U12770 ( .A(b[2146]), .B(n8672), .Z(n8673) );
  XNOR U12771 ( .A(b[2146]), .B(n8674), .Z(c[2146]) );
  XOR U12772 ( .A(n8675), .B(n8676), .Z(n8672) );
  ANDN U12773 ( .B(n8677), .A(n8678), .Z(n8675) );
  XNOR U12774 ( .A(b[2145]), .B(n8676), .Z(n8677) );
  XNOR U12775 ( .A(b[2145]), .B(n8678), .Z(c[2145]) );
  XOR U12776 ( .A(n8679), .B(n8680), .Z(n8676) );
  ANDN U12777 ( .B(n8681), .A(n8682), .Z(n8679) );
  XNOR U12778 ( .A(b[2144]), .B(n8680), .Z(n8681) );
  XNOR U12779 ( .A(b[2144]), .B(n8682), .Z(c[2144]) );
  XOR U12780 ( .A(n8683), .B(n8684), .Z(n8680) );
  ANDN U12781 ( .B(n8685), .A(n8686), .Z(n8683) );
  XNOR U12782 ( .A(b[2143]), .B(n8684), .Z(n8685) );
  XNOR U12783 ( .A(b[2143]), .B(n8686), .Z(c[2143]) );
  XOR U12784 ( .A(n8687), .B(n8688), .Z(n8684) );
  ANDN U12785 ( .B(n8689), .A(n8690), .Z(n8687) );
  XNOR U12786 ( .A(b[2142]), .B(n8688), .Z(n8689) );
  XNOR U12787 ( .A(b[2142]), .B(n8690), .Z(c[2142]) );
  XOR U12788 ( .A(n8691), .B(n8692), .Z(n8688) );
  ANDN U12789 ( .B(n8693), .A(n8694), .Z(n8691) );
  XNOR U12790 ( .A(b[2141]), .B(n8692), .Z(n8693) );
  XNOR U12791 ( .A(b[2141]), .B(n8694), .Z(c[2141]) );
  XOR U12792 ( .A(n8695), .B(n8696), .Z(n8692) );
  ANDN U12793 ( .B(n8697), .A(n8698), .Z(n8695) );
  XNOR U12794 ( .A(b[2140]), .B(n8696), .Z(n8697) );
  XNOR U12795 ( .A(b[2140]), .B(n8698), .Z(c[2140]) );
  XOR U12796 ( .A(n8699), .B(n8700), .Z(n8696) );
  ANDN U12797 ( .B(n8701), .A(n8702), .Z(n8699) );
  XNOR U12798 ( .A(b[2139]), .B(n8700), .Z(n8701) );
  XNOR U12799 ( .A(b[213]), .B(n8703), .Z(c[213]) );
  XNOR U12800 ( .A(b[2139]), .B(n8702), .Z(c[2139]) );
  XOR U12801 ( .A(n8704), .B(n8705), .Z(n8700) );
  ANDN U12802 ( .B(n8706), .A(n8707), .Z(n8704) );
  XNOR U12803 ( .A(b[2138]), .B(n8705), .Z(n8706) );
  XNOR U12804 ( .A(b[2138]), .B(n8707), .Z(c[2138]) );
  XOR U12805 ( .A(n8708), .B(n8709), .Z(n8705) );
  ANDN U12806 ( .B(n8710), .A(n8711), .Z(n8708) );
  XNOR U12807 ( .A(b[2137]), .B(n8709), .Z(n8710) );
  XNOR U12808 ( .A(b[2137]), .B(n8711), .Z(c[2137]) );
  XOR U12809 ( .A(n8712), .B(n8713), .Z(n8709) );
  ANDN U12810 ( .B(n8714), .A(n8715), .Z(n8712) );
  XNOR U12811 ( .A(b[2136]), .B(n8713), .Z(n8714) );
  XNOR U12812 ( .A(b[2136]), .B(n8715), .Z(c[2136]) );
  XOR U12813 ( .A(n8716), .B(n8717), .Z(n8713) );
  ANDN U12814 ( .B(n8718), .A(n8719), .Z(n8716) );
  XNOR U12815 ( .A(b[2135]), .B(n8717), .Z(n8718) );
  XNOR U12816 ( .A(b[2135]), .B(n8719), .Z(c[2135]) );
  XOR U12817 ( .A(n8720), .B(n8721), .Z(n8717) );
  ANDN U12818 ( .B(n8722), .A(n8723), .Z(n8720) );
  XNOR U12819 ( .A(b[2134]), .B(n8721), .Z(n8722) );
  XNOR U12820 ( .A(b[2134]), .B(n8723), .Z(c[2134]) );
  XOR U12821 ( .A(n8724), .B(n8725), .Z(n8721) );
  ANDN U12822 ( .B(n8726), .A(n8727), .Z(n8724) );
  XNOR U12823 ( .A(b[2133]), .B(n8725), .Z(n8726) );
  XNOR U12824 ( .A(b[2133]), .B(n8727), .Z(c[2133]) );
  XOR U12825 ( .A(n8728), .B(n8729), .Z(n8725) );
  ANDN U12826 ( .B(n8730), .A(n8731), .Z(n8728) );
  XNOR U12827 ( .A(b[2132]), .B(n8729), .Z(n8730) );
  XNOR U12828 ( .A(b[2132]), .B(n8731), .Z(c[2132]) );
  XOR U12829 ( .A(n8732), .B(n8733), .Z(n8729) );
  ANDN U12830 ( .B(n8734), .A(n8735), .Z(n8732) );
  XNOR U12831 ( .A(b[2131]), .B(n8733), .Z(n8734) );
  XNOR U12832 ( .A(b[2131]), .B(n8735), .Z(c[2131]) );
  XOR U12833 ( .A(n8736), .B(n8737), .Z(n8733) );
  ANDN U12834 ( .B(n8738), .A(n8739), .Z(n8736) );
  XNOR U12835 ( .A(b[2130]), .B(n8737), .Z(n8738) );
  XNOR U12836 ( .A(b[2130]), .B(n8739), .Z(c[2130]) );
  XOR U12837 ( .A(n8740), .B(n8741), .Z(n8737) );
  ANDN U12838 ( .B(n8742), .A(n8743), .Z(n8740) );
  XNOR U12839 ( .A(b[2129]), .B(n8741), .Z(n8742) );
  XNOR U12840 ( .A(b[212]), .B(n8744), .Z(c[212]) );
  XNOR U12841 ( .A(b[2129]), .B(n8743), .Z(c[2129]) );
  XOR U12842 ( .A(n8745), .B(n8746), .Z(n8741) );
  ANDN U12843 ( .B(n8747), .A(n8748), .Z(n8745) );
  XNOR U12844 ( .A(b[2128]), .B(n8746), .Z(n8747) );
  XNOR U12845 ( .A(b[2128]), .B(n8748), .Z(c[2128]) );
  XOR U12846 ( .A(n8749), .B(n8750), .Z(n8746) );
  ANDN U12847 ( .B(n8751), .A(n8752), .Z(n8749) );
  XNOR U12848 ( .A(b[2127]), .B(n8750), .Z(n8751) );
  XNOR U12849 ( .A(b[2127]), .B(n8752), .Z(c[2127]) );
  XOR U12850 ( .A(n8753), .B(n8754), .Z(n8750) );
  ANDN U12851 ( .B(n8755), .A(n8756), .Z(n8753) );
  XNOR U12852 ( .A(b[2126]), .B(n8754), .Z(n8755) );
  XNOR U12853 ( .A(b[2126]), .B(n8756), .Z(c[2126]) );
  XOR U12854 ( .A(n8757), .B(n8758), .Z(n8754) );
  ANDN U12855 ( .B(n8759), .A(n8760), .Z(n8757) );
  XNOR U12856 ( .A(b[2125]), .B(n8758), .Z(n8759) );
  XNOR U12857 ( .A(b[2125]), .B(n8760), .Z(c[2125]) );
  XOR U12858 ( .A(n8761), .B(n8762), .Z(n8758) );
  ANDN U12859 ( .B(n8763), .A(n8764), .Z(n8761) );
  XNOR U12860 ( .A(b[2124]), .B(n8762), .Z(n8763) );
  XNOR U12861 ( .A(b[2124]), .B(n8764), .Z(c[2124]) );
  XOR U12862 ( .A(n8765), .B(n8766), .Z(n8762) );
  ANDN U12863 ( .B(n8767), .A(n8768), .Z(n8765) );
  XNOR U12864 ( .A(b[2123]), .B(n8766), .Z(n8767) );
  XNOR U12865 ( .A(b[2123]), .B(n8768), .Z(c[2123]) );
  XOR U12866 ( .A(n8769), .B(n8770), .Z(n8766) );
  ANDN U12867 ( .B(n8771), .A(n8772), .Z(n8769) );
  XNOR U12868 ( .A(b[2122]), .B(n8770), .Z(n8771) );
  XNOR U12869 ( .A(b[2122]), .B(n8772), .Z(c[2122]) );
  XOR U12870 ( .A(n8773), .B(n8774), .Z(n8770) );
  ANDN U12871 ( .B(n8775), .A(n8776), .Z(n8773) );
  XNOR U12872 ( .A(b[2121]), .B(n8774), .Z(n8775) );
  XNOR U12873 ( .A(b[2121]), .B(n8776), .Z(c[2121]) );
  XOR U12874 ( .A(n8777), .B(n8778), .Z(n8774) );
  ANDN U12875 ( .B(n8779), .A(n8780), .Z(n8777) );
  XNOR U12876 ( .A(b[2120]), .B(n8778), .Z(n8779) );
  XNOR U12877 ( .A(b[2120]), .B(n8780), .Z(c[2120]) );
  XOR U12878 ( .A(n8781), .B(n8782), .Z(n8778) );
  ANDN U12879 ( .B(n8783), .A(n8784), .Z(n8781) );
  XNOR U12880 ( .A(b[2119]), .B(n8782), .Z(n8783) );
  XNOR U12881 ( .A(b[211]), .B(n8785), .Z(c[211]) );
  XNOR U12882 ( .A(b[2119]), .B(n8784), .Z(c[2119]) );
  XOR U12883 ( .A(n8786), .B(n8787), .Z(n8782) );
  ANDN U12884 ( .B(n8788), .A(n8789), .Z(n8786) );
  XNOR U12885 ( .A(b[2118]), .B(n8787), .Z(n8788) );
  XNOR U12886 ( .A(b[2118]), .B(n8789), .Z(c[2118]) );
  XOR U12887 ( .A(n8790), .B(n8791), .Z(n8787) );
  ANDN U12888 ( .B(n8792), .A(n8793), .Z(n8790) );
  XNOR U12889 ( .A(b[2117]), .B(n8791), .Z(n8792) );
  XNOR U12890 ( .A(b[2117]), .B(n8793), .Z(c[2117]) );
  XOR U12891 ( .A(n8794), .B(n8795), .Z(n8791) );
  ANDN U12892 ( .B(n8796), .A(n8797), .Z(n8794) );
  XNOR U12893 ( .A(b[2116]), .B(n8795), .Z(n8796) );
  XNOR U12894 ( .A(b[2116]), .B(n8797), .Z(c[2116]) );
  XOR U12895 ( .A(n8798), .B(n8799), .Z(n8795) );
  ANDN U12896 ( .B(n8800), .A(n8801), .Z(n8798) );
  XNOR U12897 ( .A(b[2115]), .B(n8799), .Z(n8800) );
  XNOR U12898 ( .A(b[2115]), .B(n8801), .Z(c[2115]) );
  XOR U12899 ( .A(n8802), .B(n8803), .Z(n8799) );
  ANDN U12900 ( .B(n8804), .A(n8805), .Z(n8802) );
  XNOR U12901 ( .A(b[2114]), .B(n8803), .Z(n8804) );
  XNOR U12902 ( .A(b[2114]), .B(n8805), .Z(c[2114]) );
  XOR U12903 ( .A(n8806), .B(n8807), .Z(n8803) );
  ANDN U12904 ( .B(n8808), .A(n8809), .Z(n8806) );
  XNOR U12905 ( .A(b[2113]), .B(n8807), .Z(n8808) );
  XNOR U12906 ( .A(b[2113]), .B(n8809), .Z(c[2113]) );
  XOR U12907 ( .A(n8810), .B(n8811), .Z(n8807) );
  ANDN U12908 ( .B(n8812), .A(n8813), .Z(n8810) );
  XNOR U12909 ( .A(b[2112]), .B(n8811), .Z(n8812) );
  XNOR U12910 ( .A(b[2112]), .B(n8813), .Z(c[2112]) );
  XOR U12911 ( .A(n8814), .B(n8815), .Z(n8811) );
  ANDN U12912 ( .B(n8816), .A(n8817), .Z(n8814) );
  XNOR U12913 ( .A(b[2111]), .B(n8815), .Z(n8816) );
  XNOR U12914 ( .A(b[2111]), .B(n8817), .Z(c[2111]) );
  XOR U12915 ( .A(n8818), .B(n8819), .Z(n8815) );
  ANDN U12916 ( .B(n8820), .A(n8821), .Z(n8818) );
  XNOR U12917 ( .A(b[2110]), .B(n8819), .Z(n8820) );
  XNOR U12918 ( .A(b[2110]), .B(n8821), .Z(c[2110]) );
  XOR U12919 ( .A(n8822), .B(n8823), .Z(n8819) );
  ANDN U12920 ( .B(n8824), .A(n8825), .Z(n8822) );
  XNOR U12921 ( .A(b[2109]), .B(n8823), .Z(n8824) );
  XNOR U12922 ( .A(b[210]), .B(n8826), .Z(c[210]) );
  XNOR U12923 ( .A(b[2109]), .B(n8825), .Z(c[2109]) );
  XOR U12924 ( .A(n8827), .B(n8828), .Z(n8823) );
  ANDN U12925 ( .B(n8829), .A(n8830), .Z(n8827) );
  XNOR U12926 ( .A(b[2108]), .B(n8828), .Z(n8829) );
  XNOR U12927 ( .A(b[2108]), .B(n8830), .Z(c[2108]) );
  XOR U12928 ( .A(n8831), .B(n8832), .Z(n8828) );
  ANDN U12929 ( .B(n8833), .A(n8834), .Z(n8831) );
  XNOR U12930 ( .A(b[2107]), .B(n8832), .Z(n8833) );
  XNOR U12931 ( .A(b[2107]), .B(n8834), .Z(c[2107]) );
  XOR U12932 ( .A(n8835), .B(n8836), .Z(n8832) );
  ANDN U12933 ( .B(n8837), .A(n8838), .Z(n8835) );
  XNOR U12934 ( .A(b[2106]), .B(n8836), .Z(n8837) );
  XNOR U12935 ( .A(b[2106]), .B(n8838), .Z(c[2106]) );
  XOR U12936 ( .A(n8839), .B(n8840), .Z(n8836) );
  ANDN U12937 ( .B(n8841), .A(n8842), .Z(n8839) );
  XNOR U12938 ( .A(b[2105]), .B(n8840), .Z(n8841) );
  XNOR U12939 ( .A(b[2105]), .B(n8842), .Z(c[2105]) );
  XOR U12940 ( .A(n8843), .B(n8844), .Z(n8840) );
  ANDN U12941 ( .B(n8845), .A(n8846), .Z(n8843) );
  XNOR U12942 ( .A(b[2104]), .B(n8844), .Z(n8845) );
  XNOR U12943 ( .A(b[2104]), .B(n8846), .Z(c[2104]) );
  XOR U12944 ( .A(n8847), .B(n8848), .Z(n8844) );
  ANDN U12945 ( .B(n8849), .A(n8850), .Z(n8847) );
  XNOR U12946 ( .A(b[2103]), .B(n8848), .Z(n8849) );
  XNOR U12947 ( .A(b[2103]), .B(n8850), .Z(c[2103]) );
  XOR U12948 ( .A(n8851), .B(n8852), .Z(n8848) );
  ANDN U12949 ( .B(n8853), .A(n8854), .Z(n8851) );
  XNOR U12950 ( .A(b[2102]), .B(n8852), .Z(n8853) );
  XNOR U12951 ( .A(b[2102]), .B(n8854), .Z(c[2102]) );
  XOR U12952 ( .A(n8855), .B(n8856), .Z(n8852) );
  ANDN U12953 ( .B(n8857), .A(n8858), .Z(n8855) );
  XNOR U12954 ( .A(b[2101]), .B(n8856), .Z(n8857) );
  XNOR U12955 ( .A(b[2101]), .B(n8858), .Z(c[2101]) );
  XOR U12956 ( .A(n8859), .B(n8860), .Z(n8856) );
  ANDN U12957 ( .B(n8861), .A(n8862), .Z(n8859) );
  XNOR U12958 ( .A(b[2100]), .B(n8860), .Z(n8861) );
  XNOR U12959 ( .A(b[2100]), .B(n8862), .Z(c[2100]) );
  XOR U12960 ( .A(n8863), .B(n8864), .Z(n8860) );
  ANDN U12961 ( .B(n8865), .A(n8866), .Z(n8863) );
  XNOR U12962 ( .A(b[2099]), .B(n8864), .Z(n8865) );
  XNOR U12963 ( .A(b[20]), .B(n8867), .Z(c[20]) );
  XNOR U12964 ( .A(b[209]), .B(n8868), .Z(c[209]) );
  XNOR U12965 ( .A(b[2099]), .B(n8866), .Z(c[2099]) );
  XOR U12966 ( .A(n8869), .B(n8870), .Z(n8864) );
  ANDN U12967 ( .B(n8871), .A(n8872), .Z(n8869) );
  XNOR U12968 ( .A(b[2098]), .B(n8870), .Z(n8871) );
  XNOR U12969 ( .A(b[2098]), .B(n8872), .Z(c[2098]) );
  XOR U12970 ( .A(n8873), .B(n8874), .Z(n8870) );
  ANDN U12971 ( .B(n8875), .A(n8876), .Z(n8873) );
  XNOR U12972 ( .A(b[2097]), .B(n8874), .Z(n8875) );
  XNOR U12973 ( .A(b[2097]), .B(n8876), .Z(c[2097]) );
  XOR U12974 ( .A(n8877), .B(n8878), .Z(n8874) );
  ANDN U12975 ( .B(n8879), .A(n8880), .Z(n8877) );
  XNOR U12976 ( .A(b[2096]), .B(n8878), .Z(n8879) );
  XNOR U12977 ( .A(b[2096]), .B(n8880), .Z(c[2096]) );
  XOR U12978 ( .A(n8881), .B(n8882), .Z(n8878) );
  ANDN U12979 ( .B(n8883), .A(n8884), .Z(n8881) );
  XNOR U12980 ( .A(b[2095]), .B(n8882), .Z(n8883) );
  XNOR U12981 ( .A(b[2095]), .B(n8884), .Z(c[2095]) );
  XOR U12982 ( .A(n8885), .B(n8886), .Z(n8882) );
  ANDN U12983 ( .B(n8887), .A(n8888), .Z(n8885) );
  XNOR U12984 ( .A(b[2094]), .B(n8886), .Z(n8887) );
  XNOR U12985 ( .A(b[2094]), .B(n8888), .Z(c[2094]) );
  XOR U12986 ( .A(n8889), .B(n8890), .Z(n8886) );
  ANDN U12987 ( .B(n8891), .A(n8892), .Z(n8889) );
  XNOR U12988 ( .A(b[2093]), .B(n8890), .Z(n8891) );
  XNOR U12989 ( .A(b[2093]), .B(n8892), .Z(c[2093]) );
  XOR U12990 ( .A(n8893), .B(n8894), .Z(n8890) );
  ANDN U12991 ( .B(n8895), .A(n8896), .Z(n8893) );
  XNOR U12992 ( .A(b[2092]), .B(n8894), .Z(n8895) );
  XNOR U12993 ( .A(b[2092]), .B(n8896), .Z(c[2092]) );
  XOR U12994 ( .A(n8897), .B(n8898), .Z(n8894) );
  ANDN U12995 ( .B(n8899), .A(n8900), .Z(n8897) );
  XNOR U12996 ( .A(b[2091]), .B(n8898), .Z(n8899) );
  XNOR U12997 ( .A(b[2091]), .B(n8900), .Z(c[2091]) );
  XOR U12998 ( .A(n8901), .B(n8902), .Z(n8898) );
  ANDN U12999 ( .B(n8903), .A(n8904), .Z(n8901) );
  XNOR U13000 ( .A(b[2090]), .B(n8902), .Z(n8903) );
  XNOR U13001 ( .A(b[2090]), .B(n8904), .Z(c[2090]) );
  XOR U13002 ( .A(n8905), .B(n8906), .Z(n8902) );
  ANDN U13003 ( .B(n8907), .A(n8908), .Z(n8905) );
  XNOR U13004 ( .A(b[2089]), .B(n8906), .Z(n8907) );
  XNOR U13005 ( .A(b[208]), .B(n8909), .Z(c[208]) );
  XNOR U13006 ( .A(b[2089]), .B(n8908), .Z(c[2089]) );
  XOR U13007 ( .A(n8910), .B(n8911), .Z(n8906) );
  ANDN U13008 ( .B(n8912), .A(n8913), .Z(n8910) );
  XNOR U13009 ( .A(b[2088]), .B(n8911), .Z(n8912) );
  XNOR U13010 ( .A(b[2088]), .B(n8913), .Z(c[2088]) );
  XOR U13011 ( .A(n8914), .B(n8915), .Z(n8911) );
  ANDN U13012 ( .B(n8916), .A(n8917), .Z(n8914) );
  XNOR U13013 ( .A(b[2087]), .B(n8915), .Z(n8916) );
  XNOR U13014 ( .A(b[2087]), .B(n8917), .Z(c[2087]) );
  XOR U13015 ( .A(n8918), .B(n8919), .Z(n8915) );
  ANDN U13016 ( .B(n8920), .A(n8921), .Z(n8918) );
  XNOR U13017 ( .A(b[2086]), .B(n8919), .Z(n8920) );
  XNOR U13018 ( .A(b[2086]), .B(n8921), .Z(c[2086]) );
  XOR U13019 ( .A(n8922), .B(n8923), .Z(n8919) );
  ANDN U13020 ( .B(n8924), .A(n8925), .Z(n8922) );
  XNOR U13021 ( .A(b[2085]), .B(n8923), .Z(n8924) );
  XNOR U13022 ( .A(b[2085]), .B(n8925), .Z(c[2085]) );
  XOR U13023 ( .A(n8926), .B(n8927), .Z(n8923) );
  ANDN U13024 ( .B(n8928), .A(n8929), .Z(n8926) );
  XNOR U13025 ( .A(b[2084]), .B(n8927), .Z(n8928) );
  XNOR U13026 ( .A(b[2084]), .B(n8929), .Z(c[2084]) );
  XOR U13027 ( .A(n8930), .B(n8931), .Z(n8927) );
  ANDN U13028 ( .B(n8932), .A(n8933), .Z(n8930) );
  XNOR U13029 ( .A(b[2083]), .B(n8931), .Z(n8932) );
  XNOR U13030 ( .A(b[2083]), .B(n8933), .Z(c[2083]) );
  XOR U13031 ( .A(n8934), .B(n8935), .Z(n8931) );
  ANDN U13032 ( .B(n8936), .A(n8937), .Z(n8934) );
  XNOR U13033 ( .A(b[2082]), .B(n8935), .Z(n8936) );
  XNOR U13034 ( .A(b[2082]), .B(n8937), .Z(c[2082]) );
  XOR U13035 ( .A(n8938), .B(n8939), .Z(n8935) );
  ANDN U13036 ( .B(n8940), .A(n8941), .Z(n8938) );
  XNOR U13037 ( .A(b[2081]), .B(n8939), .Z(n8940) );
  XNOR U13038 ( .A(b[2081]), .B(n8941), .Z(c[2081]) );
  XOR U13039 ( .A(n8942), .B(n8943), .Z(n8939) );
  ANDN U13040 ( .B(n8944), .A(n8945), .Z(n8942) );
  XNOR U13041 ( .A(b[2080]), .B(n8943), .Z(n8944) );
  XNOR U13042 ( .A(b[2080]), .B(n8945), .Z(c[2080]) );
  XOR U13043 ( .A(n8946), .B(n8947), .Z(n8943) );
  ANDN U13044 ( .B(n8948), .A(n8949), .Z(n8946) );
  XNOR U13045 ( .A(b[2079]), .B(n8947), .Z(n8948) );
  XNOR U13046 ( .A(b[207]), .B(n8950), .Z(c[207]) );
  XNOR U13047 ( .A(b[2079]), .B(n8949), .Z(c[2079]) );
  XOR U13048 ( .A(n8951), .B(n8952), .Z(n8947) );
  ANDN U13049 ( .B(n8953), .A(n8954), .Z(n8951) );
  XNOR U13050 ( .A(b[2078]), .B(n8952), .Z(n8953) );
  XNOR U13051 ( .A(b[2078]), .B(n8954), .Z(c[2078]) );
  XOR U13052 ( .A(n8955), .B(n8956), .Z(n8952) );
  ANDN U13053 ( .B(n8957), .A(n8958), .Z(n8955) );
  XNOR U13054 ( .A(b[2077]), .B(n8956), .Z(n8957) );
  XNOR U13055 ( .A(b[2077]), .B(n8958), .Z(c[2077]) );
  XOR U13056 ( .A(n8959), .B(n8960), .Z(n8956) );
  ANDN U13057 ( .B(n8961), .A(n8962), .Z(n8959) );
  XNOR U13058 ( .A(b[2076]), .B(n8960), .Z(n8961) );
  XNOR U13059 ( .A(b[2076]), .B(n8962), .Z(c[2076]) );
  XOR U13060 ( .A(n8963), .B(n8964), .Z(n8960) );
  ANDN U13061 ( .B(n8965), .A(n8966), .Z(n8963) );
  XNOR U13062 ( .A(b[2075]), .B(n8964), .Z(n8965) );
  XNOR U13063 ( .A(b[2075]), .B(n8966), .Z(c[2075]) );
  XOR U13064 ( .A(n8967), .B(n8968), .Z(n8964) );
  ANDN U13065 ( .B(n8969), .A(n8970), .Z(n8967) );
  XNOR U13066 ( .A(b[2074]), .B(n8968), .Z(n8969) );
  XNOR U13067 ( .A(b[2074]), .B(n8970), .Z(c[2074]) );
  XOR U13068 ( .A(n8971), .B(n8972), .Z(n8968) );
  ANDN U13069 ( .B(n8973), .A(n8974), .Z(n8971) );
  XNOR U13070 ( .A(b[2073]), .B(n8972), .Z(n8973) );
  XNOR U13071 ( .A(b[2073]), .B(n8974), .Z(c[2073]) );
  XOR U13072 ( .A(n8975), .B(n8976), .Z(n8972) );
  ANDN U13073 ( .B(n8977), .A(n8978), .Z(n8975) );
  XNOR U13074 ( .A(b[2072]), .B(n8976), .Z(n8977) );
  XNOR U13075 ( .A(b[2072]), .B(n8978), .Z(c[2072]) );
  XOR U13076 ( .A(n8979), .B(n8980), .Z(n8976) );
  ANDN U13077 ( .B(n8981), .A(n8982), .Z(n8979) );
  XNOR U13078 ( .A(b[2071]), .B(n8980), .Z(n8981) );
  XNOR U13079 ( .A(b[2071]), .B(n8982), .Z(c[2071]) );
  XOR U13080 ( .A(n8983), .B(n8984), .Z(n8980) );
  ANDN U13081 ( .B(n8985), .A(n8986), .Z(n8983) );
  XNOR U13082 ( .A(b[2070]), .B(n8984), .Z(n8985) );
  XNOR U13083 ( .A(b[2070]), .B(n8986), .Z(c[2070]) );
  XOR U13084 ( .A(n8987), .B(n8988), .Z(n8984) );
  ANDN U13085 ( .B(n8989), .A(n8990), .Z(n8987) );
  XNOR U13086 ( .A(b[2069]), .B(n8988), .Z(n8989) );
  XNOR U13087 ( .A(b[206]), .B(n8991), .Z(c[206]) );
  XNOR U13088 ( .A(b[2069]), .B(n8990), .Z(c[2069]) );
  XOR U13089 ( .A(n8992), .B(n8993), .Z(n8988) );
  ANDN U13090 ( .B(n8994), .A(n8995), .Z(n8992) );
  XNOR U13091 ( .A(b[2068]), .B(n8993), .Z(n8994) );
  XNOR U13092 ( .A(b[2068]), .B(n8995), .Z(c[2068]) );
  XOR U13093 ( .A(n8996), .B(n8997), .Z(n8993) );
  ANDN U13094 ( .B(n8998), .A(n8999), .Z(n8996) );
  XNOR U13095 ( .A(b[2067]), .B(n8997), .Z(n8998) );
  XNOR U13096 ( .A(b[2067]), .B(n8999), .Z(c[2067]) );
  XOR U13097 ( .A(n9000), .B(n9001), .Z(n8997) );
  ANDN U13098 ( .B(n9002), .A(n9003), .Z(n9000) );
  XNOR U13099 ( .A(b[2066]), .B(n9001), .Z(n9002) );
  XNOR U13100 ( .A(b[2066]), .B(n9003), .Z(c[2066]) );
  XOR U13101 ( .A(n9004), .B(n9005), .Z(n9001) );
  ANDN U13102 ( .B(n9006), .A(n9007), .Z(n9004) );
  XNOR U13103 ( .A(b[2065]), .B(n9005), .Z(n9006) );
  XNOR U13104 ( .A(b[2065]), .B(n9007), .Z(c[2065]) );
  XOR U13105 ( .A(n9008), .B(n9009), .Z(n9005) );
  ANDN U13106 ( .B(n9010), .A(n9011), .Z(n9008) );
  XNOR U13107 ( .A(b[2064]), .B(n9009), .Z(n9010) );
  XNOR U13108 ( .A(b[2064]), .B(n9011), .Z(c[2064]) );
  XOR U13109 ( .A(n9012), .B(n9013), .Z(n9009) );
  ANDN U13110 ( .B(n9014), .A(n9015), .Z(n9012) );
  XNOR U13111 ( .A(b[2063]), .B(n9013), .Z(n9014) );
  XNOR U13112 ( .A(b[2063]), .B(n9015), .Z(c[2063]) );
  XOR U13113 ( .A(n9016), .B(n9017), .Z(n9013) );
  ANDN U13114 ( .B(n9018), .A(n9019), .Z(n9016) );
  XNOR U13115 ( .A(b[2062]), .B(n9017), .Z(n9018) );
  XNOR U13116 ( .A(b[2062]), .B(n9019), .Z(c[2062]) );
  XOR U13117 ( .A(n9020), .B(n9021), .Z(n9017) );
  ANDN U13118 ( .B(n9022), .A(n9023), .Z(n9020) );
  XNOR U13119 ( .A(b[2061]), .B(n9021), .Z(n9022) );
  XNOR U13120 ( .A(b[2061]), .B(n9023), .Z(c[2061]) );
  XOR U13121 ( .A(n9024), .B(n9025), .Z(n9021) );
  ANDN U13122 ( .B(n9026), .A(n9027), .Z(n9024) );
  XNOR U13123 ( .A(b[2060]), .B(n9025), .Z(n9026) );
  XNOR U13124 ( .A(b[2060]), .B(n9027), .Z(c[2060]) );
  XOR U13125 ( .A(n9028), .B(n9029), .Z(n9025) );
  ANDN U13126 ( .B(n9030), .A(n9031), .Z(n9028) );
  XNOR U13127 ( .A(b[2059]), .B(n9029), .Z(n9030) );
  XNOR U13128 ( .A(b[205]), .B(n9032), .Z(c[205]) );
  XNOR U13129 ( .A(b[2059]), .B(n9031), .Z(c[2059]) );
  XOR U13130 ( .A(n9033), .B(n9034), .Z(n9029) );
  ANDN U13131 ( .B(n9035), .A(n9036), .Z(n9033) );
  XNOR U13132 ( .A(b[2058]), .B(n9034), .Z(n9035) );
  XNOR U13133 ( .A(b[2058]), .B(n9036), .Z(c[2058]) );
  XOR U13134 ( .A(n9037), .B(n9038), .Z(n9034) );
  ANDN U13135 ( .B(n9039), .A(n9040), .Z(n9037) );
  XNOR U13136 ( .A(b[2057]), .B(n9038), .Z(n9039) );
  XNOR U13137 ( .A(b[2057]), .B(n9040), .Z(c[2057]) );
  XOR U13138 ( .A(n9041), .B(n9042), .Z(n9038) );
  ANDN U13139 ( .B(n9043), .A(n9044), .Z(n9041) );
  XNOR U13140 ( .A(b[2056]), .B(n9042), .Z(n9043) );
  XNOR U13141 ( .A(b[2056]), .B(n9044), .Z(c[2056]) );
  XOR U13142 ( .A(n9045), .B(n9046), .Z(n9042) );
  ANDN U13143 ( .B(n9047), .A(n9048), .Z(n9045) );
  XNOR U13144 ( .A(b[2055]), .B(n9046), .Z(n9047) );
  XNOR U13145 ( .A(b[2055]), .B(n9048), .Z(c[2055]) );
  XOR U13146 ( .A(n9049), .B(n9050), .Z(n9046) );
  ANDN U13147 ( .B(n9051), .A(n9052), .Z(n9049) );
  XNOR U13148 ( .A(b[2054]), .B(n9050), .Z(n9051) );
  XNOR U13149 ( .A(b[2054]), .B(n9052), .Z(c[2054]) );
  XOR U13150 ( .A(n9053), .B(n9054), .Z(n9050) );
  ANDN U13151 ( .B(n9055), .A(n9056), .Z(n9053) );
  XNOR U13152 ( .A(b[2053]), .B(n9054), .Z(n9055) );
  XNOR U13153 ( .A(b[2053]), .B(n9056), .Z(c[2053]) );
  XOR U13154 ( .A(n9057), .B(n9058), .Z(n9054) );
  ANDN U13155 ( .B(n9059), .A(n9060), .Z(n9057) );
  XNOR U13156 ( .A(b[2052]), .B(n9058), .Z(n9059) );
  XNOR U13157 ( .A(b[2052]), .B(n9060), .Z(c[2052]) );
  XOR U13158 ( .A(n9061), .B(n9062), .Z(n9058) );
  ANDN U13159 ( .B(n9063), .A(n9064), .Z(n9061) );
  XNOR U13160 ( .A(b[2051]), .B(n9062), .Z(n9063) );
  XNOR U13161 ( .A(b[2051]), .B(n9064), .Z(c[2051]) );
  XOR U13162 ( .A(n9065), .B(n9066), .Z(n9062) );
  ANDN U13163 ( .B(n9067), .A(n9068), .Z(n9065) );
  XNOR U13164 ( .A(b[2050]), .B(n9066), .Z(n9067) );
  XNOR U13165 ( .A(b[2050]), .B(n9068), .Z(c[2050]) );
  XOR U13166 ( .A(n9069), .B(n9070), .Z(n9066) );
  ANDN U13167 ( .B(n9071), .A(n9072), .Z(n9069) );
  XNOR U13168 ( .A(b[2049]), .B(n9070), .Z(n9071) );
  XNOR U13169 ( .A(b[204]), .B(n9073), .Z(c[204]) );
  XNOR U13170 ( .A(b[2049]), .B(n9072), .Z(c[2049]) );
  XOR U13171 ( .A(n9074), .B(n9075), .Z(n9070) );
  ANDN U13172 ( .B(n9076), .A(n9077), .Z(n9074) );
  XNOR U13173 ( .A(b[2048]), .B(n9075), .Z(n9076) );
  XNOR U13174 ( .A(b[2048]), .B(n9077), .Z(c[2048]) );
  XOR U13175 ( .A(n9078), .B(n9079), .Z(n9075) );
  ANDN U13176 ( .B(n9080), .A(n9081), .Z(n9078) );
  XNOR U13177 ( .A(b[2047]), .B(n9079), .Z(n9080) );
  XNOR U13178 ( .A(b[2047]), .B(n9081), .Z(c[2047]) );
  XOR U13179 ( .A(n9082), .B(n9083), .Z(n9079) );
  ANDN U13180 ( .B(n9084), .A(n9085), .Z(n9082) );
  XNOR U13181 ( .A(b[2046]), .B(n9083), .Z(n9084) );
  XNOR U13182 ( .A(b[2046]), .B(n9085), .Z(c[2046]) );
  XOR U13183 ( .A(n9086), .B(n9087), .Z(n9083) );
  ANDN U13184 ( .B(n9088), .A(n9089), .Z(n9086) );
  XNOR U13185 ( .A(b[2045]), .B(n9087), .Z(n9088) );
  XNOR U13186 ( .A(b[2045]), .B(n9089), .Z(c[2045]) );
  XOR U13187 ( .A(n9090), .B(n9091), .Z(n9087) );
  ANDN U13188 ( .B(n9092), .A(n9093), .Z(n9090) );
  XNOR U13189 ( .A(b[2044]), .B(n9091), .Z(n9092) );
  XNOR U13190 ( .A(b[2044]), .B(n9093), .Z(c[2044]) );
  XOR U13191 ( .A(n9094), .B(n9095), .Z(n9091) );
  ANDN U13192 ( .B(n9096), .A(n9097), .Z(n9094) );
  XNOR U13193 ( .A(b[2043]), .B(n9095), .Z(n9096) );
  XNOR U13194 ( .A(b[2043]), .B(n9097), .Z(c[2043]) );
  XOR U13195 ( .A(n9098), .B(n9099), .Z(n9095) );
  ANDN U13196 ( .B(n9100), .A(n9101), .Z(n9098) );
  XNOR U13197 ( .A(b[2042]), .B(n9099), .Z(n9100) );
  XNOR U13198 ( .A(b[2042]), .B(n9101), .Z(c[2042]) );
  XOR U13199 ( .A(n9102), .B(n9103), .Z(n9099) );
  ANDN U13200 ( .B(n9104), .A(n9105), .Z(n9102) );
  XNOR U13201 ( .A(b[2041]), .B(n9103), .Z(n9104) );
  XNOR U13202 ( .A(b[2041]), .B(n9105), .Z(c[2041]) );
  XOR U13203 ( .A(n9106), .B(n9107), .Z(n9103) );
  ANDN U13204 ( .B(n9108), .A(n9109), .Z(n9106) );
  XNOR U13205 ( .A(b[2040]), .B(n9107), .Z(n9108) );
  XNOR U13206 ( .A(b[2040]), .B(n9109), .Z(c[2040]) );
  XOR U13207 ( .A(n9110), .B(n9111), .Z(n9107) );
  ANDN U13208 ( .B(n9112), .A(n9113), .Z(n9110) );
  XNOR U13209 ( .A(b[2039]), .B(n9111), .Z(n9112) );
  XNOR U13210 ( .A(b[203]), .B(n9114), .Z(c[203]) );
  XNOR U13211 ( .A(b[2039]), .B(n9113), .Z(c[2039]) );
  XOR U13212 ( .A(n9115), .B(n9116), .Z(n9111) );
  ANDN U13213 ( .B(n9117), .A(n9118), .Z(n9115) );
  XNOR U13214 ( .A(b[2038]), .B(n9116), .Z(n9117) );
  XNOR U13215 ( .A(b[2038]), .B(n9118), .Z(c[2038]) );
  XOR U13216 ( .A(n9119), .B(n9120), .Z(n9116) );
  ANDN U13217 ( .B(n9121), .A(n9122), .Z(n9119) );
  XNOR U13218 ( .A(b[2037]), .B(n9120), .Z(n9121) );
  XNOR U13219 ( .A(b[2037]), .B(n9122), .Z(c[2037]) );
  XOR U13220 ( .A(n9123), .B(n9124), .Z(n9120) );
  ANDN U13221 ( .B(n9125), .A(n9126), .Z(n9123) );
  XNOR U13222 ( .A(b[2036]), .B(n9124), .Z(n9125) );
  XNOR U13223 ( .A(b[2036]), .B(n9126), .Z(c[2036]) );
  XOR U13224 ( .A(n9127), .B(n9128), .Z(n9124) );
  ANDN U13225 ( .B(n9129), .A(n9130), .Z(n9127) );
  XNOR U13226 ( .A(b[2035]), .B(n9128), .Z(n9129) );
  XNOR U13227 ( .A(b[2035]), .B(n9130), .Z(c[2035]) );
  XOR U13228 ( .A(n9131), .B(n9132), .Z(n9128) );
  ANDN U13229 ( .B(n9133), .A(n9134), .Z(n9131) );
  XNOR U13230 ( .A(b[2034]), .B(n9132), .Z(n9133) );
  XNOR U13231 ( .A(b[2034]), .B(n9134), .Z(c[2034]) );
  XOR U13232 ( .A(n9135), .B(n9136), .Z(n9132) );
  ANDN U13233 ( .B(n9137), .A(n9138), .Z(n9135) );
  XNOR U13234 ( .A(b[2033]), .B(n9136), .Z(n9137) );
  XNOR U13235 ( .A(b[2033]), .B(n9138), .Z(c[2033]) );
  XOR U13236 ( .A(n9139), .B(n9140), .Z(n9136) );
  ANDN U13237 ( .B(n9141), .A(n9142), .Z(n9139) );
  XNOR U13238 ( .A(b[2032]), .B(n9140), .Z(n9141) );
  XNOR U13239 ( .A(b[2032]), .B(n9142), .Z(c[2032]) );
  XOR U13240 ( .A(n9143), .B(n9144), .Z(n9140) );
  ANDN U13241 ( .B(n9145), .A(n9146), .Z(n9143) );
  XNOR U13242 ( .A(b[2031]), .B(n9144), .Z(n9145) );
  XNOR U13243 ( .A(b[2031]), .B(n9146), .Z(c[2031]) );
  XOR U13244 ( .A(n9147), .B(n9148), .Z(n9144) );
  ANDN U13245 ( .B(n9149), .A(n9150), .Z(n9147) );
  XNOR U13246 ( .A(b[2030]), .B(n9148), .Z(n9149) );
  XNOR U13247 ( .A(b[2030]), .B(n9150), .Z(c[2030]) );
  XOR U13248 ( .A(n9151), .B(n9152), .Z(n9148) );
  ANDN U13249 ( .B(n9153), .A(n9154), .Z(n9151) );
  XNOR U13250 ( .A(b[2029]), .B(n9152), .Z(n9153) );
  XNOR U13251 ( .A(b[202]), .B(n9155), .Z(c[202]) );
  XNOR U13252 ( .A(b[2029]), .B(n9154), .Z(c[2029]) );
  XOR U13253 ( .A(n9156), .B(n9157), .Z(n9152) );
  ANDN U13254 ( .B(n9158), .A(n9159), .Z(n9156) );
  XNOR U13255 ( .A(b[2028]), .B(n9157), .Z(n9158) );
  XNOR U13256 ( .A(b[2028]), .B(n9159), .Z(c[2028]) );
  XOR U13257 ( .A(n9160), .B(n9161), .Z(n9157) );
  ANDN U13258 ( .B(n9162), .A(n9163), .Z(n9160) );
  XNOR U13259 ( .A(b[2027]), .B(n9161), .Z(n9162) );
  XNOR U13260 ( .A(b[2027]), .B(n9163), .Z(c[2027]) );
  XOR U13261 ( .A(n9164), .B(n9165), .Z(n9161) );
  ANDN U13262 ( .B(n9166), .A(n9167), .Z(n9164) );
  XNOR U13263 ( .A(b[2026]), .B(n9165), .Z(n9166) );
  XNOR U13264 ( .A(b[2026]), .B(n9167), .Z(c[2026]) );
  XOR U13265 ( .A(n9168), .B(n9169), .Z(n9165) );
  ANDN U13266 ( .B(n9170), .A(n9171), .Z(n9168) );
  XNOR U13267 ( .A(b[2025]), .B(n9169), .Z(n9170) );
  XNOR U13268 ( .A(b[2025]), .B(n9171), .Z(c[2025]) );
  XOR U13269 ( .A(n9172), .B(n9173), .Z(n9169) );
  ANDN U13270 ( .B(n9174), .A(n9175), .Z(n9172) );
  XNOR U13271 ( .A(b[2024]), .B(n9173), .Z(n9174) );
  XNOR U13272 ( .A(b[2024]), .B(n9175), .Z(c[2024]) );
  XOR U13273 ( .A(n9176), .B(n9177), .Z(n9173) );
  ANDN U13274 ( .B(n9178), .A(n9179), .Z(n9176) );
  XNOR U13275 ( .A(b[2023]), .B(n9177), .Z(n9178) );
  XNOR U13276 ( .A(b[2023]), .B(n9179), .Z(c[2023]) );
  XOR U13277 ( .A(n9180), .B(n9181), .Z(n9177) );
  ANDN U13278 ( .B(n9182), .A(n9183), .Z(n9180) );
  XNOR U13279 ( .A(b[2022]), .B(n9181), .Z(n9182) );
  XNOR U13280 ( .A(b[2022]), .B(n9183), .Z(c[2022]) );
  XOR U13281 ( .A(n9184), .B(n9185), .Z(n9181) );
  ANDN U13282 ( .B(n9186), .A(n9187), .Z(n9184) );
  XNOR U13283 ( .A(b[2021]), .B(n9185), .Z(n9186) );
  XNOR U13284 ( .A(b[2021]), .B(n9187), .Z(c[2021]) );
  XOR U13285 ( .A(n9188), .B(n9189), .Z(n9185) );
  ANDN U13286 ( .B(n9190), .A(n9191), .Z(n9188) );
  XNOR U13287 ( .A(b[2020]), .B(n9189), .Z(n9190) );
  XNOR U13288 ( .A(b[2020]), .B(n9191), .Z(c[2020]) );
  XOR U13289 ( .A(n9192), .B(n9193), .Z(n9189) );
  ANDN U13290 ( .B(n9194), .A(n9195), .Z(n9192) );
  XNOR U13291 ( .A(b[2019]), .B(n9193), .Z(n9194) );
  XNOR U13292 ( .A(b[201]), .B(n9196), .Z(c[201]) );
  XNOR U13293 ( .A(b[2019]), .B(n9195), .Z(c[2019]) );
  XOR U13294 ( .A(n9197), .B(n9198), .Z(n9193) );
  ANDN U13295 ( .B(n9199), .A(n9200), .Z(n9197) );
  XNOR U13296 ( .A(b[2018]), .B(n9198), .Z(n9199) );
  XNOR U13297 ( .A(b[2018]), .B(n9200), .Z(c[2018]) );
  XOR U13298 ( .A(n9201), .B(n9202), .Z(n9198) );
  ANDN U13299 ( .B(n9203), .A(n9204), .Z(n9201) );
  XNOR U13300 ( .A(b[2017]), .B(n9202), .Z(n9203) );
  XNOR U13301 ( .A(b[2017]), .B(n9204), .Z(c[2017]) );
  XOR U13302 ( .A(n9205), .B(n9206), .Z(n9202) );
  ANDN U13303 ( .B(n9207), .A(n9208), .Z(n9205) );
  XNOR U13304 ( .A(b[2016]), .B(n9206), .Z(n9207) );
  XNOR U13305 ( .A(b[2016]), .B(n9208), .Z(c[2016]) );
  XOR U13306 ( .A(n9209), .B(n9210), .Z(n9206) );
  ANDN U13307 ( .B(n9211), .A(n9212), .Z(n9209) );
  XNOR U13308 ( .A(b[2015]), .B(n9210), .Z(n9211) );
  XNOR U13309 ( .A(b[2015]), .B(n9212), .Z(c[2015]) );
  XOR U13310 ( .A(n9213), .B(n9214), .Z(n9210) );
  ANDN U13311 ( .B(n9215), .A(n9216), .Z(n9213) );
  XNOR U13312 ( .A(b[2014]), .B(n9214), .Z(n9215) );
  XNOR U13313 ( .A(b[2014]), .B(n9216), .Z(c[2014]) );
  XOR U13314 ( .A(n9217), .B(n9218), .Z(n9214) );
  ANDN U13315 ( .B(n9219), .A(n9220), .Z(n9217) );
  XNOR U13316 ( .A(b[2013]), .B(n9218), .Z(n9219) );
  XNOR U13317 ( .A(b[2013]), .B(n9220), .Z(c[2013]) );
  XOR U13318 ( .A(n9221), .B(n9222), .Z(n9218) );
  ANDN U13319 ( .B(n9223), .A(n9224), .Z(n9221) );
  XNOR U13320 ( .A(b[2012]), .B(n9222), .Z(n9223) );
  XNOR U13321 ( .A(b[2012]), .B(n9224), .Z(c[2012]) );
  XOR U13322 ( .A(n9225), .B(n9226), .Z(n9222) );
  ANDN U13323 ( .B(n9227), .A(n9228), .Z(n9225) );
  XNOR U13324 ( .A(b[2011]), .B(n9226), .Z(n9227) );
  XNOR U13325 ( .A(b[2011]), .B(n9228), .Z(c[2011]) );
  XOR U13326 ( .A(n9229), .B(n9230), .Z(n9226) );
  ANDN U13327 ( .B(n9231), .A(n9232), .Z(n9229) );
  XNOR U13328 ( .A(b[2010]), .B(n9230), .Z(n9231) );
  XNOR U13329 ( .A(b[2010]), .B(n9232), .Z(c[2010]) );
  XOR U13330 ( .A(n9233), .B(n9234), .Z(n9230) );
  ANDN U13331 ( .B(n9235), .A(n9236), .Z(n9233) );
  XNOR U13332 ( .A(b[2009]), .B(n9234), .Z(n9235) );
  XNOR U13333 ( .A(b[200]), .B(n9237), .Z(c[200]) );
  XNOR U13334 ( .A(b[2009]), .B(n9236), .Z(c[2009]) );
  XOR U13335 ( .A(n9238), .B(n9239), .Z(n9234) );
  ANDN U13336 ( .B(n9240), .A(n9241), .Z(n9238) );
  XNOR U13337 ( .A(b[2008]), .B(n9239), .Z(n9240) );
  XNOR U13338 ( .A(b[2008]), .B(n9241), .Z(c[2008]) );
  XOR U13339 ( .A(n9242), .B(n9243), .Z(n9239) );
  ANDN U13340 ( .B(n9244), .A(n9245), .Z(n9242) );
  XNOR U13341 ( .A(b[2007]), .B(n9243), .Z(n9244) );
  XNOR U13342 ( .A(b[2007]), .B(n9245), .Z(c[2007]) );
  XOR U13343 ( .A(n9246), .B(n9247), .Z(n9243) );
  ANDN U13344 ( .B(n9248), .A(n9249), .Z(n9246) );
  XNOR U13345 ( .A(b[2006]), .B(n9247), .Z(n9248) );
  XNOR U13346 ( .A(b[2006]), .B(n9249), .Z(c[2006]) );
  XOR U13347 ( .A(n9250), .B(n9251), .Z(n9247) );
  ANDN U13348 ( .B(n9252), .A(n9253), .Z(n9250) );
  XNOR U13349 ( .A(b[2005]), .B(n9251), .Z(n9252) );
  XNOR U13350 ( .A(b[2005]), .B(n9253), .Z(c[2005]) );
  XOR U13351 ( .A(n9254), .B(n9255), .Z(n9251) );
  ANDN U13352 ( .B(n9256), .A(n9257), .Z(n9254) );
  XNOR U13353 ( .A(b[2004]), .B(n9255), .Z(n9256) );
  XNOR U13354 ( .A(b[2004]), .B(n9257), .Z(c[2004]) );
  XOR U13355 ( .A(n9258), .B(n9259), .Z(n9255) );
  ANDN U13356 ( .B(n9260), .A(n9261), .Z(n9258) );
  XNOR U13357 ( .A(b[2003]), .B(n9259), .Z(n9260) );
  XNOR U13358 ( .A(b[2003]), .B(n9261), .Z(c[2003]) );
  XOR U13359 ( .A(n9262), .B(n9263), .Z(n9259) );
  ANDN U13360 ( .B(n9264), .A(n9265), .Z(n9262) );
  XNOR U13361 ( .A(b[2002]), .B(n9263), .Z(n9264) );
  XNOR U13362 ( .A(b[2002]), .B(n9265), .Z(c[2002]) );
  XOR U13363 ( .A(n9266), .B(n9267), .Z(n9263) );
  ANDN U13364 ( .B(n9268), .A(n9269), .Z(n9266) );
  XNOR U13365 ( .A(b[2001]), .B(n9267), .Z(n9268) );
  XNOR U13366 ( .A(b[2001]), .B(n9269), .Z(c[2001]) );
  XOR U13367 ( .A(n9270), .B(n9271), .Z(n9267) );
  ANDN U13368 ( .B(n9272), .A(n9273), .Z(n9270) );
  XNOR U13369 ( .A(b[2000]), .B(n9271), .Z(n9272) );
  XNOR U13370 ( .A(b[2000]), .B(n9273), .Z(c[2000]) );
  XOR U13371 ( .A(n9274), .B(n9275), .Z(n9271) );
  ANDN U13372 ( .B(n9276), .A(n9277), .Z(n9274) );
  XNOR U13373 ( .A(b[1999]), .B(n9275), .Z(n9276) );
  XNOR U13374 ( .A(b[1]), .B(n9278), .Z(c[1]) );
  XNOR U13375 ( .A(b[19]), .B(n9279), .Z(c[19]) );
  XNOR U13376 ( .A(b[199]), .B(n9280), .Z(c[199]) );
  XNOR U13377 ( .A(b[1999]), .B(n9277), .Z(c[1999]) );
  XOR U13378 ( .A(n9281), .B(n9282), .Z(n9275) );
  ANDN U13379 ( .B(n9283), .A(n9284), .Z(n9281) );
  XNOR U13380 ( .A(b[1998]), .B(n9282), .Z(n9283) );
  XNOR U13381 ( .A(b[1998]), .B(n9284), .Z(c[1998]) );
  XOR U13382 ( .A(n9285), .B(n9286), .Z(n9282) );
  ANDN U13383 ( .B(n9287), .A(n9288), .Z(n9285) );
  XNOR U13384 ( .A(b[1997]), .B(n9286), .Z(n9287) );
  XNOR U13385 ( .A(b[1997]), .B(n9288), .Z(c[1997]) );
  XOR U13386 ( .A(n9289), .B(n9290), .Z(n9286) );
  ANDN U13387 ( .B(n9291), .A(n9292), .Z(n9289) );
  XNOR U13388 ( .A(b[1996]), .B(n9290), .Z(n9291) );
  XNOR U13389 ( .A(b[1996]), .B(n9292), .Z(c[1996]) );
  XOR U13390 ( .A(n9293), .B(n9294), .Z(n9290) );
  ANDN U13391 ( .B(n9295), .A(n9296), .Z(n9293) );
  XNOR U13392 ( .A(b[1995]), .B(n9294), .Z(n9295) );
  XNOR U13393 ( .A(b[1995]), .B(n9296), .Z(c[1995]) );
  XOR U13394 ( .A(n9297), .B(n9298), .Z(n9294) );
  ANDN U13395 ( .B(n9299), .A(n9300), .Z(n9297) );
  XNOR U13396 ( .A(b[1994]), .B(n9298), .Z(n9299) );
  XNOR U13397 ( .A(b[1994]), .B(n9300), .Z(c[1994]) );
  XOR U13398 ( .A(n9301), .B(n9302), .Z(n9298) );
  ANDN U13399 ( .B(n9303), .A(n9304), .Z(n9301) );
  XNOR U13400 ( .A(b[1993]), .B(n9302), .Z(n9303) );
  XNOR U13401 ( .A(b[1993]), .B(n9304), .Z(c[1993]) );
  XOR U13402 ( .A(n9305), .B(n9306), .Z(n9302) );
  ANDN U13403 ( .B(n9307), .A(n9308), .Z(n9305) );
  XNOR U13404 ( .A(b[1992]), .B(n9306), .Z(n9307) );
  XNOR U13405 ( .A(b[1992]), .B(n9308), .Z(c[1992]) );
  XOR U13406 ( .A(n9309), .B(n9310), .Z(n9306) );
  ANDN U13407 ( .B(n9311), .A(n9312), .Z(n9309) );
  XNOR U13408 ( .A(b[1991]), .B(n9310), .Z(n9311) );
  XNOR U13409 ( .A(b[1991]), .B(n9312), .Z(c[1991]) );
  XOR U13410 ( .A(n9313), .B(n9314), .Z(n9310) );
  ANDN U13411 ( .B(n9315), .A(n9316), .Z(n9313) );
  XNOR U13412 ( .A(b[1990]), .B(n9314), .Z(n9315) );
  XNOR U13413 ( .A(b[1990]), .B(n9316), .Z(c[1990]) );
  XOR U13414 ( .A(n9317), .B(n9318), .Z(n9314) );
  ANDN U13415 ( .B(n9319), .A(n9320), .Z(n9317) );
  XNOR U13416 ( .A(b[1989]), .B(n9318), .Z(n9319) );
  XNOR U13417 ( .A(b[198]), .B(n9321), .Z(c[198]) );
  XNOR U13418 ( .A(b[1989]), .B(n9320), .Z(c[1989]) );
  XOR U13419 ( .A(n9322), .B(n9323), .Z(n9318) );
  ANDN U13420 ( .B(n9324), .A(n9325), .Z(n9322) );
  XNOR U13421 ( .A(b[1988]), .B(n9323), .Z(n9324) );
  XNOR U13422 ( .A(b[1988]), .B(n9325), .Z(c[1988]) );
  XOR U13423 ( .A(n9326), .B(n9327), .Z(n9323) );
  ANDN U13424 ( .B(n9328), .A(n9329), .Z(n9326) );
  XNOR U13425 ( .A(b[1987]), .B(n9327), .Z(n9328) );
  XNOR U13426 ( .A(b[1987]), .B(n9329), .Z(c[1987]) );
  XOR U13427 ( .A(n9330), .B(n9331), .Z(n9327) );
  ANDN U13428 ( .B(n9332), .A(n9333), .Z(n9330) );
  XNOR U13429 ( .A(b[1986]), .B(n9331), .Z(n9332) );
  XNOR U13430 ( .A(b[1986]), .B(n9333), .Z(c[1986]) );
  XOR U13431 ( .A(n9334), .B(n9335), .Z(n9331) );
  ANDN U13432 ( .B(n9336), .A(n9337), .Z(n9334) );
  XNOR U13433 ( .A(b[1985]), .B(n9335), .Z(n9336) );
  XNOR U13434 ( .A(b[1985]), .B(n9337), .Z(c[1985]) );
  XOR U13435 ( .A(n9338), .B(n9339), .Z(n9335) );
  ANDN U13436 ( .B(n9340), .A(n9341), .Z(n9338) );
  XNOR U13437 ( .A(b[1984]), .B(n9339), .Z(n9340) );
  XNOR U13438 ( .A(b[1984]), .B(n9341), .Z(c[1984]) );
  XOR U13439 ( .A(n9342), .B(n9343), .Z(n9339) );
  ANDN U13440 ( .B(n9344), .A(n9345), .Z(n9342) );
  XNOR U13441 ( .A(b[1983]), .B(n9343), .Z(n9344) );
  XNOR U13442 ( .A(b[1983]), .B(n9345), .Z(c[1983]) );
  XOR U13443 ( .A(n9346), .B(n9347), .Z(n9343) );
  ANDN U13444 ( .B(n9348), .A(n9349), .Z(n9346) );
  XNOR U13445 ( .A(b[1982]), .B(n9347), .Z(n9348) );
  XNOR U13446 ( .A(b[1982]), .B(n9349), .Z(c[1982]) );
  XOR U13447 ( .A(n9350), .B(n9351), .Z(n9347) );
  ANDN U13448 ( .B(n9352), .A(n9353), .Z(n9350) );
  XNOR U13449 ( .A(b[1981]), .B(n9351), .Z(n9352) );
  XNOR U13450 ( .A(b[1981]), .B(n9353), .Z(c[1981]) );
  XOR U13451 ( .A(n9354), .B(n9355), .Z(n9351) );
  ANDN U13452 ( .B(n9356), .A(n9357), .Z(n9354) );
  XNOR U13453 ( .A(b[1980]), .B(n9355), .Z(n9356) );
  XNOR U13454 ( .A(b[1980]), .B(n9357), .Z(c[1980]) );
  XOR U13455 ( .A(n9358), .B(n9359), .Z(n9355) );
  ANDN U13456 ( .B(n9360), .A(n9361), .Z(n9358) );
  XNOR U13457 ( .A(b[1979]), .B(n9359), .Z(n9360) );
  XNOR U13458 ( .A(b[197]), .B(n9362), .Z(c[197]) );
  XNOR U13459 ( .A(b[1979]), .B(n9361), .Z(c[1979]) );
  XOR U13460 ( .A(n9363), .B(n9364), .Z(n9359) );
  ANDN U13461 ( .B(n9365), .A(n9366), .Z(n9363) );
  XNOR U13462 ( .A(b[1978]), .B(n9364), .Z(n9365) );
  XNOR U13463 ( .A(b[1978]), .B(n9366), .Z(c[1978]) );
  XOR U13464 ( .A(n9367), .B(n9368), .Z(n9364) );
  ANDN U13465 ( .B(n9369), .A(n9370), .Z(n9367) );
  XNOR U13466 ( .A(b[1977]), .B(n9368), .Z(n9369) );
  XNOR U13467 ( .A(b[1977]), .B(n9370), .Z(c[1977]) );
  XOR U13468 ( .A(n9371), .B(n9372), .Z(n9368) );
  ANDN U13469 ( .B(n9373), .A(n9374), .Z(n9371) );
  XNOR U13470 ( .A(b[1976]), .B(n9372), .Z(n9373) );
  XNOR U13471 ( .A(b[1976]), .B(n9374), .Z(c[1976]) );
  XOR U13472 ( .A(n9375), .B(n9376), .Z(n9372) );
  ANDN U13473 ( .B(n9377), .A(n9378), .Z(n9375) );
  XNOR U13474 ( .A(b[1975]), .B(n9376), .Z(n9377) );
  XNOR U13475 ( .A(b[1975]), .B(n9378), .Z(c[1975]) );
  XOR U13476 ( .A(n9379), .B(n9380), .Z(n9376) );
  ANDN U13477 ( .B(n9381), .A(n9382), .Z(n9379) );
  XNOR U13478 ( .A(b[1974]), .B(n9380), .Z(n9381) );
  XNOR U13479 ( .A(b[1974]), .B(n9382), .Z(c[1974]) );
  XOR U13480 ( .A(n9383), .B(n9384), .Z(n9380) );
  ANDN U13481 ( .B(n9385), .A(n9386), .Z(n9383) );
  XNOR U13482 ( .A(b[1973]), .B(n9384), .Z(n9385) );
  XNOR U13483 ( .A(b[1973]), .B(n9386), .Z(c[1973]) );
  XOR U13484 ( .A(n9387), .B(n9388), .Z(n9384) );
  ANDN U13485 ( .B(n9389), .A(n9390), .Z(n9387) );
  XNOR U13486 ( .A(b[1972]), .B(n9388), .Z(n9389) );
  XNOR U13487 ( .A(b[1972]), .B(n9390), .Z(c[1972]) );
  XOR U13488 ( .A(n9391), .B(n9392), .Z(n9388) );
  ANDN U13489 ( .B(n9393), .A(n9394), .Z(n9391) );
  XNOR U13490 ( .A(b[1971]), .B(n9392), .Z(n9393) );
  XNOR U13491 ( .A(b[1971]), .B(n9394), .Z(c[1971]) );
  XOR U13492 ( .A(n9395), .B(n9396), .Z(n9392) );
  ANDN U13493 ( .B(n9397), .A(n9398), .Z(n9395) );
  XNOR U13494 ( .A(b[1970]), .B(n9396), .Z(n9397) );
  XNOR U13495 ( .A(b[1970]), .B(n9398), .Z(c[1970]) );
  XOR U13496 ( .A(n9399), .B(n9400), .Z(n9396) );
  ANDN U13497 ( .B(n9401), .A(n9402), .Z(n9399) );
  XNOR U13498 ( .A(b[1969]), .B(n9400), .Z(n9401) );
  XNOR U13499 ( .A(b[196]), .B(n9403), .Z(c[196]) );
  XNOR U13500 ( .A(b[1969]), .B(n9402), .Z(c[1969]) );
  XOR U13501 ( .A(n9404), .B(n9405), .Z(n9400) );
  ANDN U13502 ( .B(n9406), .A(n9407), .Z(n9404) );
  XNOR U13503 ( .A(b[1968]), .B(n9405), .Z(n9406) );
  XNOR U13504 ( .A(b[1968]), .B(n9407), .Z(c[1968]) );
  XOR U13505 ( .A(n9408), .B(n9409), .Z(n9405) );
  ANDN U13506 ( .B(n9410), .A(n9411), .Z(n9408) );
  XNOR U13507 ( .A(b[1967]), .B(n9409), .Z(n9410) );
  XNOR U13508 ( .A(b[1967]), .B(n9411), .Z(c[1967]) );
  XOR U13509 ( .A(n9412), .B(n9413), .Z(n9409) );
  ANDN U13510 ( .B(n9414), .A(n9415), .Z(n9412) );
  XNOR U13511 ( .A(b[1966]), .B(n9413), .Z(n9414) );
  XNOR U13512 ( .A(b[1966]), .B(n9415), .Z(c[1966]) );
  XOR U13513 ( .A(n9416), .B(n9417), .Z(n9413) );
  ANDN U13514 ( .B(n9418), .A(n9419), .Z(n9416) );
  XNOR U13515 ( .A(b[1965]), .B(n9417), .Z(n9418) );
  XNOR U13516 ( .A(b[1965]), .B(n9419), .Z(c[1965]) );
  XOR U13517 ( .A(n9420), .B(n9421), .Z(n9417) );
  ANDN U13518 ( .B(n9422), .A(n9423), .Z(n9420) );
  XNOR U13519 ( .A(b[1964]), .B(n9421), .Z(n9422) );
  XNOR U13520 ( .A(b[1964]), .B(n9423), .Z(c[1964]) );
  XOR U13521 ( .A(n9424), .B(n9425), .Z(n9421) );
  ANDN U13522 ( .B(n9426), .A(n9427), .Z(n9424) );
  XNOR U13523 ( .A(b[1963]), .B(n9425), .Z(n9426) );
  XNOR U13524 ( .A(b[1963]), .B(n9427), .Z(c[1963]) );
  XOR U13525 ( .A(n9428), .B(n9429), .Z(n9425) );
  ANDN U13526 ( .B(n9430), .A(n9431), .Z(n9428) );
  XNOR U13527 ( .A(b[1962]), .B(n9429), .Z(n9430) );
  XNOR U13528 ( .A(b[1962]), .B(n9431), .Z(c[1962]) );
  XOR U13529 ( .A(n9432), .B(n9433), .Z(n9429) );
  ANDN U13530 ( .B(n9434), .A(n9435), .Z(n9432) );
  XNOR U13531 ( .A(b[1961]), .B(n9433), .Z(n9434) );
  XNOR U13532 ( .A(b[1961]), .B(n9435), .Z(c[1961]) );
  XOR U13533 ( .A(n9436), .B(n9437), .Z(n9433) );
  ANDN U13534 ( .B(n9438), .A(n9439), .Z(n9436) );
  XNOR U13535 ( .A(b[1960]), .B(n9437), .Z(n9438) );
  XNOR U13536 ( .A(b[1960]), .B(n9439), .Z(c[1960]) );
  XOR U13537 ( .A(n9440), .B(n9441), .Z(n9437) );
  ANDN U13538 ( .B(n9442), .A(n9443), .Z(n9440) );
  XNOR U13539 ( .A(b[1959]), .B(n9441), .Z(n9442) );
  XNOR U13540 ( .A(b[195]), .B(n9444), .Z(c[195]) );
  XNOR U13541 ( .A(b[1959]), .B(n9443), .Z(c[1959]) );
  XOR U13542 ( .A(n9445), .B(n9446), .Z(n9441) );
  ANDN U13543 ( .B(n9447), .A(n9448), .Z(n9445) );
  XNOR U13544 ( .A(b[1958]), .B(n9446), .Z(n9447) );
  XNOR U13545 ( .A(b[1958]), .B(n9448), .Z(c[1958]) );
  XOR U13546 ( .A(n9449), .B(n9450), .Z(n9446) );
  ANDN U13547 ( .B(n9451), .A(n9452), .Z(n9449) );
  XNOR U13548 ( .A(b[1957]), .B(n9450), .Z(n9451) );
  XNOR U13549 ( .A(b[1957]), .B(n9452), .Z(c[1957]) );
  XOR U13550 ( .A(n9453), .B(n9454), .Z(n9450) );
  ANDN U13551 ( .B(n9455), .A(n9456), .Z(n9453) );
  XNOR U13552 ( .A(b[1956]), .B(n9454), .Z(n9455) );
  XNOR U13553 ( .A(b[1956]), .B(n9456), .Z(c[1956]) );
  XOR U13554 ( .A(n9457), .B(n9458), .Z(n9454) );
  ANDN U13555 ( .B(n9459), .A(n9460), .Z(n9457) );
  XNOR U13556 ( .A(b[1955]), .B(n9458), .Z(n9459) );
  XNOR U13557 ( .A(b[1955]), .B(n9460), .Z(c[1955]) );
  XOR U13558 ( .A(n9461), .B(n9462), .Z(n9458) );
  ANDN U13559 ( .B(n9463), .A(n9464), .Z(n9461) );
  XNOR U13560 ( .A(b[1954]), .B(n9462), .Z(n9463) );
  XNOR U13561 ( .A(b[1954]), .B(n9464), .Z(c[1954]) );
  XOR U13562 ( .A(n9465), .B(n9466), .Z(n9462) );
  ANDN U13563 ( .B(n9467), .A(n9468), .Z(n9465) );
  XNOR U13564 ( .A(b[1953]), .B(n9466), .Z(n9467) );
  XNOR U13565 ( .A(b[1953]), .B(n9468), .Z(c[1953]) );
  XOR U13566 ( .A(n9469), .B(n9470), .Z(n9466) );
  ANDN U13567 ( .B(n9471), .A(n9472), .Z(n9469) );
  XNOR U13568 ( .A(b[1952]), .B(n9470), .Z(n9471) );
  XNOR U13569 ( .A(b[1952]), .B(n9472), .Z(c[1952]) );
  XOR U13570 ( .A(n9473), .B(n9474), .Z(n9470) );
  ANDN U13571 ( .B(n9475), .A(n9476), .Z(n9473) );
  XNOR U13572 ( .A(b[1951]), .B(n9474), .Z(n9475) );
  XNOR U13573 ( .A(b[1951]), .B(n9476), .Z(c[1951]) );
  XOR U13574 ( .A(n9477), .B(n9478), .Z(n9474) );
  ANDN U13575 ( .B(n9479), .A(n9480), .Z(n9477) );
  XNOR U13576 ( .A(b[1950]), .B(n9478), .Z(n9479) );
  XNOR U13577 ( .A(b[1950]), .B(n9480), .Z(c[1950]) );
  XOR U13578 ( .A(n9481), .B(n9482), .Z(n9478) );
  ANDN U13579 ( .B(n9483), .A(n9484), .Z(n9481) );
  XNOR U13580 ( .A(b[1949]), .B(n9482), .Z(n9483) );
  XNOR U13581 ( .A(b[194]), .B(n9485), .Z(c[194]) );
  XNOR U13582 ( .A(b[1949]), .B(n9484), .Z(c[1949]) );
  XOR U13583 ( .A(n9486), .B(n9487), .Z(n9482) );
  ANDN U13584 ( .B(n9488), .A(n9489), .Z(n9486) );
  XNOR U13585 ( .A(b[1948]), .B(n9487), .Z(n9488) );
  XNOR U13586 ( .A(b[1948]), .B(n9489), .Z(c[1948]) );
  XOR U13587 ( .A(n9490), .B(n9491), .Z(n9487) );
  ANDN U13588 ( .B(n9492), .A(n9493), .Z(n9490) );
  XNOR U13589 ( .A(b[1947]), .B(n9491), .Z(n9492) );
  XNOR U13590 ( .A(b[1947]), .B(n9493), .Z(c[1947]) );
  XOR U13591 ( .A(n9494), .B(n9495), .Z(n9491) );
  ANDN U13592 ( .B(n9496), .A(n9497), .Z(n9494) );
  XNOR U13593 ( .A(b[1946]), .B(n9495), .Z(n9496) );
  XNOR U13594 ( .A(b[1946]), .B(n9497), .Z(c[1946]) );
  XOR U13595 ( .A(n9498), .B(n9499), .Z(n9495) );
  ANDN U13596 ( .B(n9500), .A(n9501), .Z(n9498) );
  XNOR U13597 ( .A(b[1945]), .B(n9499), .Z(n9500) );
  XNOR U13598 ( .A(b[1945]), .B(n9501), .Z(c[1945]) );
  XOR U13599 ( .A(n9502), .B(n9503), .Z(n9499) );
  ANDN U13600 ( .B(n9504), .A(n9505), .Z(n9502) );
  XNOR U13601 ( .A(b[1944]), .B(n9503), .Z(n9504) );
  XNOR U13602 ( .A(b[1944]), .B(n9505), .Z(c[1944]) );
  XOR U13603 ( .A(n9506), .B(n9507), .Z(n9503) );
  ANDN U13604 ( .B(n9508), .A(n9509), .Z(n9506) );
  XNOR U13605 ( .A(b[1943]), .B(n9507), .Z(n9508) );
  XNOR U13606 ( .A(b[1943]), .B(n9509), .Z(c[1943]) );
  XOR U13607 ( .A(n9510), .B(n9511), .Z(n9507) );
  ANDN U13608 ( .B(n9512), .A(n9513), .Z(n9510) );
  XNOR U13609 ( .A(b[1942]), .B(n9511), .Z(n9512) );
  XNOR U13610 ( .A(b[1942]), .B(n9513), .Z(c[1942]) );
  XOR U13611 ( .A(n9514), .B(n9515), .Z(n9511) );
  ANDN U13612 ( .B(n9516), .A(n9517), .Z(n9514) );
  XNOR U13613 ( .A(b[1941]), .B(n9515), .Z(n9516) );
  XNOR U13614 ( .A(b[1941]), .B(n9517), .Z(c[1941]) );
  XOR U13615 ( .A(n9518), .B(n9519), .Z(n9515) );
  ANDN U13616 ( .B(n9520), .A(n9521), .Z(n9518) );
  XNOR U13617 ( .A(b[1940]), .B(n9519), .Z(n9520) );
  XNOR U13618 ( .A(b[1940]), .B(n9521), .Z(c[1940]) );
  XOR U13619 ( .A(n9522), .B(n9523), .Z(n9519) );
  ANDN U13620 ( .B(n9524), .A(n9525), .Z(n9522) );
  XNOR U13621 ( .A(b[1939]), .B(n9523), .Z(n9524) );
  XNOR U13622 ( .A(b[193]), .B(n9526), .Z(c[193]) );
  XNOR U13623 ( .A(b[1939]), .B(n9525), .Z(c[1939]) );
  XOR U13624 ( .A(n9527), .B(n9528), .Z(n9523) );
  ANDN U13625 ( .B(n9529), .A(n9530), .Z(n9527) );
  XNOR U13626 ( .A(b[1938]), .B(n9528), .Z(n9529) );
  XNOR U13627 ( .A(b[1938]), .B(n9530), .Z(c[1938]) );
  XOR U13628 ( .A(n9531), .B(n9532), .Z(n9528) );
  ANDN U13629 ( .B(n9533), .A(n9534), .Z(n9531) );
  XNOR U13630 ( .A(b[1937]), .B(n9532), .Z(n9533) );
  XNOR U13631 ( .A(b[1937]), .B(n9534), .Z(c[1937]) );
  XOR U13632 ( .A(n9535), .B(n9536), .Z(n9532) );
  ANDN U13633 ( .B(n9537), .A(n9538), .Z(n9535) );
  XNOR U13634 ( .A(b[1936]), .B(n9536), .Z(n9537) );
  XNOR U13635 ( .A(b[1936]), .B(n9538), .Z(c[1936]) );
  XOR U13636 ( .A(n9539), .B(n9540), .Z(n9536) );
  ANDN U13637 ( .B(n9541), .A(n9542), .Z(n9539) );
  XNOR U13638 ( .A(b[1935]), .B(n9540), .Z(n9541) );
  XNOR U13639 ( .A(b[1935]), .B(n9542), .Z(c[1935]) );
  XOR U13640 ( .A(n9543), .B(n9544), .Z(n9540) );
  ANDN U13641 ( .B(n9545), .A(n9546), .Z(n9543) );
  XNOR U13642 ( .A(b[1934]), .B(n9544), .Z(n9545) );
  XNOR U13643 ( .A(b[1934]), .B(n9546), .Z(c[1934]) );
  XOR U13644 ( .A(n9547), .B(n9548), .Z(n9544) );
  ANDN U13645 ( .B(n9549), .A(n9550), .Z(n9547) );
  XNOR U13646 ( .A(b[1933]), .B(n9548), .Z(n9549) );
  XNOR U13647 ( .A(b[1933]), .B(n9550), .Z(c[1933]) );
  XOR U13648 ( .A(n9551), .B(n9552), .Z(n9548) );
  ANDN U13649 ( .B(n9553), .A(n9554), .Z(n9551) );
  XNOR U13650 ( .A(b[1932]), .B(n9552), .Z(n9553) );
  XNOR U13651 ( .A(b[1932]), .B(n9554), .Z(c[1932]) );
  XOR U13652 ( .A(n9555), .B(n9556), .Z(n9552) );
  ANDN U13653 ( .B(n9557), .A(n9558), .Z(n9555) );
  XNOR U13654 ( .A(b[1931]), .B(n9556), .Z(n9557) );
  XNOR U13655 ( .A(b[1931]), .B(n9558), .Z(c[1931]) );
  XOR U13656 ( .A(n9559), .B(n9560), .Z(n9556) );
  ANDN U13657 ( .B(n9561), .A(n9562), .Z(n9559) );
  XNOR U13658 ( .A(b[1930]), .B(n9560), .Z(n9561) );
  XNOR U13659 ( .A(b[1930]), .B(n9562), .Z(c[1930]) );
  XOR U13660 ( .A(n9563), .B(n9564), .Z(n9560) );
  ANDN U13661 ( .B(n9565), .A(n9566), .Z(n9563) );
  XNOR U13662 ( .A(b[1929]), .B(n9564), .Z(n9565) );
  XNOR U13663 ( .A(b[192]), .B(n9567), .Z(c[192]) );
  XNOR U13664 ( .A(b[1929]), .B(n9566), .Z(c[1929]) );
  XOR U13665 ( .A(n9568), .B(n9569), .Z(n9564) );
  ANDN U13666 ( .B(n9570), .A(n9571), .Z(n9568) );
  XNOR U13667 ( .A(b[1928]), .B(n9569), .Z(n9570) );
  XNOR U13668 ( .A(b[1928]), .B(n9571), .Z(c[1928]) );
  XOR U13669 ( .A(n9572), .B(n9573), .Z(n9569) );
  ANDN U13670 ( .B(n9574), .A(n9575), .Z(n9572) );
  XNOR U13671 ( .A(b[1927]), .B(n9573), .Z(n9574) );
  XNOR U13672 ( .A(b[1927]), .B(n9575), .Z(c[1927]) );
  XOR U13673 ( .A(n9576), .B(n9577), .Z(n9573) );
  ANDN U13674 ( .B(n9578), .A(n9579), .Z(n9576) );
  XNOR U13675 ( .A(b[1926]), .B(n9577), .Z(n9578) );
  XNOR U13676 ( .A(b[1926]), .B(n9579), .Z(c[1926]) );
  XOR U13677 ( .A(n9580), .B(n9581), .Z(n9577) );
  ANDN U13678 ( .B(n9582), .A(n9583), .Z(n9580) );
  XNOR U13679 ( .A(b[1925]), .B(n9581), .Z(n9582) );
  XNOR U13680 ( .A(b[1925]), .B(n9583), .Z(c[1925]) );
  XOR U13681 ( .A(n9584), .B(n9585), .Z(n9581) );
  ANDN U13682 ( .B(n9586), .A(n9587), .Z(n9584) );
  XNOR U13683 ( .A(b[1924]), .B(n9585), .Z(n9586) );
  XNOR U13684 ( .A(b[1924]), .B(n9587), .Z(c[1924]) );
  XOR U13685 ( .A(n9588), .B(n9589), .Z(n9585) );
  ANDN U13686 ( .B(n9590), .A(n9591), .Z(n9588) );
  XNOR U13687 ( .A(b[1923]), .B(n9589), .Z(n9590) );
  XNOR U13688 ( .A(b[1923]), .B(n9591), .Z(c[1923]) );
  XOR U13689 ( .A(n9592), .B(n9593), .Z(n9589) );
  ANDN U13690 ( .B(n9594), .A(n9595), .Z(n9592) );
  XNOR U13691 ( .A(b[1922]), .B(n9593), .Z(n9594) );
  XNOR U13692 ( .A(b[1922]), .B(n9595), .Z(c[1922]) );
  XOR U13693 ( .A(n9596), .B(n9597), .Z(n9593) );
  ANDN U13694 ( .B(n9598), .A(n9599), .Z(n9596) );
  XNOR U13695 ( .A(b[1921]), .B(n9597), .Z(n9598) );
  XNOR U13696 ( .A(b[1921]), .B(n9599), .Z(c[1921]) );
  XOR U13697 ( .A(n9600), .B(n9601), .Z(n9597) );
  ANDN U13698 ( .B(n9602), .A(n9603), .Z(n9600) );
  XNOR U13699 ( .A(b[1920]), .B(n9601), .Z(n9602) );
  XNOR U13700 ( .A(b[1920]), .B(n9603), .Z(c[1920]) );
  XOR U13701 ( .A(n9604), .B(n9605), .Z(n9601) );
  ANDN U13702 ( .B(n9606), .A(n9607), .Z(n9604) );
  XNOR U13703 ( .A(b[1919]), .B(n9605), .Z(n9606) );
  XNOR U13704 ( .A(b[191]), .B(n9608), .Z(c[191]) );
  XNOR U13705 ( .A(b[1919]), .B(n9607), .Z(c[1919]) );
  XOR U13706 ( .A(n9609), .B(n9610), .Z(n9605) );
  ANDN U13707 ( .B(n9611), .A(n9612), .Z(n9609) );
  XNOR U13708 ( .A(b[1918]), .B(n9610), .Z(n9611) );
  XNOR U13709 ( .A(b[1918]), .B(n9612), .Z(c[1918]) );
  XOR U13710 ( .A(n9613), .B(n9614), .Z(n9610) );
  ANDN U13711 ( .B(n9615), .A(n9616), .Z(n9613) );
  XNOR U13712 ( .A(b[1917]), .B(n9614), .Z(n9615) );
  XNOR U13713 ( .A(b[1917]), .B(n9616), .Z(c[1917]) );
  XOR U13714 ( .A(n9617), .B(n9618), .Z(n9614) );
  ANDN U13715 ( .B(n9619), .A(n9620), .Z(n9617) );
  XNOR U13716 ( .A(b[1916]), .B(n9618), .Z(n9619) );
  XNOR U13717 ( .A(b[1916]), .B(n9620), .Z(c[1916]) );
  XOR U13718 ( .A(n9621), .B(n9622), .Z(n9618) );
  ANDN U13719 ( .B(n9623), .A(n9624), .Z(n9621) );
  XNOR U13720 ( .A(b[1915]), .B(n9622), .Z(n9623) );
  XNOR U13721 ( .A(b[1915]), .B(n9624), .Z(c[1915]) );
  XOR U13722 ( .A(n9625), .B(n9626), .Z(n9622) );
  ANDN U13723 ( .B(n9627), .A(n9628), .Z(n9625) );
  XNOR U13724 ( .A(b[1914]), .B(n9626), .Z(n9627) );
  XNOR U13725 ( .A(b[1914]), .B(n9628), .Z(c[1914]) );
  XOR U13726 ( .A(n9629), .B(n9630), .Z(n9626) );
  ANDN U13727 ( .B(n9631), .A(n9632), .Z(n9629) );
  XNOR U13728 ( .A(b[1913]), .B(n9630), .Z(n9631) );
  XNOR U13729 ( .A(b[1913]), .B(n9632), .Z(c[1913]) );
  XOR U13730 ( .A(n9633), .B(n9634), .Z(n9630) );
  ANDN U13731 ( .B(n9635), .A(n9636), .Z(n9633) );
  XNOR U13732 ( .A(b[1912]), .B(n9634), .Z(n9635) );
  XNOR U13733 ( .A(b[1912]), .B(n9636), .Z(c[1912]) );
  XOR U13734 ( .A(n9637), .B(n9638), .Z(n9634) );
  ANDN U13735 ( .B(n9639), .A(n9640), .Z(n9637) );
  XNOR U13736 ( .A(b[1911]), .B(n9638), .Z(n9639) );
  XNOR U13737 ( .A(b[1911]), .B(n9640), .Z(c[1911]) );
  XOR U13738 ( .A(n9641), .B(n9642), .Z(n9638) );
  ANDN U13739 ( .B(n9643), .A(n9644), .Z(n9641) );
  XNOR U13740 ( .A(b[1910]), .B(n9642), .Z(n9643) );
  XNOR U13741 ( .A(b[1910]), .B(n9644), .Z(c[1910]) );
  XOR U13742 ( .A(n9645), .B(n9646), .Z(n9642) );
  ANDN U13743 ( .B(n9647), .A(n9648), .Z(n9645) );
  XNOR U13744 ( .A(b[1909]), .B(n9646), .Z(n9647) );
  XNOR U13745 ( .A(b[190]), .B(n9649), .Z(c[190]) );
  XNOR U13746 ( .A(b[1909]), .B(n9648), .Z(c[1909]) );
  XOR U13747 ( .A(n9650), .B(n9651), .Z(n9646) );
  ANDN U13748 ( .B(n9652), .A(n9653), .Z(n9650) );
  XNOR U13749 ( .A(b[1908]), .B(n9651), .Z(n9652) );
  XNOR U13750 ( .A(b[1908]), .B(n9653), .Z(c[1908]) );
  XOR U13751 ( .A(n9654), .B(n9655), .Z(n9651) );
  ANDN U13752 ( .B(n9656), .A(n9657), .Z(n9654) );
  XNOR U13753 ( .A(b[1907]), .B(n9655), .Z(n9656) );
  XNOR U13754 ( .A(b[1907]), .B(n9657), .Z(c[1907]) );
  XOR U13755 ( .A(n9658), .B(n9659), .Z(n9655) );
  ANDN U13756 ( .B(n9660), .A(n9661), .Z(n9658) );
  XNOR U13757 ( .A(b[1906]), .B(n9659), .Z(n9660) );
  XNOR U13758 ( .A(b[1906]), .B(n9661), .Z(c[1906]) );
  XOR U13759 ( .A(n9662), .B(n9663), .Z(n9659) );
  ANDN U13760 ( .B(n9664), .A(n9665), .Z(n9662) );
  XNOR U13761 ( .A(b[1905]), .B(n9663), .Z(n9664) );
  XNOR U13762 ( .A(b[1905]), .B(n9665), .Z(c[1905]) );
  XOR U13763 ( .A(n9666), .B(n9667), .Z(n9663) );
  ANDN U13764 ( .B(n9668), .A(n9669), .Z(n9666) );
  XNOR U13765 ( .A(b[1904]), .B(n9667), .Z(n9668) );
  XNOR U13766 ( .A(b[1904]), .B(n9669), .Z(c[1904]) );
  XOR U13767 ( .A(n9670), .B(n9671), .Z(n9667) );
  ANDN U13768 ( .B(n9672), .A(n9673), .Z(n9670) );
  XNOR U13769 ( .A(b[1903]), .B(n9671), .Z(n9672) );
  XNOR U13770 ( .A(b[1903]), .B(n9673), .Z(c[1903]) );
  XOR U13771 ( .A(n9674), .B(n9675), .Z(n9671) );
  ANDN U13772 ( .B(n9676), .A(n9677), .Z(n9674) );
  XNOR U13773 ( .A(b[1902]), .B(n9675), .Z(n9676) );
  XNOR U13774 ( .A(b[1902]), .B(n9677), .Z(c[1902]) );
  XOR U13775 ( .A(n9678), .B(n9679), .Z(n9675) );
  ANDN U13776 ( .B(n9680), .A(n9681), .Z(n9678) );
  XNOR U13777 ( .A(b[1901]), .B(n9679), .Z(n9680) );
  XNOR U13778 ( .A(b[1901]), .B(n9681), .Z(c[1901]) );
  XOR U13779 ( .A(n9682), .B(n9683), .Z(n9679) );
  ANDN U13780 ( .B(n9684), .A(n9685), .Z(n9682) );
  XNOR U13781 ( .A(b[1900]), .B(n9683), .Z(n9684) );
  XNOR U13782 ( .A(b[1900]), .B(n9685), .Z(c[1900]) );
  XOR U13783 ( .A(n9686), .B(n9687), .Z(n9683) );
  ANDN U13784 ( .B(n9688), .A(n9689), .Z(n9686) );
  XNOR U13785 ( .A(b[1899]), .B(n9687), .Z(n9688) );
  XNOR U13786 ( .A(b[18]), .B(n9690), .Z(c[18]) );
  XNOR U13787 ( .A(b[189]), .B(n9691), .Z(c[189]) );
  XNOR U13788 ( .A(b[1899]), .B(n9689), .Z(c[1899]) );
  XOR U13789 ( .A(n9692), .B(n9693), .Z(n9687) );
  ANDN U13790 ( .B(n9694), .A(n9695), .Z(n9692) );
  XNOR U13791 ( .A(b[1898]), .B(n9693), .Z(n9694) );
  XNOR U13792 ( .A(b[1898]), .B(n9695), .Z(c[1898]) );
  XOR U13793 ( .A(n9696), .B(n9697), .Z(n9693) );
  ANDN U13794 ( .B(n9698), .A(n9699), .Z(n9696) );
  XNOR U13795 ( .A(b[1897]), .B(n9697), .Z(n9698) );
  XNOR U13796 ( .A(b[1897]), .B(n9699), .Z(c[1897]) );
  XOR U13797 ( .A(n9700), .B(n9701), .Z(n9697) );
  ANDN U13798 ( .B(n9702), .A(n9703), .Z(n9700) );
  XNOR U13799 ( .A(b[1896]), .B(n9701), .Z(n9702) );
  XNOR U13800 ( .A(b[1896]), .B(n9703), .Z(c[1896]) );
  XOR U13801 ( .A(n9704), .B(n9705), .Z(n9701) );
  ANDN U13802 ( .B(n9706), .A(n9707), .Z(n9704) );
  XNOR U13803 ( .A(b[1895]), .B(n9705), .Z(n9706) );
  XNOR U13804 ( .A(b[1895]), .B(n9707), .Z(c[1895]) );
  XOR U13805 ( .A(n9708), .B(n9709), .Z(n9705) );
  ANDN U13806 ( .B(n9710), .A(n9711), .Z(n9708) );
  XNOR U13807 ( .A(b[1894]), .B(n9709), .Z(n9710) );
  XNOR U13808 ( .A(b[1894]), .B(n9711), .Z(c[1894]) );
  XOR U13809 ( .A(n9712), .B(n9713), .Z(n9709) );
  ANDN U13810 ( .B(n9714), .A(n9715), .Z(n9712) );
  XNOR U13811 ( .A(b[1893]), .B(n9713), .Z(n9714) );
  XNOR U13812 ( .A(b[1893]), .B(n9715), .Z(c[1893]) );
  XOR U13813 ( .A(n9716), .B(n9717), .Z(n9713) );
  ANDN U13814 ( .B(n9718), .A(n9719), .Z(n9716) );
  XNOR U13815 ( .A(b[1892]), .B(n9717), .Z(n9718) );
  XNOR U13816 ( .A(b[1892]), .B(n9719), .Z(c[1892]) );
  XOR U13817 ( .A(n9720), .B(n9721), .Z(n9717) );
  ANDN U13818 ( .B(n9722), .A(n9723), .Z(n9720) );
  XNOR U13819 ( .A(b[1891]), .B(n9721), .Z(n9722) );
  XNOR U13820 ( .A(b[1891]), .B(n9723), .Z(c[1891]) );
  XOR U13821 ( .A(n9724), .B(n9725), .Z(n9721) );
  ANDN U13822 ( .B(n9726), .A(n9727), .Z(n9724) );
  XNOR U13823 ( .A(b[1890]), .B(n9725), .Z(n9726) );
  XNOR U13824 ( .A(b[1890]), .B(n9727), .Z(c[1890]) );
  XOR U13825 ( .A(n9728), .B(n9729), .Z(n9725) );
  ANDN U13826 ( .B(n9730), .A(n9731), .Z(n9728) );
  XNOR U13827 ( .A(b[1889]), .B(n9729), .Z(n9730) );
  XNOR U13828 ( .A(b[188]), .B(n9732), .Z(c[188]) );
  XNOR U13829 ( .A(b[1889]), .B(n9731), .Z(c[1889]) );
  XOR U13830 ( .A(n9733), .B(n9734), .Z(n9729) );
  ANDN U13831 ( .B(n9735), .A(n9736), .Z(n9733) );
  XNOR U13832 ( .A(b[1888]), .B(n9734), .Z(n9735) );
  XNOR U13833 ( .A(b[1888]), .B(n9736), .Z(c[1888]) );
  XOR U13834 ( .A(n9737), .B(n9738), .Z(n9734) );
  ANDN U13835 ( .B(n9739), .A(n9740), .Z(n9737) );
  XNOR U13836 ( .A(b[1887]), .B(n9738), .Z(n9739) );
  XNOR U13837 ( .A(b[1887]), .B(n9740), .Z(c[1887]) );
  XOR U13838 ( .A(n9741), .B(n9742), .Z(n9738) );
  ANDN U13839 ( .B(n9743), .A(n9744), .Z(n9741) );
  XNOR U13840 ( .A(b[1886]), .B(n9742), .Z(n9743) );
  XNOR U13841 ( .A(b[1886]), .B(n9744), .Z(c[1886]) );
  XOR U13842 ( .A(n9745), .B(n9746), .Z(n9742) );
  ANDN U13843 ( .B(n9747), .A(n9748), .Z(n9745) );
  XNOR U13844 ( .A(b[1885]), .B(n9746), .Z(n9747) );
  XNOR U13845 ( .A(b[1885]), .B(n9748), .Z(c[1885]) );
  XOR U13846 ( .A(n9749), .B(n9750), .Z(n9746) );
  ANDN U13847 ( .B(n9751), .A(n9752), .Z(n9749) );
  XNOR U13848 ( .A(b[1884]), .B(n9750), .Z(n9751) );
  XNOR U13849 ( .A(b[1884]), .B(n9752), .Z(c[1884]) );
  XOR U13850 ( .A(n9753), .B(n9754), .Z(n9750) );
  ANDN U13851 ( .B(n9755), .A(n9756), .Z(n9753) );
  XNOR U13852 ( .A(b[1883]), .B(n9754), .Z(n9755) );
  XNOR U13853 ( .A(b[1883]), .B(n9756), .Z(c[1883]) );
  XOR U13854 ( .A(n9757), .B(n9758), .Z(n9754) );
  ANDN U13855 ( .B(n9759), .A(n9760), .Z(n9757) );
  XNOR U13856 ( .A(b[1882]), .B(n9758), .Z(n9759) );
  XNOR U13857 ( .A(b[1882]), .B(n9760), .Z(c[1882]) );
  XOR U13858 ( .A(n9761), .B(n9762), .Z(n9758) );
  ANDN U13859 ( .B(n9763), .A(n9764), .Z(n9761) );
  XNOR U13860 ( .A(b[1881]), .B(n9762), .Z(n9763) );
  XNOR U13861 ( .A(b[1881]), .B(n9764), .Z(c[1881]) );
  XOR U13862 ( .A(n9765), .B(n9766), .Z(n9762) );
  ANDN U13863 ( .B(n9767), .A(n9768), .Z(n9765) );
  XNOR U13864 ( .A(b[1880]), .B(n9766), .Z(n9767) );
  XNOR U13865 ( .A(b[1880]), .B(n9768), .Z(c[1880]) );
  XOR U13866 ( .A(n9769), .B(n9770), .Z(n9766) );
  ANDN U13867 ( .B(n9771), .A(n9772), .Z(n9769) );
  XNOR U13868 ( .A(b[1879]), .B(n9770), .Z(n9771) );
  XNOR U13869 ( .A(b[187]), .B(n9773), .Z(c[187]) );
  XNOR U13870 ( .A(b[1879]), .B(n9772), .Z(c[1879]) );
  XOR U13871 ( .A(n9774), .B(n9775), .Z(n9770) );
  ANDN U13872 ( .B(n9776), .A(n9777), .Z(n9774) );
  XNOR U13873 ( .A(b[1878]), .B(n9775), .Z(n9776) );
  XNOR U13874 ( .A(b[1878]), .B(n9777), .Z(c[1878]) );
  XOR U13875 ( .A(n9778), .B(n9779), .Z(n9775) );
  ANDN U13876 ( .B(n9780), .A(n9781), .Z(n9778) );
  XNOR U13877 ( .A(b[1877]), .B(n9779), .Z(n9780) );
  XNOR U13878 ( .A(b[1877]), .B(n9781), .Z(c[1877]) );
  XOR U13879 ( .A(n9782), .B(n9783), .Z(n9779) );
  ANDN U13880 ( .B(n9784), .A(n9785), .Z(n9782) );
  XNOR U13881 ( .A(b[1876]), .B(n9783), .Z(n9784) );
  XNOR U13882 ( .A(b[1876]), .B(n9785), .Z(c[1876]) );
  XOR U13883 ( .A(n9786), .B(n9787), .Z(n9783) );
  ANDN U13884 ( .B(n9788), .A(n9789), .Z(n9786) );
  XNOR U13885 ( .A(b[1875]), .B(n9787), .Z(n9788) );
  XNOR U13886 ( .A(b[1875]), .B(n9789), .Z(c[1875]) );
  XOR U13887 ( .A(n9790), .B(n9791), .Z(n9787) );
  ANDN U13888 ( .B(n9792), .A(n9793), .Z(n9790) );
  XNOR U13889 ( .A(b[1874]), .B(n9791), .Z(n9792) );
  XNOR U13890 ( .A(b[1874]), .B(n9793), .Z(c[1874]) );
  XOR U13891 ( .A(n9794), .B(n9795), .Z(n9791) );
  ANDN U13892 ( .B(n9796), .A(n9797), .Z(n9794) );
  XNOR U13893 ( .A(b[1873]), .B(n9795), .Z(n9796) );
  XNOR U13894 ( .A(b[1873]), .B(n9797), .Z(c[1873]) );
  XOR U13895 ( .A(n9798), .B(n9799), .Z(n9795) );
  ANDN U13896 ( .B(n9800), .A(n9801), .Z(n9798) );
  XNOR U13897 ( .A(b[1872]), .B(n9799), .Z(n9800) );
  XNOR U13898 ( .A(b[1872]), .B(n9801), .Z(c[1872]) );
  XOR U13899 ( .A(n9802), .B(n9803), .Z(n9799) );
  ANDN U13900 ( .B(n9804), .A(n9805), .Z(n9802) );
  XNOR U13901 ( .A(b[1871]), .B(n9803), .Z(n9804) );
  XNOR U13902 ( .A(b[1871]), .B(n9805), .Z(c[1871]) );
  XOR U13903 ( .A(n9806), .B(n9807), .Z(n9803) );
  ANDN U13904 ( .B(n9808), .A(n9809), .Z(n9806) );
  XNOR U13905 ( .A(b[1870]), .B(n9807), .Z(n9808) );
  XNOR U13906 ( .A(b[1870]), .B(n9809), .Z(c[1870]) );
  XOR U13907 ( .A(n9810), .B(n9811), .Z(n9807) );
  ANDN U13908 ( .B(n9812), .A(n9813), .Z(n9810) );
  XNOR U13909 ( .A(b[1869]), .B(n9811), .Z(n9812) );
  XNOR U13910 ( .A(b[186]), .B(n9814), .Z(c[186]) );
  XNOR U13911 ( .A(b[1869]), .B(n9813), .Z(c[1869]) );
  XOR U13912 ( .A(n9815), .B(n9816), .Z(n9811) );
  ANDN U13913 ( .B(n9817), .A(n9818), .Z(n9815) );
  XNOR U13914 ( .A(b[1868]), .B(n9816), .Z(n9817) );
  XNOR U13915 ( .A(b[1868]), .B(n9818), .Z(c[1868]) );
  XOR U13916 ( .A(n9819), .B(n9820), .Z(n9816) );
  ANDN U13917 ( .B(n9821), .A(n9822), .Z(n9819) );
  XNOR U13918 ( .A(b[1867]), .B(n9820), .Z(n9821) );
  XNOR U13919 ( .A(b[1867]), .B(n9822), .Z(c[1867]) );
  XOR U13920 ( .A(n9823), .B(n9824), .Z(n9820) );
  ANDN U13921 ( .B(n9825), .A(n9826), .Z(n9823) );
  XNOR U13922 ( .A(b[1866]), .B(n9824), .Z(n9825) );
  XNOR U13923 ( .A(b[1866]), .B(n9826), .Z(c[1866]) );
  XOR U13924 ( .A(n9827), .B(n9828), .Z(n9824) );
  ANDN U13925 ( .B(n9829), .A(n9830), .Z(n9827) );
  XNOR U13926 ( .A(b[1865]), .B(n9828), .Z(n9829) );
  XNOR U13927 ( .A(b[1865]), .B(n9830), .Z(c[1865]) );
  XOR U13928 ( .A(n9831), .B(n9832), .Z(n9828) );
  ANDN U13929 ( .B(n9833), .A(n9834), .Z(n9831) );
  XNOR U13930 ( .A(b[1864]), .B(n9832), .Z(n9833) );
  XNOR U13931 ( .A(b[1864]), .B(n9834), .Z(c[1864]) );
  XOR U13932 ( .A(n9835), .B(n9836), .Z(n9832) );
  ANDN U13933 ( .B(n9837), .A(n9838), .Z(n9835) );
  XNOR U13934 ( .A(b[1863]), .B(n9836), .Z(n9837) );
  XNOR U13935 ( .A(b[1863]), .B(n9838), .Z(c[1863]) );
  XOR U13936 ( .A(n9839), .B(n9840), .Z(n9836) );
  ANDN U13937 ( .B(n9841), .A(n9842), .Z(n9839) );
  XNOR U13938 ( .A(b[1862]), .B(n9840), .Z(n9841) );
  XNOR U13939 ( .A(b[1862]), .B(n9842), .Z(c[1862]) );
  XOR U13940 ( .A(n9843), .B(n9844), .Z(n9840) );
  ANDN U13941 ( .B(n9845), .A(n9846), .Z(n9843) );
  XNOR U13942 ( .A(b[1861]), .B(n9844), .Z(n9845) );
  XNOR U13943 ( .A(b[1861]), .B(n9846), .Z(c[1861]) );
  XOR U13944 ( .A(n9847), .B(n9848), .Z(n9844) );
  ANDN U13945 ( .B(n9849), .A(n9850), .Z(n9847) );
  XNOR U13946 ( .A(b[1860]), .B(n9848), .Z(n9849) );
  XNOR U13947 ( .A(b[1860]), .B(n9850), .Z(c[1860]) );
  XOR U13948 ( .A(n9851), .B(n9852), .Z(n9848) );
  ANDN U13949 ( .B(n9853), .A(n9854), .Z(n9851) );
  XNOR U13950 ( .A(b[1859]), .B(n9852), .Z(n9853) );
  XNOR U13951 ( .A(b[185]), .B(n9855), .Z(c[185]) );
  XNOR U13952 ( .A(b[1859]), .B(n9854), .Z(c[1859]) );
  XOR U13953 ( .A(n9856), .B(n9857), .Z(n9852) );
  ANDN U13954 ( .B(n9858), .A(n9859), .Z(n9856) );
  XNOR U13955 ( .A(b[1858]), .B(n9857), .Z(n9858) );
  XNOR U13956 ( .A(b[1858]), .B(n9859), .Z(c[1858]) );
  XOR U13957 ( .A(n9860), .B(n9861), .Z(n9857) );
  ANDN U13958 ( .B(n9862), .A(n9863), .Z(n9860) );
  XNOR U13959 ( .A(b[1857]), .B(n9861), .Z(n9862) );
  XNOR U13960 ( .A(b[1857]), .B(n9863), .Z(c[1857]) );
  XOR U13961 ( .A(n9864), .B(n9865), .Z(n9861) );
  ANDN U13962 ( .B(n9866), .A(n9867), .Z(n9864) );
  XNOR U13963 ( .A(b[1856]), .B(n9865), .Z(n9866) );
  XNOR U13964 ( .A(b[1856]), .B(n9867), .Z(c[1856]) );
  XOR U13965 ( .A(n9868), .B(n9869), .Z(n9865) );
  ANDN U13966 ( .B(n9870), .A(n9871), .Z(n9868) );
  XNOR U13967 ( .A(b[1855]), .B(n9869), .Z(n9870) );
  XNOR U13968 ( .A(b[1855]), .B(n9871), .Z(c[1855]) );
  XOR U13969 ( .A(n9872), .B(n9873), .Z(n9869) );
  ANDN U13970 ( .B(n9874), .A(n9875), .Z(n9872) );
  XNOR U13971 ( .A(b[1854]), .B(n9873), .Z(n9874) );
  XNOR U13972 ( .A(b[1854]), .B(n9875), .Z(c[1854]) );
  XOR U13973 ( .A(n9876), .B(n9877), .Z(n9873) );
  ANDN U13974 ( .B(n9878), .A(n9879), .Z(n9876) );
  XNOR U13975 ( .A(b[1853]), .B(n9877), .Z(n9878) );
  XNOR U13976 ( .A(b[1853]), .B(n9879), .Z(c[1853]) );
  XOR U13977 ( .A(n9880), .B(n9881), .Z(n9877) );
  ANDN U13978 ( .B(n9882), .A(n9883), .Z(n9880) );
  XNOR U13979 ( .A(b[1852]), .B(n9881), .Z(n9882) );
  XNOR U13980 ( .A(b[1852]), .B(n9883), .Z(c[1852]) );
  XOR U13981 ( .A(n9884), .B(n9885), .Z(n9881) );
  ANDN U13982 ( .B(n9886), .A(n9887), .Z(n9884) );
  XNOR U13983 ( .A(b[1851]), .B(n9885), .Z(n9886) );
  XNOR U13984 ( .A(b[1851]), .B(n9887), .Z(c[1851]) );
  XOR U13985 ( .A(n9888), .B(n9889), .Z(n9885) );
  ANDN U13986 ( .B(n9890), .A(n9891), .Z(n9888) );
  XNOR U13987 ( .A(b[1850]), .B(n9889), .Z(n9890) );
  XNOR U13988 ( .A(b[1850]), .B(n9891), .Z(c[1850]) );
  XOR U13989 ( .A(n9892), .B(n9893), .Z(n9889) );
  ANDN U13990 ( .B(n9894), .A(n9895), .Z(n9892) );
  XNOR U13991 ( .A(b[1849]), .B(n9893), .Z(n9894) );
  XNOR U13992 ( .A(b[184]), .B(n9896), .Z(c[184]) );
  XNOR U13993 ( .A(b[1849]), .B(n9895), .Z(c[1849]) );
  XOR U13994 ( .A(n9897), .B(n9898), .Z(n9893) );
  ANDN U13995 ( .B(n9899), .A(n9900), .Z(n9897) );
  XNOR U13996 ( .A(b[1848]), .B(n9898), .Z(n9899) );
  XNOR U13997 ( .A(b[1848]), .B(n9900), .Z(c[1848]) );
  XOR U13998 ( .A(n9901), .B(n9902), .Z(n9898) );
  ANDN U13999 ( .B(n9903), .A(n9904), .Z(n9901) );
  XNOR U14000 ( .A(b[1847]), .B(n9902), .Z(n9903) );
  XNOR U14001 ( .A(b[1847]), .B(n9904), .Z(c[1847]) );
  XOR U14002 ( .A(n9905), .B(n9906), .Z(n9902) );
  ANDN U14003 ( .B(n9907), .A(n9908), .Z(n9905) );
  XNOR U14004 ( .A(b[1846]), .B(n9906), .Z(n9907) );
  XNOR U14005 ( .A(b[1846]), .B(n9908), .Z(c[1846]) );
  XOR U14006 ( .A(n9909), .B(n9910), .Z(n9906) );
  ANDN U14007 ( .B(n9911), .A(n9912), .Z(n9909) );
  XNOR U14008 ( .A(b[1845]), .B(n9910), .Z(n9911) );
  XNOR U14009 ( .A(b[1845]), .B(n9912), .Z(c[1845]) );
  XOR U14010 ( .A(n9913), .B(n9914), .Z(n9910) );
  ANDN U14011 ( .B(n9915), .A(n9916), .Z(n9913) );
  XNOR U14012 ( .A(b[1844]), .B(n9914), .Z(n9915) );
  XNOR U14013 ( .A(b[1844]), .B(n9916), .Z(c[1844]) );
  XOR U14014 ( .A(n9917), .B(n9918), .Z(n9914) );
  ANDN U14015 ( .B(n9919), .A(n9920), .Z(n9917) );
  XNOR U14016 ( .A(b[1843]), .B(n9918), .Z(n9919) );
  XNOR U14017 ( .A(b[1843]), .B(n9920), .Z(c[1843]) );
  XOR U14018 ( .A(n9921), .B(n9922), .Z(n9918) );
  ANDN U14019 ( .B(n9923), .A(n9924), .Z(n9921) );
  XNOR U14020 ( .A(b[1842]), .B(n9922), .Z(n9923) );
  XNOR U14021 ( .A(b[1842]), .B(n9924), .Z(c[1842]) );
  XOR U14022 ( .A(n9925), .B(n9926), .Z(n9922) );
  ANDN U14023 ( .B(n9927), .A(n9928), .Z(n9925) );
  XNOR U14024 ( .A(b[1841]), .B(n9926), .Z(n9927) );
  XNOR U14025 ( .A(b[1841]), .B(n9928), .Z(c[1841]) );
  XOR U14026 ( .A(n9929), .B(n9930), .Z(n9926) );
  ANDN U14027 ( .B(n9931), .A(n9932), .Z(n9929) );
  XNOR U14028 ( .A(b[1840]), .B(n9930), .Z(n9931) );
  XNOR U14029 ( .A(b[1840]), .B(n9932), .Z(c[1840]) );
  XOR U14030 ( .A(n9933), .B(n9934), .Z(n9930) );
  ANDN U14031 ( .B(n9935), .A(n9936), .Z(n9933) );
  XNOR U14032 ( .A(b[1839]), .B(n9934), .Z(n9935) );
  XNOR U14033 ( .A(b[183]), .B(n9937), .Z(c[183]) );
  XNOR U14034 ( .A(b[1839]), .B(n9936), .Z(c[1839]) );
  XOR U14035 ( .A(n9938), .B(n9939), .Z(n9934) );
  ANDN U14036 ( .B(n9940), .A(n9941), .Z(n9938) );
  XNOR U14037 ( .A(b[1838]), .B(n9939), .Z(n9940) );
  XNOR U14038 ( .A(b[1838]), .B(n9941), .Z(c[1838]) );
  XOR U14039 ( .A(n9942), .B(n9943), .Z(n9939) );
  ANDN U14040 ( .B(n9944), .A(n9945), .Z(n9942) );
  XNOR U14041 ( .A(b[1837]), .B(n9943), .Z(n9944) );
  XNOR U14042 ( .A(b[1837]), .B(n9945), .Z(c[1837]) );
  XOR U14043 ( .A(n9946), .B(n9947), .Z(n9943) );
  ANDN U14044 ( .B(n9948), .A(n9949), .Z(n9946) );
  XNOR U14045 ( .A(b[1836]), .B(n9947), .Z(n9948) );
  XNOR U14046 ( .A(b[1836]), .B(n9949), .Z(c[1836]) );
  XOR U14047 ( .A(n9950), .B(n9951), .Z(n9947) );
  ANDN U14048 ( .B(n9952), .A(n9953), .Z(n9950) );
  XNOR U14049 ( .A(b[1835]), .B(n9951), .Z(n9952) );
  XNOR U14050 ( .A(b[1835]), .B(n9953), .Z(c[1835]) );
  XOR U14051 ( .A(n9954), .B(n9955), .Z(n9951) );
  ANDN U14052 ( .B(n9956), .A(n9957), .Z(n9954) );
  XNOR U14053 ( .A(b[1834]), .B(n9955), .Z(n9956) );
  XNOR U14054 ( .A(b[1834]), .B(n9957), .Z(c[1834]) );
  XOR U14055 ( .A(n9958), .B(n9959), .Z(n9955) );
  ANDN U14056 ( .B(n9960), .A(n9961), .Z(n9958) );
  XNOR U14057 ( .A(b[1833]), .B(n9959), .Z(n9960) );
  XNOR U14058 ( .A(b[1833]), .B(n9961), .Z(c[1833]) );
  XOR U14059 ( .A(n9962), .B(n9963), .Z(n9959) );
  ANDN U14060 ( .B(n9964), .A(n9965), .Z(n9962) );
  XNOR U14061 ( .A(b[1832]), .B(n9963), .Z(n9964) );
  XNOR U14062 ( .A(b[1832]), .B(n9965), .Z(c[1832]) );
  XOR U14063 ( .A(n9966), .B(n9967), .Z(n9963) );
  ANDN U14064 ( .B(n9968), .A(n9969), .Z(n9966) );
  XNOR U14065 ( .A(b[1831]), .B(n9967), .Z(n9968) );
  XNOR U14066 ( .A(b[1831]), .B(n9969), .Z(c[1831]) );
  XOR U14067 ( .A(n9970), .B(n9971), .Z(n9967) );
  ANDN U14068 ( .B(n9972), .A(n9973), .Z(n9970) );
  XNOR U14069 ( .A(b[1830]), .B(n9971), .Z(n9972) );
  XNOR U14070 ( .A(b[1830]), .B(n9973), .Z(c[1830]) );
  XOR U14071 ( .A(n9974), .B(n9975), .Z(n9971) );
  ANDN U14072 ( .B(n9976), .A(n9977), .Z(n9974) );
  XNOR U14073 ( .A(b[1829]), .B(n9975), .Z(n9976) );
  XNOR U14074 ( .A(b[182]), .B(n9978), .Z(c[182]) );
  XNOR U14075 ( .A(b[1829]), .B(n9977), .Z(c[1829]) );
  XOR U14076 ( .A(n9979), .B(n9980), .Z(n9975) );
  ANDN U14077 ( .B(n9981), .A(n9982), .Z(n9979) );
  XNOR U14078 ( .A(b[1828]), .B(n9980), .Z(n9981) );
  XNOR U14079 ( .A(b[1828]), .B(n9982), .Z(c[1828]) );
  XOR U14080 ( .A(n9983), .B(n9984), .Z(n9980) );
  ANDN U14081 ( .B(n9985), .A(n9986), .Z(n9983) );
  XNOR U14082 ( .A(b[1827]), .B(n9984), .Z(n9985) );
  XNOR U14083 ( .A(b[1827]), .B(n9986), .Z(c[1827]) );
  XOR U14084 ( .A(n9987), .B(n9988), .Z(n9984) );
  ANDN U14085 ( .B(n9989), .A(n9990), .Z(n9987) );
  XNOR U14086 ( .A(b[1826]), .B(n9988), .Z(n9989) );
  XNOR U14087 ( .A(b[1826]), .B(n9990), .Z(c[1826]) );
  XOR U14088 ( .A(n9991), .B(n9992), .Z(n9988) );
  ANDN U14089 ( .B(n9993), .A(n9994), .Z(n9991) );
  XNOR U14090 ( .A(b[1825]), .B(n9992), .Z(n9993) );
  XNOR U14091 ( .A(b[1825]), .B(n9994), .Z(c[1825]) );
  XOR U14092 ( .A(n9995), .B(n9996), .Z(n9992) );
  ANDN U14093 ( .B(n9997), .A(n9998), .Z(n9995) );
  XNOR U14094 ( .A(b[1824]), .B(n9996), .Z(n9997) );
  XNOR U14095 ( .A(b[1824]), .B(n9998), .Z(c[1824]) );
  XOR U14096 ( .A(n9999), .B(n10000), .Z(n9996) );
  ANDN U14097 ( .B(n10001), .A(n10002), .Z(n9999) );
  XNOR U14098 ( .A(b[1823]), .B(n10000), .Z(n10001) );
  XNOR U14099 ( .A(b[1823]), .B(n10002), .Z(c[1823]) );
  XOR U14100 ( .A(n10003), .B(n10004), .Z(n10000) );
  ANDN U14101 ( .B(n10005), .A(n10006), .Z(n10003) );
  XNOR U14102 ( .A(b[1822]), .B(n10004), .Z(n10005) );
  XNOR U14103 ( .A(b[1822]), .B(n10006), .Z(c[1822]) );
  XOR U14104 ( .A(n10007), .B(n10008), .Z(n10004) );
  ANDN U14105 ( .B(n10009), .A(n10010), .Z(n10007) );
  XNOR U14106 ( .A(b[1821]), .B(n10008), .Z(n10009) );
  XNOR U14107 ( .A(b[1821]), .B(n10010), .Z(c[1821]) );
  XOR U14108 ( .A(n10011), .B(n10012), .Z(n10008) );
  ANDN U14109 ( .B(n10013), .A(n10014), .Z(n10011) );
  XNOR U14110 ( .A(b[1820]), .B(n10012), .Z(n10013) );
  XNOR U14111 ( .A(b[1820]), .B(n10014), .Z(c[1820]) );
  XOR U14112 ( .A(n10015), .B(n10016), .Z(n10012) );
  ANDN U14113 ( .B(n10017), .A(n10018), .Z(n10015) );
  XNOR U14114 ( .A(b[1819]), .B(n10016), .Z(n10017) );
  XNOR U14115 ( .A(b[181]), .B(n10019), .Z(c[181]) );
  XNOR U14116 ( .A(b[1819]), .B(n10018), .Z(c[1819]) );
  XOR U14117 ( .A(n10020), .B(n10021), .Z(n10016) );
  ANDN U14118 ( .B(n10022), .A(n10023), .Z(n10020) );
  XNOR U14119 ( .A(b[1818]), .B(n10021), .Z(n10022) );
  XNOR U14120 ( .A(b[1818]), .B(n10023), .Z(c[1818]) );
  XOR U14121 ( .A(n10024), .B(n10025), .Z(n10021) );
  ANDN U14122 ( .B(n10026), .A(n10027), .Z(n10024) );
  XNOR U14123 ( .A(b[1817]), .B(n10025), .Z(n10026) );
  XNOR U14124 ( .A(b[1817]), .B(n10027), .Z(c[1817]) );
  XOR U14125 ( .A(n10028), .B(n10029), .Z(n10025) );
  ANDN U14126 ( .B(n10030), .A(n10031), .Z(n10028) );
  XNOR U14127 ( .A(b[1816]), .B(n10029), .Z(n10030) );
  XNOR U14128 ( .A(b[1816]), .B(n10031), .Z(c[1816]) );
  XOR U14129 ( .A(n10032), .B(n10033), .Z(n10029) );
  ANDN U14130 ( .B(n10034), .A(n10035), .Z(n10032) );
  XNOR U14131 ( .A(b[1815]), .B(n10033), .Z(n10034) );
  XNOR U14132 ( .A(b[1815]), .B(n10035), .Z(c[1815]) );
  XOR U14133 ( .A(n10036), .B(n10037), .Z(n10033) );
  ANDN U14134 ( .B(n10038), .A(n10039), .Z(n10036) );
  XNOR U14135 ( .A(b[1814]), .B(n10037), .Z(n10038) );
  XNOR U14136 ( .A(b[1814]), .B(n10039), .Z(c[1814]) );
  XOR U14137 ( .A(n10040), .B(n10041), .Z(n10037) );
  ANDN U14138 ( .B(n10042), .A(n10043), .Z(n10040) );
  XNOR U14139 ( .A(b[1813]), .B(n10041), .Z(n10042) );
  XNOR U14140 ( .A(b[1813]), .B(n10043), .Z(c[1813]) );
  XOR U14141 ( .A(n10044), .B(n10045), .Z(n10041) );
  ANDN U14142 ( .B(n10046), .A(n10047), .Z(n10044) );
  XNOR U14143 ( .A(b[1812]), .B(n10045), .Z(n10046) );
  XNOR U14144 ( .A(b[1812]), .B(n10047), .Z(c[1812]) );
  XOR U14145 ( .A(n10048), .B(n10049), .Z(n10045) );
  ANDN U14146 ( .B(n10050), .A(n10051), .Z(n10048) );
  XNOR U14147 ( .A(b[1811]), .B(n10049), .Z(n10050) );
  XNOR U14148 ( .A(b[1811]), .B(n10051), .Z(c[1811]) );
  XOR U14149 ( .A(n10052), .B(n10053), .Z(n10049) );
  ANDN U14150 ( .B(n10054), .A(n10055), .Z(n10052) );
  XNOR U14151 ( .A(b[1810]), .B(n10053), .Z(n10054) );
  XNOR U14152 ( .A(b[1810]), .B(n10055), .Z(c[1810]) );
  XOR U14153 ( .A(n10056), .B(n10057), .Z(n10053) );
  ANDN U14154 ( .B(n10058), .A(n10059), .Z(n10056) );
  XNOR U14155 ( .A(b[1809]), .B(n10057), .Z(n10058) );
  XNOR U14156 ( .A(b[180]), .B(n10060), .Z(c[180]) );
  XNOR U14157 ( .A(b[1809]), .B(n10059), .Z(c[1809]) );
  XOR U14158 ( .A(n10061), .B(n10062), .Z(n10057) );
  ANDN U14159 ( .B(n10063), .A(n10064), .Z(n10061) );
  XNOR U14160 ( .A(b[1808]), .B(n10062), .Z(n10063) );
  XNOR U14161 ( .A(b[1808]), .B(n10064), .Z(c[1808]) );
  XOR U14162 ( .A(n10065), .B(n10066), .Z(n10062) );
  ANDN U14163 ( .B(n10067), .A(n10068), .Z(n10065) );
  XNOR U14164 ( .A(b[1807]), .B(n10066), .Z(n10067) );
  XNOR U14165 ( .A(b[1807]), .B(n10068), .Z(c[1807]) );
  XOR U14166 ( .A(n10069), .B(n10070), .Z(n10066) );
  ANDN U14167 ( .B(n10071), .A(n10072), .Z(n10069) );
  XNOR U14168 ( .A(b[1806]), .B(n10070), .Z(n10071) );
  XNOR U14169 ( .A(b[1806]), .B(n10072), .Z(c[1806]) );
  XOR U14170 ( .A(n10073), .B(n10074), .Z(n10070) );
  ANDN U14171 ( .B(n10075), .A(n10076), .Z(n10073) );
  XNOR U14172 ( .A(b[1805]), .B(n10074), .Z(n10075) );
  XNOR U14173 ( .A(b[1805]), .B(n10076), .Z(c[1805]) );
  XOR U14174 ( .A(n10077), .B(n10078), .Z(n10074) );
  ANDN U14175 ( .B(n10079), .A(n10080), .Z(n10077) );
  XNOR U14176 ( .A(b[1804]), .B(n10078), .Z(n10079) );
  XNOR U14177 ( .A(b[1804]), .B(n10080), .Z(c[1804]) );
  XOR U14178 ( .A(n10081), .B(n10082), .Z(n10078) );
  ANDN U14179 ( .B(n10083), .A(n10084), .Z(n10081) );
  XNOR U14180 ( .A(b[1803]), .B(n10082), .Z(n10083) );
  XNOR U14181 ( .A(b[1803]), .B(n10084), .Z(c[1803]) );
  XOR U14182 ( .A(n10085), .B(n10086), .Z(n10082) );
  ANDN U14183 ( .B(n10087), .A(n10088), .Z(n10085) );
  XNOR U14184 ( .A(b[1802]), .B(n10086), .Z(n10087) );
  XNOR U14185 ( .A(b[1802]), .B(n10088), .Z(c[1802]) );
  XOR U14186 ( .A(n10089), .B(n10090), .Z(n10086) );
  ANDN U14187 ( .B(n10091), .A(n10092), .Z(n10089) );
  XNOR U14188 ( .A(b[1801]), .B(n10090), .Z(n10091) );
  XNOR U14189 ( .A(b[1801]), .B(n10092), .Z(c[1801]) );
  XOR U14190 ( .A(n10093), .B(n10094), .Z(n10090) );
  ANDN U14191 ( .B(n10095), .A(n10096), .Z(n10093) );
  XNOR U14192 ( .A(b[1800]), .B(n10094), .Z(n10095) );
  XNOR U14193 ( .A(b[1800]), .B(n10096), .Z(c[1800]) );
  XOR U14194 ( .A(n10097), .B(n10098), .Z(n10094) );
  ANDN U14195 ( .B(n10099), .A(n10100), .Z(n10097) );
  XNOR U14196 ( .A(b[1799]), .B(n10098), .Z(n10099) );
  XNOR U14197 ( .A(b[17]), .B(n10101), .Z(c[17]) );
  XNOR U14198 ( .A(b[179]), .B(n10102), .Z(c[179]) );
  XNOR U14199 ( .A(b[1799]), .B(n10100), .Z(c[1799]) );
  XOR U14200 ( .A(n10103), .B(n10104), .Z(n10098) );
  ANDN U14201 ( .B(n10105), .A(n10106), .Z(n10103) );
  XNOR U14202 ( .A(b[1798]), .B(n10104), .Z(n10105) );
  XNOR U14203 ( .A(b[1798]), .B(n10106), .Z(c[1798]) );
  XOR U14204 ( .A(n10107), .B(n10108), .Z(n10104) );
  ANDN U14205 ( .B(n10109), .A(n10110), .Z(n10107) );
  XNOR U14206 ( .A(b[1797]), .B(n10108), .Z(n10109) );
  XNOR U14207 ( .A(b[1797]), .B(n10110), .Z(c[1797]) );
  XOR U14208 ( .A(n10111), .B(n10112), .Z(n10108) );
  ANDN U14209 ( .B(n10113), .A(n10114), .Z(n10111) );
  XNOR U14210 ( .A(b[1796]), .B(n10112), .Z(n10113) );
  XNOR U14211 ( .A(b[1796]), .B(n10114), .Z(c[1796]) );
  XOR U14212 ( .A(n10115), .B(n10116), .Z(n10112) );
  ANDN U14213 ( .B(n10117), .A(n10118), .Z(n10115) );
  XNOR U14214 ( .A(b[1795]), .B(n10116), .Z(n10117) );
  XNOR U14215 ( .A(b[1795]), .B(n10118), .Z(c[1795]) );
  XOR U14216 ( .A(n10119), .B(n10120), .Z(n10116) );
  ANDN U14217 ( .B(n10121), .A(n10122), .Z(n10119) );
  XNOR U14218 ( .A(b[1794]), .B(n10120), .Z(n10121) );
  XNOR U14219 ( .A(b[1794]), .B(n10122), .Z(c[1794]) );
  XOR U14220 ( .A(n10123), .B(n10124), .Z(n10120) );
  ANDN U14221 ( .B(n10125), .A(n10126), .Z(n10123) );
  XNOR U14222 ( .A(b[1793]), .B(n10124), .Z(n10125) );
  XNOR U14223 ( .A(b[1793]), .B(n10126), .Z(c[1793]) );
  XOR U14224 ( .A(n10127), .B(n10128), .Z(n10124) );
  ANDN U14225 ( .B(n10129), .A(n10130), .Z(n10127) );
  XNOR U14226 ( .A(b[1792]), .B(n10128), .Z(n10129) );
  XNOR U14227 ( .A(b[1792]), .B(n10130), .Z(c[1792]) );
  XOR U14228 ( .A(n10131), .B(n10132), .Z(n10128) );
  ANDN U14229 ( .B(n10133), .A(n10134), .Z(n10131) );
  XNOR U14230 ( .A(b[1791]), .B(n10132), .Z(n10133) );
  XNOR U14231 ( .A(b[1791]), .B(n10134), .Z(c[1791]) );
  XOR U14232 ( .A(n10135), .B(n10136), .Z(n10132) );
  ANDN U14233 ( .B(n10137), .A(n10138), .Z(n10135) );
  XNOR U14234 ( .A(b[1790]), .B(n10136), .Z(n10137) );
  XNOR U14235 ( .A(b[1790]), .B(n10138), .Z(c[1790]) );
  XOR U14236 ( .A(n10139), .B(n10140), .Z(n10136) );
  ANDN U14237 ( .B(n10141), .A(n10142), .Z(n10139) );
  XNOR U14238 ( .A(b[1789]), .B(n10140), .Z(n10141) );
  XNOR U14239 ( .A(b[178]), .B(n10143), .Z(c[178]) );
  XNOR U14240 ( .A(b[1789]), .B(n10142), .Z(c[1789]) );
  XOR U14241 ( .A(n10144), .B(n10145), .Z(n10140) );
  ANDN U14242 ( .B(n10146), .A(n10147), .Z(n10144) );
  XNOR U14243 ( .A(b[1788]), .B(n10145), .Z(n10146) );
  XNOR U14244 ( .A(b[1788]), .B(n10147), .Z(c[1788]) );
  XOR U14245 ( .A(n10148), .B(n10149), .Z(n10145) );
  ANDN U14246 ( .B(n10150), .A(n10151), .Z(n10148) );
  XNOR U14247 ( .A(b[1787]), .B(n10149), .Z(n10150) );
  XNOR U14248 ( .A(b[1787]), .B(n10151), .Z(c[1787]) );
  XOR U14249 ( .A(n10152), .B(n10153), .Z(n10149) );
  ANDN U14250 ( .B(n10154), .A(n10155), .Z(n10152) );
  XNOR U14251 ( .A(b[1786]), .B(n10153), .Z(n10154) );
  XNOR U14252 ( .A(b[1786]), .B(n10155), .Z(c[1786]) );
  XOR U14253 ( .A(n10156), .B(n10157), .Z(n10153) );
  ANDN U14254 ( .B(n10158), .A(n10159), .Z(n10156) );
  XNOR U14255 ( .A(b[1785]), .B(n10157), .Z(n10158) );
  XNOR U14256 ( .A(b[1785]), .B(n10159), .Z(c[1785]) );
  XOR U14257 ( .A(n10160), .B(n10161), .Z(n10157) );
  ANDN U14258 ( .B(n10162), .A(n10163), .Z(n10160) );
  XNOR U14259 ( .A(b[1784]), .B(n10161), .Z(n10162) );
  XNOR U14260 ( .A(b[1784]), .B(n10163), .Z(c[1784]) );
  XOR U14261 ( .A(n10164), .B(n10165), .Z(n10161) );
  ANDN U14262 ( .B(n10166), .A(n10167), .Z(n10164) );
  XNOR U14263 ( .A(b[1783]), .B(n10165), .Z(n10166) );
  XNOR U14264 ( .A(b[1783]), .B(n10167), .Z(c[1783]) );
  XOR U14265 ( .A(n10168), .B(n10169), .Z(n10165) );
  ANDN U14266 ( .B(n10170), .A(n10171), .Z(n10168) );
  XNOR U14267 ( .A(b[1782]), .B(n10169), .Z(n10170) );
  XNOR U14268 ( .A(b[1782]), .B(n10171), .Z(c[1782]) );
  XOR U14269 ( .A(n10172), .B(n10173), .Z(n10169) );
  ANDN U14270 ( .B(n10174), .A(n10175), .Z(n10172) );
  XNOR U14271 ( .A(b[1781]), .B(n10173), .Z(n10174) );
  XNOR U14272 ( .A(b[1781]), .B(n10175), .Z(c[1781]) );
  XOR U14273 ( .A(n10176), .B(n10177), .Z(n10173) );
  ANDN U14274 ( .B(n10178), .A(n10179), .Z(n10176) );
  XNOR U14275 ( .A(b[1780]), .B(n10177), .Z(n10178) );
  XNOR U14276 ( .A(b[1780]), .B(n10179), .Z(c[1780]) );
  XOR U14277 ( .A(n10180), .B(n10181), .Z(n10177) );
  ANDN U14278 ( .B(n10182), .A(n10183), .Z(n10180) );
  XNOR U14279 ( .A(b[1779]), .B(n10181), .Z(n10182) );
  XNOR U14280 ( .A(b[177]), .B(n10184), .Z(c[177]) );
  XNOR U14281 ( .A(b[1779]), .B(n10183), .Z(c[1779]) );
  XOR U14282 ( .A(n10185), .B(n10186), .Z(n10181) );
  ANDN U14283 ( .B(n10187), .A(n10188), .Z(n10185) );
  XNOR U14284 ( .A(b[1778]), .B(n10186), .Z(n10187) );
  XNOR U14285 ( .A(b[1778]), .B(n10188), .Z(c[1778]) );
  XOR U14286 ( .A(n10189), .B(n10190), .Z(n10186) );
  ANDN U14287 ( .B(n10191), .A(n10192), .Z(n10189) );
  XNOR U14288 ( .A(b[1777]), .B(n10190), .Z(n10191) );
  XNOR U14289 ( .A(b[1777]), .B(n10192), .Z(c[1777]) );
  XOR U14290 ( .A(n10193), .B(n10194), .Z(n10190) );
  ANDN U14291 ( .B(n10195), .A(n10196), .Z(n10193) );
  XNOR U14292 ( .A(b[1776]), .B(n10194), .Z(n10195) );
  XNOR U14293 ( .A(b[1776]), .B(n10196), .Z(c[1776]) );
  XOR U14294 ( .A(n10197), .B(n10198), .Z(n10194) );
  ANDN U14295 ( .B(n10199), .A(n10200), .Z(n10197) );
  XNOR U14296 ( .A(b[1775]), .B(n10198), .Z(n10199) );
  XNOR U14297 ( .A(b[1775]), .B(n10200), .Z(c[1775]) );
  XOR U14298 ( .A(n10201), .B(n10202), .Z(n10198) );
  ANDN U14299 ( .B(n10203), .A(n10204), .Z(n10201) );
  XNOR U14300 ( .A(b[1774]), .B(n10202), .Z(n10203) );
  XNOR U14301 ( .A(b[1774]), .B(n10204), .Z(c[1774]) );
  XOR U14302 ( .A(n10205), .B(n10206), .Z(n10202) );
  ANDN U14303 ( .B(n10207), .A(n10208), .Z(n10205) );
  XNOR U14304 ( .A(b[1773]), .B(n10206), .Z(n10207) );
  XNOR U14305 ( .A(b[1773]), .B(n10208), .Z(c[1773]) );
  XOR U14306 ( .A(n10209), .B(n10210), .Z(n10206) );
  ANDN U14307 ( .B(n10211), .A(n10212), .Z(n10209) );
  XNOR U14308 ( .A(b[1772]), .B(n10210), .Z(n10211) );
  XNOR U14309 ( .A(b[1772]), .B(n10212), .Z(c[1772]) );
  XOR U14310 ( .A(n10213), .B(n10214), .Z(n10210) );
  ANDN U14311 ( .B(n10215), .A(n10216), .Z(n10213) );
  XNOR U14312 ( .A(b[1771]), .B(n10214), .Z(n10215) );
  XNOR U14313 ( .A(b[1771]), .B(n10216), .Z(c[1771]) );
  XOR U14314 ( .A(n10217), .B(n10218), .Z(n10214) );
  ANDN U14315 ( .B(n10219), .A(n10220), .Z(n10217) );
  XNOR U14316 ( .A(b[1770]), .B(n10218), .Z(n10219) );
  XNOR U14317 ( .A(b[1770]), .B(n10220), .Z(c[1770]) );
  XOR U14318 ( .A(n10221), .B(n10222), .Z(n10218) );
  ANDN U14319 ( .B(n10223), .A(n10224), .Z(n10221) );
  XNOR U14320 ( .A(b[1769]), .B(n10222), .Z(n10223) );
  XNOR U14321 ( .A(b[176]), .B(n10225), .Z(c[176]) );
  XNOR U14322 ( .A(b[1769]), .B(n10224), .Z(c[1769]) );
  XOR U14323 ( .A(n10226), .B(n10227), .Z(n10222) );
  ANDN U14324 ( .B(n10228), .A(n10229), .Z(n10226) );
  XNOR U14325 ( .A(b[1768]), .B(n10227), .Z(n10228) );
  XNOR U14326 ( .A(b[1768]), .B(n10229), .Z(c[1768]) );
  XOR U14327 ( .A(n10230), .B(n10231), .Z(n10227) );
  ANDN U14328 ( .B(n10232), .A(n10233), .Z(n10230) );
  XNOR U14329 ( .A(b[1767]), .B(n10231), .Z(n10232) );
  XNOR U14330 ( .A(b[1767]), .B(n10233), .Z(c[1767]) );
  XOR U14331 ( .A(n10234), .B(n10235), .Z(n10231) );
  ANDN U14332 ( .B(n10236), .A(n10237), .Z(n10234) );
  XNOR U14333 ( .A(b[1766]), .B(n10235), .Z(n10236) );
  XNOR U14334 ( .A(b[1766]), .B(n10237), .Z(c[1766]) );
  XOR U14335 ( .A(n10238), .B(n10239), .Z(n10235) );
  ANDN U14336 ( .B(n10240), .A(n10241), .Z(n10238) );
  XNOR U14337 ( .A(b[1765]), .B(n10239), .Z(n10240) );
  XNOR U14338 ( .A(b[1765]), .B(n10241), .Z(c[1765]) );
  XOR U14339 ( .A(n10242), .B(n10243), .Z(n10239) );
  ANDN U14340 ( .B(n10244), .A(n10245), .Z(n10242) );
  XNOR U14341 ( .A(b[1764]), .B(n10243), .Z(n10244) );
  XNOR U14342 ( .A(b[1764]), .B(n10245), .Z(c[1764]) );
  XOR U14343 ( .A(n10246), .B(n10247), .Z(n10243) );
  ANDN U14344 ( .B(n10248), .A(n10249), .Z(n10246) );
  XNOR U14345 ( .A(b[1763]), .B(n10247), .Z(n10248) );
  XNOR U14346 ( .A(b[1763]), .B(n10249), .Z(c[1763]) );
  XOR U14347 ( .A(n10250), .B(n10251), .Z(n10247) );
  ANDN U14348 ( .B(n10252), .A(n10253), .Z(n10250) );
  XNOR U14349 ( .A(b[1762]), .B(n10251), .Z(n10252) );
  XNOR U14350 ( .A(b[1762]), .B(n10253), .Z(c[1762]) );
  XOR U14351 ( .A(n10254), .B(n10255), .Z(n10251) );
  ANDN U14352 ( .B(n10256), .A(n10257), .Z(n10254) );
  XNOR U14353 ( .A(b[1761]), .B(n10255), .Z(n10256) );
  XNOR U14354 ( .A(b[1761]), .B(n10257), .Z(c[1761]) );
  XOR U14355 ( .A(n10258), .B(n10259), .Z(n10255) );
  ANDN U14356 ( .B(n10260), .A(n10261), .Z(n10258) );
  XNOR U14357 ( .A(b[1760]), .B(n10259), .Z(n10260) );
  XNOR U14358 ( .A(b[1760]), .B(n10261), .Z(c[1760]) );
  XOR U14359 ( .A(n10262), .B(n10263), .Z(n10259) );
  ANDN U14360 ( .B(n10264), .A(n10265), .Z(n10262) );
  XNOR U14361 ( .A(b[1759]), .B(n10263), .Z(n10264) );
  XNOR U14362 ( .A(b[175]), .B(n10266), .Z(c[175]) );
  XNOR U14363 ( .A(b[1759]), .B(n10265), .Z(c[1759]) );
  XOR U14364 ( .A(n10267), .B(n10268), .Z(n10263) );
  ANDN U14365 ( .B(n10269), .A(n10270), .Z(n10267) );
  XNOR U14366 ( .A(b[1758]), .B(n10268), .Z(n10269) );
  XNOR U14367 ( .A(b[1758]), .B(n10270), .Z(c[1758]) );
  XOR U14368 ( .A(n10271), .B(n10272), .Z(n10268) );
  ANDN U14369 ( .B(n10273), .A(n10274), .Z(n10271) );
  XNOR U14370 ( .A(b[1757]), .B(n10272), .Z(n10273) );
  XNOR U14371 ( .A(b[1757]), .B(n10274), .Z(c[1757]) );
  XOR U14372 ( .A(n10275), .B(n10276), .Z(n10272) );
  ANDN U14373 ( .B(n10277), .A(n10278), .Z(n10275) );
  XNOR U14374 ( .A(b[1756]), .B(n10276), .Z(n10277) );
  XNOR U14375 ( .A(b[1756]), .B(n10278), .Z(c[1756]) );
  XOR U14376 ( .A(n10279), .B(n10280), .Z(n10276) );
  ANDN U14377 ( .B(n10281), .A(n10282), .Z(n10279) );
  XNOR U14378 ( .A(b[1755]), .B(n10280), .Z(n10281) );
  XNOR U14379 ( .A(b[1755]), .B(n10282), .Z(c[1755]) );
  XOR U14380 ( .A(n10283), .B(n10284), .Z(n10280) );
  ANDN U14381 ( .B(n10285), .A(n10286), .Z(n10283) );
  XNOR U14382 ( .A(b[1754]), .B(n10284), .Z(n10285) );
  XNOR U14383 ( .A(b[1754]), .B(n10286), .Z(c[1754]) );
  XOR U14384 ( .A(n10287), .B(n10288), .Z(n10284) );
  ANDN U14385 ( .B(n10289), .A(n10290), .Z(n10287) );
  XNOR U14386 ( .A(b[1753]), .B(n10288), .Z(n10289) );
  XNOR U14387 ( .A(b[1753]), .B(n10290), .Z(c[1753]) );
  XOR U14388 ( .A(n10291), .B(n10292), .Z(n10288) );
  ANDN U14389 ( .B(n10293), .A(n10294), .Z(n10291) );
  XNOR U14390 ( .A(b[1752]), .B(n10292), .Z(n10293) );
  XNOR U14391 ( .A(b[1752]), .B(n10294), .Z(c[1752]) );
  XOR U14392 ( .A(n10295), .B(n10296), .Z(n10292) );
  ANDN U14393 ( .B(n10297), .A(n10298), .Z(n10295) );
  XNOR U14394 ( .A(b[1751]), .B(n10296), .Z(n10297) );
  XNOR U14395 ( .A(b[1751]), .B(n10298), .Z(c[1751]) );
  XOR U14396 ( .A(n10299), .B(n10300), .Z(n10296) );
  ANDN U14397 ( .B(n10301), .A(n10302), .Z(n10299) );
  XNOR U14398 ( .A(b[1750]), .B(n10300), .Z(n10301) );
  XNOR U14399 ( .A(b[1750]), .B(n10302), .Z(c[1750]) );
  XOR U14400 ( .A(n10303), .B(n10304), .Z(n10300) );
  ANDN U14401 ( .B(n10305), .A(n10306), .Z(n10303) );
  XNOR U14402 ( .A(b[1749]), .B(n10304), .Z(n10305) );
  XNOR U14403 ( .A(b[174]), .B(n10307), .Z(c[174]) );
  XNOR U14404 ( .A(b[1749]), .B(n10306), .Z(c[1749]) );
  XOR U14405 ( .A(n10308), .B(n10309), .Z(n10304) );
  ANDN U14406 ( .B(n10310), .A(n10311), .Z(n10308) );
  XNOR U14407 ( .A(b[1748]), .B(n10309), .Z(n10310) );
  XNOR U14408 ( .A(b[1748]), .B(n10311), .Z(c[1748]) );
  XOR U14409 ( .A(n10312), .B(n10313), .Z(n10309) );
  ANDN U14410 ( .B(n10314), .A(n10315), .Z(n10312) );
  XNOR U14411 ( .A(b[1747]), .B(n10313), .Z(n10314) );
  XNOR U14412 ( .A(b[1747]), .B(n10315), .Z(c[1747]) );
  XOR U14413 ( .A(n10316), .B(n10317), .Z(n10313) );
  ANDN U14414 ( .B(n10318), .A(n10319), .Z(n10316) );
  XNOR U14415 ( .A(b[1746]), .B(n10317), .Z(n10318) );
  XNOR U14416 ( .A(b[1746]), .B(n10319), .Z(c[1746]) );
  XOR U14417 ( .A(n10320), .B(n10321), .Z(n10317) );
  ANDN U14418 ( .B(n10322), .A(n10323), .Z(n10320) );
  XNOR U14419 ( .A(b[1745]), .B(n10321), .Z(n10322) );
  XNOR U14420 ( .A(b[1745]), .B(n10323), .Z(c[1745]) );
  XOR U14421 ( .A(n10324), .B(n10325), .Z(n10321) );
  ANDN U14422 ( .B(n10326), .A(n10327), .Z(n10324) );
  XNOR U14423 ( .A(b[1744]), .B(n10325), .Z(n10326) );
  XNOR U14424 ( .A(b[1744]), .B(n10327), .Z(c[1744]) );
  XOR U14425 ( .A(n10328), .B(n10329), .Z(n10325) );
  ANDN U14426 ( .B(n10330), .A(n10331), .Z(n10328) );
  XNOR U14427 ( .A(b[1743]), .B(n10329), .Z(n10330) );
  XNOR U14428 ( .A(b[1743]), .B(n10331), .Z(c[1743]) );
  XOR U14429 ( .A(n10332), .B(n10333), .Z(n10329) );
  ANDN U14430 ( .B(n10334), .A(n10335), .Z(n10332) );
  XNOR U14431 ( .A(b[1742]), .B(n10333), .Z(n10334) );
  XNOR U14432 ( .A(b[1742]), .B(n10335), .Z(c[1742]) );
  XOR U14433 ( .A(n10336), .B(n10337), .Z(n10333) );
  ANDN U14434 ( .B(n10338), .A(n10339), .Z(n10336) );
  XNOR U14435 ( .A(b[1741]), .B(n10337), .Z(n10338) );
  XNOR U14436 ( .A(b[1741]), .B(n10339), .Z(c[1741]) );
  XOR U14437 ( .A(n10340), .B(n10341), .Z(n10337) );
  ANDN U14438 ( .B(n10342), .A(n10343), .Z(n10340) );
  XNOR U14439 ( .A(b[1740]), .B(n10341), .Z(n10342) );
  XNOR U14440 ( .A(b[1740]), .B(n10343), .Z(c[1740]) );
  XOR U14441 ( .A(n10344), .B(n10345), .Z(n10341) );
  ANDN U14442 ( .B(n10346), .A(n10347), .Z(n10344) );
  XNOR U14443 ( .A(b[1739]), .B(n10345), .Z(n10346) );
  XNOR U14444 ( .A(b[173]), .B(n10348), .Z(c[173]) );
  XNOR U14445 ( .A(b[1739]), .B(n10347), .Z(c[1739]) );
  XOR U14446 ( .A(n10349), .B(n10350), .Z(n10345) );
  ANDN U14447 ( .B(n10351), .A(n10352), .Z(n10349) );
  XNOR U14448 ( .A(b[1738]), .B(n10350), .Z(n10351) );
  XNOR U14449 ( .A(b[1738]), .B(n10352), .Z(c[1738]) );
  XOR U14450 ( .A(n10353), .B(n10354), .Z(n10350) );
  ANDN U14451 ( .B(n10355), .A(n10356), .Z(n10353) );
  XNOR U14452 ( .A(b[1737]), .B(n10354), .Z(n10355) );
  XNOR U14453 ( .A(b[1737]), .B(n10356), .Z(c[1737]) );
  XOR U14454 ( .A(n10357), .B(n10358), .Z(n10354) );
  ANDN U14455 ( .B(n10359), .A(n10360), .Z(n10357) );
  XNOR U14456 ( .A(b[1736]), .B(n10358), .Z(n10359) );
  XNOR U14457 ( .A(b[1736]), .B(n10360), .Z(c[1736]) );
  XOR U14458 ( .A(n10361), .B(n10362), .Z(n10358) );
  ANDN U14459 ( .B(n10363), .A(n10364), .Z(n10361) );
  XNOR U14460 ( .A(b[1735]), .B(n10362), .Z(n10363) );
  XNOR U14461 ( .A(b[1735]), .B(n10364), .Z(c[1735]) );
  XOR U14462 ( .A(n10365), .B(n10366), .Z(n10362) );
  ANDN U14463 ( .B(n10367), .A(n10368), .Z(n10365) );
  XNOR U14464 ( .A(b[1734]), .B(n10366), .Z(n10367) );
  XNOR U14465 ( .A(b[1734]), .B(n10368), .Z(c[1734]) );
  XOR U14466 ( .A(n10369), .B(n10370), .Z(n10366) );
  ANDN U14467 ( .B(n10371), .A(n10372), .Z(n10369) );
  XNOR U14468 ( .A(b[1733]), .B(n10370), .Z(n10371) );
  XNOR U14469 ( .A(b[1733]), .B(n10372), .Z(c[1733]) );
  XOR U14470 ( .A(n10373), .B(n10374), .Z(n10370) );
  ANDN U14471 ( .B(n10375), .A(n10376), .Z(n10373) );
  XNOR U14472 ( .A(b[1732]), .B(n10374), .Z(n10375) );
  XNOR U14473 ( .A(b[1732]), .B(n10376), .Z(c[1732]) );
  XOR U14474 ( .A(n10377), .B(n10378), .Z(n10374) );
  ANDN U14475 ( .B(n10379), .A(n10380), .Z(n10377) );
  XNOR U14476 ( .A(b[1731]), .B(n10378), .Z(n10379) );
  XNOR U14477 ( .A(b[1731]), .B(n10380), .Z(c[1731]) );
  XOR U14478 ( .A(n10381), .B(n10382), .Z(n10378) );
  ANDN U14479 ( .B(n10383), .A(n10384), .Z(n10381) );
  XNOR U14480 ( .A(b[1730]), .B(n10382), .Z(n10383) );
  XNOR U14481 ( .A(b[1730]), .B(n10384), .Z(c[1730]) );
  XOR U14482 ( .A(n10385), .B(n10386), .Z(n10382) );
  ANDN U14483 ( .B(n10387), .A(n10388), .Z(n10385) );
  XNOR U14484 ( .A(b[1729]), .B(n10386), .Z(n10387) );
  XNOR U14485 ( .A(b[172]), .B(n10389), .Z(c[172]) );
  XNOR U14486 ( .A(b[1729]), .B(n10388), .Z(c[1729]) );
  XOR U14487 ( .A(n10390), .B(n10391), .Z(n10386) );
  ANDN U14488 ( .B(n10392), .A(n10393), .Z(n10390) );
  XNOR U14489 ( .A(b[1728]), .B(n10391), .Z(n10392) );
  XNOR U14490 ( .A(b[1728]), .B(n10393), .Z(c[1728]) );
  XOR U14491 ( .A(n10394), .B(n10395), .Z(n10391) );
  ANDN U14492 ( .B(n10396), .A(n10397), .Z(n10394) );
  XNOR U14493 ( .A(b[1727]), .B(n10395), .Z(n10396) );
  XNOR U14494 ( .A(b[1727]), .B(n10397), .Z(c[1727]) );
  XOR U14495 ( .A(n10398), .B(n10399), .Z(n10395) );
  ANDN U14496 ( .B(n10400), .A(n10401), .Z(n10398) );
  XNOR U14497 ( .A(b[1726]), .B(n10399), .Z(n10400) );
  XNOR U14498 ( .A(b[1726]), .B(n10401), .Z(c[1726]) );
  XOR U14499 ( .A(n10402), .B(n10403), .Z(n10399) );
  ANDN U14500 ( .B(n10404), .A(n10405), .Z(n10402) );
  XNOR U14501 ( .A(b[1725]), .B(n10403), .Z(n10404) );
  XNOR U14502 ( .A(b[1725]), .B(n10405), .Z(c[1725]) );
  XOR U14503 ( .A(n10406), .B(n10407), .Z(n10403) );
  ANDN U14504 ( .B(n10408), .A(n10409), .Z(n10406) );
  XNOR U14505 ( .A(b[1724]), .B(n10407), .Z(n10408) );
  XNOR U14506 ( .A(b[1724]), .B(n10409), .Z(c[1724]) );
  XOR U14507 ( .A(n10410), .B(n10411), .Z(n10407) );
  ANDN U14508 ( .B(n10412), .A(n10413), .Z(n10410) );
  XNOR U14509 ( .A(b[1723]), .B(n10411), .Z(n10412) );
  XNOR U14510 ( .A(b[1723]), .B(n10413), .Z(c[1723]) );
  XOR U14511 ( .A(n10414), .B(n10415), .Z(n10411) );
  ANDN U14512 ( .B(n10416), .A(n10417), .Z(n10414) );
  XNOR U14513 ( .A(b[1722]), .B(n10415), .Z(n10416) );
  XNOR U14514 ( .A(b[1722]), .B(n10417), .Z(c[1722]) );
  XOR U14515 ( .A(n10418), .B(n10419), .Z(n10415) );
  ANDN U14516 ( .B(n10420), .A(n10421), .Z(n10418) );
  XNOR U14517 ( .A(b[1721]), .B(n10419), .Z(n10420) );
  XNOR U14518 ( .A(b[1721]), .B(n10421), .Z(c[1721]) );
  XOR U14519 ( .A(n10422), .B(n10423), .Z(n10419) );
  ANDN U14520 ( .B(n10424), .A(n10425), .Z(n10422) );
  XNOR U14521 ( .A(b[1720]), .B(n10423), .Z(n10424) );
  XNOR U14522 ( .A(b[1720]), .B(n10425), .Z(c[1720]) );
  XOR U14523 ( .A(n10426), .B(n10427), .Z(n10423) );
  ANDN U14524 ( .B(n10428), .A(n10429), .Z(n10426) );
  XNOR U14525 ( .A(b[1719]), .B(n10427), .Z(n10428) );
  XNOR U14526 ( .A(b[171]), .B(n10430), .Z(c[171]) );
  XNOR U14527 ( .A(b[1719]), .B(n10429), .Z(c[1719]) );
  XOR U14528 ( .A(n10431), .B(n10432), .Z(n10427) );
  ANDN U14529 ( .B(n10433), .A(n10434), .Z(n10431) );
  XNOR U14530 ( .A(b[1718]), .B(n10432), .Z(n10433) );
  XNOR U14531 ( .A(b[1718]), .B(n10434), .Z(c[1718]) );
  XOR U14532 ( .A(n10435), .B(n10436), .Z(n10432) );
  ANDN U14533 ( .B(n10437), .A(n10438), .Z(n10435) );
  XNOR U14534 ( .A(b[1717]), .B(n10436), .Z(n10437) );
  XNOR U14535 ( .A(b[1717]), .B(n10438), .Z(c[1717]) );
  XOR U14536 ( .A(n10439), .B(n10440), .Z(n10436) );
  ANDN U14537 ( .B(n10441), .A(n10442), .Z(n10439) );
  XNOR U14538 ( .A(b[1716]), .B(n10440), .Z(n10441) );
  XNOR U14539 ( .A(b[1716]), .B(n10442), .Z(c[1716]) );
  XOR U14540 ( .A(n10443), .B(n10444), .Z(n10440) );
  ANDN U14541 ( .B(n10445), .A(n10446), .Z(n10443) );
  XNOR U14542 ( .A(b[1715]), .B(n10444), .Z(n10445) );
  XNOR U14543 ( .A(b[1715]), .B(n10446), .Z(c[1715]) );
  XOR U14544 ( .A(n10447), .B(n10448), .Z(n10444) );
  ANDN U14545 ( .B(n10449), .A(n10450), .Z(n10447) );
  XNOR U14546 ( .A(b[1714]), .B(n10448), .Z(n10449) );
  XNOR U14547 ( .A(b[1714]), .B(n10450), .Z(c[1714]) );
  XOR U14548 ( .A(n10451), .B(n10452), .Z(n10448) );
  ANDN U14549 ( .B(n10453), .A(n10454), .Z(n10451) );
  XNOR U14550 ( .A(b[1713]), .B(n10452), .Z(n10453) );
  XNOR U14551 ( .A(b[1713]), .B(n10454), .Z(c[1713]) );
  XOR U14552 ( .A(n10455), .B(n10456), .Z(n10452) );
  ANDN U14553 ( .B(n10457), .A(n10458), .Z(n10455) );
  XNOR U14554 ( .A(b[1712]), .B(n10456), .Z(n10457) );
  XNOR U14555 ( .A(b[1712]), .B(n10458), .Z(c[1712]) );
  XOR U14556 ( .A(n10459), .B(n10460), .Z(n10456) );
  ANDN U14557 ( .B(n10461), .A(n10462), .Z(n10459) );
  XNOR U14558 ( .A(b[1711]), .B(n10460), .Z(n10461) );
  XNOR U14559 ( .A(b[1711]), .B(n10462), .Z(c[1711]) );
  XOR U14560 ( .A(n10463), .B(n10464), .Z(n10460) );
  ANDN U14561 ( .B(n10465), .A(n10466), .Z(n10463) );
  XNOR U14562 ( .A(b[1710]), .B(n10464), .Z(n10465) );
  XNOR U14563 ( .A(b[1710]), .B(n10466), .Z(c[1710]) );
  XOR U14564 ( .A(n10467), .B(n10468), .Z(n10464) );
  ANDN U14565 ( .B(n10469), .A(n10470), .Z(n10467) );
  XNOR U14566 ( .A(b[1709]), .B(n10468), .Z(n10469) );
  XNOR U14567 ( .A(b[170]), .B(n10471), .Z(c[170]) );
  XNOR U14568 ( .A(b[1709]), .B(n10470), .Z(c[1709]) );
  XOR U14569 ( .A(n10472), .B(n10473), .Z(n10468) );
  ANDN U14570 ( .B(n10474), .A(n10475), .Z(n10472) );
  XNOR U14571 ( .A(b[1708]), .B(n10473), .Z(n10474) );
  XNOR U14572 ( .A(b[1708]), .B(n10475), .Z(c[1708]) );
  XOR U14573 ( .A(n10476), .B(n10477), .Z(n10473) );
  ANDN U14574 ( .B(n10478), .A(n10479), .Z(n10476) );
  XNOR U14575 ( .A(b[1707]), .B(n10477), .Z(n10478) );
  XNOR U14576 ( .A(b[1707]), .B(n10479), .Z(c[1707]) );
  XOR U14577 ( .A(n10480), .B(n10481), .Z(n10477) );
  ANDN U14578 ( .B(n10482), .A(n10483), .Z(n10480) );
  XNOR U14579 ( .A(b[1706]), .B(n10481), .Z(n10482) );
  XNOR U14580 ( .A(b[1706]), .B(n10483), .Z(c[1706]) );
  XOR U14581 ( .A(n10484), .B(n10485), .Z(n10481) );
  ANDN U14582 ( .B(n10486), .A(n10487), .Z(n10484) );
  XNOR U14583 ( .A(b[1705]), .B(n10485), .Z(n10486) );
  XNOR U14584 ( .A(b[1705]), .B(n10487), .Z(c[1705]) );
  XOR U14585 ( .A(n10488), .B(n10489), .Z(n10485) );
  ANDN U14586 ( .B(n10490), .A(n10491), .Z(n10488) );
  XNOR U14587 ( .A(b[1704]), .B(n10489), .Z(n10490) );
  XNOR U14588 ( .A(b[1704]), .B(n10491), .Z(c[1704]) );
  XOR U14589 ( .A(n10492), .B(n10493), .Z(n10489) );
  ANDN U14590 ( .B(n10494), .A(n10495), .Z(n10492) );
  XNOR U14591 ( .A(b[1703]), .B(n10493), .Z(n10494) );
  XNOR U14592 ( .A(b[1703]), .B(n10495), .Z(c[1703]) );
  XOR U14593 ( .A(n10496), .B(n10497), .Z(n10493) );
  ANDN U14594 ( .B(n10498), .A(n10499), .Z(n10496) );
  XNOR U14595 ( .A(b[1702]), .B(n10497), .Z(n10498) );
  XNOR U14596 ( .A(b[1702]), .B(n10499), .Z(c[1702]) );
  XOR U14597 ( .A(n10500), .B(n10501), .Z(n10497) );
  ANDN U14598 ( .B(n10502), .A(n10503), .Z(n10500) );
  XNOR U14599 ( .A(b[1701]), .B(n10501), .Z(n10502) );
  XNOR U14600 ( .A(b[1701]), .B(n10503), .Z(c[1701]) );
  XOR U14601 ( .A(n10504), .B(n10505), .Z(n10501) );
  ANDN U14602 ( .B(n10506), .A(n10507), .Z(n10504) );
  XNOR U14603 ( .A(b[1700]), .B(n10505), .Z(n10506) );
  XNOR U14604 ( .A(b[1700]), .B(n10507), .Z(c[1700]) );
  XOR U14605 ( .A(n10508), .B(n10509), .Z(n10505) );
  ANDN U14606 ( .B(n10510), .A(n10511), .Z(n10508) );
  XNOR U14607 ( .A(b[1699]), .B(n10509), .Z(n10510) );
  XNOR U14608 ( .A(b[16]), .B(n10512), .Z(c[16]) );
  XNOR U14609 ( .A(b[169]), .B(n10513), .Z(c[169]) );
  XNOR U14610 ( .A(b[1699]), .B(n10511), .Z(c[1699]) );
  XOR U14611 ( .A(n10514), .B(n10515), .Z(n10509) );
  ANDN U14612 ( .B(n10516), .A(n10517), .Z(n10514) );
  XNOR U14613 ( .A(b[1698]), .B(n10515), .Z(n10516) );
  XNOR U14614 ( .A(b[1698]), .B(n10517), .Z(c[1698]) );
  XOR U14615 ( .A(n10518), .B(n10519), .Z(n10515) );
  ANDN U14616 ( .B(n10520), .A(n10521), .Z(n10518) );
  XNOR U14617 ( .A(b[1697]), .B(n10519), .Z(n10520) );
  XNOR U14618 ( .A(b[1697]), .B(n10521), .Z(c[1697]) );
  XOR U14619 ( .A(n10522), .B(n10523), .Z(n10519) );
  ANDN U14620 ( .B(n10524), .A(n10525), .Z(n10522) );
  XNOR U14621 ( .A(b[1696]), .B(n10523), .Z(n10524) );
  XNOR U14622 ( .A(b[1696]), .B(n10525), .Z(c[1696]) );
  XOR U14623 ( .A(n10526), .B(n10527), .Z(n10523) );
  ANDN U14624 ( .B(n10528), .A(n10529), .Z(n10526) );
  XNOR U14625 ( .A(b[1695]), .B(n10527), .Z(n10528) );
  XNOR U14626 ( .A(b[1695]), .B(n10529), .Z(c[1695]) );
  XOR U14627 ( .A(n10530), .B(n10531), .Z(n10527) );
  ANDN U14628 ( .B(n10532), .A(n10533), .Z(n10530) );
  XNOR U14629 ( .A(b[1694]), .B(n10531), .Z(n10532) );
  XNOR U14630 ( .A(b[1694]), .B(n10533), .Z(c[1694]) );
  XOR U14631 ( .A(n10534), .B(n10535), .Z(n10531) );
  ANDN U14632 ( .B(n10536), .A(n10537), .Z(n10534) );
  XNOR U14633 ( .A(b[1693]), .B(n10535), .Z(n10536) );
  XNOR U14634 ( .A(b[1693]), .B(n10537), .Z(c[1693]) );
  XOR U14635 ( .A(n10538), .B(n10539), .Z(n10535) );
  ANDN U14636 ( .B(n10540), .A(n10541), .Z(n10538) );
  XNOR U14637 ( .A(b[1692]), .B(n10539), .Z(n10540) );
  XNOR U14638 ( .A(b[1692]), .B(n10541), .Z(c[1692]) );
  XOR U14639 ( .A(n10542), .B(n10543), .Z(n10539) );
  ANDN U14640 ( .B(n10544), .A(n10545), .Z(n10542) );
  XNOR U14641 ( .A(b[1691]), .B(n10543), .Z(n10544) );
  XNOR U14642 ( .A(b[1691]), .B(n10545), .Z(c[1691]) );
  XOR U14643 ( .A(n10546), .B(n10547), .Z(n10543) );
  ANDN U14644 ( .B(n10548), .A(n10549), .Z(n10546) );
  XNOR U14645 ( .A(b[1690]), .B(n10547), .Z(n10548) );
  XNOR U14646 ( .A(b[1690]), .B(n10549), .Z(c[1690]) );
  XOR U14647 ( .A(n10550), .B(n10551), .Z(n10547) );
  ANDN U14648 ( .B(n10552), .A(n10553), .Z(n10550) );
  XNOR U14649 ( .A(b[1689]), .B(n10551), .Z(n10552) );
  XNOR U14650 ( .A(b[168]), .B(n10554), .Z(c[168]) );
  XNOR U14651 ( .A(b[1689]), .B(n10553), .Z(c[1689]) );
  XOR U14652 ( .A(n10555), .B(n10556), .Z(n10551) );
  ANDN U14653 ( .B(n10557), .A(n10558), .Z(n10555) );
  XNOR U14654 ( .A(b[1688]), .B(n10556), .Z(n10557) );
  XNOR U14655 ( .A(b[1688]), .B(n10558), .Z(c[1688]) );
  XOR U14656 ( .A(n10559), .B(n10560), .Z(n10556) );
  ANDN U14657 ( .B(n10561), .A(n10562), .Z(n10559) );
  XNOR U14658 ( .A(b[1687]), .B(n10560), .Z(n10561) );
  XNOR U14659 ( .A(b[1687]), .B(n10562), .Z(c[1687]) );
  XOR U14660 ( .A(n10563), .B(n10564), .Z(n10560) );
  ANDN U14661 ( .B(n10565), .A(n10566), .Z(n10563) );
  XNOR U14662 ( .A(b[1686]), .B(n10564), .Z(n10565) );
  XNOR U14663 ( .A(b[1686]), .B(n10566), .Z(c[1686]) );
  XOR U14664 ( .A(n10567), .B(n10568), .Z(n10564) );
  ANDN U14665 ( .B(n10569), .A(n10570), .Z(n10567) );
  XNOR U14666 ( .A(b[1685]), .B(n10568), .Z(n10569) );
  XNOR U14667 ( .A(b[1685]), .B(n10570), .Z(c[1685]) );
  XOR U14668 ( .A(n10571), .B(n10572), .Z(n10568) );
  ANDN U14669 ( .B(n10573), .A(n10574), .Z(n10571) );
  XNOR U14670 ( .A(b[1684]), .B(n10572), .Z(n10573) );
  XNOR U14671 ( .A(b[1684]), .B(n10574), .Z(c[1684]) );
  XOR U14672 ( .A(n10575), .B(n10576), .Z(n10572) );
  ANDN U14673 ( .B(n10577), .A(n10578), .Z(n10575) );
  XNOR U14674 ( .A(b[1683]), .B(n10576), .Z(n10577) );
  XNOR U14675 ( .A(b[1683]), .B(n10578), .Z(c[1683]) );
  XOR U14676 ( .A(n10579), .B(n10580), .Z(n10576) );
  ANDN U14677 ( .B(n10581), .A(n10582), .Z(n10579) );
  XNOR U14678 ( .A(b[1682]), .B(n10580), .Z(n10581) );
  XNOR U14679 ( .A(b[1682]), .B(n10582), .Z(c[1682]) );
  XOR U14680 ( .A(n10583), .B(n10584), .Z(n10580) );
  ANDN U14681 ( .B(n10585), .A(n10586), .Z(n10583) );
  XNOR U14682 ( .A(b[1681]), .B(n10584), .Z(n10585) );
  XNOR U14683 ( .A(b[1681]), .B(n10586), .Z(c[1681]) );
  XOR U14684 ( .A(n10587), .B(n10588), .Z(n10584) );
  ANDN U14685 ( .B(n10589), .A(n10590), .Z(n10587) );
  XNOR U14686 ( .A(b[1680]), .B(n10588), .Z(n10589) );
  XNOR U14687 ( .A(b[1680]), .B(n10590), .Z(c[1680]) );
  XOR U14688 ( .A(n10591), .B(n10592), .Z(n10588) );
  ANDN U14689 ( .B(n10593), .A(n10594), .Z(n10591) );
  XNOR U14690 ( .A(b[1679]), .B(n10592), .Z(n10593) );
  XNOR U14691 ( .A(b[167]), .B(n10595), .Z(c[167]) );
  XNOR U14692 ( .A(b[1679]), .B(n10594), .Z(c[1679]) );
  XOR U14693 ( .A(n10596), .B(n10597), .Z(n10592) );
  ANDN U14694 ( .B(n10598), .A(n10599), .Z(n10596) );
  XNOR U14695 ( .A(b[1678]), .B(n10597), .Z(n10598) );
  XNOR U14696 ( .A(b[1678]), .B(n10599), .Z(c[1678]) );
  XOR U14697 ( .A(n10600), .B(n10601), .Z(n10597) );
  ANDN U14698 ( .B(n10602), .A(n10603), .Z(n10600) );
  XNOR U14699 ( .A(b[1677]), .B(n10601), .Z(n10602) );
  XNOR U14700 ( .A(b[1677]), .B(n10603), .Z(c[1677]) );
  XOR U14701 ( .A(n10604), .B(n10605), .Z(n10601) );
  ANDN U14702 ( .B(n10606), .A(n10607), .Z(n10604) );
  XNOR U14703 ( .A(b[1676]), .B(n10605), .Z(n10606) );
  XNOR U14704 ( .A(b[1676]), .B(n10607), .Z(c[1676]) );
  XOR U14705 ( .A(n10608), .B(n10609), .Z(n10605) );
  ANDN U14706 ( .B(n10610), .A(n10611), .Z(n10608) );
  XNOR U14707 ( .A(b[1675]), .B(n10609), .Z(n10610) );
  XNOR U14708 ( .A(b[1675]), .B(n10611), .Z(c[1675]) );
  XOR U14709 ( .A(n10612), .B(n10613), .Z(n10609) );
  ANDN U14710 ( .B(n10614), .A(n10615), .Z(n10612) );
  XNOR U14711 ( .A(b[1674]), .B(n10613), .Z(n10614) );
  XNOR U14712 ( .A(b[1674]), .B(n10615), .Z(c[1674]) );
  XOR U14713 ( .A(n10616), .B(n10617), .Z(n10613) );
  ANDN U14714 ( .B(n10618), .A(n10619), .Z(n10616) );
  XNOR U14715 ( .A(b[1673]), .B(n10617), .Z(n10618) );
  XNOR U14716 ( .A(b[1673]), .B(n10619), .Z(c[1673]) );
  XOR U14717 ( .A(n10620), .B(n10621), .Z(n10617) );
  ANDN U14718 ( .B(n10622), .A(n10623), .Z(n10620) );
  XNOR U14719 ( .A(b[1672]), .B(n10621), .Z(n10622) );
  XNOR U14720 ( .A(b[1672]), .B(n10623), .Z(c[1672]) );
  XOR U14721 ( .A(n10624), .B(n10625), .Z(n10621) );
  ANDN U14722 ( .B(n10626), .A(n10627), .Z(n10624) );
  XNOR U14723 ( .A(b[1671]), .B(n10625), .Z(n10626) );
  XNOR U14724 ( .A(b[1671]), .B(n10627), .Z(c[1671]) );
  XOR U14725 ( .A(n10628), .B(n10629), .Z(n10625) );
  ANDN U14726 ( .B(n10630), .A(n10631), .Z(n10628) );
  XNOR U14727 ( .A(b[1670]), .B(n10629), .Z(n10630) );
  XNOR U14728 ( .A(b[1670]), .B(n10631), .Z(c[1670]) );
  XOR U14729 ( .A(n10632), .B(n10633), .Z(n10629) );
  ANDN U14730 ( .B(n10634), .A(n10635), .Z(n10632) );
  XNOR U14731 ( .A(b[1669]), .B(n10633), .Z(n10634) );
  XNOR U14732 ( .A(b[166]), .B(n10636), .Z(c[166]) );
  XNOR U14733 ( .A(b[1669]), .B(n10635), .Z(c[1669]) );
  XOR U14734 ( .A(n10637), .B(n10638), .Z(n10633) );
  ANDN U14735 ( .B(n10639), .A(n10640), .Z(n10637) );
  XNOR U14736 ( .A(b[1668]), .B(n10638), .Z(n10639) );
  XNOR U14737 ( .A(b[1668]), .B(n10640), .Z(c[1668]) );
  XOR U14738 ( .A(n10641), .B(n10642), .Z(n10638) );
  ANDN U14739 ( .B(n10643), .A(n10644), .Z(n10641) );
  XNOR U14740 ( .A(b[1667]), .B(n10642), .Z(n10643) );
  XNOR U14741 ( .A(b[1667]), .B(n10644), .Z(c[1667]) );
  XOR U14742 ( .A(n10645), .B(n10646), .Z(n10642) );
  ANDN U14743 ( .B(n10647), .A(n10648), .Z(n10645) );
  XNOR U14744 ( .A(b[1666]), .B(n10646), .Z(n10647) );
  XNOR U14745 ( .A(b[1666]), .B(n10648), .Z(c[1666]) );
  XOR U14746 ( .A(n10649), .B(n10650), .Z(n10646) );
  ANDN U14747 ( .B(n10651), .A(n10652), .Z(n10649) );
  XNOR U14748 ( .A(b[1665]), .B(n10650), .Z(n10651) );
  XNOR U14749 ( .A(b[1665]), .B(n10652), .Z(c[1665]) );
  XOR U14750 ( .A(n10653), .B(n10654), .Z(n10650) );
  ANDN U14751 ( .B(n10655), .A(n10656), .Z(n10653) );
  XNOR U14752 ( .A(b[1664]), .B(n10654), .Z(n10655) );
  XNOR U14753 ( .A(b[1664]), .B(n10656), .Z(c[1664]) );
  XOR U14754 ( .A(n10657), .B(n10658), .Z(n10654) );
  ANDN U14755 ( .B(n10659), .A(n10660), .Z(n10657) );
  XNOR U14756 ( .A(b[1663]), .B(n10658), .Z(n10659) );
  XNOR U14757 ( .A(b[1663]), .B(n10660), .Z(c[1663]) );
  XOR U14758 ( .A(n10661), .B(n10662), .Z(n10658) );
  ANDN U14759 ( .B(n10663), .A(n10664), .Z(n10661) );
  XNOR U14760 ( .A(b[1662]), .B(n10662), .Z(n10663) );
  XNOR U14761 ( .A(b[1662]), .B(n10664), .Z(c[1662]) );
  XOR U14762 ( .A(n10665), .B(n10666), .Z(n10662) );
  ANDN U14763 ( .B(n10667), .A(n10668), .Z(n10665) );
  XNOR U14764 ( .A(b[1661]), .B(n10666), .Z(n10667) );
  XNOR U14765 ( .A(b[1661]), .B(n10668), .Z(c[1661]) );
  XOR U14766 ( .A(n10669), .B(n10670), .Z(n10666) );
  ANDN U14767 ( .B(n10671), .A(n10672), .Z(n10669) );
  XNOR U14768 ( .A(b[1660]), .B(n10670), .Z(n10671) );
  XNOR U14769 ( .A(b[1660]), .B(n10672), .Z(c[1660]) );
  XOR U14770 ( .A(n10673), .B(n10674), .Z(n10670) );
  ANDN U14771 ( .B(n10675), .A(n10676), .Z(n10673) );
  XNOR U14772 ( .A(b[1659]), .B(n10674), .Z(n10675) );
  XNOR U14773 ( .A(b[165]), .B(n10677), .Z(c[165]) );
  XNOR U14774 ( .A(b[1659]), .B(n10676), .Z(c[1659]) );
  XOR U14775 ( .A(n10678), .B(n10679), .Z(n10674) );
  ANDN U14776 ( .B(n10680), .A(n10681), .Z(n10678) );
  XNOR U14777 ( .A(b[1658]), .B(n10679), .Z(n10680) );
  XNOR U14778 ( .A(b[1658]), .B(n10681), .Z(c[1658]) );
  XOR U14779 ( .A(n10682), .B(n10683), .Z(n10679) );
  ANDN U14780 ( .B(n10684), .A(n10685), .Z(n10682) );
  XNOR U14781 ( .A(b[1657]), .B(n10683), .Z(n10684) );
  XNOR U14782 ( .A(b[1657]), .B(n10685), .Z(c[1657]) );
  XOR U14783 ( .A(n10686), .B(n10687), .Z(n10683) );
  ANDN U14784 ( .B(n10688), .A(n10689), .Z(n10686) );
  XNOR U14785 ( .A(b[1656]), .B(n10687), .Z(n10688) );
  XNOR U14786 ( .A(b[1656]), .B(n10689), .Z(c[1656]) );
  XOR U14787 ( .A(n10690), .B(n10691), .Z(n10687) );
  ANDN U14788 ( .B(n10692), .A(n10693), .Z(n10690) );
  XNOR U14789 ( .A(b[1655]), .B(n10691), .Z(n10692) );
  XNOR U14790 ( .A(b[1655]), .B(n10693), .Z(c[1655]) );
  XOR U14791 ( .A(n10694), .B(n10695), .Z(n10691) );
  ANDN U14792 ( .B(n10696), .A(n10697), .Z(n10694) );
  XNOR U14793 ( .A(b[1654]), .B(n10695), .Z(n10696) );
  XNOR U14794 ( .A(b[1654]), .B(n10697), .Z(c[1654]) );
  XOR U14795 ( .A(n10698), .B(n10699), .Z(n10695) );
  ANDN U14796 ( .B(n10700), .A(n10701), .Z(n10698) );
  XNOR U14797 ( .A(b[1653]), .B(n10699), .Z(n10700) );
  XNOR U14798 ( .A(b[1653]), .B(n10701), .Z(c[1653]) );
  XOR U14799 ( .A(n10702), .B(n10703), .Z(n10699) );
  ANDN U14800 ( .B(n10704), .A(n10705), .Z(n10702) );
  XNOR U14801 ( .A(b[1652]), .B(n10703), .Z(n10704) );
  XNOR U14802 ( .A(b[1652]), .B(n10705), .Z(c[1652]) );
  XOR U14803 ( .A(n10706), .B(n10707), .Z(n10703) );
  ANDN U14804 ( .B(n10708), .A(n10709), .Z(n10706) );
  XNOR U14805 ( .A(b[1651]), .B(n10707), .Z(n10708) );
  XNOR U14806 ( .A(b[1651]), .B(n10709), .Z(c[1651]) );
  XOR U14807 ( .A(n10710), .B(n10711), .Z(n10707) );
  ANDN U14808 ( .B(n10712), .A(n10713), .Z(n10710) );
  XNOR U14809 ( .A(b[1650]), .B(n10711), .Z(n10712) );
  XNOR U14810 ( .A(b[1650]), .B(n10713), .Z(c[1650]) );
  XOR U14811 ( .A(n10714), .B(n10715), .Z(n10711) );
  ANDN U14812 ( .B(n10716), .A(n10717), .Z(n10714) );
  XNOR U14813 ( .A(b[1649]), .B(n10715), .Z(n10716) );
  XNOR U14814 ( .A(b[164]), .B(n10718), .Z(c[164]) );
  XNOR U14815 ( .A(b[1649]), .B(n10717), .Z(c[1649]) );
  XOR U14816 ( .A(n10719), .B(n10720), .Z(n10715) );
  ANDN U14817 ( .B(n10721), .A(n10722), .Z(n10719) );
  XNOR U14818 ( .A(b[1648]), .B(n10720), .Z(n10721) );
  XNOR U14819 ( .A(b[1648]), .B(n10722), .Z(c[1648]) );
  XOR U14820 ( .A(n10723), .B(n10724), .Z(n10720) );
  ANDN U14821 ( .B(n10725), .A(n10726), .Z(n10723) );
  XNOR U14822 ( .A(b[1647]), .B(n10724), .Z(n10725) );
  XNOR U14823 ( .A(b[1647]), .B(n10726), .Z(c[1647]) );
  XOR U14824 ( .A(n10727), .B(n10728), .Z(n10724) );
  ANDN U14825 ( .B(n10729), .A(n10730), .Z(n10727) );
  XNOR U14826 ( .A(b[1646]), .B(n10728), .Z(n10729) );
  XNOR U14827 ( .A(b[1646]), .B(n10730), .Z(c[1646]) );
  XOR U14828 ( .A(n10731), .B(n10732), .Z(n10728) );
  ANDN U14829 ( .B(n10733), .A(n10734), .Z(n10731) );
  XNOR U14830 ( .A(b[1645]), .B(n10732), .Z(n10733) );
  XNOR U14831 ( .A(b[1645]), .B(n10734), .Z(c[1645]) );
  XOR U14832 ( .A(n10735), .B(n10736), .Z(n10732) );
  ANDN U14833 ( .B(n10737), .A(n10738), .Z(n10735) );
  XNOR U14834 ( .A(b[1644]), .B(n10736), .Z(n10737) );
  XNOR U14835 ( .A(b[1644]), .B(n10738), .Z(c[1644]) );
  XOR U14836 ( .A(n10739), .B(n10740), .Z(n10736) );
  ANDN U14837 ( .B(n10741), .A(n10742), .Z(n10739) );
  XNOR U14838 ( .A(b[1643]), .B(n10740), .Z(n10741) );
  XNOR U14839 ( .A(b[1643]), .B(n10742), .Z(c[1643]) );
  XOR U14840 ( .A(n10743), .B(n10744), .Z(n10740) );
  ANDN U14841 ( .B(n10745), .A(n10746), .Z(n10743) );
  XNOR U14842 ( .A(b[1642]), .B(n10744), .Z(n10745) );
  XNOR U14843 ( .A(b[1642]), .B(n10746), .Z(c[1642]) );
  XOR U14844 ( .A(n10747), .B(n10748), .Z(n10744) );
  ANDN U14845 ( .B(n10749), .A(n10750), .Z(n10747) );
  XNOR U14846 ( .A(b[1641]), .B(n10748), .Z(n10749) );
  XNOR U14847 ( .A(b[1641]), .B(n10750), .Z(c[1641]) );
  XOR U14848 ( .A(n10751), .B(n10752), .Z(n10748) );
  ANDN U14849 ( .B(n10753), .A(n10754), .Z(n10751) );
  XNOR U14850 ( .A(b[1640]), .B(n10752), .Z(n10753) );
  XNOR U14851 ( .A(b[1640]), .B(n10754), .Z(c[1640]) );
  XOR U14852 ( .A(n10755), .B(n10756), .Z(n10752) );
  ANDN U14853 ( .B(n10757), .A(n10758), .Z(n10755) );
  XNOR U14854 ( .A(b[1639]), .B(n10756), .Z(n10757) );
  XNOR U14855 ( .A(b[163]), .B(n10759), .Z(c[163]) );
  XNOR U14856 ( .A(b[1639]), .B(n10758), .Z(c[1639]) );
  XOR U14857 ( .A(n10760), .B(n10761), .Z(n10756) );
  ANDN U14858 ( .B(n10762), .A(n10763), .Z(n10760) );
  XNOR U14859 ( .A(b[1638]), .B(n10761), .Z(n10762) );
  XNOR U14860 ( .A(b[1638]), .B(n10763), .Z(c[1638]) );
  XOR U14861 ( .A(n10764), .B(n10765), .Z(n10761) );
  ANDN U14862 ( .B(n10766), .A(n10767), .Z(n10764) );
  XNOR U14863 ( .A(b[1637]), .B(n10765), .Z(n10766) );
  XNOR U14864 ( .A(b[1637]), .B(n10767), .Z(c[1637]) );
  XOR U14865 ( .A(n10768), .B(n10769), .Z(n10765) );
  ANDN U14866 ( .B(n10770), .A(n10771), .Z(n10768) );
  XNOR U14867 ( .A(b[1636]), .B(n10769), .Z(n10770) );
  XNOR U14868 ( .A(b[1636]), .B(n10771), .Z(c[1636]) );
  XOR U14869 ( .A(n10772), .B(n10773), .Z(n10769) );
  ANDN U14870 ( .B(n10774), .A(n10775), .Z(n10772) );
  XNOR U14871 ( .A(b[1635]), .B(n10773), .Z(n10774) );
  XNOR U14872 ( .A(b[1635]), .B(n10775), .Z(c[1635]) );
  XOR U14873 ( .A(n10776), .B(n10777), .Z(n10773) );
  ANDN U14874 ( .B(n10778), .A(n10779), .Z(n10776) );
  XNOR U14875 ( .A(b[1634]), .B(n10777), .Z(n10778) );
  XNOR U14876 ( .A(b[1634]), .B(n10779), .Z(c[1634]) );
  XOR U14877 ( .A(n10780), .B(n10781), .Z(n10777) );
  ANDN U14878 ( .B(n10782), .A(n10783), .Z(n10780) );
  XNOR U14879 ( .A(b[1633]), .B(n10781), .Z(n10782) );
  XNOR U14880 ( .A(b[1633]), .B(n10783), .Z(c[1633]) );
  XOR U14881 ( .A(n10784), .B(n10785), .Z(n10781) );
  ANDN U14882 ( .B(n10786), .A(n10787), .Z(n10784) );
  XNOR U14883 ( .A(b[1632]), .B(n10785), .Z(n10786) );
  XNOR U14884 ( .A(b[1632]), .B(n10787), .Z(c[1632]) );
  XOR U14885 ( .A(n10788), .B(n10789), .Z(n10785) );
  ANDN U14886 ( .B(n10790), .A(n10791), .Z(n10788) );
  XNOR U14887 ( .A(b[1631]), .B(n10789), .Z(n10790) );
  XNOR U14888 ( .A(b[1631]), .B(n10791), .Z(c[1631]) );
  XOR U14889 ( .A(n10792), .B(n10793), .Z(n10789) );
  ANDN U14890 ( .B(n10794), .A(n10795), .Z(n10792) );
  XNOR U14891 ( .A(b[1630]), .B(n10793), .Z(n10794) );
  XNOR U14892 ( .A(b[1630]), .B(n10795), .Z(c[1630]) );
  XOR U14893 ( .A(n10796), .B(n10797), .Z(n10793) );
  ANDN U14894 ( .B(n10798), .A(n10799), .Z(n10796) );
  XNOR U14895 ( .A(b[1629]), .B(n10797), .Z(n10798) );
  XNOR U14896 ( .A(b[162]), .B(n10800), .Z(c[162]) );
  XNOR U14897 ( .A(b[1629]), .B(n10799), .Z(c[1629]) );
  XOR U14898 ( .A(n10801), .B(n10802), .Z(n10797) );
  ANDN U14899 ( .B(n10803), .A(n10804), .Z(n10801) );
  XNOR U14900 ( .A(b[1628]), .B(n10802), .Z(n10803) );
  XNOR U14901 ( .A(b[1628]), .B(n10804), .Z(c[1628]) );
  XOR U14902 ( .A(n10805), .B(n10806), .Z(n10802) );
  ANDN U14903 ( .B(n10807), .A(n10808), .Z(n10805) );
  XNOR U14904 ( .A(b[1627]), .B(n10806), .Z(n10807) );
  XNOR U14905 ( .A(b[1627]), .B(n10808), .Z(c[1627]) );
  XOR U14906 ( .A(n10809), .B(n10810), .Z(n10806) );
  ANDN U14907 ( .B(n10811), .A(n10812), .Z(n10809) );
  XNOR U14908 ( .A(b[1626]), .B(n10810), .Z(n10811) );
  XNOR U14909 ( .A(b[1626]), .B(n10812), .Z(c[1626]) );
  XOR U14910 ( .A(n10813), .B(n10814), .Z(n10810) );
  ANDN U14911 ( .B(n10815), .A(n10816), .Z(n10813) );
  XNOR U14912 ( .A(b[1625]), .B(n10814), .Z(n10815) );
  XNOR U14913 ( .A(b[1625]), .B(n10816), .Z(c[1625]) );
  XOR U14914 ( .A(n10817), .B(n10818), .Z(n10814) );
  ANDN U14915 ( .B(n10819), .A(n10820), .Z(n10817) );
  XNOR U14916 ( .A(b[1624]), .B(n10818), .Z(n10819) );
  XNOR U14917 ( .A(b[1624]), .B(n10820), .Z(c[1624]) );
  XOR U14918 ( .A(n10821), .B(n10822), .Z(n10818) );
  ANDN U14919 ( .B(n10823), .A(n10824), .Z(n10821) );
  XNOR U14920 ( .A(b[1623]), .B(n10822), .Z(n10823) );
  XNOR U14921 ( .A(b[1623]), .B(n10824), .Z(c[1623]) );
  XOR U14922 ( .A(n10825), .B(n10826), .Z(n10822) );
  ANDN U14923 ( .B(n10827), .A(n10828), .Z(n10825) );
  XNOR U14924 ( .A(b[1622]), .B(n10826), .Z(n10827) );
  XNOR U14925 ( .A(b[1622]), .B(n10828), .Z(c[1622]) );
  XOR U14926 ( .A(n10829), .B(n10830), .Z(n10826) );
  ANDN U14927 ( .B(n10831), .A(n10832), .Z(n10829) );
  XNOR U14928 ( .A(b[1621]), .B(n10830), .Z(n10831) );
  XNOR U14929 ( .A(b[1621]), .B(n10832), .Z(c[1621]) );
  XOR U14930 ( .A(n10833), .B(n10834), .Z(n10830) );
  ANDN U14931 ( .B(n10835), .A(n10836), .Z(n10833) );
  XNOR U14932 ( .A(b[1620]), .B(n10834), .Z(n10835) );
  XNOR U14933 ( .A(b[1620]), .B(n10836), .Z(c[1620]) );
  XOR U14934 ( .A(n10837), .B(n10838), .Z(n10834) );
  ANDN U14935 ( .B(n10839), .A(n10840), .Z(n10837) );
  XNOR U14936 ( .A(b[1619]), .B(n10838), .Z(n10839) );
  XNOR U14937 ( .A(b[161]), .B(n10841), .Z(c[161]) );
  XNOR U14938 ( .A(b[1619]), .B(n10840), .Z(c[1619]) );
  XOR U14939 ( .A(n10842), .B(n10843), .Z(n10838) );
  ANDN U14940 ( .B(n10844), .A(n10845), .Z(n10842) );
  XNOR U14941 ( .A(b[1618]), .B(n10843), .Z(n10844) );
  XNOR U14942 ( .A(b[1618]), .B(n10845), .Z(c[1618]) );
  XOR U14943 ( .A(n10846), .B(n10847), .Z(n10843) );
  ANDN U14944 ( .B(n10848), .A(n10849), .Z(n10846) );
  XNOR U14945 ( .A(b[1617]), .B(n10847), .Z(n10848) );
  XNOR U14946 ( .A(b[1617]), .B(n10849), .Z(c[1617]) );
  XOR U14947 ( .A(n10850), .B(n10851), .Z(n10847) );
  ANDN U14948 ( .B(n10852), .A(n10853), .Z(n10850) );
  XNOR U14949 ( .A(b[1616]), .B(n10851), .Z(n10852) );
  XNOR U14950 ( .A(b[1616]), .B(n10853), .Z(c[1616]) );
  XOR U14951 ( .A(n10854), .B(n10855), .Z(n10851) );
  ANDN U14952 ( .B(n10856), .A(n10857), .Z(n10854) );
  XNOR U14953 ( .A(b[1615]), .B(n10855), .Z(n10856) );
  XNOR U14954 ( .A(b[1615]), .B(n10857), .Z(c[1615]) );
  XOR U14955 ( .A(n10858), .B(n10859), .Z(n10855) );
  ANDN U14956 ( .B(n10860), .A(n10861), .Z(n10858) );
  XNOR U14957 ( .A(b[1614]), .B(n10859), .Z(n10860) );
  XNOR U14958 ( .A(b[1614]), .B(n10861), .Z(c[1614]) );
  XOR U14959 ( .A(n10862), .B(n10863), .Z(n10859) );
  ANDN U14960 ( .B(n10864), .A(n10865), .Z(n10862) );
  XNOR U14961 ( .A(b[1613]), .B(n10863), .Z(n10864) );
  XNOR U14962 ( .A(b[1613]), .B(n10865), .Z(c[1613]) );
  XOR U14963 ( .A(n10866), .B(n10867), .Z(n10863) );
  ANDN U14964 ( .B(n10868), .A(n10869), .Z(n10866) );
  XNOR U14965 ( .A(b[1612]), .B(n10867), .Z(n10868) );
  XNOR U14966 ( .A(b[1612]), .B(n10869), .Z(c[1612]) );
  XOR U14967 ( .A(n10870), .B(n10871), .Z(n10867) );
  ANDN U14968 ( .B(n10872), .A(n10873), .Z(n10870) );
  XNOR U14969 ( .A(b[1611]), .B(n10871), .Z(n10872) );
  XNOR U14970 ( .A(b[1611]), .B(n10873), .Z(c[1611]) );
  XOR U14971 ( .A(n10874), .B(n10875), .Z(n10871) );
  ANDN U14972 ( .B(n10876), .A(n10877), .Z(n10874) );
  XNOR U14973 ( .A(b[1610]), .B(n10875), .Z(n10876) );
  XNOR U14974 ( .A(b[1610]), .B(n10877), .Z(c[1610]) );
  XOR U14975 ( .A(n10878), .B(n10879), .Z(n10875) );
  ANDN U14976 ( .B(n10880), .A(n10881), .Z(n10878) );
  XNOR U14977 ( .A(b[1609]), .B(n10879), .Z(n10880) );
  XNOR U14978 ( .A(b[160]), .B(n10882), .Z(c[160]) );
  XNOR U14979 ( .A(b[1609]), .B(n10881), .Z(c[1609]) );
  XOR U14980 ( .A(n10883), .B(n10884), .Z(n10879) );
  ANDN U14981 ( .B(n10885), .A(n10886), .Z(n10883) );
  XNOR U14982 ( .A(b[1608]), .B(n10884), .Z(n10885) );
  XNOR U14983 ( .A(b[1608]), .B(n10886), .Z(c[1608]) );
  XOR U14984 ( .A(n10887), .B(n10888), .Z(n10884) );
  ANDN U14985 ( .B(n10889), .A(n10890), .Z(n10887) );
  XNOR U14986 ( .A(b[1607]), .B(n10888), .Z(n10889) );
  XNOR U14987 ( .A(b[1607]), .B(n10890), .Z(c[1607]) );
  XOR U14988 ( .A(n10891), .B(n10892), .Z(n10888) );
  ANDN U14989 ( .B(n10893), .A(n10894), .Z(n10891) );
  XNOR U14990 ( .A(b[1606]), .B(n10892), .Z(n10893) );
  XNOR U14991 ( .A(b[1606]), .B(n10894), .Z(c[1606]) );
  XOR U14992 ( .A(n10895), .B(n10896), .Z(n10892) );
  ANDN U14993 ( .B(n10897), .A(n10898), .Z(n10895) );
  XNOR U14994 ( .A(b[1605]), .B(n10896), .Z(n10897) );
  XNOR U14995 ( .A(b[1605]), .B(n10898), .Z(c[1605]) );
  XOR U14996 ( .A(n10899), .B(n10900), .Z(n10896) );
  ANDN U14997 ( .B(n10901), .A(n10902), .Z(n10899) );
  XNOR U14998 ( .A(b[1604]), .B(n10900), .Z(n10901) );
  XNOR U14999 ( .A(b[1604]), .B(n10902), .Z(c[1604]) );
  XOR U15000 ( .A(n10903), .B(n10904), .Z(n10900) );
  ANDN U15001 ( .B(n10905), .A(n10906), .Z(n10903) );
  XNOR U15002 ( .A(b[1603]), .B(n10904), .Z(n10905) );
  XNOR U15003 ( .A(b[1603]), .B(n10906), .Z(c[1603]) );
  XOR U15004 ( .A(n10907), .B(n10908), .Z(n10904) );
  ANDN U15005 ( .B(n10909), .A(n10910), .Z(n10907) );
  XNOR U15006 ( .A(b[1602]), .B(n10908), .Z(n10909) );
  XNOR U15007 ( .A(b[1602]), .B(n10910), .Z(c[1602]) );
  XOR U15008 ( .A(n10911), .B(n10912), .Z(n10908) );
  ANDN U15009 ( .B(n10913), .A(n10914), .Z(n10911) );
  XNOR U15010 ( .A(b[1601]), .B(n10912), .Z(n10913) );
  XNOR U15011 ( .A(b[1601]), .B(n10914), .Z(c[1601]) );
  XOR U15012 ( .A(n10915), .B(n10916), .Z(n10912) );
  ANDN U15013 ( .B(n10917), .A(n10918), .Z(n10915) );
  XNOR U15014 ( .A(b[1600]), .B(n10916), .Z(n10917) );
  XNOR U15015 ( .A(b[1600]), .B(n10918), .Z(c[1600]) );
  XOR U15016 ( .A(n10919), .B(n10920), .Z(n10916) );
  ANDN U15017 ( .B(n10921), .A(n10922), .Z(n10919) );
  XNOR U15018 ( .A(b[1599]), .B(n10920), .Z(n10921) );
  XNOR U15019 ( .A(b[15]), .B(n10923), .Z(c[15]) );
  XNOR U15020 ( .A(b[159]), .B(n10924), .Z(c[159]) );
  XNOR U15021 ( .A(b[1599]), .B(n10922), .Z(c[1599]) );
  XOR U15022 ( .A(n10925), .B(n10926), .Z(n10920) );
  ANDN U15023 ( .B(n10927), .A(n10928), .Z(n10925) );
  XNOR U15024 ( .A(b[1598]), .B(n10926), .Z(n10927) );
  XNOR U15025 ( .A(b[1598]), .B(n10928), .Z(c[1598]) );
  XOR U15026 ( .A(n10929), .B(n10930), .Z(n10926) );
  ANDN U15027 ( .B(n10931), .A(n10932), .Z(n10929) );
  XNOR U15028 ( .A(b[1597]), .B(n10930), .Z(n10931) );
  XNOR U15029 ( .A(b[1597]), .B(n10932), .Z(c[1597]) );
  XOR U15030 ( .A(n10933), .B(n10934), .Z(n10930) );
  ANDN U15031 ( .B(n10935), .A(n10936), .Z(n10933) );
  XNOR U15032 ( .A(b[1596]), .B(n10934), .Z(n10935) );
  XNOR U15033 ( .A(b[1596]), .B(n10936), .Z(c[1596]) );
  XOR U15034 ( .A(n10937), .B(n10938), .Z(n10934) );
  ANDN U15035 ( .B(n10939), .A(n10940), .Z(n10937) );
  XNOR U15036 ( .A(b[1595]), .B(n10938), .Z(n10939) );
  XNOR U15037 ( .A(b[1595]), .B(n10940), .Z(c[1595]) );
  XOR U15038 ( .A(n10941), .B(n10942), .Z(n10938) );
  ANDN U15039 ( .B(n10943), .A(n10944), .Z(n10941) );
  XNOR U15040 ( .A(b[1594]), .B(n10942), .Z(n10943) );
  XNOR U15041 ( .A(b[1594]), .B(n10944), .Z(c[1594]) );
  XOR U15042 ( .A(n10945), .B(n10946), .Z(n10942) );
  ANDN U15043 ( .B(n10947), .A(n10948), .Z(n10945) );
  XNOR U15044 ( .A(b[1593]), .B(n10946), .Z(n10947) );
  XNOR U15045 ( .A(b[1593]), .B(n10948), .Z(c[1593]) );
  XOR U15046 ( .A(n10949), .B(n10950), .Z(n10946) );
  ANDN U15047 ( .B(n10951), .A(n10952), .Z(n10949) );
  XNOR U15048 ( .A(b[1592]), .B(n10950), .Z(n10951) );
  XNOR U15049 ( .A(b[1592]), .B(n10952), .Z(c[1592]) );
  XOR U15050 ( .A(n10953), .B(n10954), .Z(n10950) );
  ANDN U15051 ( .B(n10955), .A(n10956), .Z(n10953) );
  XNOR U15052 ( .A(b[1591]), .B(n10954), .Z(n10955) );
  XNOR U15053 ( .A(b[1591]), .B(n10956), .Z(c[1591]) );
  XOR U15054 ( .A(n10957), .B(n10958), .Z(n10954) );
  ANDN U15055 ( .B(n10959), .A(n10960), .Z(n10957) );
  XNOR U15056 ( .A(b[1590]), .B(n10958), .Z(n10959) );
  XNOR U15057 ( .A(b[1590]), .B(n10960), .Z(c[1590]) );
  XOR U15058 ( .A(n10961), .B(n10962), .Z(n10958) );
  ANDN U15059 ( .B(n10963), .A(n10964), .Z(n10961) );
  XNOR U15060 ( .A(b[1589]), .B(n10962), .Z(n10963) );
  XNOR U15061 ( .A(b[158]), .B(n10965), .Z(c[158]) );
  XNOR U15062 ( .A(b[1589]), .B(n10964), .Z(c[1589]) );
  XOR U15063 ( .A(n10966), .B(n10967), .Z(n10962) );
  ANDN U15064 ( .B(n10968), .A(n10969), .Z(n10966) );
  XNOR U15065 ( .A(b[1588]), .B(n10967), .Z(n10968) );
  XNOR U15066 ( .A(b[1588]), .B(n10969), .Z(c[1588]) );
  XOR U15067 ( .A(n10970), .B(n10971), .Z(n10967) );
  ANDN U15068 ( .B(n10972), .A(n10973), .Z(n10970) );
  XNOR U15069 ( .A(b[1587]), .B(n10971), .Z(n10972) );
  XNOR U15070 ( .A(b[1587]), .B(n10973), .Z(c[1587]) );
  XOR U15071 ( .A(n10974), .B(n10975), .Z(n10971) );
  ANDN U15072 ( .B(n10976), .A(n10977), .Z(n10974) );
  XNOR U15073 ( .A(b[1586]), .B(n10975), .Z(n10976) );
  XNOR U15074 ( .A(b[1586]), .B(n10977), .Z(c[1586]) );
  XOR U15075 ( .A(n10978), .B(n10979), .Z(n10975) );
  ANDN U15076 ( .B(n10980), .A(n10981), .Z(n10978) );
  XNOR U15077 ( .A(b[1585]), .B(n10979), .Z(n10980) );
  XNOR U15078 ( .A(b[1585]), .B(n10981), .Z(c[1585]) );
  XOR U15079 ( .A(n10982), .B(n10983), .Z(n10979) );
  ANDN U15080 ( .B(n10984), .A(n10985), .Z(n10982) );
  XNOR U15081 ( .A(b[1584]), .B(n10983), .Z(n10984) );
  XNOR U15082 ( .A(b[1584]), .B(n10985), .Z(c[1584]) );
  XOR U15083 ( .A(n10986), .B(n10987), .Z(n10983) );
  ANDN U15084 ( .B(n10988), .A(n10989), .Z(n10986) );
  XNOR U15085 ( .A(b[1583]), .B(n10987), .Z(n10988) );
  XNOR U15086 ( .A(b[1583]), .B(n10989), .Z(c[1583]) );
  XOR U15087 ( .A(n10990), .B(n10991), .Z(n10987) );
  ANDN U15088 ( .B(n10992), .A(n10993), .Z(n10990) );
  XNOR U15089 ( .A(b[1582]), .B(n10991), .Z(n10992) );
  XNOR U15090 ( .A(b[1582]), .B(n10993), .Z(c[1582]) );
  XOR U15091 ( .A(n10994), .B(n10995), .Z(n10991) );
  ANDN U15092 ( .B(n10996), .A(n10997), .Z(n10994) );
  XNOR U15093 ( .A(b[1581]), .B(n10995), .Z(n10996) );
  XNOR U15094 ( .A(b[1581]), .B(n10997), .Z(c[1581]) );
  XOR U15095 ( .A(n10998), .B(n10999), .Z(n10995) );
  ANDN U15096 ( .B(n11000), .A(n11001), .Z(n10998) );
  XNOR U15097 ( .A(b[1580]), .B(n10999), .Z(n11000) );
  XNOR U15098 ( .A(b[1580]), .B(n11001), .Z(c[1580]) );
  XOR U15099 ( .A(n11002), .B(n11003), .Z(n10999) );
  ANDN U15100 ( .B(n11004), .A(n11005), .Z(n11002) );
  XNOR U15101 ( .A(b[1579]), .B(n11003), .Z(n11004) );
  XNOR U15102 ( .A(b[157]), .B(n11006), .Z(c[157]) );
  XNOR U15103 ( .A(b[1579]), .B(n11005), .Z(c[1579]) );
  XOR U15104 ( .A(n11007), .B(n11008), .Z(n11003) );
  ANDN U15105 ( .B(n11009), .A(n11010), .Z(n11007) );
  XNOR U15106 ( .A(b[1578]), .B(n11008), .Z(n11009) );
  XNOR U15107 ( .A(b[1578]), .B(n11010), .Z(c[1578]) );
  XOR U15108 ( .A(n11011), .B(n11012), .Z(n11008) );
  ANDN U15109 ( .B(n11013), .A(n11014), .Z(n11011) );
  XNOR U15110 ( .A(b[1577]), .B(n11012), .Z(n11013) );
  XNOR U15111 ( .A(b[1577]), .B(n11014), .Z(c[1577]) );
  XOR U15112 ( .A(n11015), .B(n11016), .Z(n11012) );
  ANDN U15113 ( .B(n11017), .A(n11018), .Z(n11015) );
  XNOR U15114 ( .A(b[1576]), .B(n11016), .Z(n11017) );
  XNOR U15115 ( .A(b[1576]), .B(n11018), .Z(c[1576]) );
  XOR U15116 ( .A(n11019), .B(n11020), .Z(n11016) );
  ANDN U15117 ( .B(n11021), .A(n11022), .Z(n11019) );
  XNOR U15118 ( .A(b[1575]), .B(n11020), .Z(n11021) );
  XNOR U15119 ( .A(b[1575]), .B(n11022), .Z(c[1575]) );
  XOR U15120 ( .A(n11023), .B(n11024), .Z(n11020) );
  ANDN U15121 ( .B(n11025), .A(n11026), .Z(n11023) );
  XNOR U15122 ( .A(b[1574]), .B(n11024), .Z(n11025) );
  XNOR U15123 ( .A(b[1574]), .B(n11026), .Z(c[1574]) );
  XOR U15124 ( .A(n11027), .B(n11028), .Z(n11024) );
  ANDN U15125 ( .B(n11029), .A(n11030), .Z(n11027) );
  XNOR U15126 ( .A(b[1573]), .B(n11028), .Z(n11029) );
  XNOR U15127 ( .A(b[1573]), .B(n11030), .Z(c[1573]) );
  XOR U15128 ( .A(n11031), .B(n11032), .Z(n11028) );
  ANDN U15129 ( .B(n11033), .A(n11034), .Z(n11031) );
  XNOR U15130 ( .A(b[1572]), .B(n11032), .Z(n11033) );
  XNOR U15131 ( .A(b[1572]), .B(n11034), .Z(c[1572]) );
  XOR U15132 ( .A(n11035), .B(n11036), .Z(n11032) );
  ANDN U15133 ( .B(n11037), .A(n11038), .Z(n11035) );
  XNOR U15134 ( .A(b[1571]), .B(n11036), .Z(n11037) );
  XNOR U15135 ( .A(b[1571]), .B(n11038), .Z(c[1571]) );
  XOR U15136 ( .A(n11039), .B(n11040), .Z(n11036) );
  ANDN U15137 ( .B(n11041), .A(n11042), .Z(n11039) );
  XNOR U15138 ( .A(b[1570]), .B(n11040), .Z(n11041) );
  XNOR U15139 ( .A(b[1570]), .B(n11042), .Z(c[1570]) );
  XOR U15140 ( .A(n11043), .B(n11044), .Z(n11040) );
  ANDN U15141 ( .B(n11045), .A(n11046), .Z(n11043) );
  XNOR U15142 ( .A(b[1569]), .B(n11044), .Z(n11045) );
  XNOR U15143 ( .A(b[156]), .B(n11047), .Z(c[156]) );
  XNOR U15144 ( .A(b[1569]), .B(n11046), .Z(c[1569]) );
  XOR U15145 ( .A(n11048), .B(n11049), .Z(n11044) );
  ANDN U15146 ( .B(n11050), .A(n11051), .Z(n11048) );
  XNOR U15147 ( .A(b[1568]), .B(n11049), .Z(n11050) );
  XNOR U15148 ( .A(b[1568]), .B(n11051), .Z(c[1568]) );
  XOR U15149 ( .A(n11052), .B(n11053), .Z(n11049) );
  ANDN U15150 ( .B(n11054), .A(n11055), .Z(n11052) );
  XNOR U15151 ( .A(b[1567]), .B(n11053), .Z(n11054) );
  XNOR U15152 ( .A(b[1567]), .B(n11055), .Z(c[1567]) );
  XOR U15153 ( .A(n11056), .B(n11057), .Z(n11053) );
  ANDN U15154 ( .B(n11058), .A(n11059), .Z(n11056) );
  XNOR U15155 ( .A(b[1566]), .B(n11057), .Z(n11058) );
  XNOR U15156 ( .A(b[1566]), .B(n11059), .Z(c[1566]) );
  XOR U15157 ( .A(n11060), .B(n11061), .Z(n11057) );
  ANDN U15158 ( .B(n11062), .A(n11063), .Z(n11060) );
  XNOR U15159 ( .A(b[1565]), .B(n11061), .Z(n11062) );
  XNOR U15160 ( .A(b[1565]), .B(n11063), .Z(c[1565]) );
  XOR U15161 ( .A(n11064), .B(n11065), .Z(n11061) );
  ANDN U15162 ( .B(n11066), .A(n11067), .Z(n11064) );
  XNOR U15163 ( .A(b[1564]), .B(n11065), .Z(n11066) );
  XNOR U15164 ( .A(b[1564]), .B(n11067), .Z(c[1564]) );
  XOR U15165 ( .A(n11068), .B(n11069), .Z(n11065) );
  ANDN U15166 ( .B(n11070), .A(n11071), .Z(n11068) );
  XNOR U15167 ( .A(b[1563]), .B(n11069), .Z(n11070) );
  XNOR U15168 ( .A(b[1563]), .B(n11071), .Z(c[1563]) );
  XOR U15169 ( .A(n11072), .B(n11073), .Z(n11069) );
  ANDN U15170 ( .B(n11074), .A(n11075), .Z(n11072) );
  XNOR U15171 ( .A(b[1562]), .B(n11073), .Z(n11074) );
  XNOR U15172 ( .A(b[1562]), .B(n11075), .Z(c[1562]) );
  XOR U15173 ( .A(n11076), .B(n11077), .Z(n11073) );
  ANDN U15174 ( .B(n11078), .A(n11079), .Z(n11076) );
  XNOR U15175 ( .A(b[1561]), .B(n11077), .Z(n11078) );
  XNOR U15176 ( .A(b[1561]), .B(n11079), .Z(c[1561]) );
  XOR U15177 ( .A(n11080), .B(n11081), .Z(n11077) );
  ANDN U15178 ( .B(n11082), .A(n11083), .Z(n11080) );
  XNOR U15179 ( .A(b[1560]), .B(n11081), .Z(n11082) );
  XNOR U15180 ( .A(b[1560]), .B(n11083), .Z(c[1560]) );
  XOR U15181 ( .A(n11084), .B(n11085), .Z(n11081) );
  ANDN U15182 ( .B(n11086), .A(n11087), .Z(n11084) );
  XNOR U15183 ( .A(b[1559]), .B(n11085), .Z(n11086) );
  XNOR U15184 ( .A(b[155]), .B(n11088), .Z(c[155]) );
  XNOR U15185 ( .A(b[1559]), .B(n11087), .Z(c[1559]) );
  XOR U15186 ( .A(n11089), .B(n11090), .Z(n11085) );
  ANDN U15187 ( .B(n11091), .A(n11092), .Z(n11089) );
  XNOR U15188 ( .A(b[1558]), .B(n11090), .Z(n11091) );
  XNOR U15189 ( .A(b[1558]), .B(n11092), .Z(c[1558]) );
  XOR U15190 ( .A(n11093), .B(n11094), .Z(n11090) );
  ANDN U15191 ( .B(n11095), .A(n11096), .Z(n11093) );
  XNOR U15192 ( .A(b[1557]), .B(n11094), .Z(n11095) );
  XNOR U15193 ( .A(b[1557]), .B(n11096), .Z(c[1557]) );
  XOR U15194 ( .A(n11097), .B(n11098), .Z(n11094) );
  ANDN U15195 ( .B(n11099), .A(n11100), .Z(n11097) );
  XNOR U15196 ( .A(b[1556]), .B(n11098), .Z(n11099) );
  XNOR U15197 ( .A(b[1556]), .B(n11100), .Z(c[1556]) );
  XOR U15198 ( .A(n11101), .B(n11102), .Z(n11098) );
  ANDN U15199 ( .B(n11103), .A(n11104), .Z(n11101) );
  XNOR U15200 ( .A(b[1555]), .B(n11102), .Z(n11103) );
  XNOR U15201 ( .A(b[1555]), .B(n11104), .Z(c[1555]) );
  XOR U15202 ( .A(n11105), .B(n11106), .Z(n11102) );
  ANDN U15203 ( .B(n11107), .A(n11108), .Z(n11105) );
  XNOR U15204 ( .A(b[1554]), .B(n11106), .Z(n11107) );
  XNOR U15205 ( .A(b[1554]), .B(n11108), .Z(c[1554]) );
  XOR U15206 ( .A(n11109), .B(n11110), .Z(n11106) );
  ANDN U15207 ( .B(n11111), .A(n11112), .Z(n11109) );
  XNOR U15208 ( .A(b[1553]), .B(n11110), .Z(n11111) );
  XNOR U15209 ( .A(b[1553]), .B(n11112), .Z(c[1553]) );
  XOR U15210 ( .A(n11113), .B(n11114), .Z(n11110) );
  ANDN U15211 ( .B(n11115), .A(n11116), .Z(n11113) );
  XNOR U15212 ( .A(b[1552]), .B(n11114), .Z(n11115) );
  XNOR U15213 ( .A(b[1552]), .B(n11116), .Z(c[1552]) );
  XOR U15214 ( .A(n11117), .B(n11118), .Z(n11114) );
  ANDN U15215 ( .B(n11119), .A(n11120), .Z(n11117) );
  XNOR U15216 ( .A(b[1551]), .B(n11118), .Z(n11119) );
  XNOR U15217 ( .A(b[1551]), .B(n11120), .Z(c[1551]) );
  XOR U15218 ( .A(n11121), .B(n11122), .Z(n11118) );
  ANDN U15219 ( .B(n11123), .A(n11124), .Z(n11121) );
  XNOR U15220 ( .A(b[1550]), .B(n11122), .Z(n11123) );
  XNOR U15221 ( .A(b[1550]), .B(n11124), .Z(c[1550]) );
  XOR U15222 ( .A(n11125), .B(n11126), .Z(n11122) );
  ANDN U15223 ( .B(n11127), .A(n11128), .Z(n11125) );
  XNOR U15224 ( .A(b[1549]), .B(n11126), .Z(n11127) );
  XNOR U15225 ( .A(b[154]), .B(n11129), .Z(c[154]) );
  XNOR U15226 ( .A(b[1549]), .B(n11128), .Z(c[1549]) );
  XOR U15227 ( .A(n11130), .B(n11131), .Z(n11126) );
  ANDN U15228 ( .B(n11132), .A(n11133), .Z(n11130) );
  XNOR U15229 ( .A(b[1548]), .B(n11131), .Z(n11132) );
  XNOR U15230 ( .A(b[1548]), .B(n11133), .Z(c[1548]) );
  XOR U15231 ( .A(n11134), .B(n11135), .Z(n11131) );
  ANDN U15232 ( .B(n11136), .A(n11137), .Z(n11134) );
  XNOR U15233 ( .A(b[1547]), .B(n11135), .Z(n11136) );
  XNOR U15234 ( .A(b[1547]), .B(n11137), .Z(c[1547]) );
  XOR U15235 ( .A(n11138), .B(n11139), .Z(n11135) );
  ANDN U15236 ( .B(n11140), .A(n11141), .Z(n11138) );
  XNOR U15237 ( .A(b[1546]), .B(n11139), .Z(n11140) );
  XNOR U15238 ( .A(b[1546]), .B(n11141), .Z(c[1546]) );
  XOR U15239 ( .A(n11142), .B(n11143), .Z(n11139) );
  ANDN U15240 ( .B(n11144), .A(n11145), .Z(n11142) );
  XNOR U15241 ( .A(b[1545]), .B(n11143), .Z(n11144) );
  XNOR U15242 ( .A(b[1545]), .B(n11145), .Z(c[1545]) );
  XOR U15243 ( .A(n11146), .B(n11147), .Z(n11143) );
  ANDN U15244 ( .B(n11148), .A(n11149), .Z(n11146) );
  XNOR U15245 ( .A(b[1544]), .B(n11147), .Z(n11148) );
  XNOR U15246 ( .A(b[1544]), .B(n11149), .Z(c[1544]) );
  XOR U15247 ( .A(n11150), .B(n11151), .Z(n11147) );
  ANDN U15248 ( .B(n11152), .A(n11153), .Z(n11150) );
  XNOR U15249 ( .A(b[1543]), .B(n11151), .Z(n11152) );
  XNOR U15250 ( .A(b[1543]), .B(n11153), .Z(c[1543]) );
  XOR U15251 ( .A(n11154), .B(n11155), .Z(n11151) );
  ANDN U15252 ( .B(n11156), .A(n11157), .Z(n11154) );
  XNOR U15253 ( .A(b[1542]), .B(n11155), .Z(n11156) );
  XNOR U15254 ( .A(b[1542]), .B(n11157), .Z(c[1542]) );
  XOR U15255 ( .A(n11158), .B(n11159), .Z(n11155) );
  ANDN U15256 ( .B(n11160), .A(n11161), .Z(n11158) );
  XNOR U15257 ( .A(b[1541]), .B(n11159), .Z(n11160) );
  XNOR U15258 ( .A(b[1541]), .B(n11161), .Z(c[1541]) );
  XOR U15259 ( .A(n11162), .B(n11163), .Z(n11159) );
  ANDN U15260 ( .B(n11164), .A(n11165), .Z(n11162) );
  XNOR U15261 ( .A(b[1540]), .B(n11163), .Z(n11164) );
  XNOR U15262 ( .A(b[1540]), .B(n11165), .Z(c[1540]) );
  XOR U15263 ( .A(n11166), .B(n11167), .Z(n11163) );
  ANDN U15264 ( .B(n11168), .A(n11169), .Z(n11166) );
  XNOR U15265 ( .A(b[1539]), .B(n11167), .Z(n11168) );
  XNOR U15266 ( .A(b[153]), .B(n11170), .Z(c[153]) );
  XNOR U15267 ( .A(b[1539]), .B(n11169), .Z(c[1539]) );
  XOR U15268 ( .A(n11171), .B(n11172), .Z(n11167) );
  ANDN U15269 ( .B(n11173), .A(n11174), .Z(n11171) );
  XNOR U15270 ( .A(b[1538]), .B(n11172), .Z(n11173) );
  XNOR U15271 ( .A(b[1538]), .B(n11174), .Z(c[1538]) );
  XOR U15272 ( .A(n11175), .B(n11176), .Z(n11172) );
  ANDN U15273 ( .B(n11177), .A(n11178), .Z(n11175) );
  XNOR U15274 ( .A(b[1537]), .B(n11176), .Z(n11177) );
  XNOR U15275 ( .A(b[1537]), .B(n11178), .Z(c[1537]) );
  XOR U15276 ( .A(n11179), .B(n11180), .Z(n11176) );
  ANDN U15277 ( .B(n11181), .A(n11182), .Z(n11179) );
  XNOR U15278 ( .A(b[1536]), .B(n11180), .Z(n11181) );
  XNOR U15279 ( .A(b[1536]), .B(n11182), .Z(c[1536]) );
  XOR U15280 ( .A(n11183), .B(n11184), .Z(n11180) );
  ANDN U15281 ( .B(n11185), .A(n11186), .Z(n11183) );
  XNOR U15282 ( .A(b[1535]), .B(n11184), .Z(n11185) );
  XNOR U15283 ( .A(b[1535]), .B(n11186), .Z(c[1535]) );
  XOR U15284 ( .A(n11187), .B(n11188), .Z(n11184) );
  ANDN U15285 ( .B(n11189), .A(n11190), .Z(n11187) );
  XNOR U15286 ( .A(b[1534]), .B(n11188), .Z(n11189) );
  XNOR U15287 ( .A(b[1534]), .B(n11190), .Z(c[1534]) );
  XOR U15288 ( .A(n11191), .B(n11192), .Z(n11188) );
  ANDN U15289 ( .B(n11193), .A(n11194), .Z(n11191) );
  XNOR U15290 ( .A(b[1533]), .B(n11192), .Z(n11193) );
  XNOR U15291 ( .A(b[1533]), .B(n11194), .Z(c[1533]) );
  XOR U15292 ( .A(n11195), .B(n11196), .Z(n11192) );
  ANDN U15293 ( .B(n11197), .A(n11198), .Z(n11195) );
  XNOR U15294 ( .A(b[1532]), .B(n11196), .Z(n11197) );
  XNOR U15295 ( .A(b[1532]), .B(n11198), .Z(c[1532]) );
  XOR U15296 ( .A(n11199), .B(n11200), .Z(n11196) );
  ANDN U15297 ( .B(n11201), .A(n11202), .Z(n11199) );
  XNOR U15298 ( .A(b[1531]), .B(n11200), .Z(n11201) );
  XNOR U15299 ( .A(b[1531]), .B(n11202), .Z(c[1531]) );
  XOR U15300 ( .A(n11203), .B(n11204), .Z(n11200) );
  ANDN U15301 ( .B(n11205), .A(n11206), .Z(n11203) );
  XNOR U15302 ( .A(b[1530]), .B(n11204), .Z(n11205) );
  XNOR U15303 ( .A(b[1530]), .B(n11206), .Z(c[1530]) );
  XOR U15304 ( .A(n11207), .B(n11208), .Z(n11204) );
  ANDN U15305 ( .B(n11209), .A(n11210), .Z(n11207) );
  XNOR U15306 ( .A(b[1529]), .B(n11208), .Z(n11209) );
  XNOR U15307 ( .A(b[152]), .B(n11211), .Z(c[152]) );
  XNOR U15308 ( .A(b[1529]), .B(n11210), .Z(c[1529]) );
  XOR U15309 ( .A(n11212), .B(n11213), .Z(n11208) );
  ANDN U15310 ( .B(n11214), .A(n11215), .Z(n11212) );
  XNOR U15311 ( .A(b[1528]), .B(n11213), .Z(n11214) );
  XNOR U15312 ( .A(b[1528]), .B(n11215), .Z(c[1528]) );
  XOR U15313 ( .A(n11216), .B(n11217), .Z(n11213) );
  ANDN U15314 ( .B(n11218), .A(n11219), .Z(n11216) );
  XNOR U15315 ( .A(b[1527]), .B(n11217), .Z(n11218) );
  XNOR U15316 ( .A(b[1527]), .B(n11219), .Z(c[1527]) );
  XOR U15317 ( .A(n11220), .B(n11221), .Z(n11217) );
  ANDN U15318 ( .B(n11222), .A(n11223), .Z(n11220) );
  XNOR U15319 ( .A(b[1526]), .B(n11221), .Z(n11222) );
  XNOR U15320 ( .A(b[1526]), .B(n11223), .Z(c[1526]) );
  XOR U15321 ( .A(n11224), .B(n11225), .Z(n11221) );
  ANDN U15322 ( .B(n11226), .A(n11227), .Z(n11224) );
  XNOR U15323 ( .A(b[1525]), .B(n11225), .Z(n11226) );
  XNOR U15324 ( .A(b[1525]), .B(n11227), .Z(c[1525]) );
  XOR U15325 ( .A(n11228), .B(n11229), .Z(n11225) );
  ANDN U15326 ( .B(n11230), .A(n11231), .Z(n11228) );
  XNOR U15327 ( .A(b[1524]), .B(n11229), .Z(n11230) );
  XNOR U15328 ( .A(b[1524]), .B(n11231), .Z(c[1524]) );
  XOR U15329 ( .A(n11232), .B(n11233), .Z(n11229) );
  ANDN U15330 ( .B(n11234), .A(n11235), .Z(n11232) );
  XNOR U15331 ( .A(b[1523]), .B(n11233), .Z(n11234) );
  XNOR U15332 ( .A(b[1523]), .B(n11235), .Z(c[1523]) );
  XOR U15333 ( .A(n11236), .B(n11237), .Z(n11233) );
  ANDN U15334 ( .B(n11238), .A(n11239), .Z(n11236) );
  XNOR U15335 ( .A(b[1522]), .B(n11237), .Z(n11238) );
  XNOR U15336 ( .A(b[1522]), .B(n11239), .Z(c[1522]) );
  XOR U15337 ( .A(n11240), .B(n11241), .Z(n11237) );
  ANDN U15338 ( .B(n11242), .A(n11243), .Z(n11240) );
  XNOR U15339 ( .A(b[1521]), .B(n11241), .Z(n11242) );
  XNOR U15340 ( .A(b[1521]), .B(n11243), .Z(c[1521]) );
  XOR U15341 ( .A(n11244), .B(n11245), .Z(n11241) );
  ANDN U15342 ( .B(n11246), .A(n11247), .Z(n11244) );
  XNOR U15343 ( .A(b[1520]), .B(n11245), .Z(n11246) );
  XNOR U15344 ( .A(b[1520]), .B(n11247), .Z(c[1520]) );
  XOR U15345 ( .A(n11248), .B(n11249), .Z(n11245) );
  ANDN U15346 ( .B(n11250), .A(n11251), .Z(n11248) );
  XNOR U15347 ( .A(b[1519]), .B(n11249), .Z(n11250) );
  XNOR U15348 ( .A(b[151]), .B(n11252), .Z(c[151]) );
  XNOR U15349 ( .A(b[1519]), .B(n11251), .Z(c[1519]) );
  XOR U15350 ( .A(n11253), .B(n11254), .Z(n11249) );
  ANDN U15351 ( .B(n11255), .A(n11256), .Z(n11253) );
  XNOR U15352 ( .A(b[1518]), .B(n11254), .Z(n11255) );
  XNOR U15353 ( .A(b[1518]), .B(n11256), .Z(c[1518]) );
  XOR U15354 ( .A(n11257), .B(n11258), .Z(n11254) );
  ANDN U15355 ( .B(n11259), .A(n11260), .Z(n11257) );
  XNOR U15356 ( .A(b[1517]), .B(n11258), .Z(n11259) );
  XNOR U15357 ( .A(b[1517]), .B(n11260), .Z(c[1517]) );
  XOR U15358 ( .A(n11261), .B(n11262), .Z(n11258) );
  ANDN U15359 ( .B(n11263), .A(n11264), .Z(n11261) );
  XNOR U15360 ( .A(b[1516]), .B(n11262), .Z(n11263) );
  XNOR U15361 ( .A(b[1516]), .B(n11264), .Z(c[1516]) );
  XOR U15362 ( .A(n11265), .B(n11266), .Z(n11262) );
  ANDN U15363 ( .B(n11267), .A(n11268), .Z(n11265) );
  XNOR U15364 ( .A(b[1515]), .B(n11266), .Z(n11267) );
  XNOR U15365 ( .A(b[1515]), .B(n11268), .Z(c[1515]) );
  XOR U15366 ( .A(n11269), .B(n11270), .Z(n11266) );
  ANDN U15367 ( .B(n11271), .A(n11272), .Z(n11269) );
  XNOR U15368 ( .A(b[1514]), .B(n11270), .Z(n11271) );
  XNOR U15369 ( .A(b[1514]), .B(n11272), .Z(c[1514]) );
  XOR U15370 ( .A(n11273), .B(n11274), .Z(n11270) );
  ANDN U15371 ( .B(n11275), .A(n11276), .Z(n11273) );
  XNOR U15372 ( .A(b[1513]), .B(n11274), .Z(n11275) );
  XNOR U15373 ( .A(b[1513]), .B(n11276), .Z(c[1513]) );
  XOR U15374 ( .A(n11277), .B(n11278), .Z(n11274) );
  ANDN U15375 ( .B(n11279), .A(n11280), .Z(n11277) );
  XNOR U15376 ( .A(b[1512]), .B(n11278), .Z(n11279) );
  XNOR U15377 ( .A(b[1512]), .B(n11280), .Z(c[1512]) );
  XOR U15378 ( .A(n11281), .B(n11282), .Z(n11278) );
  ANDN U15379 ( .B(n11283), .A(n11284), .Z(n11281) );
  XNOR U15380 ( .A(b[1511]), .B(n11282), .Z(n11283) );
  XNOR U15381 ( .A(b[1511]), .B(n11284), .Z(c[1511]) );
  XOR U15382 ( .A(n11285), .B(n11286), .Z(n11282) );
  ANDN U15383 ( .B(n11287), .A(n11288), .Z(n11285) );
  XNOR U15384 ( .A(b[1510]), .B(n11286), .Z(n11287) );
  XNOR U15385 ( .A(b[1510]), .B(n11288), .Z(c[1510]) );
  XOR U15386 ( .A(n11289), .B(n11290), .Z(n11286) );
  ANDN U15387 ( .B(n11291), .A(n11292), .Z(n11289) );
  XNOR U15388 ( .A(b[1509]), .B(n11290), .Z(n11291) );
  XNOR U15389 ( .A(b[150]), .B(n11293), .Z(c[150]) );
  XNOR U15390 ( .A(b[1509]), .B(n11292), .Z(c[1509]) );
  XOR U15391 ( .A(n11294), .B(n11295), .Z(n11290) );
  ANDN U15392 ( .B(n11296), .A(n11297), .Z(n11294) );
  XNOR U15393 ( .A(b[1508]), .B(n11295), .Z(n11296) );
  XNOR U15394 ( .A(b[1508]), .B(n11297), .Z(c[1508]) );
  XOR U15395 ( .A(n11298), .B(n11299), .Z(n11295) );
  ANDN U15396 ( .B(n11300), .A(n11301), .Z(n11298) );
  XNOR U15397 ( .A(b[1507]), .B(n11299), .Z(n11300) );
  XNOR U15398 ( .A(b[1507]), .B(n11301), .Z(c[1507]) );
  XOR U15399 ( .A(n11302), .B(n11303), .Z(n11299) );
  ANDN U15400 ( .B(n11304), .A(n11305), .Z(n11302) );
  XNOR U15401 ( .A(b[1506]), .B(n11303), .Z(n11304) );
  XNOR U15402 ( .A(b[1506]), .B(n11305), .Z(c[1506]) );
  XOR U15403 ( .A(n11306), .B(n11307), .Z(n11303) );
  ANDN U15404 ( .B(n11308), .A(n11309), .Z(n11306) );
  XNOR U15405 ( .A(b[1505]), .B(n11307), .Z(n11308) );
  XNOR U15406 ( .A(b[1505]), .B(n11309), .Z(c[1505]) );
  XOR U15407 ( .A(n11310), .B(n11311), .Z(n11307) );
  ANDN U15408 ( .B(n11312), .A(n11313), .Z(n11310) );
  XNOR U15409 ( .A(b[1504]), .B(n11311), .Z(n11312) );
  XNOR U15410 ( .A(b[1504]), .B(n11313), .Z(c[1504]) );
  XOR U15411 ( .A(n11314), .B(n11315), .Z(n11311) );
  ANDN U15412 ( .B(n11316), .A(n11317), .Z(n11314) );
  XNOR U15413 ( .A(b[1503]), .B(n11315), .Z(n11316) );
  XNOR U15414 ( .A(b[1503]), .B(n11317), .Z(c[1503]) );
  XOR U15415 ( .A(n11318), .B(n11319), .Z(n11315) );
  ANDN U15416 ( .B(n11320), .A(n11321), .Z(n11318) );
  XNOR U15417 ( .A(b[1502]), .B(n11319), .Z(n11320) );
  XNOR U15418 ( .A(b[1502]), .B(n11321), .Z(c[1502]) );
  XOR U15419 ( .A(n11322), .B(n11323), .Z(n11319) );
  ANDN U15420 ( .B(n11324), .A(n11325), .Z(n11322) );
  XNOR U15421 ( .A(b[1501]), .B(n11323), .Z(n11324) );
  XNOR U15422 ( .A(b[1501]), .B(n11325), .Z(c[1501]) );
  XOR U15423 ( .A(n11326), .B(n11327), .Z(n11323) );
  ANDN U15424 ( .B(n11328), .A(n11329), .Z(n11326) );
  XNOR U15425 ( .A(b[1500]), .B(n11327), .Z(n11328) );
  XNOR U15426 ( .A(b[1500]), .B(n11329), .Z(c[1500]) );
  XOR U15427 ( .A(n11330), .B(n11331), .Z(n11327) );
  ANDN U15428 ( .B(n11332), .A(n11333), .Z(n11330) );
  XNOR U15429 ( .A(b[1499]), .B(n11331), .Z(n11332) );
  XNOR U15430 ( .A(b[14]), .B(n11334), .Z(c[14]) );
  XNOR U15431 ( .A(b[149]), .B(n11335), .Z(c[149]) );
  XNOR U15432 ( .A(b[1499]), .B(n11333), .Z(c[1499]) );
  XOR U15433 ( .A(n11336), .B(n11337), .Z(n11331) );
  ANDN U15434 ( .B(n11338), .A(n11339), .Z(n11336) );
  XNOR U15435 ( .A(b[1498]), .B(n11337), .Z(n11338) );
  XNOR U15436 ( .A(b[1498]), .B(n11339), .Z(c[1498]) );
  XOR U15437 ( .A(n11340), .B(n11341), .Z(n11337) );
  ANDN U15438 ( .B(n11342), .A(n11343), .Z(n11340) );
  XNOR U15439 ( .A(b[1497]), .B(n11341), .Z(n11342) );
  XNOR U15440 ( .A(b[1497]), .B(n11343), .Z(c[1497]) );
  XOR U15441 ( .A(n11344), .B(n11345), .Z(n11341) );
  ANDN U15442 ( .B(n11346), .A(n11347), .Z(n11344) );
  XNOR U15443 ( .A(b[1496]), .B(n11345), .Z(n11346) );
  XNOR U15444 ( .A(b[1496]), .B(n11347), .Z(c[1496]) );
  XOR U15445 ( .A(n11348), .B(n11349), .Z(n11345) );
  ANDN U15446 ( .B(n11350), .A(n11351), .Z(n11348) );
  XNOR U15447 ( .A(b[1495]), .B(n11349), .Z(n11350) );
  XNOR U15448 ( .A(b[1495]), .B(n11351), .Z(c[1495]) );
  XOR U15449 ( .A(n11352), .B(n11353), .Z(n11349) );
  ANDN U15450 ( .B(n11354), .A(n11355), .Z(n11352) );
  XNOR U15451 ( .A(b[1494]), .B(n11353), .Z(n11354) );
  XNOR U15452 ( .A(b[1494]), .B(n11355), .Z(c[1494]) );
  XOR U15453 ( .A(n11356), .B(n11357), .Z(n11353) );
  ANDN U15454 ( .B(n11358), .A(n11359), .Z(n11356) );
  XNOR U15455 ( .A(b[1493]), .B(n11357), .Z(n11358) );
  XNOR U15456 ( .A(b[1493]), .B(n11359), .Z(c[1493]) );
  XOR U15457 ( .A(n11360), .B(n11361), .Z(n11357) );
  ANDN U15458 ( .B(n11362), .A(n11363), .Z(n11360) );
  XNOR U15459 ( .A(b[1492]), .B(n11361), .Z(n11362) );
  XNOR U15460 ( .A(b[1492]), .B(n11363), .Z(c[1492]) );
  XOR U15461 ( .A(n11364), .B(n11365), .Z(n11361) );
  ANDN U15462 ( .B(n11366), .A(n11367), .Z(n11364) );
  XNOR U15463 ( .A(b[1491]), .B(n11365), .Z(n11366) );
  XNOR U15464 ( .A(b[1491]), .B(n11367), .Z(c[1491]) );
  XOR U15465 ( .A(n11368), .B(n11369), .Z(n11365) );
  ANDN U15466 ( .B(n11370), .A(n11371), .Z(n11368) );
  XNOR U15467 ( .A(b[1490]), .B(n11369), .Z(n11370) );
  XNOR U15468 ( .A(b[1490]), .B(n11371), .Z(c[1490]) );
  XOR U15469 ( .A(n11372), .B(n11373), .Z(n11369) );
  ANDN U15470 ( .B(n11374), .A(n11375), .Z(n11372) );
  XNOR U15471 ( .A(b[1489]), .B(n11373), .Z(n11374) );
  XNOR U15472 ( .A(b[148]), .B(n11376), .Z(c[148]) );
  XNOR U15473 ( .A(b[1489]), .B(n11375), .Z(c[1489]) );
  XOR U15474 ( .A(n11377), .B(n11378), .Z(n11373) );
  ANDN U15475 ( .B(n11379), .A(n11380), .Z(n11377) );
  XNOR U15476 ( .A(b[1488]), .B(n11378), .Z(n11379) );
  XNOR U15477 ( .A(b[1488]), .B(n11380), .Z(c[1488]) );
  XOR U15478 ( .A(n11381), .B(n11382), .Z(n11378) );
  ANDN U15479 ( .B(n11383), .A(n11384), .Z(n11381) );
  XNOR U15480 ( .A(b[1487]), .B(n11382), .Z(n11383) );
  XNOR U15481 ( .A(b[1487]), .B(n11384), .Z(c[1487]) );
  XOR U15482 ( .A(n11385), .B(n11386), .Z(n11382) );
  ANDN U15483 ( .B(n11387), .A(n11388), .Z(n11385) );
  XNOR U15484 ( .A(b[1486]), .B(n11386), .Z(n11387) );
  XNOR U15485 ( .A(b[1486]), .B(n11388), .Z(c[1486]) );
  XOR U15486 ( .A(n11389), .B(n11390), .Z(n11386) );
  ANDN U15487 ( .B(n11391), .A(n11392), .Z(n11389) );
  XNOR U15488 ( .A(b[1485]), .B(n11390), .Z(n11391) );
  XNOR U15489 ( .A(b[1485]), .B(n11392), .Z(c[1485]) );
  XOR U15490 ( .A(n11393), .B(n11394), .Z(n11390) );
  ANDN U15491 ( .B(n11395), .A(n11396), .Z(n11393) );
  XNOR U15492 ( .A(b[1484]), .B(n11394), .Z(n11395) );
  XNOR U15493 ( .A(b[1484]), .B(n11396), .Z(c[1484]) );
  XOR U15494 ( .A(n11397), .B(n11398), .Z(n11394) );
  ANDN U15495 ( .B(n11399), .A(n11400), .Z(n11397) );
  XNOR U15496 ( .A(b[1483]), .B(n11398), .Z(n11399) );
  XNOR U15497 ( .A(b[1483]), .B(n11400), .Z(c[1483]) );
  XOR U15498 ( .A(n11401), .B(n11402), .Z(n11398) );
  ANDN U15499 ( .B(n11403), .A(n11404), .Z(n11401) );
  XNOR U15500 ( .A(b[1482]), .B(n11402), .Z(n11403) );
  XNOR U15501 ( .A(b[1482]), .B(n11404), .Z(c[1482]) );
  XOR U15502 ( .A(n11405), .B(n11406), .Z(n11402) );
  ANDN U15503 ( .B(n11407), .A(n11408), .Z(n11405) );
  XNOR U15504 ( .A(b[1481]), .B(n11406), .Z(n11407) );
  XNOR U15505 ( .A(b[1481]), .B(n11408), .Z(c[1481]) );
  XOR U15506 ( .A(n11409), .B(n11410), .Z(n11406) );
  ANDN U15507 ( .B(n11411), .A(n11412), .Z(n11409) );
  XNOR U15508 ( .A(b[1480]), .B(n11410), .Z(n11411) );
  XNOR U15509 ( .A(b[1480]), .B(n11412), .Z(c[1480]) );
  XOR U15510 ( .A(n11413), .B(n11414), .Z(n11410) );
  ANDN U15511 ( .B(n11415), .A(n11416), .Z(n11413) );
  XNOR U15512 ( .A(b[1479]), .B(n11414), .Z(n11415) );
  XNOR U15513 ( .A(b[147]), .B(n11417), .Z(c[147]) );
  XNOR U15514 ( .A(b[1479]), .B(n11416), .Z(c[1479]) );
  XOR U15515 ( .A(n11418), .B(n11419), .Z(n11414) );
  ANDN U15516 ( .B(n11420), .A(n11421), .Z(n11418) );
  XNOR U15517 ( .A(b[1478]), .B(n11419), .Z(n11420) );
  XNOR U15518 ( .A(b[1478]), .B(n11421), .Z(c[1478]) );
  XOR U15519 ( .A(n11422), .B(n11423), .Z(n11419) );
  ANDN U15520 ( .B(n11424), .A(n11425), .Z(n11422) );
  XNOR U15521 ( .A(b[1477]), .B(n11423), .Z(n11424) );
  XNOR U15522 ( .A(b[1477]), .B(n11425), .Z(c[1477]) );
  XOR U15523 ( .A(n11426), .B(n11427), .Z(n11423) );
  ANDN U15524 ( .B(n11428), .A(n11429), .Z(n11426) );
  XNOR U15525 ( .A(b[1476]), .B(n11427), .Z(n11428) );
  XNOR U15526 ( .A(b[1476]), .B(n11429), .Z(c[1476]) );
  XOR U15527 ( .A(n11430), .B(n11431), .Z(n11427) );
  ANDN U15528 ( .B(n11432), .A(n11433), .Z(n11430) );
  XNOR U15529 ( .A(b[1475]), .B(n11431), .Z(n11432) );
  XNOR U15530 ( .A(b[1475]), .B(n11433), .Z(c[1475]) );
  XOR U15531 ( .A(n11434), .B(n11435), .Z(n11431) );
  ANDN U15532 ( .B(n11436), .A(n11437), .Z(n11434) );
  XNOR U15533 ( .A(b[1474]), .B(n11435), .Z(n11436) );
  XNOR U15534 ( .A(b[1474]), .B(n11437), .Z(c[1474]) );
  XOR U15535 ( .A(n11438), .B(n11439), .Z(n11435) );
  ANDN U15536 ( .B(n11440), .A(n11441), .Z(n11438) );
  XNOR U15537 ( .A(b[1473]), .B(n11439), .Z(n11440) );
  XNOR U15538 ( .A(b[1473]), .B(n11441), .Z(c[1473]) );
  XOR U15539 ( .A(n11442), .B(n11443), .Z(n11439) );
  ANDN U15540 ( .B(n11444), .A(n11445), .Z(n11442) );
  XNOR U15541 ( .A(b[1472]), .B(n11443), .Z(n11444) );
  XNOR U15542 ( .A(b[1472]), .B(n11445), .Z(c[1472]) );
  XOR U15543 ( .A(n11446), .B(n11447), .Z(n11443) );
  ANDN U15544 ( .B(n11448), .A(n11449), .Z(n11446) );
  XNOR U15545 ( .A(b[1471]), .B(n11447), .Z(n11448) );
  XNOR U15546 ( .A(b[1471]), .B(n11449), .Z(c[1471]) );
  XOR U15547 ( .A(n11450), .B(n11451), .Z(n11447) );
  ANDN U15548 ( .B(n11452), .A(n11453), .Z(n11450) );
  XNOR U15549 ( .A(b[1470]), .B(n11451), .Z(n11452) );
  XNOR U15550 ( .A(b[1470]), .B(n11453), .Z(c[1470]) );
  XOR U15551 ( .A(n11454), .B(n11455), .Z(n11451) );
  ANDN U15552 ( .B(n11456), .A(n11457), .Z(n11454) );
  XNOR U15553 ( .A(b[1469]), .B(n11455), .Z(n11456) );
  XNOR U15554 ( .A(b[146]), .B(n11458), .Z(c[146]) );
  XNOR U15555 ( .A(b[1469]), .B(n11457), .Z(c[1469]) );
  XOR U15556 ( .A(n11459), .B(n11460), .Z(n11455) );
  ANDN U15557 ( .B(n11461), .A(n11462), .Z(n11459) );
  XNOR U15558 ( .A(b[1468]), .B(n11460), .Z(n11461) );
  XNOR U15559 ( .A(b[1468]), .B(n11462), .Z(c[1468]) );
  XOR U15560 ( .A(n11463), .B(n11464), .Z(n11460) );
  ANDN U15561 ( .B(n11465), .A(n11466), .Z(n11463) );
  XNOR U15562 ( .A(b[1467]), .B(n11464), .Z(n11465) );
  XNOR U15563 ( .A(b[1467]), .B(n11466), .Z(c[1467]) );
  XOR U15564 ( .A(n11467), .B(n11468), .Z(n11464) );
  ANDN U15565 ( .B(n11469), .A(n11470), .Z(n11467) );
  XNOR U15566 ( .A(b[1466]), .B(n11468), .Z(n11469) );
  XNOR U15567 ( .A(b[1466]), .B(n11470), .Z(c[1466]) );
  XOR U15568 ( .A(n11471), .B(n11472), .Z(n11468) );
  ANDN U15569 ( .B(n11473), .A(n11474), .Z(n11471) );
  XNOR U15570 ( .A(b[1465]), .B(n11472), .Z(n11473) );
  XNOR U15571 ( .A(b[1465]), .B(n11474), .Z(c[1465]) );
  XOR U15572 ( .A(n11475), .B(n11476), .Z(n11472) );
  ANDN U15573 ( .B(n11477), .A(n11478), .Z(n11475) );
  XNOR U15574 ( .A(b[1464]), .B(n11476), .Z(n11477) );
  XNOR U15575 ( .A(b[1464]), .B(n11478), .Z(c[1464]) );
  XOR U15576 ( .A(n11479), .B(n11480), .Z(n11476) );
  ANDN U15577 ( .B(n11481), .A(n11482), .Z(n11479) );
  XNOR U15578 ( .A(b[1463]), .B(n11480), .Z(n11481) );
  XNOR U15579 ( .A(b[1463]), .B(n11482), .Z(c[1463]) );
  XOR U15580 ( .A(n11483), .B(n11484), .Z(n11480) );
  ANDN U15581 ( .B(n11485), .A(n11486), .Z(n11483) );
  XNOR U15582 ( .A(b[1462]), .B(n11484), .Z(n11485) );
  XNOR U15583 ( .A(b[1462]), .B(n11486), .Z(c[1462]) );
  XOR U15584 ( .A(n11487), .B(n11488), .Z(n11484) );
  ANDN U15585 ( .B(n11489), .A(n11490), .Z(n11487) );
  XNOR U15586 ( .A(b[1461]), .B(n11488), .Z(n11489) );
  XNOR U15587 ( .A(b[1461]), .B(n11490), .Z(c[1461]) );
  XOR U15588 ( .A(n11491), .B(n11492), .Z(n11488) );
  ANDN U15589 ( .B(n11493), .A(n11494), .Z(n11491) );
  XNOR U15590 ( .A(b[1460]), .B(n11492), .Z(n11493) );
  XNOR U15591 ( .A(b[1460]), .B(n11494), .Z(c[1460]) );
  XOR U15592 ( .A(n11495), .B(n11496), .Z(n11492) );
  ANDN U15593 ( .B(n11497), .A(n11498), .Z(n11495) );
  XNOR U15594 ( .A(b[1459]), .B(n11496), .Z(n11497) );
  XNOR U15595 ( .A(b[145]), .B(n11499), .Z(c[145]) );
  XNOR U15596 ( .A(b[1459]), .B(n11498), .Z(c[1459]) );
  XOR U15597 ( .A(n11500), .B(n11501), .Z(n11496) );
  ANDN U15598 ( .B(n11502), .A(n11503), .Z(n11500) );
  XNOR U15599 ( .A(b[1458]), .B(n11501), .Z(n11502) );
  XNOR U15600 ( .A(b[1458]), .B(n11503), .Z(c[1458]) );
  XOR U15601 ( .A(n11504), .B(n11505), .Z(n11501) );
  ANDN U15602 ( .B(n11506), .A(n11507), .Z(n11504) );
  XNOR U15603 ( .A(b[1457]), .B(n11505), .Z(n11506) );
  XNOR U15604 ( .A(b[1457]), .B(n11507), .Z(c[1457]) );
  XOR U15605 ( .A(n11508), .B(n11509), .Z(n11505) );
  ANDN U15606 ( .B(n11510), .A(n11511), .Z(n11508) );
  XNOR U15607 ( .A(b[1456]), .B(n11509), .Z(n11510) );
  XNOR U15608 ( .A(b[1456]), .B(n11511), .Z(c[1456]) );
  XOR U15609 ( .A(n11512), .B(n11513), .Z(n11509) );
  ANDN U15610 ( .B(n11514), .A(n11515), .Z(n11512) );
  XNOR U15611 ( .A(b[1455]), .B(n11513), .Z(n11514) );
  XNOR U15612 ( .A(b[1455]), .B(n11515), .Z(c[1455]) );
  XOR U15613 ( .A(n11516), .B(n11517), .Z(n11513) );
  ANDN U15614 ( .B(n11518), .A(n11519), .Z(n11516) );
  XNOR U15615 ( .A(b[1454]), .B(n11517), .Z(n11518) );
  XNOR U15616 ( .A(b[1454]), .B(n11519), .Z(c[1454]) );
  XOR U15617 ( .A(n11520), .B(n11521), .Z(n11517) );
  ANDN U15618 ( .B(n11522), .A(n11523), .Z(n11520) );
  XNOR U15619 ( .A(b[1453]), .B(n11521), .Z(n11522) );
  XNOR U15620 ( .A(b[1453]), .B(n11523), .Z(c[1453]) );
  XOR U15621 ( .A(n11524), .B(n11525), .Z(n11521) );
  ANDN U15622 ( .B(n11526), .A(n11527), .Z(n11524) );
  XNOR U15623 ( .A(b[1452]), .B(n11525), .Z(n11526) );
  XNOR U15624 ( .A(b[1452]), .B(n11527), .Z(c[1452]) );
  XOR U15625 ( .A(n11528), .B(n11529), .Z(n11525) );
  ANDN U15626 ( .B(n11530), .A(n11531), .Z(n11528) );
  XNOR U15627 ( .A(b[1451]), .B(n11529), .Z(n11530) );
  XNOR U15628 ( .A(b[1451]), .B(n11531), .Z(c[1451]) );
  XOR U15629 ( .A(n11532), .B(n11533), .Z(n11529) );
  ANDN U15630 ( .B(n11534), .A(n11535), .Z(n11532) );
  XNOR U15631 ( .A(b[1450]), .B(n11533), .Z(n11534) );
  XNOR U15632 ( .A(b[1450]), .B(n11535), .Z(c[1450]) );
  XOR U15633 ( .A(n11536), .B(n11537), .Z(n11533) );
  ANDN U15634 ( .B(n11538), .A(n11539), .Z(n11536) );
  XNOR U15635 ( .A(b[1449]), .B(n11537), .Z(n11538) );
  XNOR U15636 ( .A(b[144]), .B(n11540), .Z(c[144]) );
  XNOR U15637 ( .A(b[1449]), .B(n11539), .Z(c[1449]) );
  XOR U15638 ( .A(n11541), .B(n11542), .Z(n11537) );
  ANDN U15639 ( .B(n11543), .A(n11544), .Z(n11541) );
  XNOR U15640 ( .A(b[1448]), .B(n11542), .Z(n11543) );
  XNOR U15641 ( .A(b[1448]), .B(n11544), .Z(c[1448]) );
  XOR U15642 ( .A(n11545), .B(n11546), .Z(n11542) );
  ANDN U15643 ( .B(n11547), .A(n11548), .Z(n11545) );
  XNOR U15644 ( .A(b[1447]), .B(n11546), .Z(n11547) );
  XNOR U15645 ( .A(b[1447]), .B(n11548), .Z(c[1447]) );
  XOR U15646 ( .A(n11549), .B(n11550), .Z(n11546) );
  ANDN U15647 ( .B(n11551), .A(n11552), .Z(n11549) );
  XNOR U15648 ( .A(b[1446]), .B(n11550), .Z(n11551) );
  XNOR U15649 ( .A(b[1446]), .B(n11552), .Z(c[1446]) );
  XOR U15650 ( .A(n11553), .B(n11554), .Z(n11550) );
  ANDN U15651 ( .B(n11555), .A(n11556), .Z(n11553) );
  XNOR U15652 ( .A(b[1445]), .B(n11554), .Z(n11555) );
  XNOR U15653 ( .A(b[1445]), .B(n11556), .Z(c[1445]) );
  XOR U15654 ( .A(n11557), .B(n11558), .Z(n11554) );
  ANDN U15655 ( .B(n11559), .A(n11560), .Z(n11557) );
  XNOR U15656 ( .A(b[1444]), .B(n11558), .Z(n11559) );
  XNOR U15657 ( .A(b[1444]), .B(n11560), .Z(c[1444]) );
  XOR U15658 ( .A(n11561), .B(n11562), .Z(n11558) );
  ANDN U15659 ( .B(n11563), .A(n11564), .Z(n11561) );
  XNOR U15660 ( .A(b[1443]), .B(n11562), .Z(n11563) );
  XNOR U15661 ( .A(b[1443]), .B(n11564), .Z(c[1443]) );
  XOR U15662 ( .A(n11565), .B(n11566), .Z(n11562) );
  ANDN U15663 ( .B(n11567), .A(n11568), .Z(n11565) );
  XNOR U15664 ( .A(b[1442]), .B(n11566), .Z(n11567) );
  XNOR U15665 ( .A(b[1442]), .B(n11568), .Z(c[1442]) );
  XOR U15666 ( .A(n11569), .B(n11570), .Z(n11566) );
  ANDN U15667 ( .B(n11571), .A(n11572), .Z(n11569) );
  XNOR U15668 ( .A(b[1441]), .B(n11570), .Z(n11571) );
  XNOR U15669 ( .A(b[1441]), .B(n11572), .Z(c[1441]) );
  XOR U15670 ( .A(n11573), .B(n11574), .Z(n11570) );
  ANDN U15671 ( .B(n11575), .A(n11576), .Z(n11573) );
  XNOR U15672 ( .A(b[1440]), .B(n11574), .Z(n11575) );
  XNOR U15673 ( .A(b[1440]), .B(n11576), .Z(c[1440]) );
  XOR U15674 ( .A(n11577), .B(n11578), .Z(n11574) );
  ANDN U15675 ( .B(n11579), .A(n11580), .Z(n11577) );
  XNOR U15676 ( .A(b[1439]), .B(n11578), .Z(n11579) );
  XNOR U15677 ( .A(b[143]), .B(n11581), .Z(c[143]) );
  XNOR U15678 ( .A(b[1439]), .B(n11580), .Z(c[1439]) );
  XOR U15679 ( .A(n11582), .B(n11583), .Z(n11578) );
  ANDN U15680 ( .B(n11584), .A(n11585), .Z(n11582) );
  XNOR U15681 ( .A(b[1438]), .B(n11583), .Z(n11584) );
  XNOR U15682 ( .A(b[1438]), .B(n11585), .Z(c[1438]) );
  XOR U15683 ( .A(n11586), .B(n11587), .Z(n11583) );
  ANDN U15684 ( .B(n11588), .A(n11589), .Z(n11586) );
  XNOR U15685 ( .A(b[1437]), .B(n11587), .Z(n11588) );
  XNOR U15686 ( .A(b[1437]), .B(n11589), .Z(c[1437]) );
  XOR U15687 ( .A(n11590), .B(n11591), .Z(n11587) );
  ANDN U15688 ( .B(n11592), .A(n11593), .Z(n11590) );
  XNOR U15689 ( .A(b[1436]), .B(n11591), .Z(n11592) );
  XNOR U15690 ( .A(b[1436]), .B(n11593), .Z(c[1436]) );
  XOR U15691 ( .A(n11594), .B(n11595), .Z(n11591) );
  ANDN U15692 ( .B(n11596), .A(n11597), .Z(n11594) );
  XNOR U15693 ( .A(b[1435]), .B(n11595), .Z(n11596) );
  XNOR U15694 ( .A(b[1435]), .B(n11597), .Z(c[1435]) );
  XOR U15695 ( .A(n11598), .B(n11599), .Z(n11595) );
  ANDN U15696 ( .B(n11600), .A(n11601), .Z(n11598) );
  XNOR U15697 ( .A(b[1434]), .B(n11599), .Z(n11600) );
  XNOR U15698 ( .A(b[1434]), .B(n11601), .Z(c[1434]) );
  XOR U15699 ( .A(n11602), .B(n11603), .Z(n11599) );
  ANDN U15700 ( .B(n11604), .A(n11605), .Z(n11602) );
  XNOR U15701 ( .A(b[1433]), .B(n11603), .Z(n11604) );
  XNOR U15702 ( .A(b[1433]), .B(n11605), .Z(c[1433]) );
  XOR U15703 ( .A(n11606), .B(n11607), .Z(n11603) );
  ANDN U15704 ( .B(n11608), .A(n11609), .Z(n11606) );
  XNOR U15705 ( .A(b[1432]), .B(n11607), .Z(n11608) );
  XNOR U15706 ( .A(b[1432]), .B(n11609), .Z(c[1432]) );
  XOR U15707 ( .A(n11610), .B(n11611), .Z(n11607) );
  ANDN U15708 ( .B(n11612), .A(n11613), .Z(n11610) );
  XNOR U15709 ( .A(b[1431]), .B(n11611), .Z(n11612) );
  XNOR U15710 ( .A(b[1431]), .B(n11613), .Z(c[1431]) );
  XOR U15711 ( .A(n11614), .B(n11615), .Z(n11611) );
  ANDN U15712 ( .B(n11616), .A(n11617), .Z(n11614) );
  XNOR U15713 ( .A(b[1430]), .B(n11615), .Z(n11616) );
  XNOR U15714 ( .A(b[1430]), .B(n11617), .Z(c[1430]) );
  XOR U15715 ( .A(n11618), .B(n11619), .Z(n11615) );
  ANDN U15716 ( .B(n11620), .A(n11621), .Z(n11618) );
  XNOR U15717 ( .A(b[1429]), .B(n11619), .Z(n11620) );
  XNOR U15718 ( .A(b[142]), .B(n11622), .Z(c[142]) );
  XNOR U15719 ( .A(b[1429]), .B(n11621), .Z(c[1429]) );
  XOR U15720 ( .A(n11623), .B(n11624), .Z(n11619) );
  ANDN U15721 ( .B(n11625), .A(n11626), .Z(n11623) );
  XNOR U15722 ( .A(b[1428]), .B(n11624), .Z(n11625) );
  XNOR U15723 ( .A(b[1428]), .B(n11626), .Z(c[1428]) );
  XOR U15724 ( .A(n11627), .B(n11628), .Z(n11624) );
  ANDN U15725 ( .B(n11629), .A(n11630), .Z(n11627) );
  XNOR U15726 ( .A(b[1427]), .B(n11628), .Z(n11629) );
  XNOR U15727 ( .A(b[1427]), .B(n11630), .Z(c[1427]) );
  XOR U15728 ( .A(n11631), .B(n11632), .Z(n11628) );
  ANDN U15729 ( .B(n11633), .A(n11634), .Z(n11631) );
  XNOR U15730 ( .A(b[1426]), .B(n11632), .Z(n11633) );
  XNOR U15731 ( .A(b[1426]), .B(n11634), .Z(c[1426]) );
  XOR U15732 ( .A(n11635), .B(n11636), .Z(n11632) );
  ANDN U15733 ( .B(n11637), .A(n11638), .Z(n11635) );
  XNOR U15734 ( .A(b[1425]), .B(n11636), .Z(n11637) );
  XNOR U15735 ( .A(b[1425]), .B(n11638), .Z(c[1425]) );
  XOR U15736 ( .A(n11639), .B(n11640), .Z(n11636) );
  ANDN U15737 ( .B(n11641), .A(n11642), .Z(n11639) );
  XNOR U15738 ( .A(b[1424]), .B(n11640), .Z(n11641) );
  XNOR U15739 ( .A(b[1424]), .B(n11642), .Z(c[1424]) );
  XOR U15740 ( .A(n11643), .B(n11644), .Z(n11640) );
  ANDN U15741 ( .B(n11645), .A(n11646), .Z(n11643) );
  XNOR U15742 ( .A(b[1423]), .B(n11644), .Z(n11645) );
  XNOR U15743 ( .A(b[1423]), .B(n11646), .Z(c[1423]) );
  XOR U15744 ( .A(n11647), .B(n11648), .Z(n11644) );
  ANDN U15745 ( .B(n11649), .A(n11650), .Z(n11647) );
  XNOR U15746 ( .A(b[1422]), .B(n11648), .Z(n11649) );
  XNOR U15747 ( .A(b[1422]), .B(n11650), .Z(c[1422]) );
  XOR U15748 ( .A(n11651), .B(n11652), .Z(n11648) );
  ANDN U15749 ( .B(n11653), .A(n11654), .Z(n11651) );
  XNOR U15750 ( .A(b[1421]), .B(n11652), .Z(n11653) );
  XNOR U15751 ( .A(b[1421]), .B(n11654), .Z(c[1421]) );
  XOR U15752 ( .A(n11655), .B(n11656), .Z(n11652) );
  ANDN U15753 ( .B(n11657), .A(n11658), .Z(n11655) );
  XNOR U15754 ( .A(b[1420]), .B(n11656), .Z(n11657) );
  XNOR U15755 ( .A(b[1420]), .B(n11658), .Z(c[1420]) );
  XOR U15756 ( .A(n11659), .B(n11660), .Z(n11656) );
  ANDN U15757 ( .B(n11661), .A(n11662), .Z(n11659) );
  XNOR U15758 ( .A(b[1419]), .B(n11660), .Z(n11661) );
  XNOR U15759 ( .A(b[141]), .B(n11663), .Z(c[141]) );
  XNOR U15760 ( .A(b[1419]), .B(n11662), .Z(c[1419]) );
  XOR U15761 ( .A(n11664), .B(n11665), .Z(n11660) );
  ANDN U15762 ( .B(n11666), .A(n11667), .Z(n11664) );
  XNOR U15763 ( .A(b[1418]), .B(n11665), .Z(n11666) );
  XNOR U15764 ( .A(b[1418]), .B(n11667), .Z(c[1418]) );
  XOR U15765 ( .A(n11668), .B(n11669), .Z(n11665) );
  ANDN U15766 ( .B(n11670), .A(n11671), .Z(n11668) );
  XNOR U15767 ( .A(b[1417]), .B(n11669), .Z(n11670) );
  XNOR U15768 ( .A(b[1417]), .B(n11671), .Z(c[1417]) );
  XOR U15769 ( .A(n11672), .B(n11673), .Z(n11669) );
  ANDN U15770 ( .B(n11674), .A(n11675), .Z(n11672) );
  XNOR U15771 ( .A(b[1416]), .B(n11673), .Z(n11674) );
  XNOR U15772 ( .A(b[1416]), .B(n11675), .Z(c[1416]) );
  XOR U15773 ( .A(n11676), .B(n11677), .Z(n11673) );
  ANDN U15774 ( .B(n11678), .A(n11679), .Z(n11676) );
  XNOR U15775 ( .A(b[1415]), .B(n11677), .Z(n11678) );
  XNOR U15776 ( .A(b[1415]), .B(n11679), .Z(c[1415]) );
  XOR U15777 ( .A(n11680), .B(n11681), .Z(n11677) );
  ANDN U15778 ( .B(n11682), .A(n11683), .Z(n11680) );
  XNOR U15779 ( .A(b[1414]), .B(n11681), .Z(n11682) );
  XNOR U15780 ( .A(b[1414]), .B(n11683), .Z(c[1414]) );
  XOR U15781 ( .A(n11684), .B(n11685), .Z(n11681) );
  ANDN U15782 ( .B(n11686), .A(n11687), .Z(n11684) );
  XNOR U15783 ( .A(b[1413]), .B(n11685), .Z(n11686) );
  XNOR U15784 ( .A(b[1413]), .B(n11687), .Z(c[1413]) );
  XOR U15785 ( .A(n11688), .B(n11689), .Z(n11685) );
  ANDN U15786 ( .B(n11690), .A(n11691), .Z(n11688) );
  XNOR U15787 ( .A(b[1412]), .B(n11689), .Z(n11690) );
  XNOR U15788 ( .A(b[1412]), .B(n11691), .Z(c[1412]) );
  XOR U15789 ( .A(n11692), .B(n11693), .Z(n11689) );
  ANDN U15790 ( .B(n11694), .A(n11695), .Z(n11692) );
  XNOR U15791 ( .A(b[1411]), .B(n11693), .Z(n11694) );
  XNOR U15792 ( .A(b[1411]), .B(n11695), .Z(c[1411]) );
  XOR U15793 ( .A(n11696), .B(n11697), .Z(n11693) );
  ANDN U15794 ( .B(n11698), .A(n11699), .Z(n11696) );
  XNOR U15795 ( .A(b[1410]), .B(n11697), .Z(n11698) );
  XNOR U15796 ( .A(b[1410]), .B(n11699), .Z(c[1410]) );
  XOR U15797 ( .A(n11700), .B(n11701), .Z(n11697) );
  ANDN U15798 ( .B(n11702), .A(n11703), .Z(n11700) );
  XNOR U15799 ( .A(b[1409]), .B(n11701), .Z(n11702) );
  XNOR U15800 ( .A(b[140]), .B(n11704), .Z(c[140]) );
  XNOR U15801 ( .A(b[1409]), .B(n11703), .Z(c[1409]) );
  XOR U15802 ( .A(n11705), .B(n11706), .Z(n11701) );
  ANDN U15803 ( .B(n11707), .A(n11708), .Z(n11705) );
  XNOR U15804 ( .A(b[1408]), .B(n11706), .Z(n11707) );
  XNOR U15805 ( .A(b[1408]), .B(n11708), .Z(c[1408]) );
  XOR U15806 ( .A(n11709), .B(n11710), .Z(n11706) );
  ANDN U15807 ( .B(n11711), .A(n11712), .Z(n11709) );
  XNOR U15808 ( .A(b[1407]), .B(n11710), .Z(n11711) );
  XNOR U15809 ( .A(b[1407]), .B(n11712), .Z(c[1407]) );
  XOR U15810 ( .A(n11713), .B(n11714), .Z(n11710) );
  ANDN U15811 ( .B(n11715), .A(n11716), .Z(n11713) );
  XNOR U15812 ( .A(b[1406]), .B(n11714), .Z(n11715) );
  XNOR U15813 ( .A(b[1406]), .B(n11716), .Z(c[1406]) );
  XOR U15814 ( .A(n11717), .B(n11718), .Z(n11714) );
  ANDN U15815 ( .B(n11719), .A(n11720), .Z(n11717) );
  XNOR U15816 ( .A(b[1405]), .B(n11718), .Z(n11719) );
  XNOR U15817 ( .A(b[1405]), .B(n11720), .Z(c[1405]) );
  XOR U15818 ( .A(n11721), .B(n11722), .Z(n11718) );
  ANDN U15819 ( .B(n11723), .A(n11724), .Z(n11721) );
  XNOR U15820 ( .A(b[1404]), .B(n11722), .Z(n11723) );
  XNOR U15821 ( .A(b[1404]), .B(n11724), .Z(c[1404]) );
  XOR U15822 ( .A(n11725), .B(n11726), .Z(n11722) );
  ANDN U15823 ( .B(n11727), .A(n11728), .Z(n11725) );
  XNOR U15824 ( .A(b[1403]), .B(n11726), .Z(n11727) );
  XNOR U15825 ( .A(b[1403]), .B(n11728), .Z(c[1403]) );
  XOR U15826 ( .A(n11729), .B(n11730), .Z(n11726) );
  ANDN U15827 ( .B(n11731), .A(n11732), .Z(n11729) );
  XNOR U15828 ( .A(b[1402]), .B(n11730), .Z(n11731) );
  XNOR U15829 ( .A(b[1402]), .B(n11732), .Z(c[1402]) );
  XOR U15830 ( .A(n11733), .B(n11734), .Z(n11730) );
  ANDN U15831 ( .B(n11735), .A(n11736), .Z(n11733) );
  XNOR U15832 ( .A(b[1401]), .B(n11734), .Z(n11735) );
  XNOR U15833 ( .A(b[1401]), .B(n11736), .Z(c[1401]) );
  XOR U15834 ( .A(n11737), .B(n11738), .Z(n11734) );
  ANDN U15835 ( .B(n11739), .A(n11740), .Z(n11737) );
  XNOR U15836 ( .A(b[1400]), .B(n11738), .Z(n11739) );
  XNOR U15837 ( .A(b[1400]), .B(n11740), .Z(c[1400]) );
  XOR U15838 ( .A(n11741), .B(n11742), .Z(n11738) );
  ANDN U15839 ( .B(n11743), .A(n11744), .Z(n11741) );
  XNOR U15840 ( .A(b[1399]), .B(n11742), .Z(n11743) );
  XNOR U15841 ( .A(b[13]), .B(n11745), .Z(c[13]) );
  XNOR U15842 ( .A(b[139]), .B(n11746), .Z(c[139]) );
  XNOR U15843 ( .A(b[1399]), .B(n11744), .Z(c[1399]) );
  XOR U15844 ( .A(n11747), .B(n11748), .Z(n11742) );
  ANDN U15845 ( .B(n11749), .A(n11750), .Z(n11747) );
  XNOR U15846 ( .A(b[1398]), .B(n11748), .Z(n11749) );
  XNOR U15847 ( .A(b[1398]), .B(n11750), .Z(c[1398]) );
  XOR U15848 ( .A(n11751), .B(n11752), .Z(n11748) );
  ANDN U15849 ( .B(n11753), .A(n11754), .Z(n11751) );
  XNOR U15850 ( .A(b[1397]), .B(n11752), .Z(n11753) );
  XNOR U15851 ( .A(b[1397]), .B(n11754), .Z(c[1397]) );
  XOR U15852 ( .A(n11755), .B(n11756), .Z(n11752) );
  ANDN U15853 ( .B(n11757), .A(n11758), .Z(n11755) );
  XNOR U15854 ( .A(b[1396]), .B(n11756), .Z(n11757) );
  XNOR U15855 ( .A(b[1396]), .B(n11758), .Z(c[1396]) );
  XOR U15856 ( .A(n11759), .B(n11760), .Z(n11756) );
  ANDN U15857 ( .B(n11761), .A(n11762), .Z(n11759) );
  XNOR U15858 ( .A(b[1395]), .B(n11760), .Z(n11761) );
  XNOR U15859 ( .A(b[1395]), .B(n11762), .Z(c[1395]) );
  XOR U15860 ( .A(n11763), .B(n11764), .Z(n11760) );
  ANDN U15861 ( .B(n11765), .A(n11766), .Z(n11763) );
  XNOR U15862 ( .A(b[1394]), .B(n11764), .Z(n11765) );
  XNOR U15863 ( .A(b[1394]), .B(n11766), .Z(c[1394]) );
  XOR U15864 ( .A(n11767), .B(n11768), .Z(n11764) );
  ANDN U15865 ( .B(n11769), .A(n11770), .Z(n11767) );
  XNOR U15866 ( .A(b[1393]), .B(n11768), .Z(n11769) );
  XNOR U15867 ( .A(b[1393]), .B(n11770), .Z(c[1393]) );
  XOR U15868 ( .A(n11771), .B(n11772), .Z(n11768) );
  ANDN U15869 ( .B(n11773), .A(n11774), .Z(n11771) );
  XNOR U15870 ( .A(b[1392]), .B(n11772), .Z(n11773) );
  XNOR U15871 ( .A(b[1392]), .B(n11774), .Z(c[1392]) );
  XOR U15872 ( .A(n11775), .B(n11776), .Z(n11772) );
  ANDN U15873 ( .B(n11777), .A(n11778), .Z(n11775) );
  XNOR U15874 ( .A(b[1391]), .B(n11776), .Z(n11777) );
  XNOR U15875 ( .A(b[1391]), .B(n11778), .Z(c[1391]) );
  XOR U15876 ( .A(n11779), .B(n11780), .Z(n11776) );
  ANDN U15877 ( .B(n11781), .A(n11782), .Z(n11779) );
  XNOR U15878 ( .A(b[1390]), .B(n11780), .Z(n11781) );
  XNOR U15879 ( .A(b[1390]), .B(n11782), .Z(c[1390]) );
  XOR U15880 ( .A(n11783), .B(n11784), .Z(n11780) );
  ANDN U15881 ( .B(n11785), .A(n11786), .Z(n11783) );
  XNOR U15882 ( .A(b[1389]), .B(n11784), .Z(n11785) );
  XNOR U15883 ( .A(b[138]), .B(n11787), .Z(c[138]) );
  XNOR U15884 ( .A(b[1389]), .B(n11786), .Z(c[1389]) );
  XOR U15885 ( .A(n11788), .B(n11789), .Z(n11784) );
  ANDN U15886 ( .B(n11790), .A(n11791), .Z(n11788) );
  XNOR U15887 ( .A(b[1388]), .B(n11789), .Z(n11790) );
  XNOR U15888 ( .A(b[1388]), .B(n11791), .Z(c[1388]) );
  XOR U15889 ( .A(n11792), .B(n11793), .Z(n11789) );
  ANDN U15890 ( .B(n11794), .A(n11795), .Z(n11792) );
  XNOR U15891 ( .A(b[1387]), .B(n11793), .Z(n11794) );
  XNOR U15892 ( .A(b[1387]), .B(n11795), .Z(c[1387]) );
  XOR U15893 ( .A(n11796), .B(n11797), .Z(n11793) );
  ANDN U15894 ( .B(n11798), .A(n11799), .Z(n11796) );
  XNOR U15895 ( .A(b[1386]), .B(n11797), .Z(n11798) );
  XNOR U15896 ( .A(b[1386]), .B(n11799), .Z(c[1386]) );
  XOR U15897 ( .A(n11800), .B(n11801), .Z(n11797) );
  ANDN U15898 ( .B(n11802), .A(n11803), .Z(n11800) );
  XNOR U15899 ( .A(b[1385]), .B(n11801), .Z(n11802) );
  XNOR U15900 ( .A(b[1385]), .B(n11803), .Z(c[1385]) );
  XOR U15901 ( .A(n11804), .B(n11805), .Z(n11801) );
  ANDN U15902 ( .B(n11806), .A(n11807), .Z(n11804) );
  XNOR U15903 ( .A(b[1384]), .B(n11805), .Z(n11806) );
  XNOR U15904 ( .A(b[1384]), .B(n11807), .Z(c[1384]) );
  XOR U15905 ( .A(n11808), .B(n11809), .Z(n11805) );
  ANDN U15906 ( .B(n11810), .A(n11811), .Z(n11808) );
  XNOR U15907 ( .A(b[1383]), .B(n11809), .Z(n11810) );
  XNOR U15908 ( .A(b[1383]), .B(n11811), .Z(c[1383]) );
  XOR U15909 ( .A(n11812), .B(n11813), .Z(n11809) );
  ANDN U15910 ( .B(n11814), .A(n11815), .Z(n11812) );
  XNOR U15911 ( .A(b[1382]), .B(n11813), .Z(n11814) );
  XNOR U15912 ( .A(b[1382]), .B(n11815), .Z(c[1382]) );
  XOR U15913 ( .A(n11816), .B(n11817), .Z(n11813) );
  ANDN U15914 ( .B(n11818), .A(n11819), .Z(n11816) );
  XNOR U15915 ( .A(b[1381]), .B(n11817), .Z(n11818) );
  XNOR U15916 ( .A(b[1381]), .B(n11819), .Z(c[1381]) );
  XOR U15917 ( .A(n11820), .B(n11821), .Z(n11817) );
  ANDN U15918 ( .B(n11822), .A(n11823), .Z(n11820) );
  XNOR U15919 ( .A(b[1380]), .B(n11821), .Z(n11822) );
  XNOR U15920 ( .A(b[1380]), .B(n11823), .Z(c[1380]) );
  XOR U15921 ( .A(n11824), .B(n11825), .Z(n11821) );
  ANDN U15922 ( .B(n11826), .A(n11827), .Z(n11824) );
  XNOR U15923 ( .A(b[1379]), .B(n11825), .Z(n11826) );
  XNOR U15924 ( .A(b[137]), .B(n11828), .Z(c[137]) );
  XNOR U15925 ( .A(b[1379]), .B(n11827), .Z(c[1379]) );
  XOR U15926 ( .A(n11829), .B(n11830), .Z(n11825) );
  ANDN U15927 ( .B(n11831), .A(n11832), .Z(n11829) );
  XNOR U15928 ( .A(b[1378]), .B(n11830), .Z(n11831) );
  XNOR U15929 ( .A(b[1378]), .B(n11832), .Z(c[1378]) );
  XOR U15930 ( .A(n11833), .B(n11834), .Z(n11830) );
  ANDN U15931 ( .B(n11835), .A(n11836), .Z(n11833) );
  XNOR U15932 ( .A(b[1377]), .B(n11834), .Z(n11835) );
  XNOR U15933 ( .A(b[1377]), .B(n11836), .Z(c[1377]) );
  XOR U15934 ( .A(n11837), .B(n11838), .Z(n11834) );
  ANDN U15935 ( .B(n11839), .A(n11840), .Z(n11837) );
  XNOR U15936 ( .A(b[1376]), .B(n11838), .Z(n11839) );
  XNOR U15937 ( .A(b[1376]), .B(n11840), .Z(c[1376]) );
  XOR U15938 ( .A(n11841), .B(n11842), .Z(n11838) );
  ANDN U15939 ( .B(n11843), .A(n11844), .Z(n11841) );
  XNOR U15940 ( .A(b[1375]), .B(n11842), .Z(n11843) );
  XNOR U15941 ( .A(b[1375]), .B(n11844), .Z(c[1375]) );
  XOR U15942 ( .A(n11845), .B(n11846), .Z(n11842) );
  ANDN U15943 ( .B(n11847), .A(n11848), .Z(n11845) );
  XNOR U15944 ( .A(b[1374]), .B(n11846), .Z(n11847) );
  XNOR U15945 ( .A(b[1374]), .B(n11848), .Z(c[1374]) );
  XOR U15946 ( .A(n11849), .B(n11850), .Z(n11846) );
  ANDN U15947 ( .B(n11851), .A(n11852), .Z(n11849) );
  XNOR U15948 ( .A(b[1373]), .B(n11850), .Z(n11851) );
  XNOR U15949 ( .A(b[1373]), .B(n11852), .Z(c[1373]) );
  XOR U15950 ( .A(n11853), .B(n11854), .Z(n11850) );
  ANDN U15951 ( .B(n11855), .A(n11856), .Z(n11853) );
  XNOR U15952 ( .A(b[1372]), .B(n11854), .Z(n11855) );
  XNOR U15953 ( .A(b[1372]), .B(n11856), .Z(c[1372]) );
  XOR U15954 ( .A(n11857), .B(n11858), .Z(n11854) );
  ANDN U15955 ( .B(n11859), .A(n11860), .Z(n11857) );
  XNOR U15956 ( .A(b[1371]), .B(n11858), .Z(n11859) );
  XNOR U15957 ( .A(b[1371]), .B(n11860), .Z(c[1371]) );
  XOR U15958 ( .A(n11861), .B(n11862), .Z(n11858) );
  ANDN U15959 ( .B(n11863), .A(n11864), .Z(n11861) );
  XNOR U15960 ( .A(b[1370]), .B(n11862), .Z(n11863) );
  XNOR U15961 ( .A(b[1370]), .B(n11864), .Z(c[1370]) );
  XOR U15962 ( .A(n11865), .B(n11866), .Z(n11862) );
  ANDN U15963 ( .B(n11867), .A(n11868), .Z(n11865) );
  XNOR U15964 ( .A(b[1369]), .B(n11866), .Z(n11867) );
  XNOR U15965 ( .A(b[136]), .B(n11869), .Z(c[136]) );
  XNOR U15966 ( .A(b[1369]), .B(n11868), .Z(c[1369]) );
  XOR U15967 ( .A(n11870), .B(n11871), .Z(n11866) );
  ANDN U15968 ( .B(n11872), .A(n11873), .Z(n11870) );
  XNOR U15969 ( .A(b[1368]), .B(n11871), .Z(n11872) );
  XNOR U15970 ( .A(b[1368]), .B(n11873), .Z(c[1368]) );
  XOR U15971 ( .A(n11874), .B(n11875), .Z(n11871) );
  ANDN U15972 ( .B(n11876), .A(n11877), .Z(n11874) );
  XNOR U15973 ( .A(b[1367]), .B(n11875), .Z(n11876) );
  XNOR U15974 ( .A(b[1367]), .B(n11877), .Z(c[1367]) );
  XOR U15975 ( .A(n11878), .B(n11879), .Z(n11875) );
  ANDN U15976 ( .B(n11880), .A(n11881), .Z(n11878) );
  XNOR U15977 ( .A(b[1366]), .B(n11879), .Z(n11880) );
  XNOR U15978 ( .A(b[1366]), .B(n11881), .Z(c[1366]) );
  XOR U15979 ( .A(n11882), .B(n11883), .Z(n11879) );
  ANDN U15980 ( .B(n11884), .A(n11885), .Z(n11882) );
  XNOR U15981 ( .A(b[1365]), .B(n11883), .Z(n11884) );
  XNOR U15982 ( .A(b[1365]), .B(n11885), .Z(c[1365]) );
  XOR U15983 ( .A(n11886), .B(n11887), .Z(n11883) );
  ANDN U15984 ( .B(n11888), .A(n11889), .Z(n11886) );
  XNOR U15985 ( .A(b[1364]), .B(n11887), .Z(n11888) );
  XNOR U15986 ( .A(b[1364]), .B(n11889), .Z(c[1364]) );
  XOR U15987 ( .A(n11890), .B(n11891), .Z(n11887) );
  ANDN U15988 ( .B(n11892), .A(n11893), .Z(n11890) );
  XNOR U15989 ( .A(b[1363]), .B(n11891), .Z(n11892) );
  XNOR U15990 ( .A(b[1363]), .B(n11893), .Z(c[1363]) );
  XOR U15991 ( .A(n11894), .B(n11895), .Z(n11891) );
  ANDN U15992 ( .B(n11896), .A(n11897), .Z(n11894) );
  XNOR U15993 ( .A(b[1362]), .B(n11895), .Z(n11896) );
  XNOR U15994 ( .A(b[1362]), .B(n11897), .Z(c[1362]) );
  XOR U15995 ( .A(n11898), .B(n11899), .Z(n11895) );
  ANDN U15996 ( .B(n11900), .A(n11901), .Z(n11898) );
  XNOR U15997 ( .A(b[1361]), .B(n11899), .Z(n11900) );
  XNOR U15998 ( .A(b[1361]), .B(n11901), .Z(c[1361]) );
  XOR U15999 ( .A(n11902), .B(n11903), .Z(n11899) );
  ANDN U16000 ( .B(n11904), .A(n11905), .Z(n11902) );
  XNOR U16001 ( .A(b[1360]), .B(n11903), .Z(n11904) );
  XNOR U16002 ( .A(b[1360]), .B(n11905), .Z(c[1360]) );
  XOR U16003 ( .A(n11906), .B(n11907), .Z(n11903) );
  ANDN U16004 ( .B(n11908), .A(n11909), .Z(n11906) );
  XNOR U16005 ( .A(b[1359]), .B(n11907), .Z(n11908) );
  XNOR U16006 ( .A(b[135]), .B(n11910), .Z(c[135]) );
  XNOR U16007 ( .A(b[1359]), .B(n11909), .Z(c[1359]) );
  XOR U16008 ( .A(n11911), .B(n11912), .Z(n11907) );
  ANDN U16009 ( .B(n11913), .A(n11914), .Z(n11911) );
  XNOR U16010 ( .A(b[1358]), .B(n11912), .Z(n11913) );
  XNOR U16011 ( .A(b[1358]), .B(n11914), .Z(c[1358]) );
  XOR U16012 ( .A(n11915), .B(n11916), .Z(n11912) );
  ANDN U16013 ( .B(n11917), .A(n11918), .Z(n11915) );
  XNOR U16014 ( .A(b[1357]), .B(n11916), .Z(n11917) );
  XNOR U16015 ( .A(b[1357]), .B(n11918), .Z(c[1357]) );
  XOR U16016 ( .A(n11919), .B(n11920), .Z(n11916) );
  ANDN U16017 ( .B(n11921), .A(n11922), .Z(n11919) );
  XNOR U16018 ( .A(b[1356]), .B(n11920), .Z(n11921) );
  XNOR U16019 ( .A(b[1356]), .B(n11922), .Z(c[1356]) );
  XOR U16020 ( .A(n11923), .B(n11924), .Z(n11920) );
  ANDN U16021 ( .B(n11925), .A(n11926), .Z(n11923) );
  XNOR U16022 ( .A(b[1355]), .B(n11924), .Z(n11925) );
  XNOR U16023 ( .A(b[1355]), .B(n11926), .Z(c[1355]) );
  XOR U16024 ( .A(n11927), .B(n11928), .Z(n11924) );
  ANDN U16025 ( .B(n11929), .A(n11930), .Z(n11927) );
  XNOR U16026 ( .A(b[1354]), .B(n11928), .Z(n11929) );
  XNOR U16027 ( .A(b[1354]), .B(n11930), .Z(c[1354]) );
  XOR U16028 ( .A(n11931), .B(n11932), .Z(n11928) );
  ANDN U16029 ( .B(n11933), .A(n11934), .Z(n11931) );
  XNOR U16030 ( .A(b[1353]), .B(n11932), .Z(n11933) );
  XNOR U16031 ( .A(b[1353]), .B(n11934), .Z(c[1353]) );
  XOR U16032 ( .A(n11935), .B(n11936), .Z(n11932) );
  ANDN U16033 ( .B(n11937), .A(n11938), .Z(n11935) );
  XNOR U16034 ( .A(b[1352]), .B(n11936), .Z(n11937) );
  XNOR U16035 ( .A(b[1352]), .B(n11938), .Z(c[1352]) );
  XOR U16036 ( .A(n11939), .B(n11940), .Z(n11936) );
  ANDN U16037 ( .B(n11941), .A(n11942), .Z(n11939) );
  XNOR U16038 ( .A(b[1351]), .B(n11940), .Z(n11941) );
  XNOR U16039 ( .A(b[1351]), .B(n11942), .Z(c[1351]) );
  XOR U16040 ( .A(n11943), .B(n11944), .Z(n11940) );
  ANDN U16041 ( .B(n11945), .A(n11946), .Z(n11943) );
  XNOR U16042 ( .A(b[1350]), .B(n11944), .Z(n11945) );
  XNOR U16043 ( .A(b[1350]), .B(n11946), .Z(c[1350]) );
  XOR U16044 ( .A(n11947), .B(n11948), .Z(n11944) );
  ANDN U16045 ( .B(n11949), .A(n11950), .Z(n11947) );
  XNOR U16046 ( .A(b[1349]), .B(n11948), .Z(n11949) );
  XNOR U16047 ( .A(b[134]), .B(n11951), .Z(c[134]) );
  XNOR U16048 ( .A(b[1349]), .B(n11950), .Z(c[1349]) );
  XOR U16049 ( .A(n11952), .B(n11953), .Z(n11948) );
  ANDN U16050 ( .B(n11954), .A(n11955), .Z(n11952) );
  XNOR U16051 ( .A(b[1348]), .B(n11953), .Z(n11954) );
  XNOR U16052 ( .A(b[1348]), .B(n11955), .Z(c[1348]) );
  XOR U16053 ( .A(n11956), .B(n11957), .Z(n11953) );
  ANDN U16054 ( .B(n11958), .A(n11959), .Z(n11956) );
  XNOR U16055 ( .A(b[1347]), .B(n11957), .Z(n11958) );
  XNOR U16056 ( .A(b[1347]), .B(n11959), .Z(c[1347]) );
  XOR U16057 ( .A(n11960), .B(n11961), .Z(n11957) );
  ANDN U16058 ( .B(n11962), .A(n11963), .Z(n11960) );
  XNOR U16059 ( .A(b[1346]), .B(n11961), .Z(n11962) );
  XNOR U16060 ( .A(b[1346]), .B(n11963), .Z(c[1346]) );
  XOR U16061 ( .A(n11964), .B(n11965), .Z(n11961) );
  ANDN U16062 ( .B(n11966), .A(n11967), .Z(n11964) );
  XNOR U16063 ( .A(b[1345]), .B(n11965), .Z(n11966) );
  XNOR U16064 ( .A(b[1345]), .B(n11967), .Z(c[1345]) );
  XOR U16065 ( .A(n11968), .B(n11969), .Z(n11965) );
  ANDN U16066 ( .B(n11970), .A(n11971), .Z(n11968) );
  XNOR U16067 ( .A(b[1344]), .B(n11969), .Z(n11970) );
  XNOR U16068 ( .A(b[1344]), .B(n11971), .Z(c[1344]) );
  XOR U16069 ( .A(n11972), .B(n11973), .Z(n11969) );
  ANDN U16070 ( .B(n11974), .A(n11975), .Z(n11972) );
  XNOR U16071 ( .A(b[1343]), .B(n11973), .Z(n11974) );
  XNOR U16072 ( .A(b[1343]), .B(n11975), .Z(c[1343]) );
  XOR U16073 ( .A(n11976), .B(n11977), .Z(n11973) );
  ANDN U16074 ( .B(n11978), .A(n11979), .Z(n11976) );
  XNOR U16075 ( .A(b[1342]), .B(n11977), .Z(n11978) );
  XNOR U16076 ( .A(b[1342]), .B(n11979), .Z(c[1342]) );
  XOR U16077 ( .A(n11980), .B(n11981), .Z(n11977) );
  ANDN U16078 ( .B(n11982), .A(n11983), .Z(n11980) );
  XNOR U16079 ( .A(b[1341]), .B(n11981), .Z(n11982) );
  XNOR U16080 ( .A(b[1341]), .B(n11983), .Z(c[1341]) );
  XOR U16081 ( .A(n11984), .B(n11985), .Z(n11981) );
  ANDN U16082 ( .B(n11986), .A(n11987), .Z(n11984) );
  XNOR U16083 ( .A(b[1340]), .B(n11985), .Z(n11986) );
  XNOR U16084 ( .A(b[1340]), .B(n11987), .Z(c[1340]) );
  XOR U16085 ( .A(n11988), .B(n11989), .Z(n11985) );
  ANDN U16086 ( .B(n11990), .A(n11991), .Z(n11988) );
  XNOR U16087 ( .A(b[1339]), .B(n11989), .Z(n11990) );
  XNOR U16088 ( .A(b[133]), .B(n11992), .Z(c[133]) );
  XNOR U16089 ( .A(b[1339]), .B(n11991), .Z(c[1339]) );
  XOR U16090 ( .A(n11993), .B(n11994), .Z(n11989) );
  ANDN U16091 ( .B(n11995), .A(n11996), .Z(n11993) );
  XNOR U16092 ( .A(b[1338]), .B(n11994), .Z(n11995) );
  XNOR U16093 ( .A(b[1338]), .B(n11996), .Z(c[1338]) );
  XOR U16094 ( .A(n11997), .B(n11998), .Z(n11994) );
  ANDN U16095 ( .B(n11999), .A(n12000), .Z(n11997) );
  XNOR U16096 ( .A(b[1337]), .B(n11998), .Z(n11999) );
  XNOR U16097 ( .A(b[1337]), .B(n12000), .Z(c[1337]) );
  XOR U16098 ( .A(n12001), .B(n12002), .Z(n11998) );
  ANDN U16099 ( .B(n12003), .A(n12004), .Z(n12001) );
  XNOR U16100 ( .A(b[1336]), .B(n12002), .Z(n12003) );
  XNOR U16101 ( .A(b[1336]), .B(n12004), .Z(c[1336]) );
  XOR U16102 ( .A(n12005), .B(n12006), .Z(n12002) );
  ANDN U16103 ( .B(n12007), .A(n12008), .Z(n12005) );
  XNOR U16104 ( .A(b[1335]), .B(n12006), .Z(n12007) );
  XNOR U16105 ( .A(b[1335]), .B(n12008), .Z(c[1335]) );
  XOR U16106 ( .A(n12009), .B(n12010), .Z(n12006) );
  ANDN U16107 ( .B(n12011), .A(n12012), .Z(n12009) );
  XNOR U16108 ( .A(b[1334]), .B(n12010), .Z(n12011) );
  XNOR U16109 ( .A(b[1334]), .B(n12012), .Z(c[1334]) );
  XOR U16110 ( .A(n12013), .B(n12014), .Z(n12010) );
  ANDN U16111 ( .B(n12015), .A(n12016), .Z(n12013) );
  XNOR U16112 ( .A(b[1333]), .B(n12014), .Z(n12015) );
  XNOR U16113 ( .A(b[1333]), .B(n12016), .Z(c[1333]) );
  XOR U16114 ( .A(n12017), .B(n12018), .Z(n12014) );
  ANDN U16115 ( .B(n12019), .A(n12020), .Z(n12017) );
  XNOR U16116 ( .A(b[1332]), .B(n12018), .Z(n12019) );
  XNOR U16117 ( .A(b[1332]), .B(n12020), .Z(c[1332]) );
  XOR U16118 ( .A(n12021), .B(n12022), .Z(n12018) );
  ANDN U16119 ( .B(n12023), .A(n12024), .Z(n12021) );
  XNOR U16120 ( .A(b[1331]), .B(n12022), .Z(n12023) );
  XNOR U16121 ( .A(b[1331]), .B(n12024), .Z(c[1331]) );
  XOR U16122 ( .A(n12025), .B(n12026), .Z(n12022) );
  ANDN U16123 ( .B(n12027), .A(n12028), .Z(n12025) );
  XNOR U16124 ( .A(b[1330]), .B(n12026), .Z(n12027) );
  XNOR U16125 ( .A(b[1330]), .B(n12028), .Z(c[1330]) );
  XOR U16126 ( .A(n12029), .B(n12030), .Z(n12026) );
  ANDN U16127 ( .B(n12031), .A(n12032), .Z(n12029) );
  XNOR U16128 ( .A(b[1329]), .B(n12030), .Z(n12031) );
  XNOR U16129 ( .A(b[132]), .B(n12033), .Z(c[132]) );
  XNOR U16130 ( .A(b[1329]), .B(n12032), .Z(c[1329]) );
  XOR U16131 ( .A(n12034), .B(n12035), .Z(n12030) );
  ANDN U16132 ( .B(n12036), .A(n12037), .Z(n12034) );
  XNOR U16133 ( .A(b[1328]), .B(n12035), .Z(n12036) );
  XNOR U16134 ( .A(b[1328]), .B(n12037), .Z(c[1328]) );
  XOR U16135 ( .A(n12038), .B(n12039), .Z(n12035) );
  ANDN U16136 ( .B(n12040), .A(n12041), .Z(n12038) );
  XNOR U16137 ( .A(b[1327]), .B(n12039), .Z(n12040) );
  XNOR U16138 ( .A(b[1327]), .B(n12041), .Z(c[1327]) );
  XOR U16139 ( .A(n12042), .B(n12043), .Z(n12039) );
  ANDN U16140 ( .B(n12044), .A(n12045), .Z(n12042) );
  XNOR U16141 ( .A(b[1326]), .B(n12043), .Z(n12044) );
  XNOR U16142 ( .A(b[1326]), .B(n12045), .Z(c[1326]) );
  XOR U16143 ( .A(n12046), .B(n12047), .Z(n12043) );
  ANDN U16144 ( .B(n12048), .A(n12049), .Z(n12046) );
  XNOR U16145 ( .A(b[1325]), .B(n12047), .Z(n12048) );
  XNOR U16146 ( .A(b[1325]), .B(n12049), .Z(c[1325]) );
  XOR U16147 ( .A(n12050), .B(n12051), .Z(n12047) );
  ANDN U16148 ( .B(n12052), .A(n12053), .Z(n12050) );
  XNOR U16149 ( .A(b[1324]), .B(n12051), .Z(n12052) );
  XNOR U16150 ( .A(b[1324]), .B(n12053), .Z(c[1324]) );
  XOR U16151 ( .A(n12054), .B(n12055), .Z(n12051) );
  ANDN U16152 ( .B(n12056), .A(n12057), .Z(n12054) );
  XNOR U16153 ( .A(b[1323]), .B(n12055), .Z(n12056) );
  XNOR U16154 ( .A(b[1323]), .B(n12057), .Z(c[1323]) );
  XOR U16155 ( .A(n12058), .B(n12059), .Z(n12055) );
  ANDN U16156 ( .B(n12060), .A(n12061), .Z(n12058) );
  XNOR U16157 ( .A(b[1322]), .B(n12059), .Z(n12060) );
  XNOR U16158 ( .A(b[1322]), .B(n12061), .Z(c[1322]) );
  XOR U16159 ( .A(n12062), .B(n12063), .Z(n12059) );
  ANDN U16160 ( .B(n12064), .A(n12065), .Z(n12062) );
  XNOR U16161 ( .A(b[1321]), .B(n12063), .Z(n12064) );
  XNOR U16162 ( .A(b[1321]), .B(n12065), .Z(c[1321]) );
  XOR U16163 ( .A(n12066), .B(n12067), .Z(n12063) );
  ANDN U16164 ( .B(n12068), .A(n12069), .Z(n12066) );
  XNOR U16165 ( .A(b[1320]), .B(n12067), .Z(n12068) );
  XNOR U16166 ( .A(b[1320]), .B(n12069), .Z(c[1320]) );
  XOR U16167 ( .A(n12070), .B(n12071), .Z(n12067) );
  ANDN U16168 ( .B(n12072), .A(n12073), .Z(n12070) );
  XNOR U16169 ( .A(b[1319]), .B(n12071), .Z(n12072) );
  XNOR U16170 ( .A(b[131]), .B(n12074), .Z(c[131]) );
  XNOR U16171 ( .A(b[1319]), .B(n12073), .Z(c[1319]) );
  XOR U16172 ( .A(n12075), .B(n12076), .Z(n12071) );
  ANDN U16173 ( .B(n12077), .A(n12078), .Z(n12075) );
  XNOR U16174 ( .A(b[1318]), .B(n12076), .Z(n12077) );
  XNOR U16175 ( .A(b[1318]), .B(n12078), .Z(c[1318]) );
  XOR U16176 ( .A(n12079), .B(n12080), .Z(n12076) );
  ANDN U16177 ( .B(n12081), .A(n12082), .Z(n12079) );
  XNOR U16178 ( .A(b[1317]), .B(n12080), .Z(n12081) );
  XNOR U16179 ( .A(b[1317]), .B(n12082), .Z(c[1317]) );
  XOR U16180 ( .A(n12083), .B(n12084), .Z(n12080) );
  ANDN U16181 ( .B(n12085), .A(n12086), .Z(n12083) );
  XNOR U16182 ( .A(b[1316]), .B(n12084), .Z(n12085) );
  XNOR U16183 ( .A(b[1316]), .B(n12086), .Z(c[1316]) );
  XOR U16184 ( .A(n12087), .B(n12088), .Z(n12084) );
  ANDN U16185 ( .B(n12089), .A(n12090), .Z(n12087) );
  XNOR U16186 ( .A(b[1315]), .B(n12088), .Z(n12089) );
  XNOR U16187 ( .A(b[1315]), .B(n12090), .Z(c[1315]) );
  XOR U16188 ( .A(n12091), .B(n12092), .Z(n12088) );
  ANDN U16189 ( .B(n12093), .A(n12094), .Z(n12091) );
  XNOR U16190 ( .A(b[1314]), .B(n12092), .Z(n12093) );
  XNOR U16191 ( .A(b[1314]), .B(n12094), .Z(c[1314]) );
  XOR U16192 ( .A(n12095), .B(n12096), .Z(n12092) );
  ANDN U16193 ( .B(n12097), .A(n12098), .Z(n12095) );
  XNOR U16194 ( .A(b[1313]), .B(n12096), .Z(n12097) );
  XNOR U16195 ( .A(b[1313]), .B(n12098), .Z(c[1313]) );
  XOR U16196 ( .A(n12099), .B(n12100), .Z(n12096) );
  ANDN U16197 ( .B(n12101), .A(n12102), .Z(n12099) );
  XNOR U16198 ( .A(b[1312]), .B(n12100), .Z(n12101) );
  XNOR U16199 ( .A(b[1312]), .B(n12102), .Z(c[1312]) );
  XOR U16200 ( .A(n12103), .B(n12104), .Z(n12100) );
  ANDN U16201 ( .B(n12105), .A(n12106), .Z(n12103) );
  XNOR U16202 ( .A(b[1311]), .B(n12104), .Z(n12105) );
  XNOR U16203 ( .A(b[1311]), .B(n12106), .Z(c[1311]) );
  XOR U16204 ( .A(n12107), .B(n12108), .Z(n12104) );
  ANDN U16205 ( .B(n12109), .A(n12110), .Z(n12107) );
  XNOR U16206 ( .A(b[1310]), .B(n12108), .Z(n12109) );
  XNOR U16207 ( .A(b[1310]), .B(n12110), .Z(c[1310]) );
  XOR U16208 ( .A(n12111), .B(n12112), .Z(n12108) );
  ANDN U16209 ( .B(n12113), .A(n12114), .Z(n12111) );
  XNOR U16210 ( .A(b[1309]), .B(n12112), .Z(n12113) );
  XNOR U16211 ( .A(b[130]), .B(n12115), .Z(c[130]) );
  XNOR U16212 ( .A(b[1309]), .B(n12114), .Z(c[1309]) );
  XOR U16213 ( .A(n12116), .B(n12117), .Z(n12112) );
  ANDN U16214 ( .B(n12118), .A(n12119), .Z(n12116) );
  XNOR U16215 ( .A(b[1308]), .B(n12117), .Z(n12118) );
  XNOR U16216 ( .A(b[1308]), .B(n12119), .Z(c[1308]) );
  XOR U16217 ( .A(n12120), .B(n12121), .Z(n12117) );
  ANDN U16218 ( .B(n12122), .A(n12123), .Z(n12120) );
  XNOR U16219 ( .A(b[1307]), .B(n12121), .Z(n12122) );
  XNOR U16220 ( .A(b[1307]), .B(n12123), .Z(c[1307]) );
  XOR U16221 ( .A(n12124), .B(n12125), .Z(n12121) );
  ANDN U16222 ( .B(n12126), .A(n12127), .Z(n12124) );
  XNOR U16223 ( .A(b[1306]), .B(n12125), .Z(n12126) );
  XNOR U16224 ( .A(b[1306]), .B(n12127), .Z(c[1306]) );
  XOR U16225 ( .A(n12128), .B(n12129), .Z(n12125) );
  ANDN U16226 ( .B(n12130), .A(n12131), .Z(n12128) );
  XNOR U16227 ( .A(b[1305]), .B(n12129), .Z(n12130) );
  XNOR U16228 ( .A(b[1305]), .B(n12131), .Z(c[1305]) );
  XOR U16229 ( .A(n12132), .B(n12133), .Z(n12129) );
  ANDN U16230 ( .B(n12134), .A(n12135), .Z(n12132) );
  XNOR U16231 ( .A(b[1304]), .B(n12133), .Z(n12134) );
  XNOR U16232 ( .A(b[1304]), .B(n12135), .Z(c[1304]) );
  XOR U16233 ( .A(n12136), .B(n12137), .Z(n12133) );
  ANDN U16234 ( .B(n12138), .A(n12139), .Z(n12136) );
  XNOR U16235 ( .A(b[1303]), .B(n12137), .Z(n12138) );
  XNOR U16236 ( .A(b[1303]), .B(n12139), .Z(c[1303]) );
  XOR U16237 ( .A(n12140), .B(n12141), .Z(n12137) );
  ANDN U16238 ( .B(n12142), .A(n12143), .Z(n12140) );
  XNOR U16239 ( .A(b[1302]), .B(n12141), .Z(n12142) );
  XNOR U16240 ( .A(b[1302]), .B(n12143), .Z(c[1302]) );
  XOR U16241 ( .A(n12144), .B(n12145), .Z(n12141) );
  ANDN U16242 ( .B(n12146), .A(n12147), .Z(n12144) );
  XNOR U16243 ( .A(b[1301]), .B(n12145), .Z(n12146) );
  XNOR U16244 ( .A(b[1301]), .B(n12147), .Z(c[1301]) );
  XOR U16245 ( .A(n12148), .B(n12149), .Z(n12145) );
  ANDN U16246 ( .B(n12150), .A(n12151), .Z(n12148) );
  XNOR U16247 ( .A(b[1300]), .B(n12149), .Z(n12150) );
  XNOR U16248 ( .A(b[1300]), .B(n12151), .Z(c[1300]) );
  XOR U16249 ( .A(n12152), .B(n12153), .Z(n12149) );
  ANDN U16250 ( .B(n12154), .A(n12155), .Z(n12152) );
  XNOR U16251 ( .A(b[1299]), .B(n12153), .Z(n12154) );
  XNOR U16252 ( .A(b[12]), .B(n12156), .Z(c[12]) );
  XNOR U16253 ( .A(b[129]), .B(n12157), .Z(c[129]) );
  XNOR U16254 ( .A(b[1299]), .B(n12155), .Z(c[1299]) );
  XOR U16255 ( .A(n12158), .B(n12159), .Z(n12153) );
  ANDN U16256 ( .B(n12160), .A(n12161), .Z(n12158) );
  XNOR U16257 ( .A(b[1298]), .B(n12159), .Z(n12160) );
  XNOR U16258 ( .A(b[1298]), .B(n12161), .Z(c[1298]) );
  XOR U16259 ( .A(n12162), .B(n12163), .Z(n12159) );
  ANDN U16260 ( .B(n12164), .A(n12165), .Z(n12162) );
  XNOR U16261 ( .A(b[1297]), .B(n12163), .Z(n12164) );
  XNOR U16262 ( .A(b[1297]), .B(n12165), .Z(c[1297]) );
  XOR U16263 ( .A(n12166), .B(n12167), .Z(n12163) );
  ANDN U16264 ( .B(n12168), .A(n12169), .Z(n12166) );
  XNOR U16265 ( .A(b[1296]), .B(n12167), .Z(n12168) );
  XNOR U16266 ( .A(b[1296]), .B(n12169), .Z(c[1296]) );
  XOR U16267 ( .A(n12170), .B(n12171), .Z(n12167) );
  ANDN U16268 ( .B(n12172), .A(n12173), .Z(n12170) );
  XNOR U16269 ( .A(b[1295]), .B(n12171), .Z(n12172) );
  XNOR U16270 ( .A(b[1295]), .B(n12173), .Z(c[1295]) );
  XOR U16271 ( .A(n12174), .B(n12175), .Z(n12171) );
  ANDN U16272 ( .B(n12176), .A(n12177), .Z(n12174) );
  XNOR U16273 ( .A(b[1294]), .B(n12175), .Z(n12176) );
  XNOR U16274 ( .A(b[1294]), .B(n12177), .Z(c[1294]) );
  XOR U16275 ( .A(n12178), .B(n12179), .Z(n12175) );
  ANDN U16276 ( .B(n12180), .A(n12181), .Z(n12178) );
  XNOR U16277 ( .A(b[1293]), .B(n12179), .Z(n12180) );
  XNOR U16278 ( .A(b[1293]), .B(n12181), .Z(c[1293]) );
  XOR U16279 ( .A(n12182), .B(n12183), .Z(n12179) );
  ANDN U16280 ( .B(n12184), .A(n12185), .Z(n12182) );
  XNOR U16281 ( .A(b[1292]), .B(n12183), .Z(n12184) );
  XNOR U16282 ( .A(b[1292]), .B(n12185), .Z(c[1292]) );
  XOR U16283 ( .A(n12186), .B(n12187), .Z(n12183) );
  ANDN U16284 ( .B(n12188), .A(n12189), .Z(n12186) );
  XNOR U16285 ( .A(b[1291]), .B(n12187), .Z(n12188) );
  XNOR U16286 ( .A(b[1291]), .B(n12189), .Z(c[1291]) );
  XOR U16287 ( .A(n12190), .B(n12191), .Z(n12187) );
  ANDN U16288 ( .B(n12192), .A(n12193), .Z(n12190) );
  XNOR U16289 ( .A(b[1290]), .B(n12191), .Z(n12192) );
  XNOR U16290 ( .A(b[1290]), .B(n12193), .Z(c[1290]) );
  XOR U16291 ( .A(n12194), .B(n12195), .Z(n12191) );
  ANDN U16292 ( .B(n12196), .A(n12197), .Z(n12194) );
  XNOR U16293 ( .A(b[1289]), .B(n12195), .Z(n12196) );
  XNOR U16294 ( .A(b[128]), .B(n12198), .Z(c[128]) );
  XNOR U16295 ( .A(b[1289]), .B(n12197), .Z(c[1289]) );
  XOR U16296 ( .A(n12199), .B(n12200), .Z(n12195) );
  ANDN U16297 ( .B(n12201), .A(n12202), .Z(n12199) );
  XNOR U16298 ( .A(b[1288]), .B(n12200), .Z(n12201) );
  XNOR U16299 ( .A(b[1288]), .B(n12202), .Z(c[1288]) );
  XOR U16300 ( .A(n12203), .B(n12204), .Z(n12200) );
  ANDN U16301 ( .B(n12205), .A(n12206), .Z(n12203) );
  XNOR U16302 ( .A(b[1287]), .B(n12204), .Z(n12205) );
  XNOR U16303 ( .A(b[1287]), .B(n12206), .Z(c[1287]) );
  XOR U16304 ( .A(n12207), .B(n12208), .Z(n12204) );
  ANDN U16305 ( .B(n12209), .A(n12210), .Z(n12207) );
  XNOR U16306 ( .A(b[1286]), .B(n12208), .Z(n12209) );
  XNOR U16307 ( .A(b[1286]), .B(n12210), .Z(c[1286]) );
  XOR U16308 ( .A(n12211), .B(n12212), .Z(n12208) );
  ANDN U16309 ( .B(n12213), .A(n12214), .Z(n12211) );
  XNOR U16310 ( .A(b[1285]), .B(n12212), .Z(n12213) );
  XNOR U16311 ( .A(b[1285]), .B(n12214), .Z(c[1285]) );
  XOR U16312 ( .A(n12215), .B(n12216), .Z(n12212) );
  ANDN U16313 ( .B(n12217), .A(n12218), .Z(n12215) );
  XNOR U16314 ( .A(b[1284]), .B(n12216), .Z(n12217) );
  XNOR U16315 ( .A(b[1284]), .B(n12218), .Z(c[1284]) );
  XOR U16316 ( .A(n12219), .B(n12220), .Z(n12216) );
  ANDN U16317 ( .B(n12221), .A(n12222), .Z(n12219) );
  XNOR U16318 ( .A(b[1283]), .B(n12220), .Z(n12221) );
  XNOR U16319 ( .A(b[1283]), .B(n12222), .Z(c[1283]) );
  XOR U16320 ( .A(n12223), .B(n12224), .Z(n12220) );
  ANDN U16321 ( .B(n12225), .A(n12226), .Z(n12223) );
  XNOR U16322 ( .A(b[1282]), .B(n12224), .Z(n12225) );
  XNOR U16323 ( .A(b[1282]), .B(n12226), .Z(c[1282]) );
  XOR U16324 ( .A(n12227), .B(n12228), .Z(n12224) );
  ANDN U16325 ( .B(n12229), .A(n12230), .Z(n12227) );
  XNOR U16326 ( .A(b[1281]), .B(n12228), .Z(n12229) );
  XNOR U16327 ( .A(b[1281]), .B(n12230), .Z(c[1281]) );
  XOR U16328 ( .A(n12231), .B(n12232), .Z(n12228) );
  ANDN U16329 ( .B(n12233), .A(n12234), .Z(n12231) );
  XNOR U16330 ( .A(b[1280]), .B(n12232), .Z(n12233) );
  XNOR U16331 ( .A(b[1280]), .B(n12234), .Z(c[1280]) );
  XOR U16332 ( .A(n12235), .B(n12236), .Z(n12232) );
  ANDN U16333 ( .B(n12237), .A(n12238), .Z(n12235) );
  XNOR U16334 ( .A(b[1279]), .B(n12236), .Z(n12237) );
  XNOR U16335 ( .A(b[127]), .B(n12239), .Z(c[127]) );
  XNOR U16336 ( .A(b[1279]), .B(n12238), .Z(c[1279]) );
  XOR U16337 ( .A(n12240), .B(n12241), .Z(n12236) );
  ANDN U16338 ( .B(n12242), .A(n12243), .Z(n12240) );
  XNOR U16339 ( .A(b[1278]), .B(n12241), .Z(n12242) );
  XNOR U16340 ( .A(b[1278]), .B(n12243), .Z(c[1278]) );
  XOR U16341 ( .A(n12244), .B(n12245), .Z(n12241) );
  ANDN U16342 ( .B(n12246), .A(n12247), .Z(n12244) );
  XNOR U16343 ( .A(b[1277]), .B(n12245), .Z(n12246) );
  XNOR U16344 ( .A(b[1277]), .B(n12247), .Z(c[1277]) );
  XOR U16345 ( .A(n12248), .B(n12249), .Z(n12245) );
  ANDN U16346 ( .B(n12250), .A(n12251), .Z(n12248) );
  XNOR U16347 ( .A(b[1276]), .B(n12249), .Z(n12250) );
  XNOR U16348 ( .A(b[1276]), .B(n12251), .Z(c[1276]) );
  XOR U16349 ( .A(n12252), .B(n12253), .Z(n12249) );
  ANDN U16350 ( .B(n12254), .A(n12255), .Z(n12252) );
  XNOR U16351 ( .A(b[1275]), .B(n12253), .Z(n12254) );
  XNOR U16352 ( .A(b[1275]), .B(n12255), .Z(c[1275]) );
  XOR U16353 ( .A(n12256), .B(n12257), .Z(n12253) );
  ANDN U16354 ( .B(n12258), .A(n12259), .Z(n12256) );
  XNOR U16355 ( .A(b[1274]), .B(n12257), .Z(n12258) );
  XNOR U16356 ( .A(b[1274]), .B(n12259), .Z(c[1274]) );
  XOR U16357 ( .A(n12260), .B(n12261), .Z(n12257) );
  ANDN U16358 ( .B(n12262), .A(n12263), .Z(n12260) );
  XNOR U16359 ( .A(b[1273]), .B(n12261), .Z(n12262) );
  XNOR U16360 ( .A(b[1273]), .B(n12263), .Z(c[1273]) );
  XOR U16361 ( .A(n12264), .B(n12265), .Z(n12261) );
  ANDN U16362 ( .B(n12266), .A(n12267), .Z(n12264) );
  XNOR U16363 ( .A(b[1272]), .B(n12265), .Z(n12266) );
  XNOR U16364 ( .A(b[1272]), .B(n12267), .Z(c[1272]) );
  XOR U16365 ( .A(n12268), .B(n12269), .Z(n12265) );
  ANDN U16366 ( .B(n12270), .A(n12271), .Z(n12268) );
  XNOR U16367 ( .A(b[1271]), .B(n12269), .Z(n12270) );
  XNOR U16368 ( .A(b[1271]), .B(n12271), .Z(c[1271]) );
  XOR U16369 ( .A(n12272), .B(n12273), .Z(n12269) );
  ANDN U16370 ( .B(n12274), .A(n12275), .Z(n12272) );
  XNOR U16371 ( .A(b[1270]), .B(n12273), .Z(n12274) );
  XNOR U16372 ( .A(b[1270]), .B(n12275), .Z(c[1270]) );
  XOR U16373 ( .A(n12276), .B(n12277), .Z(n12273) );
  ANDN U16374 ( .B(n12278), .A(n12279), .Z(n12276) );
  XNOR U16375 ( .A(b[1269]), .B(n12277), .Z(n12278) );
  XNOR U16376 ( .A(b[126]), .B(n12280), .Z(c[126]) );
  XNOR U16377 ( .A(b[1269]), .B(n12279), .Z(c[1269]) );
  XOR U16378 ( .A(n12281), .B(n12282), .Z(n12277) );
  ANDN U16379 ( .B(n12283), .A(n12284), .Z(n12281) );
  XNOR U16380 ( .A(b[1268]), .B(n12282), .Z(n12283) );
  XNOR U16381 ( .A(b[1268]), .B(n12284), .Z(c[1268]) );
  XOR U16382 ( .A(n12285), .B(n12286), .Z(n12282) );
  ANDN U16383 ( .B(n12287), .A(n12288), .Z(n12285) );
  XNOR U16384 ( .A(b[1267]), .B(n12286), .Z(n12287) );
  XNOR U16385 ( .A(b[1267]), .B(n12288), .Z(c[1267]) );
  XOR U16386 ( .A(n12289), .B(n12290), .Z(n12286) );
  ANDN U16387 ( .B(n12291), .A(n12292), .Z(n12289) );
  XNOR U16388 ( .A(b[1266]), .B(n12290), .Z(n12291) );
  XNOR U16389 ( .A(b[1266]), .B(n12292), .Z(c[1266]) );
  XOR U16390 ( .A(n12293), .B(n12294), .Z(n12290) );
  ANDN U16391 ( .B(n12295), .A(n12296), .Z(n12293) );
  XNOR U16392 ( .A(b[1265]), .B(n12294), .Z(n12295) );
  XNOR U16393 ( .A(b[1265]), .B(n12296), .Z(c[1265]) );
  XOR U16394 ( .A(n12297), .B(n12298), .Z(n12294) );
  ANDN U16395 ( .B(n12299), .A(n12300), .Z(n12297) );
  XNOR U16396 ( .A(b[1264]), .B(n12298), .Z(n12299) );
  XNOR U16397 ( .A(b[1264]), .B(n12300), .Z(c[1264]) );
  XOR U16398 ( .A(n12301), .B(n12302), .Z(n12298) );
  ANDN U16399 ( .B(n12303), .A(n12304), .Z(n12301) );
  XNOR U16400 ( .A(b[1263]), .B(n12302), .Z(n12303) );
  XNOR U16401 ( .A(b[1263]), .B(n12304), .Z(c[1263]) );
  XOR U16402 ( .A(n12305), .B(n12306), .Z(n12302) );
  ANDN U16403 ( .B(n12307), .A(n12308), .Z(n12305) );
  XNOR U16404 ( .A(b[1262]), .B(n12306), .Z(n12307) );
  XNOR U16405 ( .A(b[1262]), .B(n12308), .Z(c[1262]) );
  XOR U16406 ( .A(n12309), .B(n12310), .Z(n12306) );
  ANDN U16407 ( .B(n12311), .A(n12312), .Z(n12309) );
  XNOR U16408 ( .A(b[1261]), .B(n12310), .Z(n12311) );
  XNOR U16409 ( .A(b[1261]), .B(n12312), .Z(c[1261]) );
  XOR U16410 ( .A(n12313), .B(n12314), .Z(n12310) );
  ANDN U16411 ( .B(n12315), .A(n12316), .Z(n12313) );
  XNOR U16412 ( .A(b[1260]), .B(n12314), .Z(n12315) );
  XNOR U16413 ( .A(b[1260]), .B(n12316), .Z(c[1260]) );
  XOR U16414 ( .A(n12317), .B(n12318), .Z(n12314) );
  ANDN U16415 ( .B(n12319), .A(n12320), .Z(n12317) );
  XNOR U16416 ( .A(b[1259]), .B(n12318), .Z(n12319) );
  XNOR U16417 ( .A(b[125]), .B(n12321), .Z(c[125]) );
  XNOR U16418 ( .A(b[1259]), .B(n12320), .Z(c[1259]) );
  XOR U16419 ( .A(n12322), .B(n12323), .Z(n12318) );
  ANDN U16420 ( .B(n12324), .A(n12325), .Z(n12322) );
  XNOR U16421 ( .A(b[1258]), .B(n12323), .Z(n12324) );
  XNOR U16422 ( .A(b[1258]), .B(n12325), .Z(c[1258]) );
  XOR U16423 ( .A(n12326), .B(n12327), .Z(n12323) );
  ANDN U16424 ( .B(n12328), .A(n12329), .Z(n12326) );
  XNOR U16425 ( .A(b[1257]), .B(n12327), .Z(n12328) );
  XNOR U16426 ( .A(b[1257]), .B(n12329), .Z(c[1257]) );
  XOR U16427 ( .A(n12330), .B(n12331), .Z(n12327) );
  ANDN U16428 ( .B(n12332), .A(n12333), .Z(n12330) );
  XNOR U16429 ( .A(b[1256]), .B(n12331), .Z(n12332) );
  XNOR U16430 ( .A(b[1256]), .B(n12333), .Z(c[1256]) );
  XOR U16431 ( .A(n12334), .B(n12335), .Z(n12331) );
  ANDN U16432 ( .B(n12336), .A(n12337), .Z(n12334) );
  XNOR U16433 ( .A(b[1255]), .B(n12335), .Z(n12336) );
  XNOR U16434 ( .A(b[1255]), .B(n12337), .Z(c[1255]) );
  XOR U16435 ( .A(n12338), .B(n12339), .Z(n12335) );
  ANDN U16436 ( .B(n12340), .A(n12341), .Z(n12338) );
  XNOR U16437 ( .A(b[1254]), .B(n12339), .Z(n12340) );
  XNOR U16438 ( .A(b[1254]), .B(n12341), .Z(c[1254]) );
  XOR U16439 ( .A(n12342), .B(n12343), .Z(n12339) );
  ANDN U16440 ( .B(n12344), .A(n12345), .Z(n12342) );
  XNOR U16441 ( .A(b[1253]), .B(n12343), .Z(n12344) );
  XNOR U16442 ( .A(b[1253]), .B(n12345), .Z(c[1253]) );
  XOR U16443 ( .A(n12346), .B(n12347), .Z(n12343) );
  ANDN U16444 ( .B(n12348), .A(n12349), .Z(n12346) );
  XNOR U16445 ( .A(b[1252]), .B(n12347), .Z(n12348) );
  XNOR U16446 ( .A(b[1252]), .B(n12349), .Z(c[1252]) );
  XOR U16447 ( .A(n12350), .B(n12351), .Z(n12347) );
  ANDN U16448 ( .B(n12352), .A(n12353), .Z(n12350) );
  XNOR U16449 ( .A(b[1251]), .B(n12351), .Z(n12352) );
  XNOR U16450 ( .A(b[1251]), .B(n12353), .Z(c[1251]) );
  XOR U16451 ( .A(n12354), .B(n12355), .Z(n12351) );
  ANDN U16452 ( .B(n12356), .A(n12357), .Z(n12354) );
  XNOR U16453 ( .A(b[1250]), .B(n12355), .Z(n12356) );
  XNOR U16454 ( .A(b[1250]), .B(n12357), .Z(c[1250]) );
  XOR U16455 ( .A(n12358), .B(n12359), .Z(n12355) );
  ANDN U16456 ( .B(n12360), .A(n12361), .Z(n12358) );
  XNOR U16457 ( .A(b[1249]), .B(n12359), .Z(n12360) );
  XNOR U16458 ( .A(b[124]), .B(n12362), .Z(c[124]) );
  XNOR U16459 ( .A(b[1249]), .B(n12361), .Z(c[1249]) );
  XOR U16460 ( .A(n12363), .B(n12364), .Z(n12359) );
  ANDN U16461 ( .B(n12365), .A(n12366), .Z(n12363) );
  XNOR U16462 ( .A(b[1248]), .B(n12364), .Z(n12365) );
  XNOR U16463 ( .A(b[1248]), .B(n12366), .Z(c[1248]) );
  XOR U16464 ( .A(n12367), .B(n12368), .Z(n12364) );
  ANDN U16465 ( .B(n12369), .A(n12370), .Z(n12367) );
  XNOR U16466 ( .A(b[1247]), .B(n12368), .Z(n12369) );
  XNOR U16467 ( .A(b[1247]), .B(n12370), .Z(c[1247]) );
  XOR U16468 ( .A(n12371), .B(n12372), .Z(n12368) );
  ANDN U16469 ( .B(n12373), .A(n12374), .Z(n12371) );
  XNOR U16470 ( .A(b[1246]), .B(n12372), .Z(n12373) );
  XNOR U16471 ( .A(b[1246]), .B(n12374), .Z(c[1246]) );
  XOR U16472 ( .A(n12375), .B(n12376), .Z(n12372) );
  ANDN U16473 ( .B(n12377), .A(n12378), .Z(n12375) );
  XNOR U16474 ( .A(b[1245]), .B(n12376), .Z(n12377) );
  XNOR U16475 ( .A(b[1245]), .B(n12378), .Z(c[1245]) );
  XOR U16476 ( .A(n12379), .B(n12380), .Z(n12376) );
  ANDN U16477 ( .B(n12381), .A(n12382), .Z(n12379) );
  XNOR U16478 ( .A(b[1244]), .B(n12380), .Z(n12381) );
  XNOR U16479 ( .A(b[1244]), .B(n12382), .Z(c[1244]) );
  XOR U16480 ( .A(n12383), .B(n12384), .Z(n12380) );
  ANDN U16481 ( .B(n12385), .A(n12386), .Z(n12383) );
  XNOR U16482 ( .A(b[1243]), .B(n12384), .Z(n12385) );
  XNOR U16483 ( .A(b[1243]), .B(n12386), .Z(c[1243]) );
  XOR U16484 ( .A(n12387), .B(n12388), .Z(n12384) );
  ANDN U16485 ( .B(n12389), .A(n12390), .Z(n12387) );
  XNOR U16486 ( .A(b[1242]), .B(n12388), .Z(n12389) );
  XNOR U16487 ( .A(b[1242]), .B(n12390), .Z(c[1242]) );
  XOR U16488 ( .A(n12391), .B(n12392), .Z(n12388) );
  ANDN U16489 ( .B(n12393), .A(n12394), .Z(n12391) );
  XNOR U16490 ( .A(b[1241]), .B(n12392), .Z(n12393) );
  XNOR U16491 ( .A(b[1241]), .B(n12394), .Z(c[1241]) );
  XOR U16492 ( .A(n12395), .B(n12396), .Z(n12392) );
  ANDN U16493 ( .B(n12397), .A(n12398), .Z(n12395) );
  XNOR U16494 ( .A(b[1240]), .B(n12396), .Z(n12397) );
  XNOR U16495 ( .A(b[1240]), .B(n12398), .Z(c[1240]) );
  XOR U16496 ( .A(n12399), .B(n12400), .Z(n12396) );
  ANDN U16497 ( .B(n12401), .A(n12402), .Z(n12399) );
  XNOR U16498 ( .A(b[1239]), .B(n12400), .Z(n12401) );
  XNOR U16499 ( .A(b[123]), .B(n12403), .Z(c[123]) );
  XNOR U16500 ( .A(b[1239]), .B(n12402), .Z(c[1239]) );
  XOR U16501 ( .A(n12404), .B(n12405), .Z(n12400) );
  ANDN U16502 ( .B(n12406), .A(n12407), .Z(n12404) );
  XNOR U16503 ( .A(b[1238]), .B(n12405), .Z(n12406) );
  XNOR U16504 ( .A(b[1238]), .B(n12407), .Z(c[1238]) );
  XOR U16505 ( .A(n12408), .B(n12409), .Z(n12405) );
  ANDN U16506 ( .B(n12410), .A(n12411), .Z(n12408) );
  XNOR U16507 ( .A(b[1237]), .B(n12409), .Z(n12410) );
  XNOR U16508 ( .A(b[1237]), .B(n12411), .Z(c[1237]) );
  XOR U16509 ( .A(n12412), .B(n12413), .Z(n12409) );
  ANDN U16510 ( .B(n12414), .A(n12415), .Z(n12412) );
  XNOR U16511 ( .A(b[1236]), .B(n12413), .Z(n12414) );
  XNOR U16512 ( .A(b[1236]), .B(n12415), .Z(c[1236]) );
  XOR U16513 ( .A(n12416), .B(n12417), .Z(n12413) );
  ANDN U16514 ( .B(n12418), .A(n12419), .Z(n12416) );
  XNOR U16515 ( .A(b[1235]), .B(n12417), .Z(n12418) );
  XNOR U16516 ( .A(b[1235]), .B(n12419), .Z(c[1235]) );
  XOR U16517 ( .A(n12420), .B(n12421), .Z(n12417) );
  ANDN U16518 ( .B(n12422), .A(n12423), .Z(n12420) );
  XNOR U16519 ( .A(b[1234]), .B(n12421), .Z(n12422) );
  XNOR U16520 ( .A(b[1234]), .B(n12423), .Z(c[1234]) );
  XOR U16521 ( .A(n12424), .B(n12425), .Z(n12421) );
  ANDN U16522 ( .B(n12426), .A(n12427), .Z(n12424) );
  XNOR U16523 ( .A(b[1233]), .B(n12425), .Z(n12426) );
  XNOR U16524 ( .A(b[1233]), .B(n12427), .Z(c[1233]) );
  XOR U16525 ( .A(n12428), .B(n12429), .Z(n12425) );
  ANDN U16526 ( .B(n12430), .A(n12431), .Z(n12428) );
  XNOR U16527 ( .A(b[1232]), .B(n12429), .Z(n12430) );
  XNOR U16528 ( .A(b[1232]), .B(n12431), .Z(c[1232]) );
  XOR U16529 ( .A(n12432), .B(n12433), .Z(n12429) );
  ANDN U16530 ( .B(n12434), .A(n12435), .Z(n12432) );
  XNOR U16531 ( .A(b[1231]), .B(n12433), .Z(n12434) );
  XNOR U16532 ( .A(b[1231]), .B(n12435), .Z(c[1231]) );
  XOR U16533 ( .A(n12436), .B(n12437), .Z(n12433) );
  ANDN U16534 ( .B(n12438), .A(n12439), .Z(n12436) );
  XNOR U16535 ( .A(b[1230]), .B(n12437), .Z(n12438) );
  XNOR U16536 ( .A(b[1230]), .B(n12439), .Z(c[1230]) );
  XOR U16537 ( .A(n12440), .B(n12441), .Z(n12437) );
  ANDN U16538 ( .B(n12442), .A(n12443), .Z(n12440) );
  XNOR U16539 ( .A(b[1229]), .B(n12441), .Z(n12442) );
  XNOR U16540 ( .A(b[122]), .B(n12444), .Z(c[122]) );
  XNOR U16541 ( .A(b[1229]), .B(n12443), .Z(c[1229]) );
  XOR U16542 ( .A(n12445), .B(n12446), .Z(n12441) );
  ANDN U16543 ( .B(n12447), .A(n12448), .Z(n12445) );
  XNOR U16544 ( .A(b[1228]), .B(n12446), .Z(n12447) );
  XNOR U16545 ( .A(b[1228]), .B(n12448), .Z(c[1228]) );
  XOR U16546 ( .A(n12449), .B(n12450), .Z(n12446) );
  ANDN U16547 ( .B(n12451), .A(n12452), .Z(n12449) );
  XNOR U16548 ( .A(b[1227]), .B(n12450), .Z(n12451) );
  XNOR U16549 ( .A(b[1227]), .B(n12452), .Z(c[1227]) );
  XOR U16550 ( .A(n12453), .B(n12454), .Z(n12450) );
  ANDN U16551 ( .B(n12455), .A(n12456), .Z(n12453) );
  XNOR U16552 ( .A(b[1226]), .B(n12454), .Z(n12455) );
  XNOR U16553 ( .A(b[1226]), .B(n12456), .Z(c[1226]) );
  XOR U16554 ( .A(n12457), .B(n12458), .Z(n12454) );
  ANDN U16555 ( .B(n12459), .A(n12460), .Z(n12457) );
  XNOR U16556 ( .A(b[1225]), .B(n12458), .Z(n12459) );
  XNOR U16557 ( .A(b[1225]), .B(n12460), .Z(c[1225]) );
  XOR U16558 ( .A(n12461), .B(n12462), .Z(n12458) );
  ANDN U16559 ( .B(n12463), .A(n12464), .Z(n12461) );
  XNOR U16560 ( .A(b[1224]), .B(n12462), .Z(n12463) );
  XNOR U16561 ( .A(b[1224]), .B(n12464), .Z(c[1224]) );
  XOR U16562 ( .A(n12465), .B(n12466), .Z(n12462) );
  ANDN U16563 ( .B(n12467), .A(n12468), .Z(n12465) );
  XNOR U16564 ( .A(b[1223]), .B(n12466), .Z(n12467) );
  XNOR U16565 ( .A(b[1223]), .B(n12468), .Z(c[1223]) );
  XOR U16566 ( .A(n12469), .B(n12470), .Z(n12466) );
  ANDN U16567 ( .B(n12471), .A(n12472), .Z(n12469) );
  XNOR U16568 ( .A(b[1222]), .B(n12470), .Z(n12471) );
  XNOR U16569 ( .A(b[1222]), .B(n12472), .Z(c[1222]) );
  XOR U16570 ( .A(n12473), .B(n12474), .Z(n12470) );
  ANDN U16571 ( .B(n12475), .A(n12476), .Z(n12473) );
  XNOR U16572 ( .A(b[1221]), .B(n12474), .Z(n12475) );
  XNOR U16573 ( .A(b[1221]), .B(n12476), .Z(c[1221]) );
  XOR U16574 ( .A(n12477), .B(n12478), .Z(n12474) );
  ANDN U16575 ( .B(n12479), .A(n12480), .Z(n12477) );
  XNOR U16576 ( .A(b[1220]), .B(n12478), .Z(n12479) );
  XNOR U16577 ( .A(b[1220]), .B(n12480), .Z(c[1220]) );
  XOR U16578 ( .A(n12481), .B(n12482), .Z(n12478) );
  ANDN U16579 ( .B(n12483), .A(n12484), .Z(n12481) );
  XNOR U16580 ( .A(b[1219]), .B(n12482), .Z(n12483) );
  XNOR U16581 ( .A(b[121]), .B(n12485), .Z(c[121]) );
  XNOR U16582 ( .A(b[1219]), .B(n12484), .Z(c[1219]) );
  XOR U16583 ( .A(n12486), .B(n12487), .Z(n12482) );
  ANDN U16584 ( .B(n12488), .A(n12489), .Z(n12486) );
  XNOR U16585 ( .A(b[1218]), .B(n12487), .Z(n12488) );
  XNOR U16586 ( .A(b[1218]), .B(n12489), .Z(c[1218]) );
  XOR U16587 ( .A(n12490), .B(n12491), .Z(n12487) );
  ANDN U16588 ( .B(n12492), .A(n12493), .Z(n12490) );
  XNOR U16589 ( .A(b[1217]), .B(n12491), .Z(n12492) );
  XNOR U16590 ( .A(b[1217]), .B(n12493), .Z(c[1217]) );
  XOR U16591 ( .A(n12494), .B(n12495), .Z(n12491) );
  ANDN U16592 ( .B(n12496), .A(n12497), .Z(n12494) );
  XNOR U16593 ( .A(b[1216]), .B(n12495), .Z(n12496) );
  XNOR U16594 ( .A(b[1216]), .B(n12497), .Z(c[1216]) );
  XOR U16595 ( .A(n12498), .B(n12499), .Z(n12495) );
  ANDN U16596 ( .B(n12500), .A(n12501), .Z(n12498) );
  XNOR U16597 ( .A(b[1215]), .B(n12499), .Z(n12500) );
  XNOR U16598 ( .A(b[1215]), .B(n12501), .Z(c[1215]) );
  XOR U16599 ( .A(n12502), .B(n12503), .Z(n12499) );
  ANDN U16600 ( .B(n12504), .A(n12505), .Z(n12502) );
  XNOR U16601 ( .A(b[1214]), .B(n12503), .Z(n12504) );
  XNOR U16602 ( .A(b[1214]), .B(n12505), .Z(c[1214]) );
  XOR U16603 ( .A(n12506), .B(n12507), .Z(n12503) );
  ANDN U16604 ( .B(n12508), .A(n12509), .Z(n12506) );
  XNOR U16605 ( .A(b[1213]), .B(n12507), .Z(n12508) );
  XNOR U16606 ( .A(b[1213]), .B(n12509), .Z(c[1213]) );
  XOR U16607 ( .A(n12510), .B(n12511), .Z(n12507) );
  ANDN U16608 ( .B(n12512), .A(n12513), .Z(n12510) );
  XNOR U16609 ( .A(b[1212]), .B(n12511), .Z(n12512) );
  XNOR U16610 ( .A(b[1212]), .B(n12513), .Z(c[1212]) );
  XOR U16611 ( .A(n12514), .B(n12515), .Z(n12511) );
  ANDN U16612 ( .B(n12516), .A(n12517), .Z(n12514) );
  XNOR U16613 ( .A(b[1211]), .B(n12515), .Z(n12516) );
  XNOR U16614 ( .A(b[1211]), .B(n12517), .Z(c[1211]) );
  XOR U16615 ( .A(n12518), .B(n12519), .Z(n12515) );
  ANDN U16616 ( .B(n12520), .A(n12521), .Z(n12518) );
  XNOR U16617 ( .A(b[1210]), .B(n12519), .Z(n12520) );
  XNOR U16618 ( .A(b[1210]), .B(n12521), .Z(c[1210]) );
  XOR U16619 ( .A(n12522), .B(n12523), .Z(n12519) );
  ANDN U16620 ( .B(n12524), .A(n12525), .Z(n12522) );
  XNOR U16621 ( .A(b[1209]), .B(n12523), .Z(n12524) );
  XNOR U16622 ( .A(b[120]), .B(n12526), .Z(c[120]) );
  XNOR U16623 ( .A(b[1209]), .B(n12525), .Z(c[1209]) );
  XOR U16624 ( .A(n12527), .B(n12528), .Z(n12523) );
  ANDN U16625 ( .B(n12529), .A(n12530), .Z(n12527) );
  XNOR U16626 ( .A(b[1208]), .B(n12528), .Z(n12529) );
  XNOR U16627 ( .A(b[1208]), .B(n12530), .Z(c[1208]) );
  XOR U16628 ( .A(n12531), .B(n12532), .Z(n12528) );
  ANDN U16629 ( .B(n12533), .A(n12534), .Z(n12531) );
  XNOR U16630 ( .A(b[1207]), .B(n12532), .Z(n12533) );
  XNOR U16631 ( .A(b[1207]), .B(n12534), .Z(c[1207]) );
  XOR U16632 ( .A(n12535), .B(n12536), .Z(n12532) );
  ANDN U16633 ( .B(n12537), .A(n12538), .Z(n12535) );
  XNOR U16634 ( .A(b[1206]), .B(n12536), .Z(n12537) );
  XNOR U16635 ( .A(b[1206]), .B(n12538), .Z(c[1206]) );
  XOR U16636 ( .A(n12539), .B(n12540), .Z(n12536) );
  ANDN U16637 ( .B(n12541), .A(n12542), .Z(n12539) );
  XNOR U16638 ( .A(b[1205]), .B(n12540), .Z(n12541) );
  XNOR U16639 ( .A(b[1205]), .B(n12542), .Z(c[1205]) );
  XOR U16640 ( .A(n12543), .B(n12544), .Z(n12540) );
  ANDN U16641 ( .B(n12545), .A(n12546), .Z(n12543) );
  XNOR U16642 ( .A(b[1204]), .B(n12544), .Z(n12545) );
  XNOR U16643 ( .A(b[1204]), .B(n12546), .Z(c[1204]) );
  XOR U16644 ( .A(n12547), .B(n12548), .Z(n12544) );
  ANDN U16645 ( .B(n12549), .A(n12550), .Z(n12547) );
  XNOR U16646 ( .A(b[1203]), .B(n12548), .Z(n12549) );
  XNOR U16647 ( .A(b[1203]), .B(n12550), .Z(c[1203]) );
  XOR U16648 ( .A(n12551), .B(n12552), .Z(n12548) );
  ANDN U16649 ( .B(n12553), .A(n12554), .Z(n12551) );
  XNOR U16650 ( .A(b[1202]), .B(n12552), .Z(n12553) );
  XNOR U16651 ( .A(b[1202]), .B(n12554), .Z(c[1202]) );
  XOR U16652 ( .A(n12555), .B(n12556), .Z(n12552) );
  ANDN U16653 ( .B(n12557), .A(n12558), .Z(n12555) );
  XNOR U16654 ( .A(b[1201]), .B(n12556), .Z(n12557) );
  XNOR U16655 ( .A(b[1201]), .B(n12558), .Z(c[1201]) );
  XOR U16656 ( .A(n12559), .B(n12560), .Z(n12556) );
  ANDN U16657 ( .B(n12561), .A(n12562), .Z(n12559) );
  XNOR U16658 ( .A(b[1200]), .B(n12560), .Z(n12561) );
  XNOR U16659 ( .A(b[1200]), .B(n12562), .Z(c[1200]) );
  XOR U16660 ( .A(n12563), .B(n12564), .Z(n12560) );
  ANDN U16661 ( .B(n12565), .A(n12566), .Z(n12563) );
  XNOR U16662 ( .A(b[1199]), .B(n12564), .Z(n12565) );
  XNOR U16663 ( .A(b[11]), .B(n12567), .Z(c[11]) );
  XNOR U16664 ( .A(b[119]), .B(n12568), .Z(c[119]) );
  XNOR U16665 ( .A(b[1199]), .B(n12566), .Z(c[1199]) );
  XOR U16666 ( .A(n12569), .B(n12570), .Z(n12564) );
  ANDN U16667 ( .B(n12571), .A(n12572), .Z(n12569) );
  XNOR U16668 ( .A(b[1198]), .B(n12570), .Z(n12571) );
  XNOR U16669 ( .A(b[1198]), .B(n12572), .Z(c[1198]) );
  XOR U16670 ( .A(n12573), .B(n12574), .Z(n12570) );
  ANDN U16671 ( .B(n12575), .A(n12576), .Z(n12573) );
  XNOR U16672 ( .A(b[1197]), .B(n12574), .Z(n12575) );
  XNOR U16673 ( .A(b[1197]), .B(n12576), .Z(c[1197]) );
  XOR U16674 ( .A(n12577), .B(n12578), .Z(n12574) );
  ANDN U16675 ( .B(n12579), .A(n12580), .Z(n12577) );
  XNOR U16676 ( .A(b[1196]), .B(n12578), .Z(n12579) );
  XNOR U16677 ( .A(b[1196]), .B(n12580), .Z(c[1196]) );
  XOR U16678 ( .A(n12581), .B(n12582), .Z(n12578) );
  ANDN U16679 ( .B(n12583), .A(n12584), .Z(n12581) );
  XNOR U16680 ( .A(b[1195]), .B(n12582), .Z(n12583) );
  XNOR U16681 ( .A(b[1195]), .B(n12584), .Z(c[1195]) );
  XOR U16682 ( .A(n12585), .B(n12586), .Z(n12582) );
  ANDN U16683 ( .B(n12587), .A(n12588), .Z(n12585) );
  XNOR U16684 ( .A(b[1194]), .B(n12586), .Z(n12587) );
  XNOR U16685 ( .A(b[1194]), .B(n12588), .Z(c[1194]) );
  XOR U16686 ( .A(n12589), .B(n12590), .Z(n12586) );
  ANDN U16687 ( .B(n12591), .A(n12592), .Z(n12589) );
  XNOR U16688 ( .A(b[1193]), .B(n12590), .Z(n12591) );
  XNOR U16689 ( .A(b[1193]), .B(n12592), .Z(c[1193]) );
  XOR U16690 ( .A(n12593), .B(n12594), .Z(n12590) );
  ANDN U16691 ( .B(n12595), .A(n12596), .Z(n12593) );
  XNOR U16692 ( .A(b[1192]), .B(n12594), .Z(n12595) );
  XNOR U16693 ( .A(b[1192]), .B(n12596), .Z(c[1192]) );
  XOR U16694 ( .A(n12597), .B(n12598), .Z(n12594) );
  ANDN U16695 ( .B(n12599), .A(n12600), .Z(n12597) );
  XNOR U16696 ( .A(b[1191]), .B(n12598), .Z(n12599) );
  XNOR U16697 ( .A(b[1191]), .B(n12600), .Z(c[1191]) );
  XOR U16698 ( .A(n12601), .B(n12602), .Z(n12598) );
  ANDN U16699 ( .B(n12603), .A(n12604), .Z(n12601) );
  XNOR U16700 ( .A(b[1190]), .B(n12602), .Z(n12603) );
  XNOR U16701 ( .A(b[1190]), .B(n12604), .Z(c[1190]) );
  XOR U16702 ( .A(n12605), .B(n12606), .Z(n12602) );
  ANDN U16703 ( .B(n12607), .A(n12608), .Z(n12605) );
  XNOR U16704 ( .A(b[1189]), .B(n12606), .Z(n12607) );
  XNOR U16705 ( .A(b[118]), .B(n12609), .Z(c[118]) );
  XNOR U16706 ( .A(b[1189]), .B(n12608), .Z(c[1189]) );
  XOR U16707 ( .A(n12610), .B(n12611), .Z(n12606) );
  ANDN U16708 ( .B(n12612), .A(n12613), .Z(n12610) );
  XNOR U16709 ( .A(b[1188]), .B(n12611), .Z(n12612) );
  XNOR U16710 ( .A(b[1188]), .B(n12613), .Z(c[1188]) );
  XOR U16711 ( .A(n12614), .B(n12615), .Z(n12611) );
  ANDN U16712 ( .B(n12616), .A(n12617), .Z(n12614) );
  XNOR U16713 ( .A(b[1187]), .B(n12615), .Z(n12616) );
  XNOR U16714 ( .A(b[1187]), .B(n12617), .Z(c[1187]) );
  XOR U16715 ( .A(n12618), .B(n12619), .Z(n12615) );
  ANDN U16716 ( .B(n12620), .A(n12621), .Z(n12618) );
  XNOR U16717 ( .A(b[1186]), .B(n12619), .Z(n12620) );
  XNOR U16718 ( .A(b[1186]), .B(n12621), .Z(c[1186]) );
  XOR U16719 ( .A(n12622), .B(n12623), .Z(n12619) );
  ANDN U16720 ( .B(n12624), .A(n12625), .Z(n12622) );
  XNOR U16721 ( .A(b[1185]), .B(n12623), .Z(n12624) );
  XNOR U16722 ( .A(b[1185]), .B(n12625), .Z(c[1185]) );
  XOR U16723 ( .A(n12626), .B(n12627), .Z(n12623) );
  ANDN U16724 ( .B(n12628), .A(n12629), .Z(n12626) );
  XNOR U16725 ( .A(b[1184]), .B(n12627), .Z(n12628) );
  XNOR U16726 ( .A(b[1184]), .B(n12629), .Z(c[1184]) );
  XOR U16727 ( .A(n12630), .B(n12631), .Z(n12627) );
  ANDN U16728 ( .B(n12632), .A(n12633), .Z(n12630) );
  XNOR U16729 ( .A(b[1183]), .B(n12631), .Z(n12632) );
  XNOR U16730 ( .A(b[1183]), .B(n12633), .Z(c[1183]) );
  XOR U16731 ( .A(n12634), .B(n12635), .Z(n12631) );
  ANDN U16732 ( .B(n12636), .A(n12637), .Z(n12634) );
  XNOR U16733 ( .A(b[1182]), .B(n12635), .Z(n12636) );
  XNOR U16734 ( .A(b[1182]), .B(n12637), .Z(c[1182]) );
  XOR U16735 ( .A(n12638), .B(n12639), .Z(n12635) );
  ANDN U16736 ( .B(n12640), .A(n12641), .Z(n12638) );
  XNOR U16737 ( .A(b[1181]), .B(n12639), .Z(n12640) );
  XNOR U16738 ( .A(b[1181]), .B(n12641), .Z(c[1181]) );
  XOR U16739 ( .A(n12642), .B(n12643), .Z(n12639) );
  ANDN U16740 ( .B(n12644), .A(n12645), .Z(n12642) );
  XNOR U16741 ( .A(b[1180]), .B(n12643), .Z(n12644) );
  XNOR U16742 ( .A(b[1180]), .B(n12645), .Z(c[1180]) );
  XOR U16743 ( .A(n12646), .B(n12647), .Z(n12643) );
  ANDN U16744 ( .B(n12648), .A(n12649), .Z(n12646) );
  XNOR U16745 ( .A(b[1179]), .B(n12647), .Z(n12648) );
  XNOR U16746 ( .A(b[117]), .B(n12650), .Z(c[117]) );
  XNOR U16747 ( .A(b[1179]), .B(n12649), .Z(c[1179]) );
  XOR U16748 ( .A(n12651), .B(n12652), .Z(n12647) );
  ANDN U16749 ( .B(n12653), .A(n12654), .Z(n12651) );
  XNOR U16750 ( .A(b[1178]), .B(n12652), .Z(n12653) );
  XNOR U16751 ( .A(b[1178]), .B(n12654), .Z(c[1178]) );
  XOR U16752 ( .A(n12655), .B(n12656), .Z(n12652) );
  ANDN U16753 ( .B(n12657), .A(n12658), .Z(n12655) );
  XNOR U16754 ( .A(b[1177]), .B(n12656), .Z(n12657) );
  XNOR U16755 ( .A(b[1177]), .B(n12658), .Z(c[1177]) );
  XOR U16756 ( .A(n12659), .B(n12660), .Z(n12656) );
  ANDN U16757 ( .B(n12661), .A(n12662), .Z(n12659) );
  XNOR U16758 ( .A(b[1176]), .B(n12660), .Z(n12661) );
  XNOR U16759 ( .A(b[1176]), .B(n12662), .Z(c[1176]) );
  XOR U16760 ( .A(n12663), .B(n12664), .Z(n12660) );
  ANDN U16761 ( .B(n12665), .A(n12666), .Z(n12663) );
  XNOR U16762 ( .A(b[1175]), .B(n12664), .Z(n12665) );
  XNOR U16763 ( .A(b[1175]), .B(n12666), .Z(c[1175]) );
  XOR U16764 ( .A(n12667), .B(n12668), .Z(n12664) );
  ANDN U16765 ( .B(n12669), .A(n12670), .Z(n12667) );
  XNOR U16766 ( .A(b[1174]), .B(n12668), .Z(n12669) );
  XNOR U16767 ( .A(b[1174]), .B(n12670), .Z(c[1174]) );
  XOR U16768 ( .A(n12671), .B(n12672), .Z(n12668) );
  ANDN U16769 ( .B(n12673), .A(n12674), .Z(n12671) );
  XNOR U16770 ( .A(b[1173]), .B(n12672), .Z(n12673) );
  XNOR U16771 ( .A(b[1173]), .B(n12674), .Z(c[1173]) );
  XOR U16772 ( .A(n12675), .B(n12676), .Z(n12672) );
  ANDN U16773 ( .B(n12677), .A(n12678), .Z(n12675) );
  XNOR U16774 ( .A(b[1172]), .B(n12676), .Z(n12677) );
  XNOR U16775 ( .A(b[1172]), .B(n12678), .Z(c[1172]) );
  XOR U16776 ( .A(n12679), .B(n12680), .Z(n12676) );
  ANDN U16777 ( .B(n12681), .A(n12682), .Z(n12679) );
  XNOR U16778 ( .A(b[1171]), .B(n12680), .Z(n12681) );
  XNOR U16779 ( .A(b[1171]), .B(n12682), .Z(c[1171]) );
  XOR U16780 ( .A(n12683), .B(n12684), .Z(n12680) );
  ANDN U16781 ( .B(n12685), .A(n12686), .Z(n12683) );
  XNOR U16782 ( .A(b[1170]), .B(n12684), .Z(n12685) );
  XNOR U16783 ( .A(b[1170]), .B(n12686), .Z(c[1170]) );
  XOR U16784 ( .A(n12687), .B(n12688), .Z(n12684) );
  ANDN U16785 ( .B(n12689), .A(n12690), .Z(n12687) );
  XNOR U16786 ( .A(b[1169]), .B(n12688), .Z(n12689) );
  XNOR U16787 ( .A(b[116]), .B(n12691), .Z(c[116]) );
  XNOR U16788 ( .A(b[1169]), .B(n12690), .Z(c[1169]) );
  XOR U16789 ( .A(n12692), .B(n12693), .Z(n12688) );
  ANDN U16790 ( .B(n12694), .A(n12695), .Z(n12692) );
  XNOR U16791 ( .A(b[1168]), .B(n12693), .Z(n12694) );
  XNOR U16792 ( .A(b[1168]), .B(n12695), .Z(c[1168]) );
  XOR U16793 ( .A(n12696), .B(n12697), .Z(n12693) );
  ANDN U16794 ( .B(n12698), .A(n12699), .Z(n12696) );
  XNOR U16795 ( .A(b[1167]), .B(n12697), .Z(n12698) );
  XNOR U16796 ( .A(b[1167]), .B(n12699), .Z(c[1167]) );
  XOR U16797 ( .A(n12700), .B(n12701), .Z(n12697) );
  ANDN U16798 ( .B(n12702), .A(n12703), .Z(n12700) );
  XNOR U16799 ( .A(b[1166]), .B(n12701), .Z(n12702) );
  XNOR U16800 ( .A(b[1166]), .B(n12703), .Z(c[1166]) );
  XOR U16801 ( .A(n12704), .B(n12705), .Z(n12701) );
  ANDN U16802 ( .B(n12706), .A(n12707), .Z(n12704) );
  XNOR U16803 ( .A(b[1165]), .B(n12705), .Z(n12706) );
  XNOR U16804 ( .A(b[1165]), .B(n12707), .Z(c[1165]) );
  XOR U16805 ( .A(n12708), .B(n12709), .Z(n12705) );
  ANDN U16806 ( .B(n12710), .A(n12711), .Z(n12708) );
  XNOR U16807 ( .A(b[1164]), .B(n12709), .Z(n12710) );
  XNOR U16808 ( .A(b[1164]), .B(n12711), .Z(c[1164]) );
  XOR U16809 ( .A(n12712), .B(n12713), .Z(n12709) );
  ANDN U16810 ( .B(n12714), .A(n12715), .Z(n12712) );
  XNOR U16811 ( .A(b[1163]), .B(n12713), .Z(n12714) );
  XNOR U16812 ( .A(b[1163]), .B(n12715), .Z(c[1163]) );
  XOR U16813 ( .A(n12716), .B(n12717), .Z(n12713) );
  ANDN U16814 ( .B(n12718), .A(n12719), .Z(n12716) );
  XNOR U16815 ( .A(b[1162]), .B(n12717), .Z(n12718) );
  XNOR U16816 ( .A(b[1162]), .B(n12719), .Z(c[1162]) );
  XOR U16817 ( .A(n12720), .B(n12721), .Z(n12717) );
  ANDN U16818 ( .B(n12722), .A(n12723), .Z(n12720) );
  XNOR U16819 ( .A(b[1161]), .B(n12721), .Z(n12722) );
  XNOR U16820 ( .A(b[1161]), .B(n12723), .Z(c[1161]) );
  XOR U16821 ( .A(n12724), .B(n12725), .Z(n12721) );
  ANDN U16822 ( .B(n12726), .A(n12727), .Z(n12724) );
  XNOR U16823 ( .A(b[1160]), .B(n12725), .Z(n12726) );
  XNOR U16824 ( .A(b[1160]), .B(n12727), .Z(c[1160]) );
  XOR U16825 ( .A(n12728), .B(n12729), .Z(n12725) );
  ANDN U16826 ( .B(n12730), .A(n12731), .Z(n12728) );
  XNOR U16827 ( .A(b[1159]), .B(n12729), .Z(n12730) );
  XNOR U16828 ( .A(b[115]), .B(n12732), .Z(c[115]) );
  XNOR U16829 ( .A(b[1159]), .B(n12731), .Z(c[1159]) );
  XOR U16830 ( .A(n12733), .B(n12734), .Z(n12729) );
  ANDN U16831 ( .B(n12735), .A(n12736), .Z(n12733) );
  XNOR U16832 ( .A(b[1158]), .B(n12734), .Z(n12735) );
  XNOR U16833 ( .A(b[1158]), .B(n12736), .Z(c[1158]) );
  XOR U16834 ( .A(n12737), .B(n12738), .Z(n12734) );
  ANDN U16835 ( .B(n12739), .A(n12740), .Z(n12737) );
  XNOR U16836 ( .A(b[1157]), .B(n12738), .Z(n12739) );
  XNOR U16837 ( .A(b[1157]), .B(n12740), .Z(c[1157]) );
  XOR U16838 ( .A(n12741), .B(n12742), .Z(n12738) );
  ANDN U16839 ( .B(n12743), .A(n12744), .Z(n12741) );
  XNOR U16840 ( .A(b[1156]), .B(n12742), .Z(n12743) );
  XNOR U16841 ( .A(b[1156]), .B(n12744), .Z(c[1156]) );
  XOR U16842 ( .A(n12745), .B(n12746), .Z(n12742) );
  ANDN U16843 ( .B(n12747), .A(n12748), .Z(n12745) );
  XNOR U16844 ( .A(b[1155]), .B(n12746), .Z(n12747) );
  XNOR U16845 ( .A(b[1155]), .B(n12748), .Z(c[1155]) );
  XOR U16846 ( .A(n12749), .B(n12750), .Z(n12746) );
  ANDN U16847 ( .B(n12751), .A(n12752), .Z(n12749) );
  XNOR U16848 ( .A(b[1154]), .B(n12750), .Z(n12751) );
  XNOR U16849 ( .A(b[1154]), .B(n12752), .Z(c[1154]) );
  XOR U16850 ( .A(n12753), .B(n12754), .Z(n12750) );
  ANDN U16851 ( .B(n12755), .A(n12756), .Z(n12753) );
  XNOR U16852 ( .A(b[1153]), .B(n12754), .Z(n12755) );
  XNOR U16853 ( .A(b[1153]), .B(n12756), .Z(c[1153]) );
  XOR U16854 ( .A(n12757), .B(n12758), .Z(n12754) );
  ANDN U16855 ( .B(n12759), .A(n12760), .Z(n12757) );
  XNOR U16856 ( .A(b[1152]), .B(n12758), .Z(n12759) );
  XNOR U16857 ( .A(b[1152]), .B(n12760), .Z(c[1152]) );
  XOR U16858 ( .A(n12761), .B(n12762), .Z(n12758) );
  ANDN U16859 ( .B(n12763), .A(n12764), .Z(n12761) );
  XNOR U16860 ( .A(b[1151]), .B(n12762), .Z(n12763) );
  XNOR U16861 ( .A(b[1151]), .B(n12764), .Z(c[1151]) );
  XOR U16862 ( .A(n12765), .B(n12766), .Z(n12762) );
  ANDN U16863 ( .B(n12767), .A(n12768), .Z(n12765) );
  XNOR U16864 ( .A(b[1150]), .B(n12766), .Z(n12767) );
  XNOR U16865 ( .A(b[1150]), .B(n12768), .Z(c[1150]) );
  XOR U16866 ( .A(n12769), .B(n12770), .Z(n12766) );
  ANDN U16867 ( .B(n12771), .A(n12772), .Z(n12769) );
  XNOR U16868 ( .A(b[1149]), .B(n12770), .Z(n12771) );
  XNOR U16869 ( .A(b[114]), .B(n12773), .Z(c[114]) );
  XNOR U16870 ( .A(b[1149]), .B(n12772), .Z(c[1149]) );
  XOR U16871 ( .A(n12774), .B(n12775), .Z(n12770) );
  ANDN U16872 ( .B(n12776), .A(n12777), .Z(n12774) );
  XNOR U16873 ( .A(b[1148]), .B(n12775), .Z(n12776) );
  XNOR U16874 ( .A(b[1148]), .B(n12777), .Z(c[1148]) );
  XOR U16875 ( .A(n12778), .B(n12779), .Z(n12775) );
  ANDN U16876 ( .B(n12780), .A(n12781), .Z(n12778) );
  XNOR U16877 ( .A(b[1147]), .B(n12779), .Z(n12780) );
  XNOR U16878 ( .A(b[1147]), .B(n12781), .Z(c[1147]) );
  XOR U16879 ( .A(n12782), .B(n12783), .Z(n12779) );
  ANDN U16880 ( .B(n12784), .A(n12785), .Z(n12782) );
  XNOR U16881 ( .A(b[1146]), .B(n12783), .Z(n12784) );
  XNOR U16882 ( .A(b[1146]), .B(n12785), .Z(c[1146]) );
  XOR U16883 ( .A(n12786), .B(n12787), .Z(n12783) );
  ANDN U16884 ( .B(n12788), .A(n12789), .Z(n12786) );
  XNOR U16885 ( .A(b[1145]), .B(n12787), .Z(n12788) );
  XNOR U16886 ( .A(b[1145]), .B(n12789), .Z(c[1145]) );
  XOR U16887 ( .A(n12790), .B(n12791), .Z(n12787) );
  ANDN U16888 ( .B(n12792), .A(n12793), .Z(n12790) );
  XNOR U16889 ( .A(b[1144]), .B(n12791), .Z(n12792) );
  XNOR U16890 ( .A(b[1144]), .B(n12793), .Z(c[1144]) );
  XOR U16891 ( .A(n12794), .B(n12795), .Z(n12791) );
  ANDN U16892 ( .B(n12796), .A(n12797), .Z(n12794) );
  XNOR U16893 ( .A(b[1143]), .B(n12795), .Z(n12796) );
  XNOR U16894 ( .A(b[1143]), .B(n12797), .Z(c[1143]) );
  XOR U16895 ( .A(n12798), .B(n12799), .Z(n12795) );
  ANDN U16896 ( .B(n12800), .A(n12801), .Z(n12798) );
  XNOR U16897 ( .A(b[1142]), .B(n12799), .Z(n12800) );
  XNOR U16898 ( .A(b[1142]), .B(n12801), .Z(c[1142]) );
  XOR U16899 ( .A(n12802), .B(n12803), .Z(n12799) );
  ANDN U16900 ( .B(n12804), .A(n12805), .Z(n12802) );
  XNOR U16901 ( .A(b[1141]), .B(n12803), .Z(n12804) );
  XNOR U16902 ( .A(b[1141]), .B(n12805), .Z(c[1141]) );
  XOR U16903 ( .A(n12806), .B(n12807), .Z(n12803) );
  ANDN U16904 ( .B(n12808), .A(n12809), .Z(n12806) );
  XNOR U16905 ( .A(b[1140]), .B(n12807), .Z(n12808) );
  XNOR U16906 ( .A(b[1140]), .B(n12809), .Z(c[1140]) );
  XOR U16907 ( .A(n12810), .B(n12811), .Z(n12807) );
  ANDN U16908 ( .B(n12812), .A(n12813), .Z(n12810) );
  XNOR U16909 ( .A(b[1139]), .B(n12811), .Z(n12812) );
  XNOR U16910 ( .A(b[113]), .B(n12814), .Z(c[113]) );
  XNOR U16911 ( .A(b[1139]), .B(n12813), .Z(c[1139]) );
  XOR U16912 ( .A(n12815), .B(n12816), .Z(n12811) );
  ANDN U16913 ( .B(n12817), .A(n12818), .Z(n12815) );
  XNOR U16914 ( .A(b[1138]), .B(n12816), .Z(n12817) );
  XNOR U16915 ( .A(b[1138]), .B(n12818), .Z(c[1138]) );
  XOR U16916 ( .A(n12819), .B(n12820), .Z(n12816) );
  ANDN U16917 ( .B(n12821), .A(n12822), .Z(n12819) );
  XNOR U16918 ( .A(b[1137]), .B(n12820), .Z(n12821) );
  XNOR U16919 ( .A(b[1137]), .B(n12822), .Z(c[1137]) );
  XOR U16920 ( .A(n12823), .B(n12824), .Z(n12820) );
  ANDN U16921 ( .B(n12825), .A(n12826), .Z(n12823) );
  XNOR U16922 ( .A(b[1136]), .B(n12824), .Z(n12825) );
  XNOR U16923 ( .A(b[1136]), .B(n12826), .Z(c[1136]) );
  XOR U16924 ( .A(n12827), .B(n12828), .Z(n12824) );
  ANDN U16925 ( .B(n12829), .A(n12830), .Z(n12827) );
  XNOR U16926 ( .A(b[1135]), .B(n12828), .Z(n12829) );
  XNOR U16927 ( .A(b[1135]), .B(n12830), .Z(c[1135]) );
  XOR U16928 ( .A(n12831), .B(n12832), .Z(n12828) );
  ANDN U16929 ( .B(n12833), .A(n12834), .Z(n12831) );
  XNOR U16930 ( .A(b[1134]), .B(n12832), .Z(n12833) );
  XNOR U16931 ( .A(b[1134]), .B(n12834), .Z(c[1134]) );
  XOR U16932 ( .A(n12835), .B(n12836), .Z(n12832) );
  ANDN U16933 ( .B(n12837), .A(n12838), .Z(n12835) );
  XNOR U16934 ( .A(b[1133]), .B(n12836), .Z(n12837) );
  XNOR U16935 ( .A(b[1133]), .B(n12838), .Z(c[1133]) );
  XOR U16936 ( .A(n12839), .B(n12840), .Z(n12836) );
  ANDN U16937 ( .B(n12841), .A(n12842), .Z(n12839) );
  XNOR U16938 ( .A(b[1132]), .B(n12840), .Z(n12841) );
  XNOR U16939 ( .A(b[1132]), .B(n12842), .Z(c[1132]) );
  XOR U16940 ( .A(n12843), .B(n12844), .Z(n12840) );
  ANDN U16941 ( .B(n12845), .A(n12846), .Z(n12843) );
  XNOR U16942 ( .A(b[1131]), .B(n12844), .Z(n12845) );
  XNOR U16943 ( .A(b[1131]), .B(n12846), .Z(c[1131]) );
  XOR U16944 ( .A(n12847), .B(n12848), .Z(n12844) );
  ANDN U16945 ( .B(n12849), .A(n12850), .Z(n12847) );
  XNOR U16946 ( .A(b[1130]), .B(n12848), .Z(n12849) );
  XNOR U16947 ( .A(b[1130]), .B(n12850), .Z(c[1130]) );
  XOR U16948 ( .A(n12851), .B(n12852), .Z(n12848) );
  ANDN U16949 ( .B(n12853), .A(n12854), .Z(n12851) );
  XNOR U16950 ( .A(b[1129]), .B(n12852), .Z(n12853) );
  XNOR U16951 ( .A(b[112]), .B(n12855), .Z(c[112]) );
  XNOR U16952 ( .A(b[1129]), .B(n12854), .Z(c[1129]) );
  XOR U16953 ( .A(n12856), .B(n12857), .Z(n12852) );
  ANDN U16954 ( .B(n12858), .A(n12859), .Z(n12856) );
  XNOR U16955 ( .A(b[1128]), .B(n12857), .Z(n12858) );
  XNOR U16956 ( .A(b[1128]), .B(n12859), .Z(c[1128]) );
  XOR U16957 ( .A(n12860), .B(n12861), .Z(n12857) );
  ANDN U16958 ( .B(n12862), .A(n12863), .Z(n12860) );
  XNOR U16959 ( .A(b[1127]), .B(n12861), .Z(n12862) );
  XNOR U16960 ( .A(b[1127]), .B(n12863), .Z(c[1127]) );
  XOR U16961 ( .A(n12864), .B(n12865), .Z(n12861) );
  ANDN U16962 ( .B(n12866), .A(n12867), .Z(n12864) );
  XNOR U16963 ( .A(b[1126]), .B(n12865), .Z(n12866) );
  XNOR U16964 ( .A(b[1126]), .B(n12867), .Z(c[1126]) );
  XOR U16965 ( .A(n12868), .B(n12869), .Z(n12865) );
  ANDN U16966 ( .B(n12870), .A(n12871), .Z(n12868) );
  XNOR U16967 ( .A(b[1125]), .B(n12869), .Z(n12870) );
  XNOR U16968 ( .A(b[1125]), .B(n12871), .Z(c[1125]) );
  XOR U16969 ( .A(n12872), .B(n12873), .Z(n12869) );
  ANDN U16970 ( .B(n12874), .A(n12875), .Z(n12872) );
  XNOR U16971 ( .A(b[1124]), .B(n12873), .Z(n12874) );
  XNOR U16972 ( .A(b[1124]), .B(n12875), .Z(c[1124]) );
  XOR U16973 ( .A(n12876), .B(n12877), .Z(n12873) );
  ANDN U16974 ( .B(n12878), .A(n12879), .Z(n12876) );
  XNOR U16975 ( .A(b[1123]), .B(n12877), .Z(n12878) );
  XNOR U16976 ( .A(b[1123]), .B(n12879), .Z(c[1123]) );
  XOR U16977 ( .A(n12880), .B(n12881), .Z(n12877) );
  ANDN U16978 ( .B(n12882), .A(n12883), .Z(n12880) );
  XNOR U16979 ( .A(b[1122]), .B(n12881), .Z(n12882) );
  XNOR U16980 ( .A(b[1122]), .B(n12883), .Z(c[1122]) );
  XOR U16981 ( .A(n12884), .B(n12885), .Z(n12881) );
  ANDN U16982 ( .B(n12886), .A(n12887), .Z(n12884) );
  XNOR U16983 ( .A(b[1121]), .B(n12885), .Z(n12886) );
  XNOR U16984 ( .A(b[1121]), .B(n12887), .Z(c[1121]) );
  XOR U16985 ( .A(n12888), .B(n12889), .Z(n12885) );
  ANDN U16986 ( .B(n12890), .A(n12891), .Z(n12888) );
  XNOR U16987 ( .A(b[1120]), .B(n12889), .Z(n12890) );
  XNOR U16988 ( .A(b[1120]), .B(n12891), .Z(c[1120]) );
  XOR U16989 ( .A(n12892), .B(n12893), .Z(n12889) );
  ANDN U16990 ( .B(n12894), .A(n12895), .Z(n12892) );
  XNOR U16991 ( .A(b[1119]), .B(n12893), .Z(n12894) );
  XNOR U16992 ( .A(b[111]), .B(n12896), .Z(c[111]) );
  XNOR U16993 ( .A(b[1119]), .B(n12895), .Z(c[1119]) );
  XOR U16994 ( .A(n12897), .B(n12898), .Z(n12893) );
  ANDN U16995 ( .B(n12899), .A(n12900), .Z(n12897) );
  XNOR U16996 ( .A(b[1118]), .B(n12898), .Z(n12899) );
  XNOR U16997 ( .A(b[1118]), .B(n12900), .Z(c[1118]) );
  XOR U16998 ( .A(n12901), .B(n12902), .Z(n12898) );
  ANDN U16999 ( .B(n12903), .A(n12904), .Z(n12901) );
  XNOR U17000 ( .A(b[1117]), .B(n12902), .Z(n12903) );
  XNOR U17001 ( .A(b[1117]), .B(n12904), .Z(c[1117]) );
  XOR U17002 ( .A(n12905), .B(n12906), .Z(n12902) );
  ANDN U17003 ( .B(n12907), .A(n12908), .Z(n12905) );
  XNOR U17004 ( .A(b[1116]), .B(n12906), .Z(n12907) );
  XNOR U17005 ( .A(b[1116]), .B(n12908), .Z(c[1116]) );
  XOR U17006 ( .A(n12909), .B(n12910), .Z(n12906) );
  ANDN U17007 ( .B(n12911), .A(n12912), .Z(n12909) );
  XNOR U17008 ( .A(b[1115]), .B(n12910), .Z(n12911) );
  XNOR U17009 ( .A(b[1115]), .B(n12912), .Z(c[1115]) );
  XOR U17010 ( .A(n12913), .B(n12914), .Z(n12910) );
  ANDN U17011 ( .B(n12915), .A(n12916), .Z(n12913) );
  XNOR U17012 ( .A(b[1114]), .B(n12914), .Z(n12915) );
  XNOR U17013 ( .A(b[1114]), .B(n12916), .Z(c[1114]) );
  XOR U17014 ( .A(n12917), .B(n12918), .Z(n12914) );
  ANDN U17015 ( .B(n12919), .A(n12920), .Z(n12917) );
  XNOR U17016 ( .A(b[1113]), .B(n12918), .Z(n12919) );
  XNOR U17017 ( .A(b[1113]), .B(n12920), .Z(c[1113]) );
  XOR U17018 ( .A(n12921), .B(n12922), .Z(n12918) );
  ANDN U17019 ( .B(n12923), .A(n12924), .Z(n12921) );
  XNOR U17020 ( .A(b[1112]), .B(n12922), .Z(n12923) );
  XNOR U17021 ( .A(b[1112]), .B(n12924), .Z(c[1112]) );
  XOR U17022 ( .A(n12925), .B(n12926), .Z(n12922) );
  ANDN U17023 ( .B(n12927), .A(n12928), .Z(n12925) );
  XNOR U17024 ( .A(b[1111]), .B(n12926), .Z(n12927) );
  XNOR U17025 ( .A(b[1111]), .B(n12928), .Z(c[1111]) );
  XOR U17026 ( .A(n12929), .B(n12930), .Z(n12926) );
  ANDN U17027 ( .B(n12931), .A(n12932), .Z(n12929) );
  XNOR U17028 ( .A(b[1110]), .B(n12930), .Z(n12931) );
  XNOR U17029 ( .A(b[1110]), .B(n12932), .Z(c[1110]) );
  XOR U17030 ( .A(n12933), .B(n12934), .Z(n12930) );
  ANDN U17031 ( .B(n12935), .A(n12936), .Z(n12933) );
  XNOR U17032 ( .A(b[1109]), .B(n12934), .Z(n12935) );
  XNOR U17033 ( .A(b[110]), .B(n12937), .Z(c[110]) );
  XNOR U17034 ( .A(b[1109]), .B(n12936), .Z(c[1109]) );
  XOR U17035 ( .A(n12938), .B(n12939), .Z(n12934) );
  ANDN U17036 ( .B(n12940), .A(n12941), .Z(n12938) );
  XNOR U17037 ( .A(b[1108]), .B(n12939), .Z(n12940) );
  XNOR U17038 ( .A(b[1108]), .B(n12941), .Z(c[1108]) );
  XOR U17039 ( .A(n12942), .B(n12943), .Z(n12939) );
  ANDN U17040 ( .B(n12944), .A(n12945), .Z(n12942) );
  XNOR U17041 ( .A(b[1107]), .B(n12943), .Z(n12944) );
  XNOR U17042 ( .A(b[1107]), .B(n12945), .Z(c[1107]) );
  XOR U17043 ( .A(n12946), .B(n12947), .Z(n12943) );
  ANDN U17044 ( .B(n12948), .A(n12949), .Z(n12946) );
  XNOR U17045 ( .A(b[1106]), .B(n12947), .Z(n12948) );
  XNOR U17046 ( .A(b[1106]), .B(n12949), .Z(c[1106]) );
  XOR U17047 ( .A(n12950), .B(n12951), .Z(n12947) );
  ANDN U17048 ( .B(n12952), .A(n12953), .Z(n12950) );
  XNOR U17049 ( .A(b[1105]), .B(n12951), .Z(n12952) );
  XNOR U17050 ( .A(b[1105]), .B(n12953), .Z(c[1105]) );
  XOR U17051 ( .A(n12954), .B(n12955), .Z(n12951) );
  ANDN U17052 ( .B(n12956), .A(n12957), .Z(n12954) );
  XNOR U17053 ( .A(b[1104]), .B(n12955), .Z(n12956) );
  XNOR U17054 ( .A(b[1104]), .B(n12957), .Z(c[1104]) );
  XOR U17055 ( .A(n12958), .B(n12959), .Z(n12955) );
  ANDN U17056 ( .B(n12960), .A(n12961), .Z(n12958) );
  XNOR U17057 ( .A(b[1103]), .B(n12959), .Z(n12960) );
  XNOR U17058 ( .A(b[1103]), .B(n12961), .Z(c[1103]) );
  XOR U17059 ( .A(n12962), .B(n12963), .Z(n12959) );
  ANDN U17060 ( .B(n12964), .A(n12965), .Z(n12962) );
  XNOR U17061 ( .A(b[1102]), .B(n12963), .Z(n12964) );
  XNOR U17062 ( .A(b[1102]), .B(n12965), .Z(c[1102]) );
  XOR U17063 ( .A(n12966), .B(n12967), .Z(n12963) );
  ANDN U17064 ( .B(n12968), .A(n12969), .Z(n12966) );
  XNOR U17065 ( .A(b[1101]), .B(n12967), .Z(n12968) );
  XNOR U17066 ( .A(b[1101]), .B(n12969), .Z(c[1101]) );
  XOR U17067 ( .A(n12970), .B(n12971), .Z(n12967) );
  ANDN U17068 ( .B(n12972), .A(n12973), .Z(n12970) );
  XNOR U17069 ( .A(b[1100]), .B(n12971), .Z(n12972) );
  XNOR U17070 ( .A(b[1100]), .B(n12973), .Z(c[1100]) );
  XOR U17071 ( .A(n12974), .B(n12975), .Z(n12971) );
  ANDN U17072 ( .B(n12976), .A(n12977), .Z(n12974) );
  XNOR U17073 ( .A(b[1099]), .B(n12975), .Z(n12976) );
  XNOR U17074 ( .A(b[10]), .B(n12978), .Z(c[10]) );
  XNOR U17075 ( .A(b[109]), .B(n12979), .Z(c[109]) );
  XNOR U17076 ( .A(b[1099]), .B(n12977), .Z(c[1099]) );
  XOR U17077 ( .A(n12980), .B(n12981), .Z(n12975) );
  ANDN U17078 ( .B(n12982), .A(n12983), .Z(n12980) );
  XNOR U17079 ( .A(b[1098]), .B(n12981), .Z(n12982) );
  XNOR U17080 ( .A(b[1098]), .B(n12983), .Z(c[1098]) );
  XOR U17081 ( .A(n12984), .B(n12985), .Z(n12981) );
  ANDN U17082 ( .B(n12986), .A(n12987), .Z(n12984) );
  XNOR U17083 ( .A(b[1097]), .B(n12985), .Z(n12986) );
  XNOR U17084 ( .A(b[1097]), .B(n12987), .Z(c[1097]) );
  XOR U17085 ( .A(n12988), .B(n12989), .Z(n12985) );
  ANDN U17086 ( .B(n12990), .A(n12991), .Z(n12988) );
  XNOR U17087 ( .A(b[1096]), .B(n12989), .Z(n12990) );
  XNOR U17088 ( .A(b[1096]), .B(n12991), .Z(c[1096]) );
  XOR U17089 ( .A(n12992), .B(n12993), .Z(n12989) );
  ANDN U17090 ( .B(n12994), .A(n12995), .Z(n12992) );
  XNOR U17091 ( .A(b[1095]), .B(n12993), .Z(n12994) );
  XNOR U17092 ( .A(b[1095]), .B(n12995), .Z(c[1095]) );
  XOR U17093 ( .A(n12996), .B(n12997), .Z(n12993) );
  ANDN U17094 ( .B(n12998), .A(n12999), .Z(n12996) );
  XNOR U17095 ( .A(b[1094]), .B(n12997), .Z(n12998) );
  XNOR U17096 ( .A(b[1094]), .B(n12999), .Z(c[1094]) );
  XOR U17097 ( .A(n13000), .B(n13001), .Z(n12997) );
  ANDN U17098 ( .B(n13002), .A(n13003), .Z(n13000) );
  XNOR U17099 ( .A(b[1093]), .B(n13001), .Z(n13002) );
  XNOR U17100 ( .A(b[1093]), .B(n13003), .Z(c[1093]) );
  XOR U17101 ( .A(n13004), .B(n13005), .Z(n13001) );
  ANDN U17102 ( .B(n13006), .A(n13007), .Z(n13004) );
  XNOR U17103 ( .A(b[1092]), .B(n13005), .Z(n13006) );
  XNOR U17104 ( .A(b[1092]), .B(n13007), .Z(c[1092]) );
  XOR U17105 ( .A(n13008), .B(n13009), .Z(n13005) );
  ANDN U17106 ( .B(n13010), .A(n13011), .Z(n13008) );
  XNOR U17107 ( .A(b[1091]), .B(n13009), .Z(n13010) );
  XNOR U17108 ( .A(b[1091]), .B(n13011), .Z(c[1091]) );
  XOR U17109 ( .A(n13012), .B(n13013), .Z(n13009) );
  ANDN U17110 ( .B(n13014), .A(n13015), .Z(n13012) );
  XNOR U17111 ( .A(b[1090]), .B(n13013), .Z(n13014) );
  XNOR U17112 ( .A(b[1090]), .B(n13015), .Z(c[1090]) );
  XOR U17113 ( .A(n13016), .B(n13017), .Z(n13013) );
  ANDN U17114 ( .B(n13018), .A(n13019), .Z(n13016) );
  XNOR U17115 ( .A(b[1089]), .B(n13017), .Z(n13018) );
  XNOR U17116 ( .A(b[108]), .B(n13020), .Z(c[108]) );
  XNOR U17117 ( .A(b[1089]), .B(n13019), .Z(c[1089]) );
  XOR U17118 ( .A(n13021), .B(n13022), .Z(n13017) );
  ANDN U17119 ( .B(n13023), .A(n13024), .Z(n13021) );
  XNOR U17120 ( .A(b[1088]), .B(n13022), .Z(n13023) );
  XNOR U17121 ( .A(b[1088]), .B(n13024), .Z(c[1088]) );
  XOR U17122 ( .A(n13025), .B(n13026), .Z(n13022) );
  ANDN U17123 ( .B(n13027), .A(n13028), .Z(n13025) );
  XNOR U17124 ( .A(b[1087]), .B(n13026), .Z(n13027) );
  XNOR U17125 ( .A(b[1087]), .B(n13028), .Z(c[1087]) );
  XOR U17126 ( .A(n13029), .B(n13030), .Z(n13026) );
  ANDN U17127 ( .B(n13031), .A(n13032), .Z(n13029) );
  XNOR U17128 ( .A(b[1086]), .B(n13030), .Z(n13031) );
  XNOR U17129 ( .A(b[1086]), .B(n13032), .Z(c[1086]) );
  XOR U17130 ( .A(n13033), .B(n13034), .Z(n13030) );
  ANDN U17131 ( .B(n13035), .A(n13036), .Z(n13033) );
  XNOR U17132 ( .A(b[1085]), .B(n13034), .Z(n13035) );
  XNOR U17133 ( .A(b[1085]), .B(n13036), .Z(c[1085]) );
  XOR U17134 ( .A(n13037), .B(n13038), .Z(n13034) );
  ANDN U17135 ( .B(n13039), .A(n13040), .Z(n13037) );
  XNOR U17136 ( .A(b[1084]), .B(n13038), .Z(n13039) );
  XNOR U17137 ( .A(b[1084]), .B(n13040), .Z(c[1084]) );
  XOR U17138 ( .A(n13041), .B(n13042), .Z(n13038) );
  ANDN U17139 ( .B(n13043), .A(n13044), .Z(n13041) );
  XNOR U17140 ( .A(b[1083]), .B(n13042), .Z(n13043) );
  XNOR U17141 ( .A(b[1083]), .B(n13044), .Z(c[1083]) );
  XOR U17142 ( .A(n13045), .B(n13046), .Z(n13042) );
  ANDN U17143 ( .B(n13047), .A(n13048), .Z(n13045) );
  XNOR U17144 ( .A(b[1082]), .B(n13046), .Z(n13047) );
  XNOR U17145 ( .A(b[1082]), .B(n13048), .Z(c[1082]) );
  XOR U17146 ( .A(n13049), .B(n13050), .Z(n13046) );
  ANDN U17147 ( .B(n13051), .A(n13052), .Z(n13049) );
  XNOR U17148 ( .A(b[1081]), .B(n13050), .Z(n13051) );
  XNOR U17149 ( .A(b[1081]), .B(n13052), .Z(c[1081]) );
  XOR U17150 ( .A(n13053), .B(n13054), .Z(n13050) );
  ANDN U17151 ( .B(n13055), .A(n13056), .Z(n13053) );
  XNOR U17152 ( .A(b[1080]), .B(n13054), .Z(n13055) );
  XNOR U17153 ( .A(b[1080]), .B(n13056), .Z(c[1080]) );
  XOR U17154 ( .A(n13057), .B(n13058), .Z(n13054) );
  ANDN U17155 ( .B(n13059), .A(n13060), .Z(n13057) );
  XNOR U17156 ( .A(b[1079]), .B(n13058), .Z(n13059) );
  XNOR U17157 ( .A(b[107]), .B(n13061), .Z(c[107]) );
  XNOR U17158 ( .A(b[1079]), .B(n13060), .Z(c[1079]) );
  XOR U17159 ( .A(n13062), .B(n13063), .Z(n13058) );
  ANDN U17160 ( .B(n13064), .A(n13065), .Z(n13062) );
  XNOR U17161 ( .A(b[1078]), .B(n13063), .Z(n13064) );
  XNOR U17162 ( .A(b[1078]), .B(n13065), .Z(c[1078]) );
  XOR U17163 ( .A(n13066), .B(n13067), .Z(n13063) );
  ANDN U17164 ( .B(n13068), .A(n13069), .Z(n13066) );
  XNOR U17165 ( .A(b[1077]), .B(n13067), .Z(n13068) );
  XNOR U17166 ( .A(b[1077]), .B(n13069), .Z(c[1077]) );
  XOR U17167 ( .A(n13070), .B(n13071), .Z(n13067) );
  ANDN U17168 ( .B(n13072), .A(n13073), .Z(n13070) );
  XNOR U17169 ( .A(b[1076]), .B(n13071), .Z(n13072) );
  XNOR U17170 ( .A(b[1076]), .B(n13073), .Z(c[1076]) );
  XOR U17171 ( .A(n13074), .B(n13075), .Z(n13071) );
  ANDN U17172 ( .B(n13076), .A(n13077), .Z(n13074) );
  XNOR U17173 ( .A(b[1075]), .B(n13075), .Z(n13076) );
  XNOR U17174 ( .A(b[1075]), .B(n13077), .Z(c[1075]) );
  XOR U17175 ( .A(n13078), .B(n13079), .Z(n13075) );
  ANDN U17176 ( .B(n13080), .A(n13081), .Z(n13078) );
  XNOR U17177 ( .A(b[1074]), .B(n13079), .Z(n13080) );
  XNOR U17178 ( .A(b[1074]), .B(n13081), .Z(c[1074]) );
  XOR U17179 ( .A(n13082), .B(n13083), .Z(n13079) );
  ANDN U17180 ( .B(n13084), .A(n13085), .Z(n13082) );
  XNOR U17181 ( .A(b[1073]), .B(n13083), .Z(n13084) );
  XNOR U17182 ( .A(b[1073]), .B(n13085), .Z(c[1073]) );
  XOR U17183 ( .A(n13086), .B(n13087), .Z(n13083) );
  ANDN U17184 ( .B(n13088), .A(n13089), .Z(n13086) );
  XNOR U17185 ( .A(b[1072]), .B(n13087), .Z(n13088) );
  XNOR U17186 ( .A(b[1072]), .B(n13089), .Z(c[1072]) );
  XOR U17187 ( .A(n13090), .B(n13091), .Z(n13087) );
  ANDN U17188 ( .B(n13092), .A(n13093), .Z(n13090) );
  XNOR U17189 ( .A(b[1071]), .B(n13091), .Z(n13092) );
  XNOR U17190 ( .A(b[1071]), .B(n13093), .Z(c[1071]) );
  XOR U17191 ( .A(n13094), .B(n13095), .Z(n13091) );
  ANDN U17192 ( .B(n13096), .A(n13097), .Z(n13094) );
  XNOR U17193 ( .A(b[1070]), .B(n13095), .Z(n13096) );
  XNOR U17194 ( .A(b[1070]), .B(n13097), .Z(c[1070]) );
  XOR U17195 ( .A(n13098), .B(n13099), .Z(n13095) );
  ANDN U17196 ( .B(n13100), .A(n13101), .Z(n13098) );
  XNOR U17197 ( .A(b[1069]), .B(n13099), .Z(n13100) );
  XNOR U17198 ( .A(b[106]), .B(n13102), .Z(c[106]) );
  XNOR U17199 ( .A(b[1069]), .B(n13101), .Z(c[1069]) );
  XOR U17200 ( .A(n13103), .B(n13104), .Z(n13099) );
  ANDN U17201 ( .B(n13105), .A(n13106), .Z(n13103) );
  XNOR U17202 ( .A(b[1068]), .B(n13104), .Z(n13105) );
  XNOR U17203 ( .A(b[1068]), .B(n13106), .Z(c[1068]) );
  XOR U17204 ( .A(n13107), .B(n13108), .Z(n13104) );
  ANDN U17205 ( .B(n13109), .A(n13110), .Z(n13107) );
  XNOR U17206 ( .A(b[1067]), .B(n13108), .Z(n13109) );
  XNOR U17207 ( .A(b[1067]), .B(n13110), .Z(c[1067]) );
  XOR U17208 ( .A(n13111), .B(n13112), .Z(n13108) );
  ANDN U17209 ( .B(n13113), .A(n13114), .Z(n13111) );
  XNOR U17210 ( .A(b[1066]), .B(n13112), .Z(n13113) );
  XNOR U17211 ( .A(b[1066]), .B(n13114), .Z(c[1066]) );
  XOR U17212 ( .A(n13115), .B(n13116), .Z(n13112) );
  ANDN U17213 ( .B(n13117), .A(n13118), .Z(n13115) );
  XNOR U17214 ( .A(b[1065]), .B(n13116), .Z(n13117) );
  XNOR U17215 ( .A(b[1065]), .B(n13118), .Z(c[1065]) );
  XOR U17216 ( .A(n13119), .B(n13120), .Z(n13116) );
  ANDN U17217 ( .B(n13121), .A(n13122), .Z(n13119) );
  XNOR U17218 ( .A(b[1064]), .B(n13120), .Z(n13121) );
  XNOR U17219 ( .A(b[1064]), .B(n13122), .Z(c[1064]) );
  XOR U17220 ( .A(n13123), .B(n13124), .Z(n13120) );
  ANDN U17221 ( .B(n13125), .A(n13126), .Z(n13123) );
  XNOR U17222 ( .A(b[1063]), .B(n13124), .Z(n13125) );
  XNOR U17223 ( .A(b[1063]), .B(n13126), .Z(c[1063]) );
  XOR U17224 ( .A(n13127), .B(n13128), .Z(n13124) );
  ANDN U17225 ( .B(n13129), .A(n13130), .Z(n13127) );
  XNOR U17226 ( .A(b[1062]), .B(n13128), .Z(n13129) );
  XNOR U17227 ( .A(b[1062]), .B(n13130), .Z(c[1062]) );
  XOR U17228 ( .A(n13131), .B(n13132), .Z(n13128) );
  ANDN U17229 ( .B(n13133), .A(n13134), .Z(n13131) );
  XNOR U17230 ( .A(b[1061]), .B(n13132), .Z(n13133) );
  XNOR U17231 ( .A(b[1061]), .B(n13134), .Z(c[1061]) );
  XOR U17232 ( .A(n13135), .B(n13136), .Z(n13132) );
  ANDN U17233 ( .B(n13137), .A(n13138), .Z(n13135) );
  XNOR U17234 ( .A(b[1060]), .B(n13136), .Z(n13137) );
  XNOR U17235 ( .A(b[1060]), .B(n13138), .Z(c[1060]) );
  XOR U17236 ( .A(n13139), .B(n13140), .Z(n13136) );
  ANDN U17237 ( .B(n13141), .A(n13142), .Z(n13139) );
  XNOR U17238 ( .A(b[1059]), .B(n13140), .Z(n13141) );
  XNOR U17239 ( .A(b[105]), .B(n13143), .Z(c[105]) );
  XNOR U17240 ( .A(b[1059]), .B(n13142), .Z(c[1059]) );
  XOR U17241 ( .A(n13144), .B(n13145), .Z(n13140) );
  ANDN U17242 ( .B(n13146), .A(n13147), .Z(n13144) );
  XNOR U17243 ( .A(b[1058]), .B(n13145), .Z(n13146) );
  XNOR U17244 ( .A(b[1058]), .B(n13147), .Z(c[1058]) );
  XOR U17245 ( .A(n13148), .B(n13149), .Z(n13145) );
  ANDN U17246 ( .B(n13150), .A(n13151), .Z(n13148) );
  XNOR U17247 ( .A(b[1057]), .B(n13149), .Z(n13150) );
  XNOR U17248 ( .A(b[1057]), .B(n13151), .Z(c[1057]) );
  XOR U17249 ( .A(n13152), .B(n13153), .Z(n13149) );
  ANDN U17250 ( .B(n13154), .A(n13155), .Z(n13152) );
  XNOR U17251 ( .A(b[1056]), .B(n13153), .Z(n13154) );
  XNOR U17252 ( .A(b[1056]), .B(n13155), .Z(c[1056]) );
  XOR U17253 ( .A(n13156), .B(n13157), .Z(n13153) );
  ANDN U17254 ( .B(n13158), .A(n13159), .Z(n13156) );
  XNOR U17255 ( .A(b[1055]), .B(n13157), .Z(n13158) );
  XNOR U17256 ( .A(b[1055]), .B(n13159), .Z(c[1055]) );
  XOR U17257 ( .A(n13160), .B(n13161), .Z(n13157) );
  ANDN U17258 ( .B(n13162), .A(n13163), .Z(n13160) );
  XNOR U17259 ( .A(b[1054]), .B(n13161), .Z(n13162) );
  XNOR U17260 ( .A(b[1054]), .B(n13163), .Z(c[1054]) );
  XOR U17261 ( .A(n13164), .B(n13165), .Z(n13161) );
  ANDN U17262 ( .B(n13166), .A(n13167), .Z(n13164) );
  XNOR U17263 ( .A(b[1053]), .B(n13165), .Z(n13166) );
  XNOR U17264 ( .A(b[1053]), .B(n13167), .Z(c[1053]) );
  XOR U17265 ( .A(n13168), .B(n13169), .Z(n13165) );
  ANDN U17266 ( .B(n13170), .A(n13171), .Z(n13168) );
  XNOR U17267 ( .A(b[1052]), .B(n13169), .Z(n13170) );
  XNOR U17268 ( .A(b[1052]), .B(n13171), .Z(c[1052]) );
  XOR U17269 ( .A(n13172), .B(n13173), .Z(n13169) );
  ANDN U17270 ( .B(n13174), .A(n13175), .Z(n13172) );
  XNOR U17271 ( .A(b[1051]), .B(n13173), .Z(n13174) );
  XNOR U17272 ( .A(b[1051]), .B(n13175), .Z(c[1051]) );
  XOR U17273 ( .A(n13176), .B(n13177), .Z(n13173) );
  ANDN U17274 ( .B(n13178), .A(n13179), .Z(n13176) );
  XNOR U17275 ( .A(b[1050]), .B(n13177), .Z(n13178) );
  XNOR U17276 ( .A(b[1050]), .B(n13179), .Z(c[1050]) );
  XOR U17277 ( .A(n13180), .B(n13181), .Z(n13177) );
  ANDN U17278 ( .B(n13182), .A(n13183), .Z(n13180) );
  XNOR U17279 ( .A(b[1049]), .B(n13181), .Z(n13182) );
  XNOR U17280 ( .A(b[104]), .B(n13184), .Z(c[104]) );
  XNOR U17281 ( .A(b[1049]), .B(n13183), .Z(c[1049]) );
  XOR U17282 ( .A(n13185), .B(n13186), .Z(n13181) );
  ANDN U17283 ( .B(n13187), .A(n13188), .Z(n13185) );
  XNOR U17284 ( .A(b[1048]), .B(n13186), .Z(n13187) );
  XNOR U17285 ( .A(b[1048]), .B(n13188), .Z(c[1048]) );
  XOR U17286 ( .A(n13189), .B(n13190), .Z(n13186) );
  ANDN U17287 ( .B(n13191), .A(n13192), .Z(n13189) );
  XNOR U17288 ( .A(b[1047]), .B(n13190), .Z(n13191) );
  XNOR U17289 ( .A(b[1047]), .B(n13192), .Z(c[1047]) );
  XOR U17290 ( .A(n13193), .B(n13194), .Z(n13190) );
  ANDN U17291 ( .B(n13195), .A(n13196), .Z(n13193) );
  XNOR U17292 ( .A(b[1046]), .B(n13194), .Z(n13195) );
  XNOR U17293 ( .A(b[1046]), .B(n13196), .Z(c[1046]) );
  XOR U17294 ( .A(n13197), .B(n13198), .Z(n13194) );
  ANDN U17295 ( .B(n13199), .A(n13200), .Z(n13197) );
  XNOR U17296 ( .A(b[1045]), .B(n13198), .Z(n13199) );
  XNOR U17297 ( .A(b[1045]), .B(n13200), .Z(c[1045]) );
  XOR U17298 ( .A(n13201), .B(n13202), .Z(n13198) );
  ANDN U17299 ( .B(n13203), .A(n13204), .Z(n13201) );
  XNOR U17300 ( .A(b[1044]), .B(n13202), .Z(n13203) );
  XNOR U17301 ( .A(b[1044]), .B(n13204), .Z(c[1044]) );
  XOR U17302 ( .A(n13205), .B(n13206), .Z(n13202) );
  ANDN U17303 ( .B(n13207), .A(n13208), .Z(n13205) );
  XNOR U17304 ( .A(b[1043]), .B(n13206), .Z(n13207) );
  XNOR U17305 ( .A(b[1043]), .B(n13208), .Z(c[1043]) );
  XOR U17306 ( .A(n13209), .B(n13210), .Z(n13206) );
  ANDN U17307 ( .B(n13211), .A(n13212), .Z(n13209) );
  XNOR U17308 ( .A(b[1042]), .B(n13210), .Z(n13211) );
  XNOR U17309 ( .A(b[1042]), .B(n13212), .Z(c[1042]) );
  XOR U17310 ( .A(n13213), .B(n13214), .Z(n13210) );
  ANDN U17311 ( .B(n13215), .A(n13216), .Z(n13213) );
  XNOR U17312 ( .A(b[1041]), .B(n13214), .Z(n13215) );
  XNOR U17313 ( .A(b[1041]), .B(n13216), .Z(c[1041]) );
  XOR U17314 ( .A(n13217), .B(n13218), .Z(n13214) );
  ANDN U17315 ( .B(n13219), .A(n13220), .Z(n13217) );
  XNOR U17316 ( .A(b[1040]), .B(n13218), .Z(n13219) );
  XNOR U17317 ( .A(b[1040]), .B(n13220), .Z(c[1040]) );
  XOR U17318 ( .A(n13221), .B(n13222), .Z(n13218) );
  ANDN U17319 ( .B(n13223), .A(n13224), .Z(n13221) );
  XNOR U17320 ( .A(b[1039]), .B(n13222), .Z(n13223) );
  XNOR U17321 ( .A(b[103]), .B(n13225), .Z(c[103]) );
  XNOR U17322 ( .A(b[1039]), .B(n13224), .Z(c[1039]) );
  XOR U17323 ( .A(n13226), .B(n13227), .Z(n13222) );
  ANDN U17324 ( .B(n13228), .A(n13229), .Z(n13226) );
  XNOR U17325 ( .A(b[1038]), .B(n13227), .Z(n13228) );
  XNOR U17326 ( .A(b[1038]), .B(n13229), .Z(c[1038]) );
  XOR U17327 ( .A(n13230), .B(n13231), .Z(n13227) );
  ANDN U17328 ( .B(n13232), .A(n13233), .Z(n13230) );
  XNOR U17329 ( .A(b[1037]), .B(n13231), .Z(n13232) );
  XNOR U17330 ( .A(b[1037]), .B(n13233), .Z(c[1037]) );
  XOR U17331 ( .A(n13234), .B(n13235), .Z(n13231) );
  ANDN U17332 ( .B(n13236), .A(n13237), .Z(n13234) );
  XNOR U17333 ( .A(b[1036]), .B(n13235), .Z(n13236) );
  XNOR U17334 ( .A(b[1036]), .B(n13237), .Z(c[1036]) );
  XOR U17335 ( .A(n13238), .B(n13239), .Z(n13235) );
  ANDN U17336 ( .B(n13240), .A(n13241), .Z(n13238) );
  XNOR U17337 ( .A(b[1035]), .B(n13239), .Z(n13240) );
  XNOR U17338 ( .A(b[1035]), .B(n13241), .Z(c[1035]) );
  XOR U17339 ( .A(n13242), .B(n13243), .Z(n13239) );
  ANDN U17340 ( .B(n13244), .A(n13245), .Z(n13242) );
  XNOR U17341 ( .A(b[1034]), .B(n13243), .Z(n13244) );
  XNOR U17342 ( .A(b[1034]), .B(n13245), .Z(c[1034]) );
  XOR U17343 ( .A(n13246), .B(n13247), .Z(n13243) );
  ANDN U17344 ( .B(n13248), .A(n13249), .Z(n13246) );
  XNOR U17345 ( .A(b[1033]), .B(n13247), .Z(n13248) );
  XNOR U17346 ( .A(b[1033]), .B(n13249), .Z(c[1033]) );
  XOR U17347 ( .A(n13250), .B(n13251), .Z(n13247) );
  ANDN U17348 ( .B(n13252), .A(n13253), .Z(n13250) );
  XNOR U17349 ( .A(b[1032]), .B(n13251), .Z(n13252) );
  XNOR U17350 ( .A(b[1032]), .B(n13253), .Z(c[1032]) );
  XOR U17351 ( .A(n13254), .B(n13255), .Z(n13251) );
  ANDN U17352 ( .B(n13256), .A(n13257), .Z(n13254) );
  XNOR U17353 ( .A(b[1031]), .B(n13255), .Z(n13256) );
  XNOR U17354 ( .A(b[1031]), .B(n13257), .Z(c[1031]) );
  XOR U17355 ( .A(n13258), .B(n13259), .Z(n13255) );
  ANDN U17356 ( .B(n13260), .A(n13261), .Z(n13258) );
  XNOR U17357 ( .A(b[1030]), .B(n13259), .Z(n13260) );
  XNOR U17358 ( .A(b[1030]), .B(n13261), .Z(c[1030]) );
  XOR U17359 ( .A(n13262), .B(n13263), .Z(n13259) );
  ANDN U17360 ( .B(n13264), .A(n13265), .Z(n13262) );
  XNOR U17361 ( .A(b[1029]), .B(n13263), .Z(n13264) );
  XNOR U17362 ( .A(b[102]), .B(n13266), .Z(c[102]) );
  XNOR U17363 ( .A(b[1029]), .B(n13265), .Z(c[1029]) );
  XOR U17364 ( .A(n13267), .B(n13268), .Z(n13263) );
  ANDN U17365 ( .B(n13269), .A(n13270), .Z(n13267) );
  XNOR U17366 ( .A(b[1028]), .B(n13268), .Z(n13269) );
  XNOR U17367 ( .A(b[1028]), .B(n13270), .Z(c[1028]) );
  XOR U17368 ( .A(n13271), .B(n13272), .Z(n13268) );
  ANDN U17369 ( .B(n13273), .A(n13274), .Z(n13271) );
  XNOR U17370 ( .A(b[1027]), .B(n13272), .Z(n13273) );
  XNOR U17371 ( .A(b[1027]), .B(n13274), .Z(c[1027]) );
  XOR U17372 ( .A(n13275), .B(n13276), .Z(n13272) );
  ANDN U17373 ( .B(n13277), .A(n13278), .Z(n13275) );
  XNOR U17374 ( .A(b[1026]), .B(n13276), .Z(n13277) );
  XNOR U17375 ( .A(b[1026]), .B(n13278), .Z(c[1026]) );
  XOR U17376 ( .A(n13279), .B(n13280), .Z(n13276) );
  ANDN U17377 ( .B(n13281), .A(n13282), .Z(n13279) );
  XNOR U17378 ( .A(b[1025]), .B(n13280), .Z(n13281) );
  XNOR U17379 ( .A(b[1025]), .B(n13282), .Z(c[1025]) );
  XOR U17380 ( .A(n13283), .B(n13284), .Z(n13280) );
  ANDN U17381 ( .B(n13285), .A(n13286), .Z(n13283) );
  XNOR U17382 ( .A(b[1024]), .B(n13284), .Z(n13285) );
  XNOR U17383 ( .A(b[1024]), .B(n13286), .Z(c[1024]) );
  XOR U17384 ( .A(n13287), .B(n13288), .Z(n13284) );
  ANDN U17385 ( .B(n13289), .A(n13290), .Z(n13287) );
  XNOR U17386 ( .A(b[1023]), .B(n13288), .Z(n13289) );
  XNOR U17387 ( .A(b[1023]), .B(n13290), .Z(c[1023]) );
  XOR U17388 ( .A(n13291), .B(n13292), .Z(n13288) );
  ANDN U17389 ( .B(n13293), .A(n13294), .Z(n13291) );
  XNOR U17390 ( .A(b[1022]), .B(n13292), .Z(n13293) );
  XNOR U17391 ( .A(b[1022]), .B(n13294), .Z(c[1022]) );
  XOR U17392 ( .A(n13295), .B(n13296), .Z(n13292) );
  ANDN U17393 ( .B(n13297), .A(n13298), .Z(n13295) );
  XNOR U17394 ( .A(b[1021]), .B(n13296), .Z(n13297) );
  XNOR U17395 ( .A(b[1021]), .B(n13298), .Z(c[1021]) );
  XOR U17396 ( .A(n13299), .B(n13300), .Z(n13296) );
  ANDN U17397 ( .B(n13301), .A(n13302), .Z(n13299) );
  XNOR U17398 ( .A(b[1020]), .B(n13300), .Z(n13301) );
  XNOR U17399 ( .A(b[1020]), .B(n13302), .Z(c[1020]) );
  XOR U17400 ( .A(n13303), .B(n13304), .Z(n13300) );
  ANDN U17401 ( .B(n13305), .A(n13306), .Z(n13303) );
  XNOR U17402 ( .A(b[1019]), .B(n13304), .Z(n13305) );
  XNOR U17403 ( .A(b[101]), .B(n13307), .Z(c[101]) );
  XNOR U17404 ( .A(b[1019]), .B(n13306), .Z(c[1019]) );
  XOR U17405 ( .A(n13308), .B(n13309), .Z(n13304) );
  ANDN U17406 ( .B(n13310), .A(n13311), .Z(n13308) );
  XNOR U17407 ( .A(b[1018]), .B(n13309), .Z(n13310) );
  XNOR U17408 ( .A(b[1018]), .B(n13311), .Z(c[1018]) );
  XOR U17409 ( .A(n13312), .B(n13313), .Z(n13309) );
  ANDN U17410 ( .B(n13314), .A(n13315), .Z(n13312) );
  XNOR U17411 ( .A(b[1017]), .B(n13313), .Z(n13314) );
  XNOR U17412 ( .A(b[1017]), .B(n13315), .Z(c[1017]) );
  XOR U17413 ( .A(n13316), .B(n13317), .Z(n13313) );
  ANDN U17414 ( .B(n13318), .A(n13319), .Z(n13316) );
  XNOR U17415 ( .A(b[1016]), .B(n13317), .Z(n13318) );
  XNOR U17416 ( .A(b[1016]), .B(n13319), .Z(c[1016]) );
  XOR U17417 ( .A(n13320), .B(n13321), .Z(n13317) );
  ANDN U17418 ( .B(n13322), .A(n13323), .Z(n13320) );
  XNOR U17419 ( .A(b[1015]), .B(n13321), .Z(n13322) );
  XNOR U17420 ( .A(b[1015]), .B(n13323), .Z(c[1015]) );
  XOR U17421 ( .A(n13324), .B(n13325), .Z(n13321) );
  ANDN U17422 ( .B(n13326), .A(n13327), .Z(n13324) );
  XNOR U17423 ( .A(b[1014]), .B(n13325), .Z(n13326) );
  XNOR U17424 ( .A(b[1014]), .B(n13327), .Z(c[1014]) );
  XOR U17425 ( .A(n13328), .B(n13329), .Z(n13325) );
  ANDN U17426 ( .B(n13330), .A(n13331), .Z(n13328) );
  XNOR U17427 ( .A(b[1013]), .B(n13329), .Z(n13330) );
  XNOR U17428 ( .A(b[1013]), .B(n13331), .Z(c[1013]) );
  XOR U17429 ( .A(n13332), .B(n13333), .Z(n13329) );
  ANDN U17430 ( .B(n13334), .A(n13335), .Z(n13332) );
  XNOR U17431 ( .A(b[1012]), .B(n13333), .Z(n13334) );
  XNOR U17432 ( .A(b[1012]), .B(n13335), .Z(c[1012]) );
  XOR U17433 ( .A(n13336), .B(n13337), .Z(n13333) );
  ANDN U17434 ( .B(n13338), .A(n13339), .Z(n13336) );
  XNOR U17435 ( .A(b[1011]), .B(n13337), .Z(n13338) );
  XNOR U17436 ( .A(b[1011]), .B(n13339), .Z(c[1011]) );
  XOR U17437 ( .A(n13340), .B(n13341), .Z(n13337) );
  ANDN U17438 ( .B(n13342), .A(n13343), .Z(n13340) );
  XNOR U17439 ( .A(b[1010]), .B(n13341), .Z(n13342) );
  XNOR U17440 ( .A(b[1010]), .B(n13343), .Z(c[1010]) );
  XOR U17441 ( .A(n13344), .B(n13345), .Z(n13341) );
  ANDN U17442 ( .B(n13346), .A(n13347), .Z(n13344) );
  XNOR U17443 ( .A(b[1009]), .B(n13345), .Z(n13346) );
  XNOR U17444 ( .A(b[100]), .B(n13348), .Z(c[100]) );
  XNOR U17445 ( .A(b[1009]), .B(n13347), .Z(c[1009]) );
  XOR U17446 ( .A(n13349), .B(n13350), .Z(n13345) );
  ANDN U17447 ( .B(n13351), .A(n13352), .Z(n13349) );
  XNOR U17448 ( .A(b[1008]), .B(n13350), .Z(n13351) );
  XNOR U17449 ( .A(b[1008]), .B(n13352), .Z(c[1008]) );
  XOR U17450 ( .A(n13353), .B(n13354), .Z(n13350) );
  ANDN U17451 ( .B(n13355), .A(n13356), .Z(n13353) );
  XNOR U17452 ( .A(b[1007]), .B(n13354), .Z(n13355) );
  XNOR U17453 ( .A(b[1007]), .B(n13356), .Z(c[1007]) );
  XOR U17454 ( .A(n13357), .B(n13358), .Z(n13354) );
  ANDN U17455 ( .B(n13359), .A(n13360), .Z(n13357) );
  XNOR U17456 ( .A(b[1006]), .B(n13358), .Z(n13359) );
  XNOR U17457 ( .A(b[1006]), .B(n13360), .Z(c[1006]) );
  XOR U17458 ( .A(n13361), .B(n13362), .Z(n13358) );
  ANDN U17459 ( .B(n13363), .A(n13364), .Z(n13361) );
  XNOR U17460 ( .A(b[1005]), .B(n13362), .Z(n13363) );
  XNOR U17461 ( .A(b[1005]), .B(n13364), .Z(c[1005]) );
  XOR U17462 ( .A(n13365), .B(n13366), .Z(n13362) );
  ANDN U17463 ( .B(n13367), .A(n13368), .Z(n13365) );
  XNOR U17464 ( .A(b[1004]), .B(n13366), .Z(n13367) );
  XNOR U17465 ( .A(b[1004]), .B(n13368), .Z(c[1004]) );
  XOR U17466 ( .A(n13369), .B(n13370), .Z(n13366) );
  ANDN U17467 ( .B(n13371), .A(n13372), .Z(n13369) );
  XNOR U17468 ( .A(b[1003]), .B(n13370), .Z(n13371) );
  XNOR U17469 ( .A(b[1003]), .B(n13372), .Z(c[1003]) );
  XOR U17470 ( .A(n13373), .B(n13374), .Z(n13370) );
  ANDN U17471 ( .B(n13375), .A(n13376), .Z(n13373) );
  XNOR U17472 ( .A(b[1002]), .B(n13374), .Z(n13375) );
  XNOR U17473 ( .A(b[1002]), .B(n13376), .Z(c[1002]) );
  XOR U17474 ( .A(n13377), .B(n13378), .Z(n13374) );
  ANDN U17475 ( .B(n13379), .A(n13380), .Z(n13377) );
  XNOR U17476 ( .A(b[1001]), .B(n13378), .Z(n13379) );
  XNOR U17477 ( .A(b[1001]), .B(n13380), .Z(c[1001]) );
  XOR U17478 ( .A(n13381), .B(n13382), .Z(n13378) );
  ANDN U17479 ( .B(n13383), .A(n13384), .Z(n13381) );
  XNOR U17480 ( .A(b[1000]), .B(n13382), .Z(n13383) );
  XNOR U17481 ( .A(b[1000]), .B(n13384), .Z(c[1000]) );
  XOR U17482 ( .A(n13385), .B(n13386), .Z(n13382) );
  ANDN U17483 ( .B(n13387), .A(n8), .Z(n13385) );
  XNOR U17484 ( .A(b[999]), .B(n13386), .Z(n13387) );
  XOR U17485 ( .A(n13388), .B(n13389), .Z(n13386) );
  ANDN U17486 ( .B(n13390), .A(n9), .Z(n13388) );
  XNOR U17487 ( .A(b[998]), .B(n13389), .Z(n13390) );
  XOR U17488 ( .A(n13391), .B(n13392), .Z(n13389) );
  ANDN U17489 ( .B(n13393), .A(n10), .Z(n13391) );
  XNOR U17490 ( .A(b[997]), .B(n13392), .Z(n13393) );
  XOR U17491 ( .A(n13394), .B(n13395), .Z(n13392) );
  ANDN U17492 ( .B(n13396), .A(n11), .Z(n13394) );
  XNOR U17493 ( .A(b[996]), .B(n13395), .Z(n13396) );
  XOR U17494 ( .A(n13397), .B(n13398), .Z(n13395) );
  ANDN U17495 ( .B(n13399), .A(n12), .Z(n13397) );
  XNOR U17496 ( .A(b[995]), .B(n13398), .Z(n13399) );
  XOR U17497 ( .A(n13400), .B(n13401), .Z(n13398) );
  ANDN U17498 ( .B(n13402), .A(n13), .Z(n13400) );
  XNOR U17499 ( .A(b[994]), .B(n13401), .Z(n13402) );
  XOR U17500 ( .A(n13403), .B(n13404), .Z(n13401) );
  ANDN U17501 ( .B(n13405), .A(n14), .Z(n13403) );
  XNOR U17502 ( .A(b[993]), .B(n13404), .Z(n13405) );
  XOR U17503 ( .A(n13406), .B(n13407), .Z(n13404) );
  ANDN U17504 ( .B(n13408), .A(n15), .Z(n13406) );
  XNOR U17505 ( .A(b[992]), .B(n13407), .Z(n13408) );
  XOR U17506 ( .A(n13409), .B(n13410), .Z(n13407) );
  ANDN U17507 ( .B(n13411), .A(n16), .Z(n13409) );
  XNOR U17508 ( .A(b[991]), .B(n13410), .Z(n13411) );
  XOR U17509 ( .A(n13412), .B(n13413), .Z(n13410) );
  ANDN U17510 ( .B(n13414), .A(n17), .Z(n13412) );
  XNOR U17511 ( .A(b[990]), .B(n13413), .Z(n13414) );
  XOR U17512 ( .A(n13415), .B(n13416), .Z(n13413) );
  ANDN U17513 ( .B(n13417), .A(n19), .Z(n13415) );
  XNOR U17514 ( .A(b[989]), .B(n13416), .Z(n13417) );
  XOR U17515 ( .A(n13418), .B(n13419), .Z(n13416) );
  ANDN U17516 ( .B(n13420), .A(n20), .Z(n13418) );
  XNOR U17517 ( .A(b[988]), .B(n13419), .Z(n13420) );
  XOR U17518 ( .A(n13421), .B(n13422), .Z(n13419) );
  ANDN U17519 ( .B(n13423), .A(n21), .Z(n13421) );
  XNOR U17520 ( .A(b[987]), .B(n13422), .Z(n13423) );
  XOR U17521 ( .A(n13424), .B(n13425), .Z(n13422) );
  ANDN U17522 ( .B(n13426), .A(n22), .Z(n13424) );
  XNOR U17523 ( .A(b[986]), .B(n13425), .Z(n13426) );
  XOR U17524 ( .A(n13427), .B(n13428), .Z(n13425) );
  ANDN U17525 ( .B(n13429), .A(n23), .Z(n13427) );
  XNOR U17526 ( .A(b[985]), .B(n13428), .Z(n13429) );
  XOR U17527 ( .A(n13430), .B(n13431), .Z(n13428) );
  ANDN U17528 ( .B(n13432), .A(n24), .Z(n13430) );
  XNOR U17529 ( .A(b[984]), .B(n13431), .Z(n13432) );
  XOR U17530 ( .A(n13433), .B(n13434), .Z(n13431) );
  ANDN U17531 ( .B(n13435), .A(n25), .Z(n13433) );
  XNOR U17532 ( .A(b[983]), .B(n13434), .Z(n13435) );
  XOR U17533 ( .A(n13436), .B(n13437), .Z(n13434) );
  ANDN U17534 ( .B(n13438), .A(n26), .Z(n13436) );
  XNOR U17535 ( .A(b[982]), .B(n13437), .Z(n13438) );
  XOR U17536 ( .A(n13439), .B(n13440), .Z(n13437) );
  ANDN U17537 ( .B(n13441), .A(n27), .Z(n13439) );
  XNOR U17538 ( .A(b[981]), .B(n13440), .Z(n13441) );
  XOR U17539 ( .A(n13442), .B(n13443), .Z(n13440) );
  ANDN U17540 ( .B(n13444), .A(n28), .Z(n13442) );
  XNOR U17541 ( .A(b[980]), .B(n13443), .Z(n13444) );
  XOR U17542 ( .A(n13445), .B(n13446), .Z(n13443) );
  ANDN U17543 ( .B(n13447), .A(n30), .Z(n13445) );
  XNOR U17544 ( .A(b[979]), .B(n13446), .Z(n13447) );
  XOR U17545 ( .A(n13448), .B(n13449), .Z(n13446) );
  ANDN U17546 ( .B(n13450), .A(n31), .Z(n13448) );
  XNOR U17547 ( .A(b[978]), .B(n13449), .Z(n13450) );
  XOR U17548 ( .A(n13451), .B(n13452), .Z(n13449) );
  ANDN U17549 ( .B(n13453), .A(n32), .Z(n13451) );
  XNOR U17550 ( .A(b[977]), .B(n13452), .Z(n13453) );
  XOR U17551 ( .A(n13454), .B(n13455), .Z(n13452) );
  ANDN U17552 ( .B(n13456), .A(n33), .Z(n13454) );
  XNOR U17553 ( .A(b[976]), .B(n13455), .Z(n13456) );
  XOR U17554 ( .A(n13457), .B(n13458), .Z(n13455) );
  ANDN U17555 ( .B(n13459), .A(n34), .Z(n13457) );
  XNOR U17556 ( .A(b[975]), .B(n13458), .Z(n13459) );
  XOR U17557 ( .A(n13460), .B(n13461), .Z(n13458) );
  ANDN U17558 ( .B(n13462), .A(n35), .Z(n13460) );
  XNOR U17559 ( .A(b[974]), .B(n13461), .Z(n13462) );
  XOR U17560 ( .A(n13463), .B(n13464), .Z(n13461) );
  ANDN U17561 ( .B(n13465), .A(n36), .Z(n13463) );
  XNOR U17562 ( .A(b[973]), .B(n13464), .Z(n13465) );
  XOR U17563 ( .A(n13466), .B(n13467), .Z(n13464) );
  ANDN U17564 ( .B(n13468), .A(n37), .Z(n13466) );
  XNOR U17565 ( .A(b[972]), .B(n13467), .Z(n13468) );
  XOR U17566 ( .A(n13469), .B(n13470), .Z(n13467) );
  ANDN U17567 ( .B(n13471), .A(n38), .Z(n13469) );
  XNOR U17568 ( .A(b[971]), .B(n13470), .Z(n13471) );
  XOR U17569 ( .A(n13472), .B(n13473), .Z(n13470) );
  ANDN U17570 ( .B(n13474), .A(n39), .Z(n13472) );
  XNOR U17571 ( .A(b[970]), .B(n13473), .Z(n13474) );
  XOR U17572 ( .A(n13475), .B(n13476), .Z(n13473) );
  ANDN U17573 ( .B(n13477), .A(n41), .Z(n13475) );
  XNOR U17574 ( .A(b[969]), .B(n13476), .Z(n13477) );
  XOR U17575 ( .A(n13478), .B(n13479), .Z(n13476) );
  ANDN U17576 ( .B(n13480), .A(n42), .Z(n13478) );
  XNOR U17577 ( .A(b[968]), .B(n13479), .Z(n13480) );
  XOR U17578 ( .A(n13481), .B(n13482), .Z(n13479) );
  ANDN U17579 ( .B(n13483), .A(n43), .Z(n13481) );
  XNOR U17580 ( .A(b[967]), .B(n13482), .Z(n13483) );
  XOR U17581 ( .A(n13484), .B(n13485), .Z(n13482) );
  ANDN U17582 ( .B(n13486), .A(n44), .Z(n13484) );
  XNOR U17583 ( .A(b[966]), .B(n13485), .Z(n13486) );
  XOR U17584 ( .A(n13487), .B(n13488), .Z(n13485) );
  ANDN U17585 ( .B(n13489), .A(n45), .Z(n13487) );
  XNOR U17586 ( .A(b[965]), .B(n13488), .Z(n13489) );
  XOR U17587 ( .A(n13490), .B(n13491), .Z(n13488) );
  ANDN U17588 ( .B(n13492), .A(n46), .Z(n13490) );
  XNOR U17589 ( .A(b[964]), .B(n13491), .Z(n13492) );
  XOR U17590 ( .A(n13493), .B(n13494), .Z(n13491) );
  ANDN U17591 ( .B(n13495), .A(n47), .Z(n13493) );
  XNOR U17592 ( .A(b[963]), .B(n13494), .Z(n13495) );
  XOR U17593 ( .A(n13496), .B(n13497), .Z(n13494) );
  ANDN U17594 ( .B(n13498), .A(n48), .Z(n13496) );
  XNOR U17595 ( .A(b[962]), .B(n13497), .Z(n13498) );
  XOR U17596 ( .A(n13499), .B(n13500), .Z(n13497) );
  ANDN U17597 ( .B(n13501), .A(n49), .Z(n13499) );
  XNOR U17598 ( .A(b[961]), .B(n13500), .Z(n13501) );
  XOR U17599 ( .A(n13502), .B(n13503), .Z(n13500) );
  ANDN U17600 ( .B(n13504), .A(n50), .Z(n13502) );
  XNOR U17601 ( .A(b[960]), .B(n13503), .Z(n13504) );
  XOR U17602 ( .A(n13505), .B(n13506), .Z(n13503) );
  ANDN U17603 ( .B(n13507), .A(n52), .Z(n13505) );
  XNOR U17604 ( .A(b[959]), .B(n13506), .Z(n13507) );
  XOR U17605 ( .A(n13508), .B(n13509), .Z(n13506) );
  ANDN U17606 ( .B(n13510), .A(n53), .Z(n13508) );
  XNOR U17607 ( .A(b[958]), .B(n13509), .Z(n13510) );
  XOR U17608 ( .A(n13511), .B(n13512), .Z(n13509) );
  ANDN U17609 ( .B(n13513), .A(n54), .Z(n13511) );
  XNOR U17610 ( .A(b[957]), .B(n13512), .Z(n13513) );
  XOR U17611 ( .A(n13514), .B(n13515), .Z(n13512) );
  ANDN U17612 ( .B(n13516), .A(n55), .Z(n13514) );
  XNOR U17613 ( .A(b[956]), .B(n13515), .Z(n13516) );
  XOR U17614 ( .A(n13517), .B(n13518), .Z(n13515) );
  ANDN U17615 ( .B(n13519), .A(n56), .Z(n13517) );
  XNOR U17616 ( .A(b[955]), .B(n13518), .Z(n13519) );
  XOR U17617 ( .A(n13520), .B(n13521), .Z(n13518) );
  ANDN U17618 ( .B(n13522), .A(n57), .Z(n13520) );
  XNOR U17619 ( .A(b[954]), .B(n13521), .Z(n13522) );
  XOR U17620 ( .A(n13523), .B(n13524), .Z(n13521) );
  ANDN U17621 ( .B(n13525), .A(n58), .Z(n13523) );
  XNOR U17622 ( .A(b[953]), .B(n13524), .Z(n13525) );
  XOR U17623 ( .A(n13526), .B(n13527), .Z(n13524) );
  ANDN U17624 ( .B(n13528), .A(n59), .Z(n13526) );
  XNOR U17625 ( .A(b[952]), .B(n13527), .Z(n13528) );
  XOR U17626 ( .A(n13529), .B(n13530), .Z(n13527) );
  ANDN U17627 ( .B(n13531), .A(n60), .Z(n13529) );
  XNOR U17628 ( .A(b[951]), .B(n13530), .Z(n13531) );
  XOR U17629 ( .A(n13532), .B(n13533), .Z(n13530) );
  ANDN U17630 ( .B(n13534), .A(n61), .Z(n13532) );
  XNOR U17631 ( .A(b[950]), .B(n13533), .Z(n13534) );
  XOR U17632 ( .A(n13535), .B(n13536), .Z(n13533) );
  ANDN U17633 ( .B(n13537), .A(n63), .Z(n13535) );
  XNOR U17634 ( .A(b[949]), .B(n13536), .Z(n13537) );
  XOR U17635 ( .A(n13538), .B(n13539), .Z(n13536) );
  ANDN U17636 ( .B(n13540), .A(n64), .Z(n13538) );
  XNOR U17637 ( .A(b[948]), .B(n13539), .Z(n13540) );
  XOR U17638 ( .A(n13541), .B(n13542), .Z(n13539) );
  ANDN U17639 ( .B(n13543), .A(n65), .Z(n13541) );
  XNOR U17640 ( .A(b[947]), .B(n13542), .Z(n13543) );
  XOR U17641 ( .A(n13544), .B(n13545), .Z(n13542) );
  ANDN U17642 ( .B(n13546), .A(n66), .Z(n13544) );
  XNOR U17643 ( .A(b[946]), .B(n13545), .Z(n13546) );
  XOR U17644 ( .A(n13547), .B(n13548), .Z(n13545) );
  ANDN U17645 ( .B(n13549), .A(n67), .Z(n13547) );
  XNOR U17646 ( .A(b[945]), .B(n13548), .Z(n13549) );
  XOR U17647 ( .A(n13550), .B(n13551), .Z(n13548) );
  ANDN U17648 ( .B(n13552), .A(n68), .Z(n13550) );
  XNOR U17649 ( .A(b[944]), .B(n13551), .Z(n13552) );
  XOR U17650 ( .A(n13553), .B(n13554), .Z(n13551) );
  ANDN U17651 ( .B(n13555), .A(n69), .Z(n13553) );
  XNOR U17652 ( .A(b[943]), .B(n13554), .Z(n13555) );
  XOR U17653 ( .A(n13556), .B(n13557), .Z(n13554) );
  ANDN U17654 ( .B(n13558), .A(n70), .Z(n13556) );
  XNOR U17655 ( .A(b[942]), .B(n13557), .Z(n13558) );
  XOR U17656 ( .A(n13559), .B(n13560), .Z(n13557) );
  ANDN U17657 ( .B(n13561), .A(n71), .Z(n13559) );
  XNOR U17658 ( .A(b[941]), .B(n13560), .Z(n13561) );
  XOR U17659 ( .A(n13562), .B(n13563), .Z(n13560) );
  ANDN U17660 ( .B(n13564), .A(n72), .Z(n13562) );
  XNOR U17661 ( .A(b[940]), .B(n13563), .Z(n13564) );
  XOR U17662 ( .A(n13565), .B(n13566), .Z(n13563) );
  ANDN U17663 ( .B(n13567), .A(n74), .Z(n13565) );
  XNOR U17664 ( .A(b[939]), .B(n13566), .Z(n13567) );
  XOR U17665 ( .A(n13568), .B(n13569), .Z(n13566) );
  ANDN U17666 ( .B(n13570), .A(n75), .Z(n13568) );
  XNOR U17667 ( .A(b[938]), .B(n13569), .Z(n13570) );
  XOR U17668 ( .A(n13571), .B(n13572), .Z(n13569) );
  ANDN U17669 ( .B(n13573), .A(n76), .Z(n13571) );
  XNOR U17670 ( .A(b[937]), .B(n13572), .Z(n13573) );
  XOR U17671 ( .A(n13574), .B(n13575), .Z(n13572) );
  ANDN U17672 ( .B(n13576), .A(n77), .Z(n13574) );
  XNOR U17673 ( .A(b[936]), .B(n13575), .Z(n13576) );
  XOR U17674 ( .A(n13577), .B(n13578), .Z(n13575) );
  ANDN U17675 ( .B(n13579), .A(n78), .Z(n13577) );
  XNOR U17676 ( .A(b[935]), .B(n13578), .Z(n13579) );
  XOR U17677 ( .A(n13580), .B(n13581), .Z(n13578) );
  ANDN U17678 ( .B(n13582), .A(n79), .Z(n13580) );
  XNOR U17679 ( .A(b[934]), .B(n13581), .Z(n13582) );
  XOR U17680 ( .A(n13583), .B(n13584), .Z(n13581) );
  ANDN U17681 ( .B(n13585), .A(n80), .Z(n13583) );
  XNOR U17682 ( .A(b[933]), .B(n13584), .Z(n13585) );
  XOR U17683 ( .A(n13586), .B(n13587), .Z(n13584) );
  ANDN U17684 ( .B(n13588), .A(n81), .Z(n13586) );
  XNOR U17685 ( .A(b[932]), .B(n13587), .Z(n13588) );
  XOR U17686 ( .A(n13589), .B(n13590), .Z(n13587) );
  ANDN U17687 ( .B(n13591), .A(n82), .Z(n13589) );
  XNOR U17688 ( .A(b[931]), .B(n13590), .Z(n13591) );
  XOR U17689 ( .A(n13592), .B(n13593), .Z(n13590) );
  ANDN U17690 ( .B(n13594), .A(n83), .Z(n13592) );
  XNOR U17691 ( .A(b[930]), .B(n13593), .Z(n13594) );
  XOR U17692 ( .A(n13595), .B(n13596), .Z(n13593) );
  ANDN U17693 ( .B(n13597), .A(n85), .Z(n13595) );
  XNOR U17694 ( .A(b[929]), .B(n13596), .Z(n13597) );
  XOR U17695 ( .A(n13598), .B(n13599), .Z(n13596) );
  ANDN U17696 ( .B(n13600), .A(n86), .Z(n13598) );
  XNOR U17697 ( .A(b[928]), .B(n13599), .Z(n13600) );
  XOR U17698 ( .A(n13601), .B(n13602), .Z(n13599) );
  ANDN U17699 ( .B(n13603), .A(n87), .Z(n13601) );
  XNOR U17700 ( .A(b[927]), .B(n13602), .Z(n13603) );
  XOR U17701 ( .A(n13604), .B(n13605), .Z(n13602) );
  ANDN U17702 ( .B(n13606), .A(n88), .Z(n13604) );
  XNOR U17703 ( .A(b[926]), .B(n13605), .Z(n13606) );
  XOR U17704 ( .A(n13607), .B(n13608), .Z(n13605) );
  ANDN U17705 ( .B(n13609), .A(n89), .Z(n13607) );
  XNOR U17706 ( .A(b[925]), .B(n13608), .Z(n13609) );
  XOR U17707 ( .A(n13610), .B(n13611), .Z(n13608) );
  ANDN U17708 ( .B(n13612), .A(n90), .Z(n13610) );
  XNOR U17709 ( .A(b[924]), .B(n13611), .Z(n13612) );
  XOR U17710 ( .A(n13613), .B(n13614), .Z(n13611) );
  ANDN U17711 ( .B(n13615), .A(n91), .Z(n13613) );
  XNOR U17712 ( .A(b[923]), .B(n13614), .Z(n13615) );
  XOR U17713 ( .A(n13616), .B(n13617), .Z(n13614) );
  ANDN U17714 ( .B(n13618), .A(n92), .Z(n13616) );
  XNOR U17715 ( .A(b[922]), .B(n13617), .Z(n13618) );
  XOR U17716 ( .A(n13619), .B(n13620), .Z(n13617) );
  ANDN U17717 ( .B(n13621), .A(n93), .Z(n13619) );
  XNOR U17718 ( .A(b[921]), .B(n13620), .Z(n13621) );
  XOR U17719 ( .A(n13622), .B(n13623), .Z(n13620) );
  ANDN U17720 ( .B(n13624), .A(n94), .Z(n13622) );
  XNOR U17721 ( .A(b[920]), .B(n13623), .Z(n13624) );
  XOR U17722 ( .A(n13625), .B(n13626), .Z(n13623) );
  ANDN U17723 ( .B(n13627), .A(n96), .Z(n13625) );
  XNOR U17724 ( .A(b[919]), .B(n13626), .Z(n13627) );
  XOR U17725 ( .A(n13628), .B(n13629), .Z(n13626) );
  ANDN U17726 ( .B(n13630), .A(n97), .Z(n13628) );
  XNOR U17727 ( .A(b[918]), .B(n13629), .Z(n13630) );
  XOR U17728 ( .A(n13631), .B(n13632), .Z(n13629) );
  ANDN U17729 ( .B(n13633), .A(n98), .Z(n13631) );
  XNOR U17730 ( .A(b[917]), .B(n13632), .Z(n13633) );
  XOR U17731 ( .A(n13634), .B(n13635), .Z(n13632) );
  ANDN U17732 ( .B(n13636), .A(n99), .Z(n13634) );
  XNOR U17733 ( .A(b[916]), .B(n13635), .Z(n13636) );
  XOR U17734 ( .A(n13637), .B(n13638), .Z(n13635) );
  ANDN U17735 ( .B(n13639), .A(n100), .Z(n13637) );
  XNOR U17736 ( .A(b[915]), .B(n13638), .Z(n13639) );
  XOR U17737 ( .A(n13640), .B(n13641), .Z(n13638) );
  ANDN U17738 ( .B(n13642), .A(n101), .Z(n13640) );
  XNOR U17739 ( .A(b[914]), .B(n13641), .Z(n13642) );
  XOR U17740 ( .A(n13643), .B(n13644), .Z(n13641) );
  ANDN U17741 ( .B(n13645), .A(n102), .Z(n13643) );
  XNOR U17742 ( .A(b[913]), .B(n13644), .Z(n13645) );
  XOR U17743 ( .A(n13646), .B(n13647), .Z(n13644) );
  ANDN U17744 ( .B(n13648), .A(n103), .Z(n13646) );
  XNOR U17745 ( .A(b[912]), .B(n13647), .Z(n13648) );
  XOR U17746 ( .A(n13649), .B(n13650), .Z(n13647) );
  ANDN U17747 ( .B(n13651), .A(n104), .Z(n13649) );
  XNOR U17748 ( .A(b[911]), .B(n13650), .Z(n13651) );
  XOR U17749 ( .A(n13652), .B(n13653), .Z(n13650) );
  ANDN U17750 ( .B(n13654), .A(n105), .Z(n13652) );
  XNOR U17751 ( .A(b[910]), .B(n13653), .Z(n13654) );
  XOR U17752 ( .A(n13655), .B(n13656), .Z(n13653) );
  ANDN U17753 ( .B(n13657), .A(n107), .Z(n13655) );
  XNOR U17754 ( .A(b[909]), .B(n13656), .Z(n13657) );
  XOR U17755 ( .A(n13658), .B(n13659), .Z(n13656) );
  ANDN U17756 ( .B(n13660), .A(n108), .Z(n13658) );
  XNOR U17757 ( .A(b[908]), .B(n13659), .Z(n13660) );
  XOR U17758 ( .A(n13661), .B(n13662), .Z(n13659) );
  ANDN U17759 ( .B(n13663), .A(n109), .Z(n13661) );
  XNOR U17760 ( .A(b[907]), .B(n13662), .Z(n13663) );
  XOR U17761 ( .A(n13664), .B(n13665), .Z(n13662) );
  ANDN U17762 ( .B(n13666), .A(n110), .Z(n13664) );
  XNOR U17763 ( .A(b[906]), .B(n13665), .Z(n13666) );
  XOR U17764 ( .A(n13667), .B(n13668), .Z(n13665) );
  ANDN U17765 ( .B(n13669), .A(n111), .Z(n13667) );
  XNOR U17766 ( .A(b[905]), .B(n13668), .Z(n13669) );
  XOR U17767 ( .A(n13670), .B(n13671), .Z(n13668) );
  ANDN U17768 ( .B(n13672), .A(n112), .Z(n13670) );
  XNOR U17769 ( .A(b[904]), .B(n13671), .Z(n13672) );
  XOR U17770 ( .A(n13673), .B(n13674), .Z(n13671) );
  ANDN U17771 ( .B(n13675), .A(n113), .Z(n13673) );
  XNOR U17772 ( .A(b[903]), .B(n13674), .Z(n13675) );
  XOR U17773 ( .A(n13676), .B(n13677), .Z(n13674) );
  ANDN U17774 ( .B(n13678), .A(n114), .Z(n13676) );
  XNOR U17775 ( .A(b[902]), .B(n13677), .Z(n13678) );
  XOR U17776 ( .A(n13679), .B(n13680), .Z(n13677) );
  ANDN U17777 ( .B(n13681), .A(n115), .Z(n13679) );
  XNOR U17778 ( .A(b[901]), .B(n13680), .Z(n13681) );
  XOR U17779 ( .A(n13682), .B(n13683), .Z(n13680) );
  ANDN U17780 ( .B(n13684), .A(n116), .Z(n13682) );
  XNOR U17781 ( .A(b[900]), .B(n13683), .Z(n13684) );
  XOR U17782 ( .A(n13685), .B(n13686), .Z(n13683) );
  ANDN U17783 ( .B(n13687), .A(n119), .Z(n13685) );
  XNOR U17784 ( .A(b[899]), .B(n13686), .Z(n13687) );
  XOR U17785 ( .A(n13688), .B(n13689), .Z(n13686) );
  ANDN U17786 ( .B(n13690), .A(n120), .Z(n13688) );
  XNOR U17787 ( .A(b[898]), .B(n13689), .Z(n13690) );
  XOR U17788 ( .A(n13691), .B(n13692), .Z(n13689) );
  ANDN U17789 ( .B(n13693), .A(n121), .Z(n13691) );
  XNOR U17790 ( .A(b[897]), .B(n13692), .Z(n13693) );
  XOR U17791 ( .A(n13694), .B(n13695), .Z(n13692) );
  ANDN U17792 ( .B(n13696), .A(n122), .Z(n13694) );
  XNOR U17793 ( .A(b[896]), .B(n13695), .Z(n13696) );
  XOR U17794 ( .A(n13697), .B(n13698), .Z(n13695) );
  ANDN U17795 ( .B(n13699), .A(n123), .Z(n13697) );
  XNOR U17796 ( .A(b[895]), .B(n13698), .Z(n13699) );
  XOR U17797 ( .A(n13700), .B(n13701), .Z(n13698) );
  ANDN U17798 ( .B(n13702), .A(n124), .Z(n13700) );
  XNOR U17799 ( .A(b[894]), .B(n13701), .Z(n13702) );
  XOR U17800 ( .A(n13703), .B(n13704), .Z(n13701) );
  ANDN U17801 ( .B(n13705), .A(n125), .Z(n13703) );
  XNOR U17802 ( .A(b[893]), .B(n13704), .Z(n13705) );
  XOR U17803 ( .A(n13706), .B(n13707), .Z(n13704) );
  ANDN U17804 ( .B(n13708), .A(n126), .Z(n13706) );
  XNOR U17805 ( .A(b[892]), .B(n13707), .Z(n13708) );
  XOR U17806 ( .A(n13709), .B(n13710), .Z(n13707) );
  ANDN U17807 ( .B(n13711), .A(n127), .Z(n13709) );
  XNOR U17808 ( .A(b[891]), .B(n13710), .Z(n13711) );
  XOR U17809 ( .A(n13712), .B(n13713), .Z(n13710) );
  ANDN U17810 ( .B(n13714), .A(n128), .Z(n13712) );
  XNOR U17811 ( .A(b[890]), .B(n13713), .Z(n13714) );
  XOR U17812 ( .A(n13715), .B(n13716), .Z(n13713) );
  ANDN U17813 ( .B(n13717), .A(n130), .Z(n13715) );
  XNOR U17814 ( .A(b[889]), .B(n13716), .Z(n13717) );
  XOR U17815 ( .A(n13718), .B(n13719), .Z(n13716) );
  ANDN U17816 ( .B(n13720), .A(n131), .Z(n13718) );
  XNOR U17817 ( .A(b[888]), .B(n13719), .Z(n13720) );
  XOR U17818 ( .A(n13721), .B(n13722), .Z(n13719) );
  ANDN U17819 ( .B(n13723), .A(n132), .Z(n13721) );
  XNOR U17820 ( .A(b[887]), .B(n13722), .Z(n13723) );
  XOR U17821 ( .A(n13724), .B(n13725), .Z(n13722) );
  ANDN U17822 ( .B(n13726), .A(n133), .Z(n13724) );
  XNOR U17823 ( .A(b[886]), .B(n13725), .Z(n13726) );
  XOR U17824 ( .A(n13727), .B(n13728), .Z(n13725) );
  ANDN U17825 ( .B(n13729), .A(n134), .Z(n13727) );
  XNOR U17826 ( .A(b[885]), .B(n13728), .Z(n13729) );
  XOR U17827 ( .A(n13730), .B(n13731), .Z(n13728) );
  ANDN U17828 ( .B(n13732), .A(n135), .Z(n13730) );
  XNOR U17829 ( .A(b[884]), .B(n13731), .Z(n13732) );
  XOR U17830 ( .A(n13733), .B(n13734), .Z(n13731) );
  ANDN U17831 ( .B(n13735), .A(n136), .Z(n13733) );
  XNOR U17832 ( .A(b[883]), .B(n13734), .Z(n13735) );
  XOR U17833 ( .A(n13736), .B(n13737), .Z(n13734) );
  ANDN U17834 ( .B(n13738), .A(n137), .Z(n13736) );
  XNOR U17835 ( .A(b[882]), .B(n13737), .Z(n13738) );
  XOR U17836 ( .A(n13739), .B(n13740), .Z(n13737) );
  ANDN U17837 ( .B(n13741), .A(n138), .Z(n13739) );
  XNOR U17838 ( .A(b[881]), .B(n13740), .Z(n13741) );
  XOR U17839 ( .A(n13742), .B(n13743), .Z(n13740) );
  ANDN U17840 ( .B(n13744), .A(n139), .Z(n13742) );
  XNOR U17841 ( .A(b[880]), .B(n13743), .Z(n13744) );
  XOR U17842 ( .A(n13745), .B(n13746), .Z(n13743) );
  ANDN U17843 ( .B(n13747), .A(n141), .Z(n13745) );
  XNOR U17844 ( .A(b[879]), .B(n13746), .Z(n13747) );
  XOR U17845 ( .A(n13748), .B(n13749), .Z(n13746) );
  ANDN U17846 ( .B(n13750), .A(n142), .Z(n13748) );
  XNOR U17847 ( .A(b[878]), .B(n13749), .Z(n13750) );
  XOR U17848 ( .A(n13751), .B(n13752), .Z(n13749) );
  ANDN U17849 ( .B(n13753), .A(n143), .Z(n13751) );
  XNOR U17850 ( .A(b[877]), .B(n13752), .Z(n13753) );
  XOR U17851 ( .A(n13754), .B(n13755), .Z(n13752) );
  ANDN U17852 ( .B(n13756), .A(n144), .Z(n13754) );
  XNOR U17853 ( .A(b[876]), .B(n13755), .Z(n13756) );
  XOR U17854 ( .A(n13757), .B(n13758), .Z(n13755) );
  ANDN U17855 ( .B(n13759), .A(n145), .Z(n13757) );
  XNOR U17856 ( .A(b[875]), .B(n13758), .Z(n13759) );
  XOR U17857 ( .A(n13760), .B(n13761), .Z(n13758) );
  ANDN U17858 ( .B(n13762), .A(n146), .Z(n13760) );
  XNOR U17859 ( .A(b[874]), .B(n13761), .Z(n13762) );
  XOR U17860 ( .A(n13763), .B(n13764), .Z(n13761) );
  ANDN U17861 ( .B(n13765), .A(n147), .Z(n13763) );
  XNOR U17862 ( .A(b[873]), .B(n13764), .Z(n13765) );
  XOR U17863 ( .A(n13766), .B(n13767), .Z(n13764) );
  ANDN U17864 ( .B(n13768), .A(n148), .Z(n13766) );
  XNOR U17865 ( .A(b[872]), .B(n13767), .Z(n13768) );
  XOR U17866 ( .A(n13769), .B(n13770), .Z(n13767) );
  ANDN U17867 ( .B(n13771), .A(n149), .Z(n13769) );
  XNOR U17868 ( .A(b[871]), .B(n13770), .Z(n13771) );
  XOR U17869 ( .A(n13772), .B(n13773), .Z(n13770) );
  ANDN U17870 ( .B(n13774), .A(n150), .Z(n13772) );
  XNOR U17871 ( .A(b[870]), .B(n13773), .Z(n13774) );
  XOR U17872 ( .A(n13775), .B(n13776), .Z(n13773) );
  ANDN U17873 ( .B(n13777), .A(n152), .Z(n13775) );
  XNOR U17874 ( .A(b[869]), .B(n13776), .Z(n13777) );
  XOR U17875 ( .A(n13778), .B(n13779), .Z(n13776) );
  ANDN U17876 ( .B(n13780), .A(n153), .Z(n13778) );
  XNOR U17877 ( .A(b[868]), .B(n13779), .Z(n13780) );
  XOR U17878 ( .A(n13781), .B(n13782), .Z(n13779) );
  ANDN U17879 ( .B(n13783), .A(n154), .Z(n13781) );
  XNOR U17880 ( .A(b[867]), .B(n13782), .Z(n13783) );
  XOR U17881 ( .A(n13784), .B(n13785), .Z(n13782) );
  ANDN U17882 ( .B(n13786), .A(n155), .Z(n13784) );
  XNOR U17883 ( .A(b[866]), .B(n13785), .Z(n13786) );
  XOR U17884 ( .A(n13787), .B(n13788), .Z(n13785) );
  ANDN U17885 ( .B(n13789), .A(n156), .Z(n13787) );
  XNOR U17886 ( .A(b[865]), .B(n13788), .Z(n13789) );
  XOR U17887 ( .A(n13790), .B(n13791), .Z(n13788) );
  ANDN U17888 ( .B(n13792), .A(n157), .Z(n13790) );
  XNOR U17889 ( .A(b[864]), .B(n13791), .Z(n13792) );
  XOR U17890 ( .A(n13793), .B(n13794), .Z(n13791) );
  ANDN U17891 ( .B(n13795), .A(n158), .Z(n13793) );
  XNOR U17892 ( .A(b[863]), .B(n13794), .Z(n13795) );
  XOR U17893 ( .A(n13796), .B(n13797), .Z(n13794) );
  ANDN U17894 ( .B(n13798), .A(n159), .Z(n13796) );
  XNOR U17895 ( .A(b[862]), .B(n13797), .Z(n13798) );
  XOR U17896 ( .A(n13799), .B(n13800), .Z(n13797) );
  ANDN U17897 ( .B(n13801), .A(n160), .Z(n13799) );
  XNOR U17898 ( .A(b[861]), .B(n13800), .Z(n13801) );
  XOR U17899 ( .A(n13802), .B(n13803), .Z(n13800) );
  ANDN U17900 ( .B(n13804), .A(n161), .Z(n13802) );
  XNOR U17901 ( .A(b[860]), .B(n13803), .Z(n13804) );
  XOR U17902 ( .A(n13805), .B(n13806), .Z(n13803) );
  ANDN U17903 ( .B(n13807), .A(n163), .Z(n13805) );
  XNOR U17904 ( .A(b[859]), .B(n13806), .Z(n13807) );
  XOR U17905 ( .A(n13808), .B(n13809), .Z(n13806) );
  ANDN U17906 ( .B(n13810), .A(n164), .Z(n13808) );
  XNOR U17907 ( .A(b[858]), .B(n13809), .Z(n13810) );
  XOR U17908 ( .A(n13811), .B(n13812), .Z(n13809) );
  ANDN U17909 ( .B(n13813), .A(n165), .Z(n13811) );
  XNOR U17910 ( .A(b[857]), .B(n13812), .Z(n13813) );
  XOR U17911 ( .A(n13814), .B(n13815), .Z(n13812) );
  ANDN U17912 ( .B(n13816), .A(n166), .Z(n13814) );
  XNOR U17913 ( .A(b[856]), .B(n13815), .Z(n13816) );
  XOR U17914 ( .A(n13817), .B(n13818), .Z(n13815) );
  ANDN U17915 ( .B(n13819), .A(n167), .Z(n13817) );
  XNOR U17916 ( .A(b[855]), .B(n13818), .Z(n13819) );
  XOR U17917 ( .A(n13820), .B(n13821), .Z(n13818) );
  ANDN U17918 ( .B(n13822), .A(n168), .Z(n13820) );
  XNOR U17919 ( .A(b[854]), .B(n13821), .Z(n13822) );
  XOR U17920 ( .A(n13823), .B(n13824), .Z(n13821) );
  ANDN U17921 ( .B(n13825), .A(n169), .Z(n13823) );
  XNOR U17922 ( .A(b[853]), .B(n13824), .Z(n13825) );
  XOR U17923 ( .A(n13826), .B(n13827), .Z(n13824) );
  ANDN U17924 ( .B(n13828), .A(n170), .Z(n13826) );
  XNOR U17925 ( .A(b[852]), .B(n13827), .Z(n13828) );
  XOR U17926 ( .A(n13829), .B(n13830), .Z(n13827) );
  ANDN U17927 ( .B(n13831), .A(n171), .Z(n13829) );
  XNOR U17928 ( .A(b[851]), .B(n13830), .Z(n13831) );
  XOR U17929 ( .A(n13832), .B(n13833), .Z(n13830) );
  ANDN U17930 ( .B(n13834), .A(n172), .Z(n13832) );
  XNOR U17931 ( .A(b[850]), .B(n13833), .Z(n13834) );
  XOR U17932 ( .A(n13835), .B(n13836), .Z(n13833) );
  ANDN U17933 ( .B(n13837), .A(n174), .Z(n13835) );
  XNOR U17934 ( .A(b[849]), .B(n13836), .Z(n13837) );
  XOR U17935 ( .A(n13838), .B(n13839), .Z(n13836) );
  ANDN U17936 ( .B(n13840), .A(n175), .Z(n13838) );
  XNOR U17937 ( .A(b[848]), .B(n13839), .Z(n13840) );
  XOR U17938 ( .A(n13841), .B(n13842), .Z(n13839) );
  ANDN U17939 ( .B(n13843), .A(n176), .Z(n13841) );
  XNOR U17940 ( .A(b[847]), .B(n13842), .Z(n13843) );
  XOR U17941 ( .A(n13844), .B(n13845), .Z(n13842) );
  ANDN U17942 ( .B(n13846), .A(n177), .Z(n13844) );
  XNOR U17943 ( .A(b[846]), .B(n13845), .Z(n13846) );
  XOR U17944 ( .A(n13847), .B(n13848), .Z(n13845) );
  ANDN U17945 ( .B(n13849), .A(n178), .Z(n13847) );
  XNOR U17946 ( .A(b[845]), .B(n13848), .Z(n13849) );
  XOR U17947 ( .A(n13850), .B(n13851), .Z(n13848) );
  ANDN U17948 ( .B(n13852), .A(n179), .Z(n13850) );
  XNOR U17949 ( .A(b[844]), .B(n13851), .Z(n13852) );
  XOR U17950 ( .A(n13853), .B(n13854), .Z(n13851) );
  ANDN U17951 ( .B(n13855), .A(n180), .Z(n13853) );
  XNOR U17952 ( .A(b[843]), .B(n13854), .Z(n13855) );
  XOR U17953 ( .A(n13856), .B(n13857), .Z(n13854) );
  ANDN U17954 ( .B(n13858), .A(n181), .Z(n13856) );
  XNOR U17955 ( .A(b[842]), .B(n13857), .Z(n13858) );
  XOR U17956 ( .A(n13859), .B(n13860), .Z(n13857) );
  ANDN U17957 ( .B(n13861), .A(n182), .Z(n13859) );
  XNOR U17958 ( .A(b[841]), .B(n13860), .Z(n13861) );
  XOR U17959 ( .A(n13862), .B(n13863), .Z(n13860) );
  ANDN U17960 ( .B(n13864), .A(n183), .Z(n13862) );
  XNOR U17961 ( .A(b[840]), .B(n13863), .Z(n13864) );
  XOR U17962 ( .A(n13865), .B(n13866), .Z(n13863) );
  ANDN U17963 ( .B(n13867), .A(n185), .Z(n13865) );
  XNOR U17964 ( .A(b[839]), .B(n13866), .Z(n13867) );
  XOR U17965 ( .A(n13868), .B(n13869), .Z(n13866) );
  ANDN U17966 ( .B(n13870), .A(n186), .Z(n13868) );
  XNOR U17967 ( .A(b[838]), .B(n13869), .Z(n13870) );
  XOR U17968 ( .A(n13871), .B(n13872), .Z(n13869) );
  ANDN U17969 ( .B(n13873), .A(n187), .Z(n13871) );
  XNOR U17970 ( .A(b[837]), .B(n13872), .Z(n13873) );
  XOR U17971 ( .A(n13874), .B(n13875), .Z(n13872) );
  ANDN U17972 ( .B(n13876), .A(n188), .Z(n13874) );
  XNOR U17973 ( .A(b[836]), .B(n13875), .Z(n13876) );
  XOR U17974 ( .A(n13877), .B(n13878), .Z(n13875) );
  ANDN U17975 ( .B(n13879), .A(n189), .Z(n13877) );
  XNOR U17976 ( .A(b[835]), .B(n13878), .Z(n13879) );
  XOR U17977 ( .A(n13880), .B(n13881), .Z(n13878) );
  ANDN U17978 ( .B(n13882), .A(n190), .Z(n13880) );
  XNOR U17979 ( .A(b[834]), .B(n13881), .Z(n13882) );
  XOR U17980 ( .A(n13883), .B(n13884), .Z(n13881) );
  ANDN U17981 ( .B(n13885), .A(n191), .Z(n13883) );
  XNOR U17982 ( .A(b[833]), .B(n13884), .Z(n13885) );
  XOR U17983 ( .A(n13886), .B(n13887), .Z(n13884) );
  ANDN U17984 ( .B(n13888), .A(n192), .Z(n13886) );
  XNOR U17985 ( .A(b[832]), .B(n13887), .Z(n13888) );
  XOR U17986 ( .A(n13889), .B(n13890), .Z(n13887) );
  ANDN U17987 ( .B(n13891), .A(n193), .Z(n13889) );
  XNOR U17988 ( .A(b[831]), .B(n13890), .Z(n13891) );
  XOR U17989 ( .A(n13892), .B(n13893), .Z(n13890) );
  ANDN U17990 ( .B(n13894), .A(n194), .Z(n13892) );
  XNOR U17991 ( .A(b[830]), .B(n13893), .Z(n13894) );
  XOR U17992 ( .A(n13895), .B(n13896), .Z(n13893) );
  ANDN U17993 ( .B(n13897), .A(n196), .Z(n13895) );
  XNOR U17994 ( .A(b[829]), .B(n13896), .Z(n13897) );
  XOR U17995 ( .A(n13898), .B(n13899), .Z(n13896) );
  ANDN U17996 ( .B(n13900), .A(n197), .Z(n13898) );
  XNOR U17997 ( .A(b[828]), .B(n13899), .Z(n13900) );
  XOR U17998 ( .A(n13901), .B(n13902), .Z(n13899) );
  ANDN U17999 ( .B(n13903), .A(n198), .Z(n13901) );
  XNOR U18000 ( .A(b[827]), .B(n13902), .Z(n13903) );
  XOR U18001 ( .A(n13904), .B(n13905), .Z(n13902) );
  ANDN U18002 ( .B(n13906), .A(n199), .Z(n13904) );
  XNOR U18003 ( .A(b[826]), .B(n13905), .Z(n13906) );
  XOR U18004 ( .A(n13907), .B(n13908), .Z(n13905) );
  ANDN U18005 ( .B(n13909), .A(n200), .Z(n13907) );
  XNOR U18006 ( .A(b[825]), .B(n13908), .Z(n13909) );
  XOR U18007 ( .A(n13910), .B(n13911), .Z(n13908) );
  ANDN U18008 ( .B(n13912), .A(n201), .Z(n13910) );
  XNOR U18009 ( .A(b[824]), .B(n13911), .Z(n13912) );
  XOR U18010 ( .A(n13913), .B(n13914), .Z(n13911) );
  ANDN U18011 ( .B(n13915), .A(n202), .Z(n13913) );
  XNOR U18012 ( .A(b[823]), .B(n13914), .Z(n13915) );
  XOR U18013 ( .A(n13916), .B(n13917), .Z(n13914) );
  ANDN U18014 ( .B(n13918), .A(n203), .Z(n13916) );
  XNOR U18015 ( .A(b[822]), .B(n13917), .Z(n13918) );
  XOR U18016 ( .A(n13919), .B(n13920), .Z(n13917) );
  ANDN U18017 ( .B(n13921), .A(n204), .Z(n13919) );
  XNOR U18018 ( .A(b[821]), .B(n13920), .Z(n13921) );
  XOR U18019 ( .A(n13922), .B(n13923), .Z(n13920) );
  ANDN U18020 ( .B(n13924), .A(n205), .Z(n13922) );
  XNOR U18021 ( .A(b[820]), .B(n13923), .Z(n13924) );
  XOR U18022 ( .A(n13925), .B(n13926), .Z(n13923) );
  ANDN U18023 ( .B(n13927), .A(n207), .Z(n13925) );
  XNOR U18024 ( .A(b[819]), .B(n13926), .Z(n13927) );
  XOR U18025 ( .A(n13928), .B(n13929), .Z(n13926) );
  ANDN U18026 ( .B(n13930), .A(n208), .Z(n13928) );
  XNOR U18027 ( .A(b[818]), .B(n13929), .Z(n13930) );
  XOR U18028 ( .A(n13931), .B(n13932), .Z(n13929) );
  ANDN U18029 ( .B(n13933), .A(n209), .Z(n13931) );
  XNOR U18030 ( .A(b[817]), .B(n13932), .Z(n13933) );
  XOR U18031 ( .A(n13934), .B(n13935), .Z(n13932) );
  ANDN U18032 ( .B(n13936), .A(n210), .Z(n13934) );
  XNOR U18033 ( .A(b[816]), .B(n13935), .Z(n13936) );
  XOR U18034 ( .A(n13937), .B(n13938), .Z(n13935) );
  ANDN U18035 ( .B(n13939), .A(n211), .Z(n13937) );
  XNOR U18036 ( .A(b[815]), .B(n13938), .Z(n13939) );
  XOR U18037 ( .A(n13940), .B(n13941), .Z(n13938) );
  ANDN U18038 ( .B(n13942), .A(n212), .Z(n13940) );
  XNOR U18039 ( .A(b[814]), .B(n13941), .Z(n13942) );
  XOR U18040 ( .A(n13943), .B(n13944), .Z(n13941) );
  ANDN U18041 ( .B(n13945), .A(n213), .Z(n13943) );
  XNOR U18042 ( .A(b[813]), .B(n13944), .Z(n13945) );
  XOR U18043 ( .A(n13946), .B(n13947), .Z(n13944) );
  ANDN U18044 ( .B(n13948), .A(n214), .Z(n13946) );
  XNOR U18045 ( .A(b[812]), .B(n13947), .Z(n13948) );
  XOR U18046 ( .A(n13949), .B(n13950), .Z(n13947) );
  ANDN U18047 ( .B(n13951), .A(n215), .Z(n13949) );
  XNOR U18048 ( .A(b[811]), .B(n13950), .Z(n13951) );
  XOR U18049 ( .A(n13952), .B(n13953), .Z(n13950) );
  ANDN U18050 ( .B(n13954), .A(n216), .Z(n13952) );
  XNOR U18051 ( .A(b[810]), .B(n13953), .Z(n13954) );
  XOR U18052 ( .A(n13955), .B(n13956), .Z(n13953) );
  ANDN U18053 ( .B(n13957), .A(n218), .Z(n13955) );
  XNOR U18054 ( .A(b[809]), .B(n13956), .Z(n13957) );
  XOR U18055 ( .A(n13958), .B(n13959), .Z(n13956) );
  ANDN U18056 ( .B(n13960), .A(n219), .Z(n13958) );
  XNOR U18057 ( .A(b[808]), .B(n13959), .Z(n13960) );
  XOR U18058 ( .A(n13961), .B(n13962), .Z(n13959) );
  ANDN U18059 ( .B(n13963), .A(n220), .Z(n13961) );
  XNOR U18060 ( .A(b[807]), .B(n13962), .Z(n13963) );
  XOR U18061 ( .A(n13964), .B(n13965), .Z(n13962) );
  ANDN U18062 ( .B(n13966), .A(n221), .Z(n13964) );
  XNOR U18063 ( .A(b[806]), .B(n13965), .Z(n13966) );
  XOR U18064 ( .A(n13967), .B(n13968), .Z(n13965) );
  ANDN U18065 ( .B(n13969), .A(n222), .Z(n13967) );
  XNOR U18066 ( .A(b[805]), .B(n13968), .Z(n13969) );
  XOR U18067 ( .A(n13970), .B(n13971), .Z(n13968) );
  ANDN U18068 ( .B(n13972), .A(n223), .Z(n13970) );
  XNOR U18069 ( .A(b[804]), .B(n13971), .Z(n13972) );
  XOR U18070 ( .A(n13973), .B(n13974), .Z(n13971) );
  ANDN U18071 ( .B(n13975), .A(n224), .Z(n13973) );
  XNOR U18072 ( .A(b[803]), .B(n13974), .Z(n13975) );
  XOR U18073 ( .A(n13976), .B(n13977), .Z(n13974) );
  ANDN U18074 ( .B(n13978), .A(n225), .Z(n13976) );
  XNOR U18075 ( .A(b[802]), .B(n13977), .Z(n13978) );
  XOR U18076 ( .A(n13979), .B(n13980), .Z(n13977) );
  ANDN U18077 ( .B(n13981), .A(n226), .Z(n13979) );
  XNOR U18078 ( .A(b[801]), .B(n13980), .Z(n13981) );
  XOR U18079 ( .A(n13982), .B(n13983), .Z(n13980) );
  ANDN U18080 ( .B(n13984), .A(n227), .Z(n13982) );
  XNOR U18081 ( .A(b[800]), .B(n13983), .Z(n13984) );
  XOR U18082 ( .A(n13985), .B(n13986), .Z(n13983) );
  ANDN U18083 ( .B(n13987), .A(n230), .Z(n13985) );
  XNOR U18084 ( .A(b[799]), .B(n13986), .Z(n13987) );
  XOR U18085 ( .A(n13988), .B(n13989), .Z(n13986) );
  ANDN U18086 ( .B(n13990), .A(n231), .Z(n13988) );
  XNOR U18087 ( .A(b[798]), .B(n13989), .Z(n13990) );
  XOR U18088 ( .A(n13991), .B(n13992), .Z(n13989) );
  ANDN U18089 ( .B(n13993), .A(n232), .Z(n13991) );
  XNOR U18090 ( .A(b[797]), .B(n13992), .Z(n13993) );
  XOR U18091 ( .A(n13994), .B(n13995), .Z(n13992) );
  ANDN U18092 ( .B(n13996), .A(n233), .Z(n13994) );
  XNOR U18093 ( .A(b[796]), .B(n13995), .Z(n13996) );
  XOR U18094 ( .A(n13997), .B(n13998), .Z(n13995) );
  ANDN U18095 ( .B(n13999), .A(n234), .Z(n13997) );
  XNOR U18096 ( .A(b[795]), .B(n13998), .Z(n13999) );
  XOR U18097 ( .A(n14000), .B(n14001), .Z(n13998) );
  ANDN U18098 ( .B(n14002), .A(n235), .Z(n14000) );
  XNOR U18099 ( .A(b[794]), .B(n14001), .Z(n14002) );
  XOR U18100 ( .A(n14003), .B(n14004), .Z(n14001) );
  ANDN U18101 ( .B(n14005), .A(n236), .Z(n14003) );
  XNOR U18102 ( .A(b[793]), .B(n14004), .Z(n14005) );
  XOR U18103 ( .A(n14006), .B(n14007), .Z(n14004) );
  ANDN U18104 ( .B(n14008), .A(n237), .Z(n14006) );
  XNOR U18105 ( .A(b[792]), .B(n14007), .Z(n14008) );
  XOR U18106 ( .A(n14009), .B(n14010), .Z(n14007) );
  ANDN U18107 ( .B(n14011), .A(n238), .Z(n14009) );
  XNOR U18108 ( .A(b[791]), .B(n14010), .Z(n14011) );
  XOR U18109 ( .A(n14012), .B(n14013), .Z(n14010) );
  ANDN U18110 ( .B(n14014), .A(n239), .Z(n14012) );
  XNOR U18111 ( .A(b[790]), .B(n14013), .Z(n14014) );
  XOR U18112 ( .A(n14015), .B(n14016), .Z(n14013) );
  ANDN U18113 ( .B(n14017), .A(n241), .Z(n14015) );
  XNOR U18114 ( .A(b[789]), .B(n14016), .Z(n14017) );
  XOR U18115 ( .A(n14018), .B(n14019), .Z(n14016) );
  ANDN U18116 ( .B(n14020), .A(n242), .Z(n14018) );
  XNOR U18117 ( .A(b[788]), .B(n14019), .Z(n14020) );
  XOR U18118 ( .A(n14021), .B(n14022), .Z(n14019) );
  ANDN U18119 ( .B(n14023), .A(n243), .Z(n14021) );
  XNOR U18120 ( .A(b[787]), .B(n14022), .Z(n14023) );
  XOR U18121 ( .A(n14024), .B(n14025), .Z(n14022) );
  ANDN U18122 ( .B(n14026), .A(n244), .Z(n14024) );
  XNOR U18123 ( .A(b[786]), .B(n14025), .Z(n14026) );
  XOR U18124 ( .A(n14027), .B(n14028), .Z(n14025) );
  ANDN U18125 ( .B(n14029), .A(n245), .Z(n14027) );
  XNOR U18126 ( .A(b[785]), .B(n14028), .Z(n14029) );
  XOR U18127 ( .A(n14030), .B(n14031), .Z(n14028) );
  ANDN U18128 ( .B(n14032), .A(n246), .Z(n14030) );
  XNOR U18129 ( .A(b[784]), .B(n14031), .Z(n14032) );
  XOR U18130 ( .A(n14033), .B(n14034), .Z(n14031) );
  ANDN U18131 ( .B(n14035), .A(n247), .Z(n14033) );
  XNOR U18132 ( .A(b[783]), .B(n14034), .Z(n14035) );
  XOR U18133 ( .A(n14036), .B(n14037), .Z(n14034) );
  ANDN U18134 ( .B(n14038), .A(n248), .Z(n14036) );
  XNOR U18135 ( .A(b[782]), .B(n14037), .Z(n14038) );
  XOR U18136 ( .A(n14039), .B(n14040), .Z(n14037) );
  ANDN U18137 ( .B(n14041), .A(n249), .Z(n14039) );
  XNOR U18138 ( .A(b[781]), .B(n14040), .Z(n14041) );
  XOR U18139 ( .A(n14042), .B(n14043), .Z(n14040) );
  ANDN U18140 ( .B(n14044), .A(n250), .Z(n14042) );
  XNOR U18141 ( .A(b[780]), .B(n14043), .Z(n14044) );
  XOR U18142 ( .A(n14045), .B(n14046), .Z(n14043) );
  ANDN U18143 ( .B(n14047), .A(n252), .Z(n14045) );
  XNOR U18144 ( .A(b[779]), .B(n14046), .Z(n14047) );
  XOR U18145 ( .A(n14048), .B(n14049), .Z(n14046) );
  ANDN U18146 ( .B(n14050), .A(n253), .Z(n14048) );
  XNOR U18147 ( .A(b[778]), .B(n14049), .Z(n14050) );
  XOR U18148 ( .A(n14051), .B(n14052), .Z(n14049) );
  ANDN U18149 ( .B(n14053), .A(n254), .Z(n14051) );
  XNOR U18150 ( .A(b[777]), .B(n14052), .Z(n14053) );
  XOR U18151 ( .A(n14054), .B(n14055), .Z(n14052) );
  ANDN U18152 ( .B(n14056), .A(n255), .Z(n14054) );
  XNOR U18153 ( .A(b[776]), .B(n14055), .Z(n14056) );
  XOR U18154 ( .A(n14057), .B(n14058), .Z(n14055) );
  ANDN U18155 ( .B(n14059), .A(n256), .Z(n14057) );
  XNOR U18156 ( .A(b[775]), .B(n14058), .Z(n14059) );
  XOR U18157 ( .A(n14060), .B(n14061), .Z(n14058) );
  ANDN U18158 ( .B(n14062), .A(n257), .Z(n14060) );
  XNOR U18159 ( .A(b[774]), .B(n14061), .Z(n14062) );
  XOR U18160 ( .A(n14063), .B(n14064), .Z(n14061) );
  ANDN U18161 ( .B(n14065), .A(n258), .Z(n14063) );
  XNOR U18162 ( .A(b[773]), .B(n14064), .Z(n14065) );
  XOR U18163 ( .A(n14066), .B(n14067), .Z(n14064) );
  ANDN U18164 ( .B(n14068), .A(n259), .Z(n14066) );
  XNOR U18165 ( .A(b[772]), .B(n14067), .Z(n14068) );
  XOR U18166 ( .A(n14069), .B(n14070), .Z(n14067) );
  ANDN U18167 ( .B(n14071), .A(n260), .Z(n14069) );
  XNOR U18168 ( .A(b[771]), .B(n14070), .Z(n14071) );
  XOR U18169 ( .A(n14072), .B(n14073), .Z(n14070) );
  ANDN U18170 ( .B(n14074), .A(n261), .Z(n14072) );
  XNOR U18171 ( .A(b[770]), .B(n14073), .Z(n14074) );
  XOR U18172 ( .A(n14075), .B(n14076), .Z(n14073) );
  ANDN U18173 ( .B(n14077), .A(n263), .Z(n14075) );
  XNOR U18174 ( .A(b[769]), .B(n14076), .Z(n14077) );
  XOR U18175 ( .A(n14078), .B(n14079), .Z(n14076) );
  ANDN U18176 ( .B(n14080), .A(n264), .Z(n14078) );
  XNOR U18177 ( .A(b[768]), .B(n14079), .Z(n14080) );
  XOR U18178 ( .A(n14081), .B(n14082), .Z(n14079) );
  ANDN U18179 ( .B(n14083), .A(n265), .Z(n14081) );
  XNOR U18180 ( .A(b[767]), .B(n14082), .Z(n14083) );
  XOR U18181 ( .A(n14084), .B(n14085), .Z(n14082) );
  ANDN U18182 ( .B(n14086), .A(n266), .Z(n14084) );
  XNOR U18183 ( .A(b[766]), .B(n14085), .Z(n14086) );
  XOR U18184 ( .A(n14087), .B(n14088), .Z(n14085) );
  ANDN U18185 ( .B(n14089), .A(n267), .Z(n14087) );
  XNOR U18186 ( .A(b[765]), .B(n14088), .Z(n14089) );
  XOR U18187 ( .A(n14090), .B(n14091), .Z(n14088) );
  ANDN U18188 ( .B(n14092), .A(n268), .Z(n14090) );
  XNOR U18189 ( .A(b[764]), .B(n14091), .Z(n14092) );
  XOR U18190 ( .A(n14093), .B(n14094), .Z(n14091) );
  ANDN U18191 ( .B(n14095), .A(n269), .Z(n14093) );
  XNOR U18192 ( .A(b[763]), .B(n14094), .Z(n14095) );
  XOR U18193 ( .A(n14096), .B(n14097), .Z(n14094) );
  ANDN U18194 ( .B(n14098), .A(n270), .Z(n14096) );
  XNOR U18195 ( .A(b[762]), .B(n14097), .Z(n14098) );
  XOR U18196 ( .A(n14099), .B(n14100), .Z(n14097) );
  ANDN U18197 ( .B(n14101), .A(n271), .Z(n14099) );
  XNOR U18198 ( .A(b[761]), .B(n14100), .Z(n14101) );
  XOR U18199 ( .A(n14102), .B(n14103), .Z(n14100) );
  ANDN U18200 ( .B(n14104), .A(n272), .Z(n14102) );
  XNOR U18201 ( .A(b[760]), .B(n14103), .Z(n14104) );
  XOR U18202 ( .A(n14105), .B(n14106), .Z(n14103) );
  ANDN U18203 ( .B(n14107), .A(n274), .Z(n14105) );
  XNOR U18204 ( .A(b[759]), .B(n14106), .Z(n14107) );
  XOR U18205 ( .A(n14108), .B(n14109), .Z(n14106) );
  ANDN U18206 ( .B(n14110), .A(n275), .Z(n14108) );
  XNOR U18207 ( .A(b[758]), .B(n14109), .Z(n14110) );
  XOR U18208 ( .A(n14111), .B(n14112), .Z(n14109) );
  ANDN U18209 ( .B(n14113), .A(n276), .Z(n14111) );
  XNOR U18210 ( .A(b[757]), .B(n14112), .Z(n14113) );
  XOR U18211 ( .A(n14114), .B(n14115), .Z(n14112) );
  ANDN U18212 ( .B(n14116), .A(n277), .Z(n14114) );
  XNOR U18213 ( .A(b[756]), .B(n14115), .Z(n14116) );
  XOR U18214 ( .A(n14117), .B(n14118), .Z(n14115) );
  ANDN U18215 ( .B(n14119), .A(n278), .Z(n14117) );
  XNOR U18216 ( .A(b[755]), .B(n14118), .Z(n14119) );
  XOR U18217 ( .A(n14120), .B(n14121), .Z(n14118) );
  ANDN U18218 ( .B(n14122), .A(n279), .Z(n14120) );
  XNOR U18219 ( .A(b[754]), .B(n14121), .Z(n14122) );
  XOR U18220 ( .A(n14123), .B(n14124), .Z(n14121) );
  ANDN U18221 ( .B(n14125), .A(n280), .Z(n14123) );
  XNOR U18222 ( .A(b[753]), .B(n14124), .Z(n14125) );
  XOR U18223 ( .A(n14126), .B(n14127), .Z(n14124) );
  ANDN U18224 ( .B(n14128), .A(n281), .Z(n14126) );
  XNOR U18225 ( .A(b[752]), .B(n14127), .Z(n14128) );
  XOR U18226 ( .A(n14129), .B(n14130), .Z(n14127) );
  ANDN U18227 ( .B(n14131), .A(n282), .Z(n14129) );
  XNOR U18228 ( .A(b[751]), .B(n14130), .Z(n14131) );
  XOR U18229 ( .A(n14132), .B(n14133), .Z(n14130) );
  ANDN U18230 ( .B(n14134), .A(n283), .Z(n14132) );
  XNOR U18231 ( .A(b[750]), .B(n14133), .Z(n14134) );
  XOR U18232 ( .A(n14135), .B(n14136), .Z(n14133) );
  ANDN U18233 ( .B(n14137), .A(n285), .Z(n14135) );
  XNOR U18234 ( .A(b[749]), .B(n14136), .Z(n14137) );
  XOR U18235 ( .A(n14138), .B(n14139), .Z(n14136) );
  ANDN U18236 ( .B(n14140), .A(n286), .Z(n14138) );
  XNOR U18237 ( .A(b[748]), .B(n14139), .Z(n14140) );
  XOR U18238 ( .A(n14141), .B(n14142), .Z(n14139) );
  ANDN U18239 ( .B(n14143), .A(n287), .Z(n14141) );
  XNOR U18240 ( .A(b[747]), .B(n14142), .Z(n14143) );
  XOR U18241 ( .A(n14144), .B(n14145), .Z(n14142) );
  ANDN U18242 ( .B(n14146), .A(n288), .Z(n14144) );
  XNOR U18243 ( .A(b[746]), .B(n14145), .Z(n14146) );
  XOR U18244 ( .A(n14147), .B(n14148), .Z(n14145) );
  ANDN U18245 ( .B(n14149), .A(n289), .Z(n14147) );
  XNOR U18246 ( .A(b[745]), .B(n14148), .Z(n14149) );
  XOR U18247 ( .A(n14150), .B(n14151), .Z(n14148) );
  ANDN U18248 ( .B(n14152), .A(n290), .Z(n14150) );
  XNOR U18249 ( .A(b[744]), .B(n14151), .Z(n14152) );
  XOR U18250 ( .A(n14153), .B(n14154), .Z(n14151) );
  ANDN U18251 ( .B(n14155), .A(n291), .Z(n14153) );
  XNOR U18252 ( .A(b[743]), .B(n14154), .Z(n14155) );
  XOR U18253 ( .A(n14156), .B(n14157), .Z(n14154) );
  ANDN U18254 ( .B(n14158), .A(n292), .Z(n14156) );
  XNOR U18255 ( .A(b[742]), .B(n14157), .Z(n14158) );
  XOR U18256 ( .A(n14159), .B(n14160), .Z(n14157) );
  ANDN U18257 ( .B(n14161), .A(n293), .Z(n14159) );
  XNOR U18258 ( .A(b[741]), .B(n14160), .Z(n14161) );
  XOR U18259 ( .A(n14162), .B(n14163), .Z(n14160) );
  ANDN U18260 ( .B(n14164), .A(n294), .Z(n14162) );
  XNOR U18261 ( .A(b[740]), .B(n14163), .Z(n14164) );
  XOR U18262 ( .A(n14165), .B(n14166), .Z(n14163) );
  ANDN U18263 ( .B(n14167), .A(n296), .Z(n14165) );
  XNOR U18264 ( .A(b[739]), .B(n14166), .Z(n14167) );
  XOR U18265 ( .A(n14168), .B(n14169), .Z(n14166) );
  ANDN U18266 ( .B(n14170), .A(n297), .Z(n14168) );
  XNOR U18267 ( .A(b[738]), .B(n14169), .Z(n14170) );
  XOR U18268 ( .A(n14171), .B(n14172), .Z(n14169) );
  ANDN U18269 ( .B(n14173), .A(n298), .Z(n14171) );
  XNOR U18270 ( .A(b[737]), .B(n14172), .Z(n14173) );
  XOR U18271 ( .A(n14174), .B(n14175), .Z(n14172) );
  ANDN U18272 ( .B(n14176), .A(n299), .Z(n14174) );
  XNOR U18273 ( .A(b[736]), .B(n14175), .Z(n14176) );
  XOR U18274 ( .A(n14177), .B(n14178), .Z(n14175) );
  ANDN U18275 ( .B(n14179), .A(n300), .Z(n14177) );
  XNOR U18276 ( .A(b[735]), .B(n14178), .Z(n14179) );
  XOR U18277 ( .A(n14180), .B(n14181), .Z(n14178) );
  ANDN U18278 ( .B(n14182), .A(n301), .Z(n14180) );
  XNOR U18279 ( .A(b[734]), .B(n14181), .Z(n14182) );
  XOR U18280 ( .A(n14183), .B(n14184), .Z(n14181) );
  ANDN U18281 ( .B(n14185), .A(n302), .Z(n14183) );
  XNOR U18282 ( .A(b[733]), .B(n14184), .Z(n14185) );
  XOR U18283 ( .A(n14186), .B(n14187), .Z(n14184) );
  ANDN U18284 ( .B(n14188), .A(n303), .Z(n14186) );
  XNOR U18285 ( .A(b[732]), .B(n14187), .Z(n14188) );
  XOR U18286 ( .A(n14189), .B(n14190), .Z(n14187) );
  ANDN U18287 ( .B(n14191), .A(n304), .Z(n14189) );
  XNOR U18288 ( .A(b[731]), .B(n14190), .Z(n14191) );
  XOR U18289 ( .A(n14192), .B(n14193), .Z(n14190) );
  ANDN U18290 ( .B(n14194), .A(n305), .Z(n14192) );
  XNOR U18291 ( .A(b[730]), .B(n14193), .Z(n14194) );
  XOR U18292 ( .A(n14195), .B(n14196), .Z(n14193) );
  ANDN U18293 ( .B(n14197), .A(n307), .Z(n14195) );
  XNOR U18294 ( .A(b[729]), .B(n14196), .Z(n14197) );
  XOR U18295 ( .A(n14198), .B(n14199), .Z(n14196) );
  ANDN U18296 ( .B(n14200), .A(n308), .Z(n14198) );
  XNOR U18297 ( .A(b[728]), .B(n14199), .Z(n14200) );
  XOR U18298 ( .A(n14201), .B(n14202), .Z(n14199) );
  ANDN U18299 ( .B(n14203), .A(n309), .Z(n14201) );
  XNOR U18300 ( .A(b[727]), .B(n14202), .Z(n14203) );
  XOR U18301 ( .A(n14204), .B(n14205), .Z(n14202) );
  ANDN U18302 ( .B(n14206), .A(n310), .Z(n14204) );
  XNOR U18303 ( .A(b[726]), .B(n14205), .Z(n14206) );
  XOR U18304 ( .A(n14207), .B(n14208), .Z(n14205) );
  ANDN U18305 ( .B(n14209), .A(n311), .Z(n14207) );
  XNOR U18306 ( .A(b[725]), .B(n14208), .Z(n14209) );
  XOR U18307 ( .A(n14210), .B(n14211), .Z(n14208) );
  ANDN U18308 ( .B(n14212), .A(n312), .Z(n14210) );
  XNOR U18309 ( .A(b[724]), .B(n14211), .Z(n14212) );
  XOR U18310 ( .A(n14213), .B(n14214), .Z(n14211) );
  ANDN U18311 ( .B(n14215), .A(n313), .Z(n14213) );
  XNOR U18312 ( .A(b[723]), .B(n14214), .Z(n14215) );
  XOR U18313 ( .A(n14216), .B(n14217), .Z(n14214) );
  ANDN U18314 ( .B(n14218), .A(n314), .Z(n14216) );
  XNOR U18315 ( .A(b[722]), .B(n14217), .Z(n14218) );
  XOR U18316 ( .A(n14219), .B(n14220), .Z(n14217) );
  ANDN U18317 ( .B(n14221), .A(n315), .Z(n14219) );
  XNOR U18318 ( .A(b[721]), .B(n14220), .Z(n14221) );
  XOR U18319 ( .A(n14222), .B(n14223), .Z(n14220) );
  ANDN U18320 ( .B(n14224), .A(n316), .Z(n14222) );
  XNOR U18321 ( .A(b[720]), .B(n14223), .Z(n14224) );
  XOR U18322 ( .A(n14225), .B(n14226), .Z(n14223) );
  ANDN U18323 ( .B(n14227), .A(n318), .Z(n14225) );
  XNOR U18324 ( .A(b[719]), .B(n14226), .Z(n14227) );
  XOR U18325 ( .A(n14228), .B(n14229), .Z(n14226) );
  ANDN U18326 ( .B(n14230), .A(n319), .Z(n14228) );
  XNOR U18327 ( .A(b[718]), .B(n14229), .Z(n14230) );
  XOR U18328 ( .A(n14231), .B(n14232), .Z(n14229) );
  ANDN U18329 ( .B(n14233), .A(n320), .Z(n14231) );
  XNOR U18330 ( .A(b[717]), .B(n14232), .Z(n14233) );
  XOR U18331 ( .A(n14234), .B(n14235), .Z(n14232) );
  ANDN U18332 ( .B(n14236), .A(n321), .Z(n14234) );
  XNOR U18333 ( .A(b[716]), .B(n14235), .Z(n14236) );
  XOR U18334 ( .A(n14237), .B(n14238), .Z(n14235) );
  ANDN U18335 ( .B(n14239), .A(n322), .Z(n14237) );
  XNOR U18336 ( .A(b[715]), .B(n14238), .Z(n14239) );
  XOR U18337 ( .A(n14240), .B(n14241), .Z(n14238) );
  ANDN U18338 ( .B(n14242), .A(n323), .Z(n14240) );
  XNOR U18339 ( .A(b[714]), .B(n14241), .Z(n14242) );
  XOR U18340 ( .A(n14243), .B(n14244), .Z(n14241) );
  ANDN U18341 ( .B(n14245), .A(n324), .Z(n14243) );
  XNOR U18342 ( .A(b[713]), .B(n14244), .Z(n14245) );
  XOR U18343 ( .A(n14246), .B(n14247), .Z(n14244) );
  ANDN U18344 ( .B(n14248), .A(n325), .Z(n14246) );
  XNOR U18345 ( .A(b[712]), .B(n14247), .Z(n14248) );
  XOR U18346 ( .A(n14249), .B(n14250), .Z(n14247) );
  ANDN U18347 ( .B(n14251), .A(n326), .Z(n14249) );
  XNOR U18348 ( .A(b[711]), .B(n14250), .Z(n14251) );
  XOR U18349 ( .A(n14252), .B(n14253), .Z(n14250) );
  ANDN U18350 ( .B(n14254), .A(n327), .Z(n14252) );
  XNOR U18351 ( .A(b[710]), .B(n14253), .Z(n14254) );
  XOR U18352 ( .A(n14255), .B(n14256), .Z(n14253) );
  ANDN U18353 ( .B(n14257), .A(n329), .Z(n14255) );
  XNOR U18354 ( .A(b[709]), .B(n14256), .Z(n14257) );
  XOR U18355 ( .A(n14258), .B(n14259), .Z(n14256) );
  ANDN U18356 ( .B(n14260), .A(n330), .Z(n14258) );
  XNOR U18357 ( .A(b[708]), .B(n14259), .Z(n14260) );
  XOR U18358 ( .A(n14261), .B(n14262), .Z(n14259) );
  ANDN U18359 ( .B(n14263), .A(n331), .Z(n14261) );
  XNOR U18360 ( .A(b[707]), .B(n14262), .Z(n14263) );
  XOR U18361 ( .A(n14264), .B(n14265), .Z(n14262) );
  ANDN U18362 ( .B(n14266), .A(n332), .Z(n14264) );
  XNOR U18363 ( .A(b[706]), .B(n14265), .Z(n14266) );
  XOR U18364 ( .A(n14267), .B(n14268), .Z(n14265) );
  ANDN U18365 ( .B(n14269), .A(n333), .Z(n14267) );
  XNOR U18366 ( .A(b[705]), .B(n14268), .Z(n14269) );
  XOR U18367 ( .A(n14270), .B(n14271), .Z(n14268) );
  ANDN U18368 ( .B(n14272), .A(n334), .Z(n14270) );
  XNOR U18369 ( .A(b[704]), .B(n14271), .Z(n14272) );
  XOR U18370 ( .A(n14273), .B(n14274), .Z(n14271) );
  ANDN U18371 ( .B(n14275), .A(n335), .Z(n14273) );
  XNOR U18372 ( .A(b[703]), .B(n14274), .Z(n14275) );
  XOR U18373 ( .A(n14276), .B(n14277), .Z(n14274) );
  ANDN U18374 ( .B(n14278), .A(n336), .Z(n14276) );
  XNOR U18375 ( .A(b[702]), .B(n14277), .Z(n14278) );
  XOR U18376 ( .A(n14279), .B(n14280), .Z(n14277) );
  ANDN U18377 ( .B(n14281), .A(n337), .Z(n14279) );
  XNOR U18378 ( .A(b[701]), .B(n14280), .Z(n14281) );
  XOR U18379 ( .A(n14282), .B(n14283), .Z(n14280) );
  ANDN U18380 ( .B(n14284), .A(n338), .Z(n14282) );
  XNOR U18381 ( .A(b[700]), .B(n14283), .Z(n14284) );
  XOR U18382 ( .A(n14285), .B(n14286), .Z(n14283) );
  ANDN U18383 ( .B(n14287), .A(n341), .Z(n14285) );
  XNOR U18384 ( .A(b[699]), .B(n14286), .Z(n14287) );
  XOR U18385 ( .A(n14288), .B(n14289), .Z(n14286) );
  ANDN U18386 ( .B(n14290), .A(n342), .Z(n14288) );
  XNOR U18387 ( .A(b[698]), .B(n14289), .Z(n14290) );
  XOR U18388 ( .A(n14291), .B(n14292), .Z(n14289) );
  ANDN U18389 ( .B(n14293), .A(n343), .Z(n14291) );
  XNOR U18390 ( .A(b[697]), .B(n14292), .Z(n14293) );
  XOR U18391 ( .A(n14294), .B(n14295), .Z(n14292) );
  ANDN U18392 ( .B(n14296), .A(n344), .Z(n14294) );
  XNOR U18393 ( .A(b[696]), .B(n14295), .Z(n14296) );
  XOR U18394 ( .A(n14297), .B(n14298), .Z(n14295) );
  ANDN U18395 ( .B(n14299), .A(n345), .Z(n14297) );
  XNOR U18396 ( .A(b[695]), .B(n14298), .Z(n14299) );
  XOR U18397 ( .A(n14300), .B(n14301), .Z(n14298) );
  ANDN U18398 ( .B(n14302), .A(n346), .Z(n14300) );
  XNOR U18399 ( .A(b[694]), .B(n14301), .Z(n14302) );
  XOR U18400 ( .A(n14303), .B(n14304), .Z(n14301) );
  ANDN U18401 ( .B(n14305), .A(n347), .Z(n14303) );
  XNOR U18402 ( .A(b[693]), .B(n14304), .Z(n14305) );
  XOR U18403 ( .A(n14306), .B(n14307), .Z(n14304) );
  ANDN U18404 ( .B(n14308), .A(n348), .Z(n14306) );
  XNOR U18405 ( .A(b[692]), .B(n14307), .Z(n14308) );
  XOR U18406 ( .A(n14309), .B(n14310), .Z(n14307) );
  ANDN U18407 ( .B(n14311), .A(n349), .Z(n14309) );
  XNOR U18408 ( .A(b[691]), .B(n14310), .Z(n14311) );
  XOR U18409 ( .A(n14312), .B(n14313), .Z(n14310) );
  ANDN U18410 ( .B(n14314), .A(n350), .Z(n14312) );
  XNOR U18411 ( .A(b[690]), .B(n14313), .Z(n14314) );
  XOR U18412 ( .A(n14315), .B(n14316), .Z(n14313) );
  ANDN U18413 ( .B(n14317), .A(n352), .Z(n14315) );
  XNOR U18414 ( .A(b[689]), .B(n14316), .Z(n14317) );
  XOR U18415 ( .A(n14318), .B(n14319), .Z(n14316) );
  ANDN U18416 ( .B(n14320), .A(n353), .Z(n14318) );
  XNOR U18417 ( .A(b[688]), .B(n14319), .Z(n14320) );
  XOR U18418 ( .A(n14321), .B(n14322), .Z(n14319) );
  ANDN U18419 ( .B(n14323), .A(n354), .Z(n14321) );
  XNOR U18420 ( .A(b[687]), .B(n14322), .Z(n14323) );
  XOR U18421 ( .A(n14324), .B(n14325), .Z(n14322) );
  ANDN U18422 ( .B(n14326), .A(n355), .Z(n14324) );
  XNOR U18423 ( .A(b[686]), .B(n14325), .Z(n14326) );
  XOR U18424 ( .A(n14327), .B(n14328), .Z(n14325) );
  ANDN U18425 ( .B(n14329), .A(n356), .Z(n14327) );
  XNOR U18426 ( .A(b[685]), .B(n14328), .Z(n14329) );
  XOR U18427 ( .A(n14330), .B(n14331), .Z(n14328) );
  ANDN U18428 ( .B(n14332), .A(n357), .Z(n14330) );
  XNOR U18429 ( .A(b[684]), .B(n14331), .Z(n14332) );
  XOR U18430 ( .A(n14333), .B(n14334), .Z(n14331) );
  ANDN U18431 ( .B(n14335), .A(n358), .Z(n14333) );
  XNOR U18432 ( .A(b[683]), .B(n14334), .Z(n14335) );
  XOR U18433 ( .A(n14336), .B(n14337), .Z(n14334) );
  ANDN U18434 ( .B(n14338), .A(n359), .Z(n14336) );
  XNOR U18435 ( .A(b[682]), .B(n14337), .Z(n14338) );
  XOR U18436 ( .A(n14339), .B(n14340), .Z(n14337) );
  ANDN U18437 ( .B(n14341), .A(n360), .Z(n14339) );
  XNOR U18438 ( .A(b[681]), .B(n14340), .Z(n14341) );
  XOR U18439 ( .A(n14342), .B(n14343), .Z(n14340) );
  ANDN U18440 ( .B(n14344), .A(n361), .Z(n14342) );
  XNOR U18441 ( .A(b[680]), .B(n14343), .Z(n14344) );
  XOR U18442 ( .A(n14345), .B(n14346), .Z(n14343) );
  ANDN U18443 ( .B(n14347), .A(n363), .Z(n14345) );
  XNOR U18444 ( .A(b[679]), .B(n14346), .Z(n14347) );
  XOR U18445 ( .A(n14348), .B(n14349), .Z(n14346) );
  ANDN U18446 ( .B(n14350), .A(n364), .Z(n14348) );
  XNOR U18447 ( .A(b[678]), .B(n14349), .Z(n14350) );
  XOR U18448 ( .A(n14351), .B(n14352), .Z(n14349) );
  ANDN U18449 ( .B(n14353), .A(n365), .Z(n14351) );
  XNOR U18450 ( .A(b[677]), .B(n14352), .Z(n14353) );
  XOR U18451 ( .A(n14354), .B(n14355), .Z(n14352) );
  ANDN U18452 ( .B(n14356), .A(n366), .Z(n14354) );
  XNOR U18453 ( .A(b[676]), .B(n14355), .Z(n14356) );
  XOR U18454 ( .A(n14357), .B(n14358), .Z(n14355) );
  ANDN U18455 ( .B(n14359), .A(n367), .Z(n14357) );
  XNOR U18456 ( .A(b[675]), .B(n14358), .Z(n14359) );
  XOR U18457 ( .A(n14360), .B(n14361), .Z(n14358) );
  ANDN U18458 ( .B(n14362), .A(n368), .Z(n14360) );
  XNOR U18459 ( .A(b[674]), .B(n14361), .Z(n14362) );
  XOR U18460 ( .A(n14363), .B(n14364), .Z(n14361) );
  ANDN U18461 ( .B(n14365), .A(n369), .Z(n14363) );
  XNOR U18462 ( .A(b[673]), .B(n14364), .Z(n14365) );
  XOR U18463 ( .A(n14366), .B(n14367), .Z(n14364) );
  ANDN U18464 ( .B(n14368), .A(n370), .Z(n14366) );
  XNOR U18465 ( .A(b[672]), .B(n14367), .Z(n14368) );
  XOR U18466 ( .A(n14369), .B(n14370), .Z(n14367) );
  ANDN U18467 ( .B(n14371), .A(n371), .Z(n14369) );
  XNOR U18468 ( .A(b[671]), .B(n14370), .Z(n14371) );
  XOR U18469 ( .A(n14372), .B(n14373), .Z(n14370) );
  ANDN U18470 ( .B(n14374), .A(n372), .Z(n14372) );
  XNOR U18471 ( .A(b[670]), .B(n14373), .Z(n14374) );
  XOR U18472 ( .A(n14375), .B(n14376), .Z(n14373) );
  ANDN U18473 ( .B(n14377), .A(n374), .Z(n14375) );
  XNOR U18474 ( .A(b[669]), .B(n14376), .Z(n14377) );
  XOR U18475 ( .A(n14378), .B(n14379), .Z(n14376) );
  ANDN U18476 ( .B(n14380), .A(n375), .Z(n14378) );
  XNOR U18477 ( .A(b[668]), .B(n14379), .Z(n14380) );
  XOR U18478 ( .A(n14381), .B(n14382), .Z(n14379) );
  ANDN U18479 ( .B(n14383), .A(n376), .Z(n14381) );
  XNOR U18480 ( .A(b[667]), .B(n14382), .Z(n14383) );
  XOR U18481 ( .A(n14384), .B(n14385), .Z(n14382) );
  ANDN U18482 ( .B(n14386), .A(n377), .Z(n14384) );
  XNOR U18483 ( .A(b[666]), .B(n14385), .Z(n14386) );
  XOR U18484 ( .A(n14387), .B(n14388), .Z(n14385) );
  ANDN U18485 ( .B(n14389), .A(n378), .Z(n14387) );
  XNOR U18486 ( .A(b[665]), .B(n14388), .Z(n14389) );
  XOR U18487 ( .A(n14390), .B(n14391), .Z(n14388) );
  ANDN U18488 ( .B(n14392), .A(n379), .Z(n14390) );
  XNOR U18489 ( .A(b[664]), .B(n14391), .Z(n14392) );
  XOR U18490 ( .A(n14393), .B(n14394), .Z(n14391) );
  ANDN U18491 ( .B(n14395), .A(n380), .Z(n14393) );
  XNOR U18492 ( .A(b[663]), .B(n14394), .Z(n14395) );
  XOR U18493 ( .A(n14396), .B(n14397), .Z(n14394) );
  ANDN U18494 ( .B(n14398), .A(n381), .Z(n14396) );
  XNOR U18495 ( .A(b[662]), .B(n14397), .Z(n14398) );
  XOR U18496 ( .A(n14399), .B(n14400), .Z(n14397) );
  ANDN U18497 ( .B(n14401), .A(n382), .Z(n14399) );
  XNOR U18498 ( .A(b[661]), .B(n14400), .Z(n14401) );
  XOR U18499 ( .A(n14402), .B(n14403), .Z(n14400) );
  ANDN U18500 ( .B(n14404), .A(n383), .Z(n14402) );
  XNOR U18501 ( .A(b[660]), .B(n14403), .Z(n14404) );
  XOR U18502 ( .A(n14405), .B(n14406), .Z(n14403) );
  ANDN U18503 ( .B(n14407), .A(n385), .Z(n14405) );
  XNOR U18504 ( .A(b[659]), .B(n14406), .Z(n14407) );
  XOR U18505 ( .A(n14408), .B(n14409), .Z(n14406) );
  ANDN U18506 ( .B(n14410), .A(n386), .Z(n14408) );
  XNOR U18507 ( .A(b[658]), .B(n14409), .Z(n14410) );
  XOR U18508 ( .A(n14411), .B(n14412), .Z(n14409) );
  ANDN U18509 ( .B(n14413), .A(n387), .Z(n14411) );
  XNOR U18510 ( .A(b[657]), .B(n14412), .Z(n14413) );
  XOR U18511 ( .A(n14414), .B(n14415), .Z(n14412) );
  ANDN U18512 ( .B(n14416), .A(n388), .Z(n14414) );
  XNOR U18513 ( .A(b[656]), .B(n14415), .Z(n14416) );
  XOR U18514 ( .A(n14417), .B(n14418), .Z(n14415) );
  ANDN U18515 ( .B(n14419), .A(n389), .Z(n14417) );
  XNOR U18516 ( .A(b[655]), .B(n14418), .Z(n14419) );
  XOR U18517 ( .A(n14420), .B(n14421), .Z(n14418) );
  ANDN U18518 ( .B(n14422), .A(n390), .Z(n14420) );
  XNOR U18519 ( .A(b[654]), .B(n14421), .Z(n14422) );
  XOR U18520 ( .A(n14423), .B(n14424), .Z(n14421) );
  ANDN U18521 ( .B(n14425), .A(n391), .Z(n14423) );
  XNOR U18522 ( .A(b[653]), .B(n14424), .Z(n14425) );
  XOR U18523 ( .A(n14426), .B(n14427), .Z(n14424) );
  ANDN U18524 ( .B(n14428), .A(n392), .Z(n14426) );
  XNOR U18525 ( .A(b[652]), .B(n14427), .Z(n14428) );
  XOR U18526 ( .A(n14429), .B(n14430), .Z(n14427) );
  ANDN U18527 ( .B(n14431), .A(n393), .Z(n14429) );
  XNOR U18528 ( .A(b[651]), .B(n14430), .Z(n14431) );
  XOR U18529 ( .A(n14432), .B(n14433), .Z(n14430) );
  ANDN U18530 ( .B(n14434), .A(n394), .Z(n14432) );
  XNOR U18531 ( .A(b[650]), .B(n14433), .Z(n14434) );
  XOR U18532 ( .A(n14435), .B(n14436), .Z(n14433) );
  ANDN U18533 ( .B(n14437), .A(n396), .Z(n14435) );
  XNOR U18534 ( .A(b[649]), .B(n14436), .Z(n14437) );
  XOR U18535 ( .A(n14438), .B(n14439), .Z(n14436) );
  ANDN U18536 ( .B(n14440), .A(n397), .Z(n14438) );
  XNOR U18537 ( .A(b[648]), .B(n14439), .Z(n14440) );
  XOR U18538 ( .A(n14441), .B(n14442), .Z(n14439) );
  ANDN U18539 ( .B(n14443), .A(n398), .Z(n14441) );
  XNOR U18540 ( .A(b[647]), .B(n14442), .Z(n14443) );
  XOR U18541 ( .A(n14444), .B(n14445), .Z(n14442) );
  ANDN U18542 ( .B(n14446), .A(n399), .Z(n14444) );
  XNOR U18543 ( .A(b[646]), .B(n14445), .Z(n14446) );
  XOR U18544 ( .A(n14447), .B(n14448), .Z(n14445) );
  ANDN U18545 ( .B(n14449), .A(n400), .Z(n14447) );
  XNOR U18546 ( .A(b[645]), .B(n14448), .Z(n14449) );
  XOR U18547 ( .A(n14450), .B(n14451), .Z(n14448) );
  ANDN U18548 ( .B(n14452), .A(n401), .Z(n14450) );
  XNOR U18549 ( .A(b[644]), .B(n14451), .Z(n14452) );
  XOR U18550 ( .A(n14453), .B(n14454), .Z(n14451) );
  ANDN U18551 ( .B(n14455), .A(n402), .Z(n14453) );
  XNOR U18552 ( .A(b[643]), .B(n14454), .Z(n14455) );
  XOR U18553 ( .A(n14456), .B(n14457), .Z(n14454) );
  ANDN U18554 ( .B(n14458), .A(n403), .Z(n14456) );
  XNOR U18555 ( .A(b[642]), .B(n14457), .Z(n14458) );
  XOR U18556 ( .A(n14459), .B(n14460), .Z(n14457) );
  ANDN U18557 ( .B(n14461), .A(n404), .Z(n14459) );
  XNOR U18558 ( .A(b[641]), .B(n14460), .Z(n14461) );
  XOR U18559 ( .A(n14462), .B(n14463), .Z(n14460) );
  ANDN U18560 ( .B(n14464), .A(n405), .Z(n14462) );
  XNOR U18561 ( .A(b[640]), .B(n14463), .Z(n14464) );
  XOR U18562 ( .A(n14465), .B(n14466), .Z(n14463) );
  ANDN U18563 ( .B(n14467), .A(n407), .Z(n14465) );
  XNOR U18564 ( .A(b[639]), .B(n14466), .Z(n14467) );
  XOR U18565 ( .A(n14468), .B(n14469), .Z(n14466) );
  ANDN U18566 ( .B(n14470), .A(n408), .Z(n14468) );
  XNOR U18567 ( .A(b[638]), .B(n14469), .Z(n14470) );
  XOR U18568 ( .A(n14471), .B(n14472), .Z(n14469) );
  ANDN U18569 ( .B(n14473), .A(n409), .Z(n14471) );
  XNOR U18570 ( .A(b[637]), .B(n14472), .Z(n14473) );
  XOR U18571 ( .A(n14474), .B(n14475), .Z(n14472) );
  ANDN U18572 ( .B(n14476), .A(n410), .Z(n14474) );
  XNOR U18573 ( .A(b[636]), .B(n14475), .Z(n14476) );
  XOR U18574 ( .A(n14477), .B(n14478), .Z(n14475) );
  ANDN U18575 ( .B(n14479), .A(n411), .Z(n14477) );
  XNOR U18576 ( .A(b[635]), .B(n14478), .Z(n14479) );
  XOR U18577 ( .A(n14480), .B(n14481), .Z(n14478) );
  ANDN U18578 ( .B(n14482), .A(n412), .Z(n14480) );
  XNOR U18579 ( .A(b[634]), .B(n14481), .Z(n14482) );
  XOR U18580 ( .A(n14483), .B(n14484), .Z(n14481) );
  ANDN U18581 ( .B(n14485), .A(n413), .Z(n14483) );
  XNOR U18582 ( .A(b[633]), .B(n14484), .Z(n14485) );
  XOR U18583 ( .A(n14486), .B(n14487), .Z(n14484) );
  ANDN U18584 ( .B(n14488), .A(n414), .Z(n14486) );
  XNOR U18585 ( .A(b[632]), .B(n14487), .Z(n14488) );
  XOR U18586 ( .A(n14489), .B(n14490), .Z(n14487) );
  ANDN U18587 ( .B(n14491), .A(n415), .Z(n14489) );
  XNOR U18588 ( .A(b[631]), .B(n14490), .Z(n14491) );
  XOR U18589 ( .A(n14492), .B(n14493), .Z(n14490) );
  ANDN U18590 ( .B(n14494), .A(n416), .Z(n14492) );
  XNOR U18591 ( .A(b[630]), .B(n14493), .Z(n14494) );
  XOR U18592 ( .A(n14495), .B(n14496), .Z(n14493) );
  ANDN U18593 ( .B(n14497), .A(n418), .Z(n14495) );
  XNOR U18594 ( .A(b[629]), .B(n14496), .Z(n14497) );
  XOR U18595 ( .A(n14498), .B(n14499), .Z(n14496) );
  ANDN U18596 ( .B(n14500), .A(n419), .Z(n14498) );
  XNOR U18597 ( .A(b[628]), .B(n14499), .Z(n14500) );
  XOR U18598 ( .A(n14501), .B(n14502), .Z(n14499) );
  ANDN U18599 ( .B(n14503), .A(n420), .Z(n14501) );
  XNOR U18600 ( .A(b[627]), .B(n14502), .Z(n14503) );
  XOR U18601 ( .A(n14504), .B(n14505), .Z(n14502) );
  ANDN U18602 ( .B(n14506), .A(n421), .Z(n14504) );
  XNOR U18603 ( .A(b[626]), .B(n14505), .Z(n14506) );
  XOR U18604 ( .A(n14507), .B(n14508), .Z(n14505) );
  ANDN U18605 ( .B(n14509), .A(n422), .Z(n14507) );
  XNOR U18606 ( .A(b[625]), .B(n14508), .Z(n14509) );
  XOR U18607 ( .A(n14510), .B(n14511), .Z(n14508) );
  ANDN U18608 ( .B(n14512), .A(n423), .Z(n14510) );
  XNOR U18609 ( .A(b[624]), .B(n14511), .Z(n14512) );
  XOR U18610 ( .A(n14513), .B(n14514), .Z(n14511) );
  ANDN U18611 ( .B(n14515), .A(n424), .Z(n14513) );
  XNOR U18612 ( .A(b[623]), .B(n14514), .Z(n14515) );
  XOR U18613 ( .A(n14516), .B(n14517), .Z(n14514) );
  ANDN U18614 ( .B(n14518), .A(n425), .Z(n14516) );
  XNOR U18615 ( .A(b[622]), .B(n14517), .Z(n14518) );
  XOR U18616 ( .A(n14519), .B(n14520), .Z(n14517) );
  ANDN U18617 ( .B(n14521), .A(n426), .Z(n14519) );
  XNOR U18618 ( .A(b[621]), .B(n14520), .Z(n14521) );
  XOR U18619 ( .A(n14522), .B(n14523), .Z(n14520) );
  ANDN U18620 ( .B(n14524), .A(n427), .Z(n14522) );
  XNOR U18621 ( .A(b[620]), .B(n14523), .Z(n14524) );
  XOR U18622 ( .A(n14525), .B(n14526), .Z(n14523) );
  ANDN U18623 ( .B(n14527), .A(n429), .Z(n14525) );
  XNOR U18624 ( .A(b[619]), .B(n14526), .Z(n14527) );
  XOR U18625 ( .A(n14528), .B(n14529), .Z(n14526) );
  ANDN U18626 ( .B(n14530), .A(n430), .Z(n14528) );
  XNOR U18627 ( .A(b[618]), .B(n14529), .Z(n14530) );
  XOR U18628 ( .A(n14531), .B(n14532), .Z(n14529) );
  ANDN U18629 ( .B(n14533), .A(n431), .Z(n14531) );
  XNOR U18630 ( .A(b[617]), .B(n14532), .Z(n14533) );
  XOR U18631 ( .A(n14534), .B(n14535), .Z(n14532) );
  ANDN U18632 ( .B(n14536), .A(n432), .Z(n14534) );
  XNOR U18633 ( .A(b[616]), .B(n14535), .Z(n14536) );
  XOR U18634 ( .A(n14537), .B(n14538), .Z(n14535) );
  ANDN U18635 ( .B(n14539), .A(n433), .Z(n14537) );
  XNOR U18636 ( .A(b[615]), .B(n14538), .Z(n14539) );
  XOR U18637 ( .A(n14540), .B(n14541), .Z(n14538) );
  ANDN U18638 ( .B(n14542), .A(n434), .Z(n14540) );
  XNOR U18639 ( .A(b[614]), .B(n14541), .Z(n14542) );
  XOR U18640 ( .A(n14543), .B(n14544), .Z(n14541) );
  ANDN U18641 ( .B(n14545), .A(n435), .Z(n14543) );
  XNOR U18642 ( .A(b[613]), .B(n14544), .Z(n14545) );
  XOR U18643 ( .A(n14546), .B(n14547), .Z(n14544) );
  ANDN U18644 ( .B(n14548), .A(n436), .Z(n14546) );
  XNOR U18645 ( .A(b[612]), .B(n14547), .Z(n14548) );
  XOR U18646 ( .A(n14549), .B(n14550), .Z(n14547) );
  ANDN U18647 ( .B(n14551), .A(n437), .Z(n14549) );
  XNOR U18648 ( .A(b[611]), .B(n14550), .Z(n14551) );
  XOR U18649 ( .A(n14552), .B(n14553), .Z(n14550) );
  ANDN U18650 ( .B(n14554), .A(n438), .Z(n14552) );
  XNOR U18651 ( .A(b[610]), .B(n14553), .Z(n14554) );
  XOR U18652 ( .A(n14555), .B(n14556), .Z(n14553) );
  ANDN U18653 ( .B(n14557), .A(n440), .Z(n14555) );
  XNOR U18654 ( .A(b[609]), .B(n14556), .Z(n14557) );
  XOR U18655 ( .A(n14558), .B(n14559), .Z(n14556) );
  ANDN U18656 ( .B(n14560), .A(n441), .Z(n14558) );
  XNOR U18657 ( .A(b[608]), .B(n14559), .Z(n14560) );
  XOR U18658 ( .A(n14561), .B(n14562), .Z(n14559) );
  ANDN U18659 ( .B(n14563), .A(n442), .Z(n14561) );
  XNOR U18660 ( .A(b[607]), .B(n14562), .Z(n14563) );
  XOR U18661 ( .A(n14564), .B(n14565), .Z(n14562) );
  ANDN U18662 ( .B(n14566), .A(n443), .Z(n14564) );
  XNOR U18663 ( .A(b[606]), .B(n14565), .Z(n14566) );
  XOR U18664 ( .A(n14567), .B(n14568), .Z(n14565) );
  ANDN U18665 ( .B(n14569), .A(n444), .Z(n14567) );
  XNOR U18666 ( .A(b[605]), .B(n14568), .Z(n14569) );
  XOR U18667 ( .A(n14570), .B(n14571), .Z(n14568) );
  ANDN U18668 ( .B(n14572), .A(n445), .Z(n14570) );
  XNOR U18669 ( .A(b[604]), .B(n14571), .Z(n14572) );
  XOR U18670 ( .A(n14573), .B(n14574), .Z(n14571) );
  ANDN U18671 ( .B(n14575), .A(n446), .Z(n14573) );
  XNOR U18672 ( .A(b[603]), .B(n14574), .Z(n14575) );
  XOR U18673 ( .A(n14576), .B(n14577), .Z(n14574) );
  ANDN U18674 ( .B(n14578), .A(n447), .Z(n14576) );
  XNOR U18675 ( .A(b[602]), .B(n14577), .Z(n14578) );
  XOR U18676 ( .A(n14579), .B(n14580), .Z(n14577) );
  ANDN U18677 ( .B(n14581), .A(n448), .Z(n14579) );
  XNOR U18678 ( .A(b[601]), .B(n14580), .Z(n14581) );
  XOR U18679 ( .A(n14582), .B(n14583), .Z(n14580) );
  ANDN U18680 ( .B(n14584), .A(n449), .Z(n14582) );
  XNOR U18681 ( .A(b[600]), .B(n14583), .Z(n14584) );
  XOR U18682 ( .A(n14585), .B(n14586), .Z(n14583) );
  ANDN U18683 ( .B(n14587), .A(n452), .Z(n14585) );
  XNOR U18684 ( .A(b[599]), .B(n14586), .Z(n14587) );
  XOR U18685 ( .A(n14588), .B(n14589), .Z(n14586) );
  ANDN U18686 ( .B(n14590), .A(n453), .Z(n14588) );
  XNOR U18687 ( .A(b[598]), .B(n14589), .Z(n14590) );
  XOR U18688 ( .A(n14591), .B(n14592), .Z(n14589) );
  ANDN U18689 ( .B(n14593), .A(n454), .Z(n14591) );
  XNOR U18690 ( .A(b[597]), .B(n14592), .Z(n14593) );
  XOR U18691 ( .A(n14594), .B(n14595), .Z(n14592) );
  ANDN U18692 ( .B(n14596), .A(n455), .Z(n14594) );
  XNOR U18693 ( .A(b[596]), .B(n14595), .Z(n14596) );
  XOR U18694 ( .A(n14597), .B(n14598), .Z(n14595) );
  ANDN U18695 ( .B(n14599), .A(n456), .Z(n14597) );
  XNOR U18696 ( .A(b[595]), .B(n14598), .Z(n14599) );
  XOR U18697 ( .A(n14600), .B(n14601), .Z(n14598) );
  ANDN U18698 ( .B(n14602), .A(n457), .Z(n14600) );
  XNOR U18699 ( .A(b[594]), .B(n14601), .Z(n14602) );
  XOR U18700 ( .A(n14603), .B(n14604), .Z(n14601) );
  ANDN U18701 ( .B(n14605), .A(n458), .Z(n14603) );
  XNOR U18702 ( .A(b[593]), .B(n14604), .Z(n14605) );
  XOR U18703 ( .A(n14606), .B(n14607), .Z(n14604) );
  ANDN U18704 ( .B(n14608), .A(n459), .Z(n14606) );
  XNOR U18705 ( .A(b[592]), .B(n14607), .Z(n14608) );
  XOR U18706 ( .A(n14609), .B(n14610), .Z(n14607) );
  ANDN U18707 ( .B(n14611), .A(n460), .Z(n14609) );
  XNOR U18708 ( .A(b[591]), .B(n14610), .Z(n14611) );
  XOR U18709 ( .A(n14612), .B(n14613), .Z(n14610) );
  ANDN U18710 ( .B(n14614), .A(n461), .Z(n14612) );
  XNOR U18711 ( .A(b[590]), .B(n14613), .Z(n14614) );
  XOR U18712 ( .A(n14615), .B(n14616), .Z(n14613) );
  ANDN U18713 ( .B(n14617), .A(n463), .Z(n14615) );
  XNOR U18714 ( .A(b[589]), .B(n14616), .Z(n14617) );
  XOR U18715 ( .A(n14618), .B(n14619), .Z(n14616) );
  ANDN U18716 ( .B(n14620), .A(n464), .Z(n14618) );
  XNOR U18717 ( .A(b[588]), .B(n14619), .Z(n14620) );
  XOR U18718 ( .A(n14621), .B(n14622), .Z(n14619) );
  ANDN U18719 ( .B(n14623), .A(n465), .Z(n14621) );
  XNOR U18720 ( .A(b[587]), .B(n14622), .Z(n14623) );
  XOR U18721 ( .A(n14624), .B(n14625), .Z(n14622) );
  ANDN U18722 ( .B(n14626), .A(n466), .Z(n14624) );
  XNOR U18723 ( .A(b[586]), .B(n14625), .Z(n14626) );
  XOR U18724 ( .A(n14627), .B(n14628), .Z(n14625) );
  ANDN U18725 ( .B(n14629), .A(n467), .Z(n14627) );
  XNOR U18726 ( .A(b[585]), .B(n14628), .Z(n14629) );
  XOR U18727 ( .A(n14630), .B(n14631), .Z(n14628) );
  ANDN U18728 ( .B(n14632), .A(n468), .Z(n14630) );
  XNOR U18729 ( .A(b[584]), .B(n14631), .Z(n14632) );
  XOR U18730 ( .A(n14633), .B(n14634), .Z(n14631) );
  ANDN U18731 ( .B(n14635), .A(n469), .Z(n14633) );
  XNOR U18732 ( .A(b[583]), .B(n14634), .Z(n14635) );
  XOR U18733 ( .A(n14636), .B(n14637), .Z(n14634) );
  ANDN U18734 ( .B(n14638), .A(n470), .Z(n14636) );
  XNOR U18735 ( .A(b[582]), .B(n14637), .Z(n14638) );
  XOR U18736 ( .A(n14639), .B(n14640), .Z(n14637) );
  ANDN U18737 ( .B(n14641), .A(n471), .Z(n14639) );
  XNOR U18738 ( .A(b[581]), .B(n14640), .Z(n14641) );
  XOR U18739 ( .A(n14642), .B(n14643), .Z(n14640) );
  ANDN U18740 ( .B(n14644), .A(n472), .Z(n14642) );
  XNOR U18741 ( .A(b[580]), .B(n14643), .Z(n14644) );
  XOR U18742 ( .A(n14645), .B(n14646), .Z(n14643) );
  ANDN U18743 ( .B(n14647), .A(n474), .Z(n14645) );
  XNOR U18744 ( .A(b[579]), .B(n14646), .Z(n14647) );
  XOR U18745 ( .A(n14648), .B(n14649), .Z(n14646) );
  ANDN U18746 ( .B(n14650), .A(n475), .Z(n14648) );
  XNOR U18747 ( .A(b[578]), .B(n14649), .Z(n14650) );
  XOR U18748 ( .A(n14651), .B(n14652), .Z(n14649) );
  ANDN U18749 ( .B(n14653), .A(n476), .Z(n14651) );
  XNOR U18750 ( .A(b[577]), .B(n14652), .Z(n14653) );
  XOR U18751 ( .A(n14654), .B(n14655), .Z(n14652) );
  ANDN U18752 ( .B(n14656), .A(n477), .Z(n14654) );
  XNOR U18753 ( .A(b[576]), .B(n14655), .Z(n14656) );
  XOR U18754 ( .A(n14657), .B(n14658), .Z(n14655) );
  ANDN U18755 ( .B(n14659), .A(n478), .Z(n14657) );
  XNOR U18756 ( .A(b[575]), .B(n14658), .Z(n14659) );
  XOR U18757 ( .A(n14660), .B(n14661), .Z(n14658) );
  ANDN U18758 ( .B(n14662), .A(n479), .Z(n14660) );
  XNOR U18759 ( .A(b[574]), .B(n14661), .Z(n14662) );
  XOR U18760 ( .A(n14663), .B(n14664), .Z(n14661) );
  ANDN U18761 ( .B(n14665), .A(n480), .Z(n14663) );
  XNOR U18762 ( .A(b[573]), .B(n14664), .Z(n14665) );
  XOR U18763 ( .A(n14666), .B(n14667), .Z(n14664) );
  ANDN U18764 ( .B(n14668), .A(n481), .Z(n14666) );
  XNOR U18765 ( .A(b[572]), .B(n14667), .Z(n14668) );
  XOR U18766 ( .A(n14669), .B(n14670), .Z(n14667) );
  ANDN U18767 ( .B(n14671), .A(n482), .Z(n14669) );
  XNOR U18768 ( .A(b[571]), .B(n14670), .Z(n14671) );
  XOR U18769 ( .A(n14672), .B(n14673), .Z(n14670) );
  ANDN U18770 ( .B(n14674), .A(n483), .Z(n14672) );
  XNOR U18771 ( .A(b[570]), .B(n14673), .Z(n14674) );
  XOR U18772 ( .A(n14675), .B(n14676), .Z(n14673) );
  ANDN U18773 ( .B(n14677), .A(n485), .Z(n14675) );
  XNOR U18774 ( .A(b[569]), .B(n14676), .Z(n14677) );
  XOR U18775 ( .A(n14678), .B(n14679), .Z(n14676) );
  ANDN U18776 ( .B(n14680), .A(n486), .Z(n14678) );
  XNOR U18777 ( .A(b[568]), .B(n14679), .Z(n14680) );
  XOR U18778 ( .A(n14681), .B(n14682), .Z(n14679) );
  ANDN U18779 ( .B(n14683), .A(n487), .Z(n14681) );
  XNOR U18780 ( .A(b[567]), .B(n14682), .Z(n14683) );
  XOR U18781 ( .A(n14684), .B(n14685), .Z(n14682) );
  ANDN U18782 ( .B(n14686), .A(n488), .Z(n14684) );
  XNOR U18783 ( .A(b[566]), .B(n14685), .Z(n14686) );
  XOR U18784 ( .A(n14687), .B(n14688), .Z(n14685) );
  ANDN U18785 ( .B(n14689), .A(n489), .Z(n14687) );
  XNOR U18786 ( .A(b[565]), .B(n14688), .Z(n14689) );
  XOR U18787 ( .A(n14690), .B(n14691), .Z(n14688) );
  ANDN U18788 ( .B(n14692), .A(n490), .Z(n14690) );
  XNOR U18789 ( .A(b[564]), .B(n14691), .Z(n14692) );
  XOR U18790 ( .A(n14693), .B(n14694), .Z(n14691) );
  ANDN U18791 ( .B(n14695), .A(n491), .Z(n14693) );
  XNOR U18792 ( .A(b[563]), .B(n14694), .Z(n14695) );
  XOR U18793 ( .A(n14696), .B(n14697), .Z(n14694) );
  ANDN U18794 ( .B(n14698), .A(n492), .Z(n14696) );
  XNOR U18795 ( .A(b[562]), .B(n14697), .Z(n14698) );
  XOR U18796 ( .A(n14699), .B(n14700), .Z(n14697) );
  ANDN U18797 ( .B(n14701), .A(n493), .Z(n14699) );
  XNOR U18798 ( .A(b[561]), .B(n14700), .Z(n14701) );
  XOR U18799 ( .A(n14702), .B(n14703), .Z(n14700) );
  ANDN U18800 ( .B(n14704), .A(n494), .Z(n14702) );
  XNOR U18801 ( .A(b[560]), .B(n14703), .Z(n14704) );
  XOR U18802 ( .A(n14705), .B(n14706), .Z(n14703) );
  ANDN U18803 ( .B(n14707), .A(n496), .Z(n14705) );
  XNOR U18804 ( .A(b[559]), .B(n14706), .Z(n14707) );
  XOR U18805 ( .A(n14708), .B(n14709), .Z(n14706) );
  ANDN U18806 ( .B(n14710), .A(n497), .Z(n14708) );
  XNOR U18807 ( .A(b[558]), .B(n14709), .Z(n14710) );
  XOR U18808 ( .A(n14711), .B(n14712), .Z(n14709) );
  ANDN U18809 ( .B(n14713), .A(n498), .Z(n14711) );
  XNOR U18810 ( .A(b[557]), .B(n14712), .Z(n14713) );
  XOR U18811 ( .A(n14714), .B(n14715), .Z(n14712) );
  ANDN U18812 ( .B(n14716), .A(n499), .Z(n14714) );
  XNOR U18813 ( .A(b[556]), .B(n14715), .Z(n14716) );
  XOR U18814 ( .A(n14717), .B(n14718), .Z(n14715) );
  ANDN U18815 ( .B(n14719), .A(n500), .Z(n14717) );
  XNOR U18816 ( .A(b[555]), .B(n14718), .Z(n14719) );
  XOR U18817 ( .A(n14720), .B(n14721), .Z(n14718) );
  ANDN U18818 ( .B(n14722), .A(n501), .Z(n14720) );
  XNOR U18819 ( .A(b[554]), .B(n14721), .Z(n14722) );
  XOR U18820 ( .A(n14723), .B(n14724), .Z(n14721) );
  ANDN U18821 ( .B(n14725), .A(n502), .Z(n14723) );
  XNOR U18822 ( .A(b[553]), .B(n14724), .Z(n14725) );
  XOR U18823 ( .A(n14726), .B(n14727), .Z(n14724) );
  ANDN U18824 ( .B(n14728), .A(n503), .Z(n14726) );
  XNOR U18825 ( .A(b[552]), .B(n14727), .Z(n14728) );
  XOR U18826 ( .A(n14729), .B(n14730), .Z(n14727) );
  ANDN U18827 ( .B(n14731), .A(n504), .Z(n14729) );
  XNOR U18828 ( .A(b[551]), .B(n14730), .Z(n14731) );
  XOR U18829 ( .A(n14732), .B(n14733), .Z(n14730) );
  ANDN U18830 ( .B(n14734), .A(n505), .Z(n14732) );
  XNOR U18831 ( .A(b[550]), .B(n14733), .Z(n14734) );
  XOR U18832 ( .A(n14735), .B(n14736), .Z(n14733) );
  ANDN U18833 ( .B(n14737), .A(n507), .Z(n14735) );
  XNOR U18834 ( .A(b[549]), .B(n14736), .Z(n14737) );
  XOR U18835 ( .A(n14738), .B(n14739), .Z(n14736) );
  ANDN U18836 ( .B(n14740), .A(n508), .Z(n14738) );
  XNOR U18837 ( .A(b[548]), .B(n14739), .Z(n14740) );
  XOR U18838 ( .A(n14741), .B(n14742), .Z(n14739) );
  ANDN U18839 ( .B(n14743), .A(n509), .Z(n14741) );
  XNOR U18840 ( .A(b[547]), .B(n14742), .Z(n14743) );
  XOR U18841 ( .A(n14744), .B(n14745), .Z(n14742) );
  ANDN U18842 ( .B(n14746), .A(n510), .Z(n14744) );
  XNOR U18843 ( .A(b[546]), .B(n14745), .Z(n14746) );
  XOR U18844 ( .A(n14747), .B(n14748), .Z(n14745) );
  ANDN U18845 ( .B(n14749), .A(n511), .Z(n14747) );
  XNOR U18846 ( .A(b[545]), .B(n14748), .Z(n14749) );
  XOR U18847 ( .A(n14750), .B(n14751), .Z(n14748) );
  ANDN U18848 ( .B(n14752), .A(n512), .Z(n14750) );
  XNOR U18849 ( .A(b[544]), .B(n14751), .Z(n14752) );
  XOR U18850 ( .A(n14753), .B(n14754), .Z(n14751) );
  ANDN U18851 ( .B(n14755), .A(n513), .Z(n14753) );
  XNOR U18852 ( .A(b[543]), .B(n14754), .Z(n14755) );
  XOR U18853 ( .A(n14756), .B(n14757), .Z(n14754) );
  ANDN U18854 ( .B(n14758), .A(n514), .Z(n14756) );
  XNOR U18855 ( .A(b[542]), .B(n14757), .Z(n14758) );
  XOR U18856 ( .A(n14759), .B(n14760), .Z(n14757) );
  ANDN U18857 ( .B(n14761), .A(n515), .Z(n14759) );
  XNOR U18858 ( .A(b[541]), .B(n14760), .Z(n14761) );
  XOR U18859 ( .A(n14762), .B(n14763), .Z(n14760) );
  ANDN U18860 ( .B(n14764), .A(n516), .Z(n14762) );
  XNOR U18861 ( .A(b[540]), .B(n14763), .Z(n14764) );
  XOR U18862 ( .A(n14765), .B(n14766), .Z(n14763) );
  ANDN U18863 ( .B(n14767), .A(n518), .Z(n14765) );
  XNOR U18864 ( .A(b[539]), .B(n14766), .Z(n14767) );
  XOR U18865 ( .A(n14768), .B(n14769), .Z(n14766) );
  ANDN U18866 ( .B(n14770), .A(n519), .Z(n14768) );
  XNOR U18867 ( .A(b[538]), .B(n14769), .Z(n14770) );
  XOR U18868 ( .A(n14771), .B(n14772), .Z(n14769) );
  ANDN U18869 ( .B(n14773), .A(n520), .Z(n14771) );
  XNOR U18870 ( .A(b[537]), .B(n14772), .Z(n14773) );
  XOR U18871 ( .A(n14774), .B(n14775), .Z(n14772) );
  ANDN U18872 ( .B(n14776), .A(n521), .Z(n14774) );
  XNOR U18873 ( .A(b[536]), .B(n14775), .Z(n14776) );
  XOR U18874 ( .A(n14777), .B(n14778), .Z(n14775) );
  ANDN U18875 ( .B(n14779), .A(n522), .Z(n14777) );
  XNOR U18876 ( .A(b[535]), .B(n14778), .Z(n14779) );
  XOR U18877 ( .A(n14780), .B(n14781), .Z(n14778) );
  ANDN U18878 ( .B(n14782), .A(n523), .Z(n14780) );
  XNOR U18879 ( .A(b[534]), .B(n14781), .Z(n14782) );
  XOR U18880 ( .A(n14783), .B(n14784), .Z(n14781) );
  ANDN U18881 ( .B(n14785), .A(n524), .Z(n14783) );
  XNOR U18882 ( .A(b[533]), .B(n14784), .Z(n14785) );
  XOR U18883 ( .A(n14786), .B(n14787), .Z(n14784) );
  ANDN U18884 ( .B(n14788), .A(n525), .Z(n14786) );
  XNOR U18885 ( .A(b[532]), .B(n14787), .Z(n14788) );
  XOR U18886 ( .A(n14789), .B(n14790), .Z(n14787) );
  ANDN U18887 ( .B(n14791), .A(n526), .Z(n14789) );
  XNOR U18888 ( .A(b[531]), .B(n14790), .Z(n14791) );
  XOR U18889 ( .A(n14792), .B(n14793), .Z(n14790) );
  ANDN U18890 ( .B(n14794), .A(n527), .Z(n14792) );
  XNOR U18891 ( .A(b[530]), .B(n14793), .Z(n14794) );
  XOR U18892 ( .A(n14795), .B(n14796), .Z(n14793) );
  ANDN U18893 ( .B(n14797), .A(n529), .Z(n14795) );
  XNOR U18894 ( .A(b[529]), .B(n14796), .Z(n14797) );
  XOR U18895 ( .A(n14798), .B(n14799), .Z(n14796) );
  ANDN U18896 ( .B(n14800), .A(n530), .Z(n14798) );
  XNOR U18897 ( .A(b[528]), .B(n14799), .Z(n14800) );
  XOR U18898 ( .A(n14801), .B(n14802), .Z(n14799) );
  ANDN U18899 ( .B(n14803), .A(n531), .Z(n14801) );
  XNOR U18900 ( .A(b[527]), .B(n14802), .Z(n14803) );
  XOR U18901 ( .A(n14804), .B(n14805), .Z(n14802) );
  ANDN U18902 ( .B(n14806), .A(n532), .Z(n14804) );
  XNOR U18903 ( .A(b[526]), .B(n14805), .Z(n14806) );
  XOR U18904 ( .A(n14807), .B(n14808), .Z(n14805) );
  ANDN U18905 ( .B(n14809), .A(n533), .Z(n14807) );
  XNOR U18906 ( .A(b[525]), .B(n14808), .Z(n14809) );
  XOR U18907 ( .A(n14810), .B(n14811), .Z(n14808) );
  ANDN U18908 ( .B(n14812), .A(n534), .Z(n14810) );
  XNOR U18909 ( .A(b[524]), .B(n14811), .Z(n14812) );
  XOR U18910 ( .A(n14813), .B(n14814), .Z(n14811) );
  ANDN U18911 ( .B(n14815), .A(n535), .Z(n14813) );
  XNOR U18912 ( .A(b[523]), .B(n14814), .Z(n14815) );
  XOR U18913 ( .A(n14816), .B(n14817), .Z(n14814) );
  ANDN U18914 ( .B(n14818), .A(n536), .Z(n14816) );
  XNOR U18915 ( .A(b[522]), .B(n14817), .Z(n14818) );
  XOR U18916 ( .A(n14819), .B(n14820), .Z(n14817) );
  ANDN U18917 ( .B(n14821), .A(n537), .Z(n14819) );
  XNOR U18918 ( .A(b[521]), .B(n14820), .Z(n14821) );
  XOR U18919 ( .A(n14822), .B(n14823), .Z(n14820) );
  ANDN U18920 ( .B(n14824), .A(n538), .Z(n14822) );
  XNOR U18921 ( .A(b[520]), .B(n14823), .Z(n14824) );
  XOR U18922 ( .A(n14825), .B(n14826), .Z(n14823) );
  ANDN U18923 ( .B(n14827), .A(n540), .Z(n14825) );
  XNOR U18924 ( .A(b[519]), .B(n14826), .Z(n14827) );
  XOR U18925 ( .A(n14828), .B(n14829), .Z(n14826) );
  ANDN U18926 ( .B(n14830), .A(n541), .Z(n14828) );
  XNOR U18927 ( .A(b[518]), .B(n14829), .Z(n14830) );
  XOR U18928 ( .A(n14831), .B(n14832), .Z(n14829) );
  ANDN U18929 ( .B(n14833), .A(n542), .Z(n14831) );
  XNOR U18930 ( .A(b[517]), .B(n14832), .Z(n14833) );
  XOR U18931 ( .A(n14834), .B(n14835), .Z(n14832) );
  ANDN U18932 ( .B(n14836), .A(n543), .Z(n14834) );
  XNOR U18933 ( .A(b[516]), .B(n14835), .Z(n14836) );
  XOR U18934 ( .A(n14837), .B(n14838), .Z(n14835) );
  ANDN U18935 ( .B(n14839), .A(n544), .Z(n14837) );
  XNOR U18936 ( .A(b[515]), .B(n14838), .Z(n14839) );
  XOR U18937 ( .A(n14840), .B(n14841), .Z(n14838) );
  ANDN U18938 ( .B(n14842), .A(n545), .Z(n14840) );
  XNOR U18939 ( .A(b[514]), .B(n14841), .Z(n14842) );
  XOR U18940 ( .A(n14843), .B(n14844), .Z(n14841) );
  ANDN U18941 ( .B(n14845), .A(n546), .Z(n14843) );
  XNOR U18942 ( .A(b[513]), .B(n14844), .Z(n14845) );
  XOR U18943 ( .A(n14846), .B(n14847), .Z(n14844) );
  ANDN U18944 ( .B(n14848), .A(n547), .Z(n14846) );
  XNOR U18945 ( .A(b[512]), .B(n14847), .Z(n14848) );
  XOR U18946 ( .A(n14849), .B(n14850), .Z(n14847) );
  ANDN U18947 ( .B(n14851), .A(n548), .Z(n14849) );
  XNOR U18948 ( .A(b[511]), .B(n14850), .Z(n14851) );
  XOR U18949 ( .A(n14852), .B(n14853), .Z(n14850) );
  ANDN U18950 ( .B(n14854), .A(n549), .Z(n14852) );
  XNOR U18951 ( .A(b[510]), .B(n14853), .Z(n14854) );
  XOR U18952 ( .A(n14855), .B(n14856), .Z(n14853) );
  ANDN U18953 ( .B(n14857), .A(n551), .Z(n14855) );
  XNOR U18954 ( .A(b[509]), .B(n14856), .Z(n14857) );
  XOR U18955 ( .A(n14858), .B(n14859), .Z(n14856) );
  ANDN U18956 ( .B(n14860), .A(n552), .Z(n14858) );
  XNOR U18957 ( .A(b[508]), .B(n14859), .Z(n14860) );
  XOR U18958 ( .A(n14861), .B(n14862), .Z(n14859) );
  ANDN U18959 ( .B(n14863), .A(n553), .Z(n14861) );
  XNOR U18960 ( .A(b[507]), .B(n14862), .Z(n14863) );
  XOR U18961 ( .A(n14864), .B(n14865), .Z(n14862) );
  ANDN U18962 ( .B(n14866), .A(n554), .Z(n14864) );
  XNOR U18963 ( .A(b[506]), .B(n14865), .Z(n14866) );
  XOR U18964 ( .A(n14867), .B(n14868), .Z(n14865) );
  ANDN U18965 ( .B(n14869), .A(n555), .Z(n14867) );
  XNOR U18966 ( .A(b[505]), .B(n14868), .Z(n14869) );
  XOR U18967 ( .A(n14870), .B(n14871), .Z(n14868) );
  ANDN U18968 ( .B(n14872), .A(n556), .Z(n14870) );
  XNOR U18969 ( .A(b[504]), .B(n14871), .Z(n14872) );
  XOR U18970 ( .A(n14873), .B(n14874), .Z(n14871) );
  ANDN U18971 ( .B(n14875), .A(n557), .Z(n14873) );
  XNOR U18972 ( .A(b[503]), .B(n14874), .Z(n14875) );
  XOR U18973 ( .A(n14876), .B(n14877), .Z(n14874) );
  ANDN U18974 ( .B(n14878), .A(n558), .Z(n14876) );
  XNOR U18975 ( .A(b[502]), .B(n14877), .Z(n14878) );
  XOR U18976 ( .A(n14879), .B(n14880), .Z(n14877) );
  ANDN U18977 ( .B(n14881), .A(n559), .Z(n14879) );
  XNOR U18978 ( .A(b[501]), .B(n14880), .Z(n14881) );
  XOR U18979 ( .A(n14882), .B(n14883), .Z(n14880) );
  ANDN U18980 ( .B(n14884), .A(n560), .Z(n14882) );
  XNOR U18981 ( .A(b[500]), .B(n14883), .Z(n14884) );
  XOR U18982 ( .A(n14885), .B(n14886), .Z(n14883) );
  ANDN U18983 ( .B(n14887), .A(n563), .Z(n14885) );
  XNOR U18984 ( .A(b[499]), .B(n14886), .Z(n14887) );
  XOR U18985 ( .A(n14888), .B(n14889), .Z(n14886) );
  ANDN U18986 ( .B(n14890), .A(n564), .Z(n14888) );
  XNOR U18987 ( .A(b[498]), .B(n14889), .Z(n14890) );
  XOR U18988 ( .A(n14891), .B(n14892), .Z(n14889) );
  ANDN U18989 ( .B(n14893), .A(n565), .Z(n14891) );
  XNOR U18990 ( .A(b[497]), .B(n14892), .Z(n14893) );
  XOR U18991 ( .A(n14894), .B(n14895), .Z(n14892) );
  ANDN U18992 ( .B(n14896), .A(n566), .Z(n14894) );
  XNOR U18993 ( .A(b[496]), .B(n14895), .Z(n14896) );
  XOR U18994 ( .A(n14897), .B(n14898), .Z(n14895) );
  ANDN U18995 ( .B(n14899), .A(n567), .Z(n14897) );
  XNOR U18996 ( .A(b[495]), .B(n14898), .Z(n14899) );
  XOR U18997 ( .A(n14900), .B(n14901), .Z(n14898) );
  ANDN U18998 ( .B(n14902), .A(n568), .Z(n14900) );
  XNOR U18999 ( .A(b[494]), .B(n14901), .Z(n14902) );
  XOR U19000 ( .A(n14903), .B(n14904), .Z(n14901) );
  ANDN U19001 ( .B(n14905), .A(n569), .Z(n14903) );
  XNOR U19002 ( .A(b[493]), .B(n14904), .Z(n14905) );
  XOR U19003 ( .A(n14906), .B(n14907), .Z(n14904) );
  ANDN U19004 ( .B(n14908), .A(n570), .Z(n14906) );
  XNOR U19005 ( .A(b[492]), .B(n14907), .Z(n14908) );
  XOR U19006 ( .A(n14909), .B(n14910), .Z(n14907) );
  ANDN U19007 ( .B(n14911), .A(n571), .Z(n14909) );
  XNOR U19008 ( .A(b[491]), .B(n14910), .Z(n14911) );
  XOR U19009 ( .A(n14912), .B(n14913), .Z(n14910) );
  ANDN U19010 ( .B(n14914), .A(n572), .Z(n14912) );
  XNOR U19011 ( .A(b[490]), .B(n14913), .Z(n14914) );
  XOR U19012 ( .A(n14915), .B(n14916), .Z(n14913) );
  ANDN U19013 ( .B(n14917), .A(n574), .Z(n14915) );
  XNOR U19014 ( .A(b[489]), .B(n14916), .Z(n14917) );
  XOR U19015 ( .A(n14918), .B(n14919), .Z(n14916) );
  ANDN U19016 ( .B(n14920), .A(n575), .Z(n14918) );
  XNOR U19017 ( .A(b[488]), .B(n14919), .Z(n14920) );
  XOR U19018 ( .A(n14921), .B(n14922), .Z(n14919) );
  ANDN U19019 ( .B(n14923), .A(n576), .Z(n14921) );
  XNOR U19020 ( .A(b[487]), .B(n14922), .Z(n14923) );
  XOR U19021 ( .A(n14924), .B(n14925), .Z(n14922) );
  ANDN U19022 ( .B(n14926), .A(n577), .Z(n14924) );
  XNOR U19023 ( .A(b[486]), .B(n14925), .Z(n14926) );
  XOR U19024 ( .A(n14927), .B(n14928), .Z(n14925) );
  ANDN U19025 ( .B(n14929), .A(n578), .Z(n14927) );
  XNOR U19026 ( .A(b[485]), .B(n14928), .Z(n14929) );
  XOR U19027 ( .A(n14930), .B(n14931), .Z(n14928) );
  ANDN U19028 ( .B(n14932), .A(n579), .Z(n14930) );
  XNOR U19029 ( .A(b[484]), .B(n14931), .Z(n14932) );
  XOR U19030 ( .A(n14933), .B(n14934), .Z(n14931) );
  ANDN U19031 ( .B(n14935), .A(n580), .Z(n14933) );
  XNOR U19032 ( .A(b[483]), .B(n14934), .Z(n14935) );
  XOR U19033 ( .A(n14936), .B(n14937), .Z(n14934) );
  ANDN U19034 ( .B(n14938), .A(n581), .Z(n14936) );
  XNOR U19035 ( .A(b[482]), .B(n14937), .Z(n14938) );
  XOR U19036 ( .A(n14939), .B(n14940), .Z(n14937) );
  ANDN U19037 ( .B(n14941), .A(n582), .Z(n14939) );
  XNOR U19038 ( .A(b[481]), .B(n14940), .Z(n14941) );
  XOR U19039 ( .A(n14942), .B(n14943), .Z(n14940) );
  ANDN U19040 ( .B(n14944), .A(n583), .Z(n14942) );
  XNOR U19041 ( .A(b[480]), .B(n14943), .Z(n14944) );
  XOR U19042 ( .A(n14945), .B(n14946), .Z(n14943) );
  ANDN U19043 ( .B(n14947), .A(n585), .Z(n14945) );
  XNOR U19044 ( .A(b[479]), .B(n14946), .Z(n14947) );
  XOR U19045 ( .A(n14948), .B(n14949), .Z(n14946) );
  ANDN U19046 ( .B(n14950), .A(n586), .Z(n14948) );
  XNOR U19047 ( .A(b[478]), .B(n14949), .Z(n14950) );
  XOR U19048 ( .A(n14951), .B(n14952), .Z(n14949) );
  ANDN U19049 ( .B(n14953), .A(n587), .Z(n14951) );
  XNOR U19050 ( .A(b[477]), .B(n14952), .Z(n14953) );
  XOR U19051 ( .A(n14954), .B(n14955), .Z(n14952) );
  ANDN U19052 ( .B(n14956), .A(n588), .Z(n14954) );
  XNOR U19053 ( .A(b[476]), .B(n14955), .Z(n14956) );
  XOR U19054 ( .A(n14957), .B(n14958), .Z(n14955) );
  ANDN U19055 ( .B(n14959), .A(n589), .Z(n14957) );
  XNOR U19056 ( .A(b[475]), .B(n14958), .Z(n14959) );
  XOR U19057 ( .A(n14960), .B(n14961), .Z(n14958) );
  ANDN U19058 ( .B(n14962), .A(n590), .Z(n14960) );
  XNOR U19059 ( .A(b[474]), .B(n14961), .Z(n14962) );
  XOR U19060 ( .A(n14963), .B(n14964), .Z(n14961) );
  ANDN U19061 ( .B(n14965), .A(n591), .Z(n14963) );
  XNOR U19062 ( .A(b[473]), .B(n14964), .Z(n14965) );
  XOR U19063 ( .A(n14966), .B(n14967), .Z(n14964) );
  ANDN U19064 ( .B(n14968), .A(n592), .Z(n14966) );
  XNOR U19065 ( .A(b[472]), .B(n14967), .Z(n14968) );
  XOR U19066 ( .A(n14969), .B(n14970), .Z(n14967) );
  ANDN U19067 ( .B(n14971), .A(n593), .Z(n14969) );
  XNOR U19068 ( .A(b[471]), .B(n14970), .Z(n14971) );
  XOR U19069 ( .A(n14972), .B(n14973), .Z(n14970) );
  ANDN U19070 ( .B(n14974), .A(n594), .Z(n14972) );
  XNOR U19071 ( .A(b[470]), .B(n14973), .Z(n14974) );
  XOR U19072 ( .A(n14975), .B(n14976), .Z(n14973) );
  ANDN U19073 ( .B(n14977), .A(n596), .Z(n14975) );
  XNOR U19074 ( .A(b[469]), .B(n14976), .Z(n14977) );
  XOR U19075 ( .A(n14978), .B(n14979), .Z(n14976) );
  ANDN U19076 ( .B(n14980), .A(n597), .Z(n14978) );
  XNOR U19077 ( .A(b[468]), .B(n14979), .Z(n14980) );
  XOR U19078 ( .A(n14981), .B(n14982), .Z(n14979) );
  ANDN U19079 ( .B(n14983), .A(n598), .Z(n14981) );
  XNOR U19080 ( .A(b[467]), .B(n14982), .Z(n14983) );
  XOR U19081 ( .A(n14984), .B(n14985), .Z(n14982) );
  ANDN U19082 ( .B(n14986), .A(n599), .Z(n14984) );
  XNOR U19083 ( .A(b[466]), .B(n14985), .Z(n14986) );
  XOR U19084 ( .A(n14987), .B(n14988), .Z(n14985) );
  ANDN U19085 ( .B(n14989), .A(n600), .Z(n14987) );
  XNOR U19086 ( .A(b[465]), .B(n14988), .Z(n14989) );
  XOR U19087 ( .A(n14990), .B(n14991), .Z(n14988) );
  ANDN U19088 ( .B(n14992), .A(n601), .Z(n14990) );
  XNOR U19089 ( .A(b[464]), .B(n14991), .Z(n14992) );
  XOR U19090 ( .A(n14993), .B(n14994), .Z(n14991) );
  ANDN U19091 ( .B(n14995), .A(n602), .Z(n14993) );
  XNOR U19092 ( .A(b[463]), .B(n14994), .Z(n14995) );
  XOR U19093 ( .A(n14996), .B(n14997), .Z(n14994) );
  ANDN U19094 ( .B(n14998), .A(n603), .Z(n14996) );
  XNOR U19095 ( .A(b[462]), .B(n14997), .Z(n14998) );
  XOR U19096 ( .A(n14999), .B(n15000), .Z(n14997) );
  ANDN U19097 ( .B(n15001), .A(n604), .Z(n14999) );
  XNOR U19098 ( .A(b[461]), .B(n15000), .Z(n15001) );
  XOR U19099 ( .A(n15002), .B(n15003), .Z(n15000) );
  ANDN U19100 ( .B(n15004), .A(n605), .Z(n15002) );
  XNOR U19101 ( .A(b[460]), .B(n15003), .Z(n15004) );
  XOR U19102 ( .A(n15005), .B(n15006), .Z(n15003) );
  ANDN U19103 ( .B(n15007), .A(n607), .Z(n15005) );
  XNOR U19104 ( .A(b[459]), .B(n15006), .Z(n15007) );
  XOR U19105 ( .A(n15008), .B(n15009), .Z(n15006) );
  ANDN U19106 ( .B(n15010), .A(n608), .Z(n15008) );
  XNOR U19107 ( .A(b[458]), .B(n15009), .Z(n15010) );
  XOR U19108 ( .A(n15011), .B(n15012), .Z(n15009) );
  ANDN U19109 ( .B(n15013), .A(n609), .Z(n15011) );
  XNOR U19110 ( .A(b[457]), .B(n15012), .Z(n15013) );
  XOR U19111 ( .A(n15014), .B(n15015), .Z(n15012) );
  ANDN U19112 ( .B(n15016), .A(n610), .Z(n15014) );
  XNOR U19113 ( .A(b[456]), .B(n15015), .Z(n15016) );
  XOR U19114 ( .A(n15017), .B(n15018), .Z(n15015) );
  ANDN U19115 ( .B(n15019), .A(n611), .Z(n15017) );
  XNOR U19116 ( .A(b[455]), .B(n15018), .Z(n15019) );
  XOR U19117 ( .A(n15020), .B(n15021), .Z(n15018) );
  ANDN U19118 ( .B(n15022), .A(n612), .Z(n15020) );
  XNOR U19119 ( .A(b[454]), .B(n15021), .Z(n15022) );
  XOR U19120 ( .A(n15023), .B(n15024), .Z(n15021) );
  ANDN U19121 ( .B(n15025), .A(n613), .Z(n15023) );
  XNOR U19122 ( .A(b[453]), .B(n15024), .Z(n15025) );
  XOR U19123 ( .A(n15026), .B(n15027), .Z(n15024) );
  ANDN U19124 ( .B(n15028), .A(n614), .Z(n15026) );
  XNOR U19125 ( .A(b[452]), .B(n15027), .Z(n15028) );
  XOR U19126 ( .A(n15029), .B(n15030), .Z(n15027) );
  ANDN U19127 ( .B(n15031), .A(n615), .Z(n15029) );
  XNOR U19128 ( .A(b[451]), .B(n15030), .Z(n15031) );
  XOR U19129 ( .A(n15032), .B(n15033), .Z(n15030) );
  ANDN U19130 ( .B(n15034), .A(n616), .Z(n15032) );
  XNOR U19131 ( .A(b[450]), .B(n15033), .Z(n15034) );
  XOR U19132 ( .A(n15035), .B(n15036), .Z(n15033) );
  ANDN U19133 ( .B(n15037), .A(n618), .Z(n15035) );
  XNOR U19134 ( .A(b[449]), .B(n15036), .Z(n15037) );
  XOR U19135 ( .A(n15038), .B(n15039), .Z(n15036) );
  ANDN U19136 ( .B(n15040), .A(n619), .Z(n15038) );
  XNOR U19137 ( .A(b[448]), .B(n15039), .Z(n15040) );
  XOR U19138 ( .A(n15041), .B(n15042), .Z(n15039) );
  ANDN U19139 ( .B(n15043), .A(n620), .Z(n15041) );
  XNOR U19140 ( .A(b[447]), .B(n15042), .Z(n15043) );
  XOR U19141 ( .A(n15044), .B(n15045), .Z(n15042) );
  ANDN U19142 ( .B(n15046), .A(n621), .Z(n15044) );
  XNOR U19143 ( .A(b[446]), .B(n15045), .Z(n15046) );
  XOR U19144 ( .A(n15047), .B(n15048), .Z(n15045) );
  ANDN U19145 ( .B(n15049), .A(n622), .Z(n15047) );
  XNOR U19146 ( .A(b[445]), .B(n15048), .Z(n15049) );
  XOR U19147 ( .A(n15050), .B(n15051), .Z(n15048) );
  ANDN U19148 ( .B(n15052), .A(n623), .Z(n15050) );
  XNOR U19149 ( .A(b[444]), .B(n15051), .Z(n15052) );
  XOR U19150 ( .A(n15053), .B(n15054), .Z(n15051) );
  ANDN U19151 ( .B(n15055), .A(n624), .Z(n15053) );
  XNOR U19152 ( .A(b[443]), .B(n15054), .Z(n15055) );
  XOR U19153 ( .A(n15056), .B(n15057), .Z(n15054) );
  ANDN U19154 ( .B(n15058), .A(n625), .Z(n15056) );
  XNOR U19155 ( .A(b[442]), .B(n15057), .Z(n15058) );
  XOR U19156 ( .A(n15059), .B(n15060), .Z(n15057) );
  ANDN U19157 ( .B(n15061), .A(n626), .Z(n15059) );
  XNOR U19158 ( .A(b[441]), .B(n15060), .Z(n15061) );
  XOR U19159 ( .A(n15062), .B(n15063), .Z(n15060) );
  ANDN U19160 ( .B(n15064), .A(n627), .Z(n15062) );
  XNOR U19161 ( .A(b[440]), .B(n15063), .Z(n15064) );
  XOR U19162 ( .A(n15065), .B(n15066), .Z(n15063) );
  ANDN U19163 ( .B(n15067), .A(n629), .Z(n15065) );
  XNOR U19164 ( .A(b[439]), .B(n15066), .Z(n15067) );
  XOR U19165 ( .A(n15068), .B(n15069), .Z(n15066) );
  ANDN U19166 ( .B(n15070), .A(n630), .Z(n15068) );
  XNOR U19167 ( .A(b[438]), .B(n15069), .Z(n15070) );
  XOR U19168 ( .A(n15071), .B(n15072), .Z(n15069) );
  ANDN U19169 ( .B(n15073), .A(n631), .Z(n15071) );
  XNOR U19170 ( .A(b[437]), .B(n15072), .Z(n15073) );
  XOR U19171 ( .A(n15074), .B(n15075), .Z(n15072) );
  ANDN U19172 ( .B(n15076), .A(n632), .Z(n15074) );
  XNOR U19173 ( .A(b[436]), .B(n15075), .Z(n15076) );
  XOR U19174 ( .A(n15077), .B(n15078), .Z(n15075) );
  ANDN U19175 ( .B(n15079), .A(n633), .Z(n15077) );
  XNOR U19176 ( .A(b[435]), .B(n15078), .Z(n15079) );
  XOR U19177 ( .A(n15080), .B(n15081), .Z(n15078) );
  ANDN U19178 ( .B(n15082), .A(n634), .Z(n15080) );
  XNOR U19179 ( .A(b[434]), .B(n15081), .Z(n15082) );
  XOR U19180 ( .A(n15083), .B(n15084), .Z(n15081) );
  ANDN U19181 ( .B(n15085), .A(n635), .Z(n15083) );
  XNOR U19182 ( .A(b[433]), .B(n15084), .Z(n15085) );
  XOR U19183 ( .A(n15086), .B(n15087), .Z(n15084) );
  ANDN U19184 ( .B(n15088), .A(n636), .Z(n15086) );
  XNOR U19185 ( .A(b[432]), .B(n15087), .Z(n15088) );
  XOR U19186 ( .A(n15089), .B(n15090), .Z(n15087) );
  ANDN U19187 ( .B(n15091), .A(n637), .Z(n15089) );
  XNOR U19188 ( .A(b[431]), .B(n15090), .Z(n15091) );
  XOR U19189 ( .A(n15092), .B(n15093), .Z(n15090) );
  ANDN U19190 ( .B(n15094), .A(n638), .Z(n15092) );
  XNOR U19191 ( .A(b[430]), .B(n15093), .Z(n15094) );
  XOR U19192 ( .A(n15095), .B(n15096), .Z(n15093) );
  ANDN U19193 ( .B(n15097), .A(n640), .Z(n15095) );
  XNOR U19194 ( .A(b[429]), .B(n15096), .Z(n15097) );
  XOR U19195 ( .A(n15098), .B(n15099), .Z(n15096) );
  ANDN U19196 ( .B(n15100), .A(n641), .Z(n15098) );
  XNOR U19197 ( .A(b[428]), .B(n15099), .Z(n15100) );
  XOR U19198 ( .A(n15101), .B(n15102), .Z(n15099) );
  ANDN U19199 ( .B(n15103), .A(n642), .Z(n15101) );
  XNOR U19200 ( .A(b[427]), .B(n15102), .Z(n15103) );
  XOR U19201 ( .A(n15104), .B(n15105), .Z(n15102) );
  ANDN U19202 ( .B(n15106), .A(n643), .Z(n15104) );
  XNOR U19203 ( .A(b[426]), .B(n15105), .Z(n15106) );
  XOR U19204 ( .A(n15107), .B(n15108), .Z(n15105) );
  ANDN U19205 ( .B(n15109), .A(n644), .Z(n15107) );
  XNOR U19206 ( .A(b[425]), .B(n15108), .Z(n15109) );
  XOR U19207 ( .A(n15110), .B(n15111), .Z(n15108) );
  ANDN U19208 ( .B(n15112), .A(n645), .Z(n15110) );
  XNOR U19209 ( .A(b[424]), .B(n15111), .Z(n15112) );
  XOR U19210 ( .A(n15113), .B(n15114), .Z(n15111) );
  ANDN U19211 ( .B(n15115), .A(n646), .Z(n15113) );
  XNOR U19212 ( .A(b[423]), .B(n15114), .Z(n15115) );
  XOR U19213 ( .A(n15116), .B(n15117), .Z(n15114) );
  ANDN U19214 ( .B(n15118), .A(n647), .Z(n15116) );
  XNOR U19215 ( .A(b[422]), .B(n15117), .Z(n15118) );
  XOR U19216 ( .A(n15119), .B(n15120), .Z(n15117) );
  ANDN U19217 ( .B(n15121), .A(n648), .Z(n15119) );
  XNOR U19218 ( .A(b[421]), .B(n15120), .Z(n15121) );
  XOR U19219 ( .A(n15122), .B(n15123), .Z(n15120) );
  ANDN U19220 ( .B(n15124), .A(n649), .Z(n15122) );
  XNOR U19221 ( .A(b[420]), .B(n15123), .Z(n15124) );
  XOR U19222 ( .A(n15125), .B(n15126), .Z(n15123) );
  ANDN U19223 ( .B(n15127), .A(n651), .Z(n15125) );
  XNOR U19224 ( .A(b[419]), .B(n15126), .Z(n15127) );
  XOR U19225 ( .A(n15128), .B(n15129), .Z(n15126) );
  ANDN U19226 ( .B(n15130), .A(n652), .Z(n15128) );
  XNOR U19227 ( .A(b[418]), .B(n15129), .Z(n15130) );
  XOR U19228 ( .A(n15131), .B(n15132), .Z(n15129) );
  ANDN U19229 ( .B(n15133), .A(n653), .Z(n15131) );
  XNOR U19230 ( .A(b[417]), .B(n15132), .Z(n15133) );
  XOR U19231 ( .A(n15134), .B(n15135), .Z(n15132) );
  ANDN U19232 ( .B(n15136), .A(n654), .Z(n15134) );
  XNOR U19233 ( .A(b[416]), .B(n15135), .Z(n15136) );
  XOR U19234 ( .A(n15137), .B(n15138), .Z(n15135) );
  ANDN U19235 ( .B(n15139), .A(n655), .Z(n15137) );
  XNOR U19236 ( .A(b[415]), .B(n15138), .Z(n15139) );
  XOR U19237 ( .A(n15140), .B(n15141), .Z(n15138) );
  ANDN U19238 ( .B(n15142), .A(n656), .Z(n15140) );
  XNOR U19239 ( .A(b[414]), .B(n15141), .Z(n15142) );
  XOR U19240 ( .A(n15143), .B(n15144), .Z(n15141) );
  ANDN U19241 ( .B(n15145), .A(n657), .Z(n15143) );
  XNOR U19242 ( .A(b[413]), .B(n15144), .Z(n15145) );
  XOR U19243 ( .A(n15146), .B(n15147), .Z(n15144) );
  ANDN U19244 ( .B(n15148), .A(n658), .Z(n15146) );
  XNOR U19245 ( .A(b[412]), .B(n15147), .Z(n15148) );
  XOR U19246 ( .A(n15149), .B(n15150), .Z(n15147) );
  ANDN U19247 ( .B(n15151), .A(n659), .Z(n15149) );
  XNOR U19248 ( .A(b[411]), .B(n15150), .Z(n15151) );
  XOR U19249 ( .A(n15152), .B(n15153), .Z(n15150) );
  ANDN U19250 ( .B(n15154), .A(n660), .Z(n15152) );
  XNOR U19251 ( .A(b[410]), .B(n15153), .Z(n15154) );
  XOR U19252 ( .A(n15155), .B(n15156), .Z(n15153) );
  ANDN U19253 ( .B(n15157), .A(n662), .Z(n15155) );
  XNOR U19254 ( .A(b[409]), .B(n15156), .Z(n15157) );
  XOR U19255 ( .A(n15158), .B(n15159), .Z(n15156) );
  ANDN U19256 ( .B(n15160), .A(n687), .Z(n15158) );
  XNOR U19257 ( .A(b[408]), .B(n15159), .Z(n15160) );
  XOR U19258 ( .A(n15161), .B(n15162), .Z(n15159) );
  ANDN U19259 ( .B(n15163), .A(n728), .Z(n15161) );
  XNOR U19260 ( .A(b[407]), .B(n15162), .Z(n15163) );
  XOR U19261 ( .A(n15164), .B(n15165), .Z(n15162) );
  ANDN U19262 ( .B(n15166), .A(n769), .Z(n15164) );
  XNOR U19263 ( .A(b[406]), .B(n15165), .Z(n15166) );
  XOR U19264 ( .A(n15167), .B(n15168), .Z(n15165) );
  ANDN U19265 ( .B(n15169), .A(n810), .Z(n15167) );
  XNOR U19266 ( .A(b[405]), .B(n15168), .Z(n15169) );
  XOR U19267 ( .A(n15170), .B(n15171), .Z(n15168) );
  ANDN U19268 ( .B(n15172), .A(n851), .Z(n15170) );
  XNOR U19269 ( .A(b[404]), .B(n15171), .Z(n15172) );
  XOR U19270 ( .A(n15173), .B(n15174), .Z(n15171) );
  ANDN U19271 ( .B(n15175), .A(n892), .Z(n15173) );
  XNOR U19272 ( .A(b[403]), .B(n15174), .Z(n15175) );
  XOR U19273 ( .A(n15176), .B(n15177), .Z(n15174) );
  ANDN U19274 ( .B(n15178), .A(n933), .Z(n15176) );
  XNOR U19275 ( .A(b[402]), .B(n15177), .Z(n15178) );
  XOR U19276 ( .A(n15179), .B(n15180), .Z(n15177) );
  ANDN U19277 ( .B(n15181), .A(n974), .Z(n15179) );
  XNOR U19278 ( .A(b[401]), .B(n15180), .Z(n15181) );
  XOR U19279 ( .A(n15182), .B(n15183), .Z(n15180) );
  ANDN U19280 ( .B(n15184), .A(n1015), .Z(n15182) );
  XNOR U19281 ( .A(b[400]), .B(n15183), .Z(n15184) );
  XOR U19282 ( .A(n15185), .B(n15186), .Z(n15183) );
  ANDN U19283 ( .B(n15187), .A(n1058), .Z(n15185) );
  XNOR U19284 ( .A(b[399]), .B(n15186), .Z(n15187) );
  XOR U19285 ( .A(n15188), .B(n15189), .Z(n15186) );
  ANDN U19286 ( .B(n15190), .A(n1099), .Z(n15188) );
  XNOR U19287 ( .A(b[398]), .B(n15189), .Z(n15190) );
  XOR U19288 ( .A(n15191), .B(n15192), .Z(n15189) );
  ANDN U19289 ( .B(n15193), .A(n1140), .Z(n15191) );
  XNOR U19290 ( .A(b[397]), .B(n15192), .Z(n15193) );
  XOR U19291 ( .A(n15194), .B(n15195), .Z(n15192) );
  ANDN U19292 ( .B(n15196), .A(n1181), .Z(n15194) );
  XNOR U19293 ( .A(b[396]), .B(n15195), .Z(n15196) );
  XOR U19294 ( .A(n15197), .B(n15198), .Z(n15195) );
  ANDN U19295 ( .B(n15199), .A(n1222), .Z(n15197) );
  XNOR U19296 ( .A(b[395]), .B(n15198), .Z(n15199) );
  XOR U19297 ( .A(n15200), .B(n15201), .Z(n15198) );
  ANDN U19298 ( .B(n15202), .A(n1263), .Z(n15200) );
  XNOR U19299 ( .A(b[394]), .B(n15201), .Z(n15202) );
  XOR U19300 ( .A(n15203), .B(n15204), .Z(n15201) );
  ANDN U19301 ( .B(n15205), .A(n1304), .Z(n15203) );
  XNOR U19302 ( .A(b[393]), .B(n15204), .Z(n15205) );
  XOR U19303 ( .A(n15206), .B(n15207), .Z(n15204) );
  ANDN U19304 ( .B(n15208), .A(n1345), .Z(n15206) );
  XNOR U19305 ( .A(b[392]), .B(n15207), .Z(n15208) );
  XOR U19306 ( .A(n15209), .B(n15210), .Z(n15207) );
  ANDN U19307 ( .B(n15211), .A(n1386), .Z(n15209) );
  XNOR U19308 ( .A(b[391]), .B(n15210), .Z(n15211) );
  XOR U19309 ( .A(n15212), .B(n15213), .Z(n15210) );
  ANDN U19310 ( .B(n15214), .A(n1427), .Z(n15212) );
  XNOR U19311 ( .A(b[390]), .B(n15213), .Z(n15214) );
  XOR U19312 ( .A(n15215), .B(n15216), .Z(n15213) );
  ANDN U19313 ( .B(n15217), .A(n1469), .Z(n15215) );
  XNOR U19314 ( .A(b[389]), .B(n15216), .Z(n15217) );
  XOR U19315 ( .A(n15218), .B(n15219), .Z(n15216) );
  ANDN U19316 ( .B(n15220), .A(n1510), .Z(n15218) );
  XNOR U19317 ( .A(b[388]), .B(n15219), .Z(n15220) );
  XOR U19318 ( .A(n15221), .B(n15222), .Z(n15219) );
  ANDN U19319 ( .B(n15223), .A(n1551), .Z(n15221) );
  XNOR U19320 ( .A(b[387]), .B(n15222), .Z(n15223) );
  XOR U19321 ( .A(n15224), .B(n15225), .Z(n15222) );
  ANDN U19322 ( .B(n15226), .A(n1592), .Z(n15224) );
  XNOR U19323 ( .A(b[386]), .B(n15225), .Z(n15226) );
  XOR U19324 ( .A(n15227), .B(n15228), .Z(n15225) );
  ANDN U19325 ( .B(n15229), .A(n1633), .Z(n15227) );
  XNOR U19326 ( .A(b[385]), .B(n15228), .Z(n15229) );
  XOR U19327 ( .A(n15230), .B(n15231), .Z(n15228) );
  ANDN U19328 ( .B(n15232), .A(n1674), .Z(n15230) );
  XNOR U19329 ( .A(b[384]), .B(n15231), .Z(n15232) );
  XOR U19330 ( .A(n15233), .B(n15234), .Z(n15231) );
  ANDN U19331 ( .B(n15235), .A(n1715), .Z(n15233) );
  XNOR U19332 ( .A(b[383]), .B(n15234), .Z(n15235) );
  XOR U19333 ( .A(n15236), .B(n15237), .Z(n15234) );
  ANDN U19334 ( .B(n15238), .A(n1756), .Z(n15236) );
  XNOR U19335 ( .A(b[382]), .B(n15237), .Z(n15238) );
  XOR U19336 ( .A(n15239), .B(n15240), .Z(n15237) );
  ANDN U19337 ( .B(n15241), .A(n1797), .Z(n15239) );
  XNOR U19338 ( .A(b[381]), .B(n15240), .Z(n15241) );
  XOR U19339 ( .A(n15242), .B(n15243), .Z(n15240) );
  ANDN U19340 ( .B(n15244), .A(n1838), .Z(n15242) );
  XNOR U19341 ( .A(b[380]), .B(n15243), .Z(n15244) );
  XOR U19342 ( .A(n15245), .B(n15246), .Z(n15243) );
  ANDN U19343 ( .B(n15247), .A(n1880), .Z(n15245) );
  XNOR U19344 ( .A(b[379]), .B(n15246), .Z(n15247) );
  XOR U19345 ( .A(n15248), .B(n15249), .Z(n15246) );
  ANDN U19346 ( .B(n15250), .A(n1921), .Z(n15248) );
  XNOR U19347 ( .A(b[378]), .B(n15249), .Z(n15250) );
  XOR U19348 ( .A(n15251), .B(n15252), .Z(n15249) );
  ANDN U19349 ( .B(n15253), .A(n1962), .Z(n15251) );
  XNOR U19350 ( .A(b[377]), .B(n15252), .Z(n15253) );
  XOR U19351 ( .A(n15254), .B(n15255), .Z(n15252) );
  ANDN U19352 ( .B(n15256), .A(n2003), .Z(n15254) );
  XNOR U19353 ( .A(b[376]), .B(n15255), .Z(n15256) );
  XOR U19354 ( .A(n15257), .B(n15258), .Z(n15255) );
  ANDN U19355 ( .B(n15259), .A(n2044), .Z(n15257) );
  XNOR U19356 ( .A(b[375]), .B(n15258), .Z(n15259) );
  XOR U19357 ( .A(n15260), .B(n15261), .Z(n15258) );
  ANDN U19358 ( .B(n15262), .A(n2085), .Z(n15260) );
  XNOR U19359 ( .A(b[374]), .B(n15261), .Z(n15262) );
  XOR U19360 ( .A(n15263), .B(n15264), .Z(n15261) );
  ANDN U19361 ( .B(n15265), .A(n2126), .Z(n15263) );
  XNOR U19362 ( .A(b[373]), .B(n15264), .Z(n15265) );
  XOR U19363 ( .A(n15266), .B(n15267), .Z(n15264) );
  ANDN U19364 ( .B(n15268), .A(n2167), .Z(n15266) );
  XNOR U19365 ( .A(b[372]), .B(n15267), .Z(n15268) );
  XOR U19366 ( .A(n15269), .B(n15270), .Z(n15267) );
  ANDN U19367 ( .B(n15271), .A(n2208), .Z(n15269) );
  XNOR U19368 ( .A(b[371]), .B(n15270), .Z(n15271) );
  XOR U19369 ( .A(n15272), .B(n15273), .Z(n15270) );
  ANDN U19370 ( .B(n15274), .A(n2249), .Z(n15272) );
  XNOR U19371 ( .A(b[370]), .B(n15273), .Z(n15274) );
  XOR U19372 ( .A(n15275), .B(n15276), .Z(n15273) );
  ANDN U19373 ( .B(n15277), .A(n2291), .Z(n15275) );
  XNOR U19374 ( .A(b[369]), .B(n15276), .Z(n15277) );
  XOR U19375 ( .A(n15278), .B(n15279), .Z(n15276) );
  ANDN U19376 ( .B(n15280), .A(n2332), .Z(n15278) );
  XNOR U19377 ( .A(b[368]), .B(n15279), .Z(n15280) );
  XOR U19378 ( .A(n15281), .B(n15282), .Z(n15279) );
  ANDN U19379 ( .B(n15283), .A(n2373), .Z(n15281) );
  XNOR U19380 ( .A(b[367]), .B(n15282), .Z(n15283) );
  XOR U19381 ( .A(n15284), .B(n15285), .Z(n15282) );
  ANDN U19382 ( .B(n15286), .A(n2414), .Z(n15284) );
  XNOR U19383 ( .A(b[366]), .B(n15285), .Z(n15286) );
  XOR U19384 ( .A(n15287), .B(n15288), .Z(n15285) );
  ANDN U19385 ( .B(n15289), .A(n2455), .Z(n15287) );
  XNOR U19386 ( .A(b[365]), .B(n15288), .Z(n15289) );
  XOR U19387 ( .A(n15290), .B(n15291), .Z(n15288) );
  ANDN U19388 ( .B(n15292), .A(n2496), .Z(n15290) );
  XNOR U19389 ( .A(b[364]), .B(n15291), .Z(n15292) );
  XOR U19390 ( .A(n15293), .B(n15294), .Z(n15291) );
  ANDN U19391 ( .B(n15295), .A(n2537), .Z(n15293) );
  XNOR U19392 ( .A(b[363]), .B(n15294), .Z(n15295) );
  XOR U19393 ( .A(n15296), .B(n15297), .Z(n15294) );
  ANDN U19394 ( .B(n15298), .A(n2578), .Z(n15296) );
  XNOR U19395 ( .A(b[362]), .B(n15297), .Z(n15298) );
  XOR U19396 ( .A(n15299), .B(n15300), .Z(n15297) );
  ANDN U19397 ( .B(n15301), .A(n2619), .Z(n15299) );
  XNOR U19398 ( .A(b[361]), .B(n15300), .Z(n15301) );
  XOR U19399 ( .A(n15302), .B(n15303), .Z(n15300) );
  ANDN U19400 ( .B(n15304), .A(n2660), .Z(n15302) );
  XNOR U19401 ( .A(b[360]), .B(n15303), .Z(n15304) );
  XOR U19402 ( .A(n15305), .B(n15306), .Z(n15303) );
  ANDN U19403 ( .B(n15307), .A(n2702), .Z(n15305) );
  XNOR U19404 ( .A(b[359]), .B(n15306), .Z(n15307) );
  XOR U19405 ( .A(n15308), .B(n15309), .Z(n15306) );
  ANDN U19406 ( .B(n15310), .A(n2743), .Z(n15308) );
  XNOR U19407 ( .A(b[358]), .B(n15309), .Z(n15310) );
  XOR U19408 ( .A(n15311), .B(n15312), .Z(n15309) );
  ANDN U19409 ( .B(n15313), .A(n2784), .Z(n15311) );
  XNOR U19410 ( .A(b[357]), .B(n15312), .Z(n15313) );
  XOR U19411 ( .A(n15314), .B(n15315), .Z(n15312) );
  ANDN U19412 ( .B(n15316), .A(n2825), .Z(n15314) );
  XNOR U19413 ( .A(b[356]), .B(n15315), .Z(n15316) );
  XOR U19414 ( .A(n15317), .B(n15318), .Z(n15315) );
  ANDN U19415 ( .B(n15319), .A(n2866), .Z(n15317) );
  XNOR U19416 ( .A(b[355]), .B(n15318), .Z(n15319) );
  XOR U19417 ( .A(n15320), .B(n15321), .Z(n15318) );
  ANDN U19418 ( .B(n15322), .A(n2907), .Z(n15320) );
  XNOR U19419 ( .A(b[354]), .B(n15321), .Z(n15322) );
  XOR U19420 ( .A(n15323), .B(n15324), .Z(n15321) );
  ANDN U19421 ( .B(n15325), .A(n2948), .Z(n15323) );
  XNOR U19422 ( .A(b[353]), .B(n15324), .Z(n15325) );
  XOR U19423 ( .A(n15326), .B(n15327), .Z(n15324) );
  ANDN U19424 ( .B(n15328), .A(n2989), .Z(n15326) );
  XNOR U19425 ( .A(b[352]), .B(n15327), .Z(n15328) );
  XOR U19426 ( .A(n15329), .B(n15330), .Z(n15327) );
  ANDN U19427 ( .B(n15331), .A(n3030), .Z(n15329) );
  XNOR U19428 ( .A(b[351]), .B(n15330), .Z(n15331) );
  XOR U19429 ( .A(n15332), .B(n15333), .Z(n15330) );
  ANDN U19430 ( .B(n15334), .A(n3071), .Z(n15332) );
  XNOR U19431 ( .A(b[350]), .B(n15333), .Z(n15334) );
  XOR U19432 ( .A(n15335), .B(n15336), .Z(n15333) );
  ANDN U19433 ( .B(n15337), .A(n3113), .Z(n15335) );
  XNOR U19434 ( .A(b[349]), .B(n15336), .Z(n15337) );
  XOR U19435 ( .A(n15338), .B(n15339), .Z(n15336) );
  ANDN U19436 ( .B(n15340), .A(n3154), .Z(n15338) );
  XNOR U19437 ( .A(b[348]), .B(n15339), .Z(n15340) );
  XOR U19438 ( .A(n15341), .B(n15342), .Z(n15339) );
  ANDN U19439 ( .B(n15343), .A(n3195), .Z(n15341) );
  XNOR U19440 ( .A(b[347]), .B(n15342), .Z(n15343) );
  XOR U19441 ( .A(n15344), .B(n15345), .Z(n15342) );
  ANDN U19442 ( .B(n15346), .A(n3236), .Z(n15344) );
  XNOR U19443 ( .A(b[346]), .B(n15345), .Z(n15346) );
  XOR U19444 ( .A(n15347), .B(n15348), .Z(n15345) );
  ANDN U19445 ( .B(n15349), .A(n3277), .Z(n15347) );
  XNOR U19446 ( .A(b[345]), .B(n15348), .Z(n15349) );
  XOR U19447 ( .A(n15350), .B(n15351), .Z(n15348) );
  ANDN U19448 ( .B(n15352), .A(n3318), .Z(n15350) );
  XNOR U19449 ( .A(b[344]), .B(n15351), .Z(n15352) );
  XOR U19450 ( .A(n15353), .B(n15354), .Z(n15351) );
  ANDN U19451 ( .B(n15355), .A(n3359), .Z(n15353) );
  XNOR U19452 ( .A(b[343]), .B(n15354), .Z(n15355) );
  XOR U19453 ( .A(n15356), .B(n15357), .Z(n15354) );
  ANDN U19454 ( .B(n15358), .A(n3400), .Z(n15356) );
  XNOR U19455 ( .A(b[342]), .B(n15357), .Z(n15358) );
  XOR U19456 ( .A(n15359), .B(n15360), .Z(n15357) );
  ANDN U19457 ( .B(n15361), .A(n3441), .Z(n15359) );
  XNOR U19458 ( .A(b[341]), .B(n15360), .Z(n15361) );
  XOR U19459 ( .A(n15362), .B(n15363), .Z(n15360) );
  ANDN U19460 ( .B(n15364), .A(n3482), .Z(n15362) );
  XNOR U19461 ( .A(b[340]), .B(n15363), .Z(n15364) );
  XOR U19462 ( .A(n15365), .B(n15366), .Z(n15363) );
  ANDN U19463 ( .B(n15367), .A(n3524), .Z(n15365) );
  XNOR U19464 ( .A(b[339]), .B(n15366), .Z(n15367) );
  XOR U19465 ( .A(n15368), .B(n15369), .Z(n15366) );
  ANDN U19466 ( .B(n15370), .A(n3565), .Z(n15368) );
  XNOR U19467 ( .A(b[338]), .B(n15369), .Z(n15370) );
  XOR U19468 ( .A(n15371), .B(n15372), .Z(n15369) );
  ANDN U19469 ( .B(n15373), .A(n3606), .Z(n15371) );
  XNOR U19470 ( .A(b[337]), .B(n15372), .Z(n15373) );
  XOR U19471 ( .A(n15374), .B(n15375), .Z(n15372) );
  ANDN U19472 ( .B(n15376), .A(n3647), .Z(n15374) );
  XNOR U19473 ( .A(b[336]), .B(n15375), .Z(n15376) );
  XOR U19474 ( .A(n15377), .B(n15378), .Z(n15375) );
  ANDN U19475 ( .B(n15379), .A(n3688), .Z(n15377) );
  XNOR U19476 ( .A(b[335]), .B(n15378), .Z(n15379) );
  XOR U19477 ( .A(n15380), .B(n15381), .Z(n15378) );
  ANDN U19478 ( .B(n15382), .A(n3729), .Z(n15380) );
  XNOR U19479 ( .A(b[334]), .B(n15381), .Z(n15382) );
  XOR U19480 ( .A(n15383), .B(n15384), .Z(n15381) );
  ANDN U19481 ( .B(n15385), .A(n3770), .Z(n15383) );
  XNOR U19482 ( .A(b[333]), .B(n15384), .Z(n15385) );
  XOR U19483 ( .A(n15386), .B(n15387), .Z(n15384) );
  ANDN U19484 ( .B(n15388), .A(n3811), .Z(n15386) );
  XNOR U19485 ( .A(b[332]), .B(n15387), .Z(n15388) );
  XOR U19486 ( .A(n15389), .B(n15390), .Z(n15387) );
  ANDN U19487 ( .B(n15391), .A(n3852), .Z(n15389) );
  XNOR U19488 ( .A(b[331]), .B(n15390), .Z(n15391) );
  XOR U19489 ( .A(n15392), .B(n15393), .Z(n15390) );
  ANDN U19490 ( .B(n15394), .A(n3893), .Z(n15392) );
  XNOR U19491 ( .A(b[330]), .B(n15393), .Z(n15394) );
  XOR U19492 ( .A(n15395), .B(n15396), .Z(n15393) );
  ANDN U19493 ( .B(n15397), .A(n3935), .Z(n15395) );
  XNOR U19494 ( .A(b[329]), .B(n15396), .Z(n15397) );
  XOR U19495 ( .A(n15398), .B(n15399), .Z(n15396) );
  ANDN U19496 ( .B(n15400), .A(n3976), .Z(n15398) );
  XNOR U19497 ( .A(b[328]), .B(n15399), .Z(n15400) );
  XOR U19498 ( .A(n15401), .B(n15402), .Z(n15399) );
  ANDN U19499 ( .B(n15403), .A(n4017), .Z(n15401) );
  XNOR U19500 ( .A(b[327]), .B(n15402), .Z(n15403) );
  XOR U19501 ( .A(n15404), .B(n15405), .Z(n15402) );
  ANDN U19502 ( .B(n15406), .A(n4058), .Z(n15404) );
  XNOR U19503 ( .A(b[326]), .B(n15405), .Z(n15406) );
  XOR U19504 ( .A(n15407), .B(n15408), .Z(n15405) );
  ANDN U19505 ( .B(n15409), .A(n4099), .Z(n15407) );
  XNOR U19506 ( .A(b[325]), .B(n15408), .Z(n15409) );
  XOR U19507 ( .A(n15410), .B(n15411), .Z(n15408) );
  ANDN U19508 ( .B(n15412), .A(n4140), .Z(n15410) );
  XNOR U19509 ( .A(b[324]), .B(n15411), .Z(n15412) );
  XOR U19510 ( .A(n15413), .B(n15414), .Z(n15411) );
  ANDN U19511 ( .B(n15415), .A(n4181), .Z(n15413) );
  XNOR U19512 ( .A(b[323]), .B(n15414), .Z(n15415) );
  XOR U19513 ( .A(n15416), .B(n15417), .Z(n15414) );
  ANDN U19514 ( .B(n15418), .A(n4222), .Z(n15416) );
  XNOR U19515 ( .A(b[322]), .B(n15417), .Z(n15418) );
  XOR U19516 ( .A(n15419), .B(n15420), .Z(n15417) );
  ANDN U19517 ( .B(n15421), .A(n4263), .Z(n15419) );
  XNOR U19518 ( .A(b[321]), .B(n15420), .Z(n15421) );
  XOR U19519 ( .A(n15422), .B(n15423), .Z(n15420) );
  ANDN U19520 ( .B(n15424), .A(n4304), .Z(n15422) );
  XNOR U19521 ( .A(b[320]), .B(n15423), .Z(n15424) );
  XOR U19522 ( .A(n15425), .B(n15426), .Z(n15423) );
  ANDN U19523 ( .B(n15427), .A(n4346), .Z(n15425) );
  XNOR U19524 ( .A(b[319]), .B(n15426), .Z(n15427) );
  XOR U19525 ( .A(n15428), .B(n15429), .Z(n15426) );
  ANDN U19526 ( .B(n15430), .A(n4387), .Z(n15428) );
  XNOR U19527 ( .A(b[318]), .B(n15429), .Z(n15430) );
  XOR U19528 ( .A(n15431), .B(n15432), .Z(n15429) );
  ANDN U19529 ( .B(n15433), .A(n4428), .Z(n15431) );
  XNOR U19530 ( .A(b[317]), .B(n15432), .Z(n15433) );
  XOR U19531 ( .A(n15434), .B(n15435), .Z(n15432) );
  ANDN U19532 ( .B(n15436), .A(n4469), .Z(n15434) );
  XNOR U19533 ( .A(b[316]), .B(n15435), .Z(n15436) );
  XOR U19534 ( .A(n15437), .B(n15438), .Z(n15435) );
  ANDN U19535 ( .B(n15439), .A(n4510), .Z(n15437) );
  XNOR U19536 ( .A(b[315]), .B(n15438), .Z(n15439) );
  XOR U19537 ( .A(n15440), .B(n15441), .Z(n15438) );
  ANDN U19538 ( .B(n15442), .A(n4551), .Z(n15440) );
  XNOR U19539 ( .A(b[314]), .B(n15441), .Z(n15442) );
  XOR U19540 ( .A(n15443), .B(n15444), .Z(n15441) );
  ANDN U19541 ( .B(n15445), .A(n4592), .Z(n15443) );
  XNOR U19542 ( .A(b[313]), .B(n15444), .Z(n15445) );
  XOR U19543 ( .A(n15446), .B(n15447), .Z(n15444) );
  ANDN U19544 ( .B(n15448), .A(n4633), .Z(n15446) );
  XNOR U19545 ( .A(b[312]), .B(n15447), .Z(n15448) );
  XOR U19546 ( .A(n15449), .B(n15450), .Z(n15447) );
  ANDN U19547 ( .B(n15451), .A(n4674), .Z(n15449) );
  XNOR U19548 ( .A(b[311]), .B(n15450), .Z(n15451) );
  XOR U19549 ( .A(n15452), .B(n15453), .Z(n15450) );
  ANDN U19550 ( .B(n15454), .A(n4715), .Z(n15452) );
  XNOR U19551 ( .A(b[310]), .B(n15453), .Z(n15454) );
  XOR U19552 ( .A(n15455), .B(n15456), .Z(n15453) );
  ANDN U19553 ( .B(n15457), .A(n4757), .Z(n15455) );
  XNOR U19554 ( .A(b[309]), .B(n15456), .Z(n15457) );
  XOR U19555 ( .A(n15458), .B(n15459), .Z(n15456) );
  ANDN U19556 ( .B(n15460), .A(n4798), .Z(n15458) );
  XNOR U19557 ( .A(b[308]), .B(n15459), .Z(n15460) );
  XOR U19558 ( .A(n15461), .B(n15462), .Z(n15459) );
  ANDN U19559 ( .B(n15463), .A(n4839), .Z(n15461) );
  XNOR U19560 ( .A(b[307]), .B(n15462), .Z(n15463) );
  XOR U19561 ( .A(n15464), .B(n15465), .Z(n15462) );
  ANDN U19562 ( .B(n15466), .A(n4880), .Z(n15464) );
  XNOR U19563 ( .A(b[306]), .B(n15465), .Z(n15466) );
  XOR U19564 ( .A(n15467), .B(n15468), .Z(n15465) );
  ANDN U19565 ( .B(n15469), .A(n4921), .Z(n15467) );
  XNOR U19566 ( .A(b[305]), .B(n15468), .Z(n15469) );
  XOR U19567 ( .A(n15470), .B(n15471), .Z(n15468) );
  ANDN U19568 ( .B(n15472), .A(n4962), .Z(n15470) );
  XNOR U19569 ( .A(b[304]), .B(n15471), .Z(n15472) );
  XOR U19570 ( .A(n15473), .B(n15474), .Z(n15471) );
  ANDN U19571 ( .B(n15475), .A(n5003), .Z(n15473) );
  XNOR U19572 ( .A(b[303]), .B(n15474), .Z(n15475) );
  XOR U19573 ( .A(n15476), .B(n15477), .Z(n15474) );
  ANDN U19574 ( .B(n15478), .A(n5044), .Z(n15476) );
  XNOR U19575 ( .A(b[302]), .B(n15477), .Z(n15478) );
  XOR U19576 ( .A(n15479), .B(n15480), .Z(n15477) );
  ANDN U19577 ( .B(n15481), .A(n5085), .Z(n15479) );
  XNOR U19578 ( .A(b[301]), .B(n15480), .Z(n15481) );
  XOR U19579 ( .A(n15482), .B(n15483), .Z(n15480) );
  ANDN U19580 ( .B(n15484), .A(n5126), .Z(n15482) );
  XNOR U19581 ( .A(b[300]), .B(n15483), .Z(n15484) );
  XOR U19582 ( .A(n15485), .B(n15486), .Z(n15483) );
  ANDN U19583 ( .B(n15487), .A(n5169), .Z(n15485) );
  XNOR U19584 ( .A(b[299]), .B(n15486), .Z(n15487) );
  XOR U19585 ( .A(n15488), .B(n15489), .Z(n15486) );
  ANDN U19586 ( .B(n15490), .A(n5210), .Z(n15488) );
  XNOR U19587 ( .A(b[298]), .B(n15489), .Z(n15490) );
  XOR U19588 ( .A(n15491), .B(n15492), .Z(n15489) );
  ANDN U19589 ( .B(n15493), .A(n5251), .Z(n15491) );
  XNOR U19590 ( .A(b[297]), .B(n15492), .Z(n15493) );
  XOR U19591 ( .A(n15494), .B(n15495), .Z(n15492) );
  ANDN U19592 ( .B(n15496), .A(n5292), .Z(n15494) );
  XNOR U19593 ( .A(b[296]), .B(n15495), .Z(n15496) );
  XOR U19594 ( .A(n15497), .B(n15498), .Z(n15495) );
  ANDN U19595 ( .B(n15499), .A(n5333), .Z(n15497) );
  XNOR U19596 ( .A(b[295]), .B(n15498), .Z(n15499) );
  XOR U19597 ( .A(n15500), .B(n15501), .Z(n15498) );
  ANDN U19598 ( .B(n15502), .A(n5374), .Z(n15500) );
  XNOR U19599 ( .A(b[294]), .B(n15501), .Z(n15502) );
  XOR U19600 ( .A(n15503), .B(n15504), .Z(n15501) );
  ANDN U19601 ( .B(n15505), .A(n5415), .Z(n15503) );
  XNOR U19602 ( .A(b[293]), .B(n15504), .Z(n15505) );
  XOR U19603 ( .A(n15506), .B(n15507), .Z(n15504) );
  ANDN U19604 ( .B(n15508), .A(n5456), .Z(n15506) );
  XNOR U19605 ( .A(b[292]), .B(n15507), .Z(n15508) );
  XOR U19606 ( .A(n15509), .B(n15510), .Z(n15507) );
  ANDN U19607 ( .B(n15511), .A(n5497), .Z(n15509) );
  XNOR U19608 ( .A(b[291]), .B(n15510), .Z(n15511) );
  XOR U19609 ( .A(n15512), .B(n15513), .Z(n15510) );
  ANDN U19610 ( .B(n15514), .A(n5538), .Z(n15512) );
  XNOR U19611 ( .A(b[290]), .B(n15513), .Z(n15514) );
  XOR U19612 ( .A(n15515), .B(n15516), .Z(n15513) );
  ANDN U19613 ( .B(n15517), .A(n5580), .Z(n15515) );
  XNOR U19614 ( .A(b[289]), .B(n15516), .Z(n15517) );
  XOR U19615 ( .A(n15518), .B(n15519), .Z(n15516) );
  ANDN U19616 ( .B(n15520), .A(n5621), .Z(n15518) );
  XNOR U19617 ( .A(b[288]), .B(n15519), .Z(n15520) );
  XOR U19618 ( .A(n15521), .B(n15522), .Z(n15519) );
  ANDN U19619 ( .B(n15523), .A(n5662), .Z(n15521) );
  XNOR U19620 ( .A(b[287]), .B(n15522), .Z(n15523) );
  XOR U19621 ( .A(n15524), .B(n15525), .Z(n15522) );
  ANDN U19622 ( .B(n15526), .A(n5703), .Z(n15524) );
  XNOR U19623 ( .A(b[286]), .B(n15525), .Z(n15526) );
  XOR U19624 ( .A(n15527), .B(n15528), .Z(n15525) );
  ANDN U19625 ( .B(n15529), .A(n5744), .Z(n15527) );
  XNOR U19626 ( .A(b[285]), .B(n15528), .Z(n15529) );
  XOR U19627 ( .A(n15530), .B(n15531), .Z(n15528) );
  ANDN U19628 ( .B(n15532), .A(n5785), .Z(n15530) );
  XNOR U19629 ( .A(b[284]), .B(n15531), .Z(n15532) );
  XOR U19630 ( .A(n15533), .B(n15534), .Z(n15531) );
  ANDN U19631 ( .B(n15535), .A(n5826), .Z(n15533) );
  XNOR U19632 ( .A(b[283]), .B(n15534), .Z(n15535) );
  XOR U19633 ( .A(n15536), .B(n15537), .Z(n15534) );
  ANDN U19634 ( .B(n15538), .A(n5867), .Z(n15536) );
  XNOR U19635 ( .A(b[282]), .B(n15537), .Z(n15538) );
  XOR U19636 ( .A(n15539), .B(n15540), .Z(n15537) );
  ANDN U19637 ( .B(n15541), .A(n5908), .Z(n15539) );
  XNOR U19638 ( .A(b[281]), .B(n15540), .Z(n15541) );
  XOR U19639 ( .A(n15542), .B(n15543), .Z(n15540) );
  ANDN U19640 ( .B(n15544), .A(n5949), .Z(n15542) );
  XNOR U19641 ( .A(b[280]), .B(n15543), .Z(n15544) );
  XOR U19642 ( .A(n15545), .B(n15546), .Z(n15543) );
  ANDN U19643 ( .B(n15547), .A(n5991), .Z(n15545) );
  XNOR U19644 ( .A(b[279]), .B(n15546), .Z(n15547) );
  XOR U19645 ( .A(n15548), .B(n15549), .Z(n15546) );
  ANDN U19646 ( .B(n15550), .A(n6032), .Z(n15548) );
  XNOR U19647 ( .A(b[278]), .B(n15549), .Z(n15550) );
  XOR U19648 ( .A(n15551), .B(n15552), .Z(n15549) );
  ANDN U19649 ( .B(n15553), .A(n6073), .Z(n15551) );
  XNOR U19650 ( .A(b[277]), .B(n15552), .Z(n15553) );
  XOR U19651 ( .A(n15554), .B(n15555), .Z(n15552) );
  ANDN U19652 ( .B(n15556), .A(n6114), .Z(n15554) );
  XNOR U19653 ( .A(b[276]), .B(n15555), .Z(n15556) );
  XOR U19654 ( .A(n15557), .B(n15558), .Z(n15555) );
  ANDN U19655 ( .B(n15559), .A(n6155), .Z(n15557) );
  XNOR U19656 ( .A(b[275]), .B(n15558), .Z(n15559) );
  XOR U19657 ( .A(n15560), .B(n15561), .Z(n15558) );
  ANDN U19658 ( .B(n15562), .A(n6196), .Z(n15560) );
  XNOR U19659 ( .A(b[274]), .B(n15561), .Z(n15562) );
  XOR U19660 ( .A(n15563), .B(n15564), .Z(n15561) );
  ANDN U19661 ( .B(n15565), .A(n6237), .Z(n15563) );
  XNOR U19662 ( .A(b[273]), .B(n15564), .Z(n15565) );
  XOR U19663 ( .A(n15566), .B(n15567), .Z(n15564) );
  ANDN U19664 ( .B(n15568), .A(n6278), .Z(n15566) );
  XNOR U19665 ( .A(b[272]), .B(n15567), .Z(n15568) );
  XOR U19666 ( .A(n15569), .B(n15570), .Z(n15567) );
  ANDN U19667 ( .B(n15571), .A(n6319), .Z(n15569) );
  XNOR U19668 ( .A(b[271]), .B(n15570), .Z(n15571) );
  XOR U19669 ( .A(n15572), .B(n15573), .Z(n15570) );
  ANDN U19670 ( .B(n15574), .A(n6360), .Z(n15572) );
  XNOR U19671 ( .A(b[270]), .B(n15573), .Z(n15574) );
  XOR U19672 ( .A(n15575), .B(n15576), .Z(n15573) );
  ANDN U19673 ( .B(n15577), .A(n6402), .Z(n15575) );
  XNOR U19674 ( .A(b[269]), .B(n15576), .Z(n15577) );
  XOR U19675 ( .A(n15578), .B(n15579), .Z(n15576) );
  ANDN U19676 ( .B(n15580), .A(n6443), .Z(n15578) );
  XNOR U19677 ( .A(b[268]), .B(n15579), .Z(n15580) );
  XOR U19678 ( .A(n15581), .B(n15582), .Z(n15579) );
  ANDN U19679 ( .B(n15583), .A(n6484), .Z(n15581) );
  XNOR U19680 ( .A(b[267]), .B(n15582), .Z(n15583) );
  XOR U19681 ( .A(n15584), .B(n15585), .Z(n15582) );
  ANDN U19682 ( .B(n15586), .A(n6525), .Z(n15584) );
  XNOR U19683 ( .A(b[266]), .B(n15585), .Z(n15586) );
  XOR U19684 ( .A(n15587), .B(n15588), .Z(n15585) );
  ANDN U19685 ( .B(n15589), .A(n6566), .Z(n15587) );
  XNOR U19686 ( .A(b[265]), .B(n15588), .Z(n15589) );
  XOR U19687 ( .A(n15590), .B(n15591), .Z(n15588) );
  ANDN U19688 ( .B(n15592), .A(n6607), .Z(n15590) );
  XNOR U19689 ( .A(b[264]), .B(n15591), .Z(n15592) );
  XOR U19690 ( .A(n15593), .B(n15594), .Z(n15591) );
  ANDN U19691 ( .B(n15595), .A(n6648), .Z(n15593) );
  XNOR U19692 ( .A(b[263]), .B(n15594), .Z(n15595) );
  XOR U19693 ( .A(n15596), .B(n15597), .Z(n15594) );
  ANDN U19694 ( .B(n15598), .A(n6689), .Z(n15596) );
  XNOR U19695 ( .A(b[262]), .B(n15597), .Z(n15598) );
  XOR U19696 ( .A(n15599), .B(n15600), .Z(n15597) );
  ANDN U19697 ( .B(n15601), .A(n6730), .Z(n15599) );
  XNOR U19698 ( .A(b[261]), .B(n15600), .Z(n15601) );
  XOR U19699 ( .A(n15602), .B(n15603), .Z(n15600) );
  ANDN U19700 ( .B(n15604), .A(n6771), .Z(n15602) );
  XNOR U19701 ( .A(b[260]), .B(n15603), .Z(n15604) );
  XOR U19702 ( .A(n15605), .B(n15606), .Z(n15603) );
  ANDN U19703 ( .B(n15607), .A(n6813), .Z(n15605) );
  XNOR U19704 ( .A(b[259]), .B(n15606), .Z(n15607) );
  XOR U19705 ( .A(n15608), .B(n15609), .Z(n15606) );
  ANDN U19706 ( .B(n15610), .A(n6854), .Z(n15608) );
  XNOR U19707 ( .A(b[258]), .B(n15609), .Z(n15610) );
  XOR U19708 ( .A(n15611), .B(n15612), .Z(n15609) );
  ANDN U19709 ( .B(n15613), .A(n6895), .Z(n15611) );
  XNOR U19710 ( .A(b[257]), .B(n15612), .Z(n15613) );
  XOR U19711 ( .A(n15614), .B(n15615), .Z(n15612) );
  ANDN U19712 ( .B(n15616), .A(n6936), .Z(n15614) );
  XNOR U19713 ( .A(b[256]), .B(n15615), .Z(n15616) );
  XOR U19714 ( .A(n15617), .B(n15618), .Z(n15615) );
  ANDN U19715 ( .B(n15619), .A(n6977), .Z(n15617) );
  XNOR U19716 ( .A(b[255]), .B(n15618), .Z(n15619) );
  XOR U19717 ( .A(n15620), .B(n15621), .Z(n15618) );
  ANDN U19718 ( .B(n15622), .A(n7018), .Z(n15620) );
  XNOR U19719 ( .A(b[254]), .B(n15621), .Z(n15622) );
  XOR U19720 ( .A(n15623), .B(n15624), .Z(n15621) );
  ANDN U19721 ( .B(n15625), .A(n7059), .Z(n15623) );
  XNOR U19722 ( .A(b[253]), .B(n15624), .Z(n15625) );
  XOR U19723 ( .A(n15626), .B(n15627), .Z(n15624) );
  ANDN U19724 ( .B(n15628), .A(n7100), .Z(n15626) );
  XNOR U19725 ( .A(b[252]), .B(n15627), .Z(n15628) );
  XOR U19726 ( .A(n15629), .B(n15630), .Z(n15627) );
  ANDN U19727 ( .B(n15631), .A(n7141), .Z(n15629) );
  XNOR U19728 ( .A(b[251]), .B(n15630), .Z(n15631) );
  XOR U19729 ( .A(n15632), .B(n15633), .Z(n15630) );
  ANDN U19730 ( .B(n15634), .A(n7182), .Z(n15632) );
  XNOR U19731 ( .A(b[250]), .B(n15633), .Z(n15634) );
  XOR U19732 ( .A(n15635), .B(n15636), .Z(n15633) );
  ANDN U19733 ( .B(n15637), .A(n7224), .Z(n15635) );
  XNOR U19734 ( .A(b[249]), .B(n15636), .Z(n15637) );
  XOR U19735 ( .A(n15638), .B(n15639), .Z(n15636) );
  ANDN U19736 ( .B(n15640), .A(n7265), .Z(n15638) );
  XNOR U19737 ( .A(b[248]), .B(n15639), .Z(n15640) );
  XOR U19738 ( .A(n15641), .B(n15642), .Z(n15639) );
  ANDN U19739 ( .B(n15643), .A(n7306), .Z(n15641) );
  XNOR U19740 ( .A(b[247]), .B(n15642), .Z(n15643) );
  XOR U19741 ( .A(n15644), .B(n15645), .Z(n15642) );
  ANDN U19742 ( .B(n15646), .A(n7347), .Z(n15644) );
  XNOR U19743 ( .A(b[246]), .B(n15645), .Z(n15646) );
  XOR U19744 ( .A(n15647), .B(n15648), .Z(n15645) );
  ANDN U19745 ( .B(n15649), .A(n7388), .Z(n15647) );
  XNOR U19746 ( .A(b[245]), .B(n15648), .Z(n15649) );
  XOR U19747 ( .A(n15650), .B(n15651), .Z(n15648) );
  ANDN U19748 ( .B(n15652), .A(n7429), .Z(n15650) );
  XNOR U19749 ( .A(b[244]), .B(n15651), .Z(n15652) );
  XOR U19750 ( .A(n15653), .B(n15654), .Z(n15651) );
  ANDN U19751 ( .B(n15655), .A(n7470), .Z(n15653) );
  XNOR U19752 ( .A(b[243]), .B(n15654), .Z(n15655) );
  XOR U19753 ( .A(n15656), .B(n15657), .Z(n15654) );
  ANDN U19754 ( .B(n15658), .A(n7511), .Z(n15656) );
  XNOR U19755 ( .A(b[242]), .B(n15657), .Z(n15658) );
  XOR U19756 ( .A(n15659), .B(n15660), .Z(n15657) );
  ANDN U19757 ( .B(n15661), .A(n7552), .Z(n15659) );
  XNOR U19758 ( .A(b[241]), .B(n15660), .Z(n15661) );
  XOR U19759 ( .A(n15662), .B(n15663), .Z(n15660) );
  ANDN U19760 ( .B(n15664), .A(n7593), .Z(n15662) );
  XNOR U19761 ( .A(b[240]), .B(n15663), .Z(n15664) );
  XOR U19762 ( .A(n15665), .B(n15666), .Z(n15663) );
  ANDN U19763 ( .B(n15667), .A(n7635), .Z(n15665) );
  XNOR U19764 ( .A(b[239]), .B(n15666), .Z(n15667) );
  XOR U19765 ( .A(n15668), .B(n15669), .Z(n15666) );
  ANDN U19766 ( .B(n15670), .A(n7676), .Z(n15668) );
  XNOR U19767 ( .A(b[238]), .B(n15669), .Z(n15670) );
  XOR U19768 ( .A(n15671), .B(n15672), .Z(n15669) );
  ANDN U19769 ( .B(n15673), .A(n7717), .Z(n15671) );
  XNOR U19770 ( .A(b[237]), .B(n15672), .Z(n15673) );
  XOR U19771 ( .A(n15674), .B(n15675), .Z(n15672) );
  ANDN U19772 ( .B(n15676), .A(n7758), .Z(n15674) );
  XNOR U19773 ( .A(b[236]), .B(n15675), .Z(n15676) );
  XOR U19774 ( .A(n15677), .B(n15678), .Z(n15675) );
  ANDN U19775 ( .B(n15679), .A(n7799), .Z(n15677) );
  XNOR U19776 ( .A(b[235]), .B(n15678), .Z(n15679) );
  XOR U19777 ( .A(n15680), .B(n15681), .Z(n15678) );
  ANDN U19778 ( .B(n15682), .A(n7840), .Z(n15680) );
  XNOR U19779 ( .A(b[234]), .B(n15681), .Z(n15682) );
  XOR U19780 ( .A(n15683), .B(n15684), .Z(n15681) );
  ANDN U19781 ( .B(n15685), .A(n7881), .Z(n15683) );
  XNOR U19782 ( .A(b[233]), .B(n15684), .Z(n15685) );
  XOR U19783 ( .A(n15686), .B(n15687), .Z(n15684) );
  ANDN U19784 ( .B(n15688), .A(n7922), .Z(n15686) );
  XNOR U19785 ( .A(b[232]), .B(n15687), .Z(n15688) );
  XOR U19786 ( .A(n15689), .B(n15690), .Z(n15687) );
  ANDN U19787 ( .B(n15691), .A(n7963), .Z(n15689) );
  XNOR U19788 ( .A(b[231]), .B(n15690), .Z(n15691) );
  XOR U19789 ( .A(n15692), .B(n15693), .Z(n15690) );
  ANDN U19790 ( .B(n15694), .A(n8004), .Z(n15692) );
  XNOR U19791 ( .A(b[230]), .B(n15693), .Z(n15694) );
  XOR U19792 ( .A(n15695), .B(n15696), .Z(n15693) );
  ANDN U19793 ( .B(n15697), .A(n8046), .Z(n15695) );
  XNOR U19794 ( .A(b[229]), .B(n15696), .Z(n15697) );
  XOR U19795 ( .A(n15698), .B(n15699), .Z(n15696) );
  ANDN U19796 ( .B(n15700), .A(n8087), .Z(n15698) );
  XNOR U19797 ( .A(b[228]), .B(n15699), .Z(n15700) );
  XOR U19798 ( .A(n15701), .B(n15702), .Z(n15699) );
  ANDN U19799 ( .B(n15703), .A(n8128), .Z(n15701) );
  XNOR U19800 ( .A(b[227]), .B(n15702), .Z(n15703) );
  XOR U19801 ( .A(n15704), .B(n15705), .Z(n15702) );
  ANDN U19802 ( .B(n15706), .A(n8169), .Z(n15704) );
  XNOR U19803 ( .A(b[226]), .B(n15705), .Z(n15706) );
  XOR U19804 ( .A(n15707), .B(n15708), .Z(n15705) );
  ANDN U19805 ( .B(n15709), .A(n8210), .Z(n15707) );
  XNOR U19806 ( .A(b[225]), .B(n15708), .Z(n15709) );
  XOR U19807 ( .A(n15710), .B(n15711), .Z(n15708) );
  ANDN U19808 ( .B(n15712), .A(n8251), .Z(n15710) );
  XNOR U19809 ( .A(b[224]), .B(n15711), .Z(n15712) );
  XOR U19810 ( .A(n15713), .B(n15714), .Z(n15711) );
  ANDN U19811 ( .B(n15715), .A(n8292), .Z(n15713) );
  XNOR U19812 ( .A(b[223]), .B(n15714), .Z(n15715) );
  XOR U19813 ( .A(n15716), .B(n15717), .Z(n15714) );
  ANDN U19814 ( .B(n15718), .A(n8333), .Z(n15716) );
  XNOR U19815 ( .A(b[222]), .B(n15717), .Z(n15718) );
  XOR U19816 ( .A(n15719), .B(n15720), .Z(n15717) );
  ANDN U19817 ( .B(n15721), .A(n8374), .Z(n15719) );
  XNOR U19818 ( .A(b[221]), .B(n15720), .Z(n15721) );
  XOR U19819 ( .A(n15722), .B(n15723), .Z(n15720) );
  ANDN U19820 ( .B(n15724), .A(n8415), .Z(n15722) );
  XNOR U19821 ( .A(b[220]), .B(n15723), .Z(n15724) );
  XOR U19822 ( .A(n15725), .B(n15726), .Z(n15723) );
  ANDN U19823 ( .B(n15727), .A(n8457), .Z(n15725) );
  XNOR U19824 ( .A(b[219]), .B(n15726), .Z(n15727) );
  XOR U19825 ( .A(n15728), .B(n15729), .Z(n15726) );
  ANDN U19826 ( .B(n15730), .A(n8498), .Z(n15728) );
  XNOR U19827 ( .A(b[218]), .B(n15729), .Z(n15730) );
  XOR U19828 ( .A(n15731), .B(n15732), .Z(n15729) );
  ANDN U19829 ( .B(n15733), .A(n8539), .Z(n15731) );
  XNOR U19830 ( .A(b[217]), .B(n15732), .Z(n15733) );
  XOR U19831 ( .A(n15734), .B(n15735), .Z(n15732) );
  ANDN U19832 ( .B(n15736), .A(n8580), .Z(n15734) );
  XNOR U19833 ( .A(b[216]), .B(n15735), .Z(n15736) );
  XOR U19834 ( .A(n15737), .B(n15738), .Z(n15735) );
  ANDN U19835 ( .B(n15739), .A(n8621), .Z(n15737) );
  XNOR U19836 ( .A(b[215]), .B(n15738), .Z(n15739) );
  XOR U19837 ( .A(n15740), .B(n15741), .Z(n15738) );
  ANDN U19838 ( .B(n15742), .A(n8662), .Z(n15740) );
  XNOR U19839 ( .A(b[214]), .B(n15741), .Z(n15742) );
  XOR U19840 ( .A(n15743), .B(n15744), .Z(n15741) );
  ANDN U19841 ( .B(n15745), .A(n8703), .Z(n15743) );
  XNOR U19842 ( .A(b[213]), .B(n15744), .Z(n15745) );
  XOR U19843 ( .A(n15746), .B(n15747), .Z(n15744) );
  ANDN U19844 ( .B(n15748), .A(n8744), .Z(n15746) );
  XNOR U19845 ( .A(b[212]), .B(n15747), .Z(n15748) );
  XOR U19846 ( .A(n15749), .B(n15750), .Z(n15747) );
  ANDN U19847 ( .B(n15751), .A(n8785), .Z(n15749) );
  XNOR U19848 ( .A(b[211]), .B(n15750), .Z(n15751) );
  XOR U19849 ( .A(n15752), .B(n15753), .Z(n15750) );
  ANDN U19850 ( .B(n15754), .A(n8826), .Z(n15752) );
  XNOR U19851 ( .A(b[210]), .B(n15753), .Z(n15754) );
  XOR U19852 ( .A(n15755), .B(n15756), .Z(n15753) );
  ANDN U19853 ( .B(n15757), .A(n8868), .Z(n15755) );
  XNOR U19854 ( .A(b[209]), .B(n15756), .Z(n15757) );
  XOR U19855 ( .A(n15758), .B(n15759), .Z(n15756) );
  ANDN U19856 ( .B(n15760), .A(n8909), .Z(n15758) );
  XNOR U19857 ( .A(b[208]), .B(n15759), .Z(n15760) );
  XOR U19858 ( .A(n15761), .B(n15762), .Z(n15759) );
  ANDN U19859 ( .B(n15763), .A(n8950), .Z(n15761) );
  XNOR U19860 ( .A(b[207]), .B(n15762), .Z(n15763) );
  XOR U19861 ( .A(n15764), .B(n15765), .Z(n15762) );
  ANDN U19862 ( .B(n15766), .A(n8991), .Z(n15764) );
  XNOR U19863 ( .A(b[206]), .B(n15765), .Z(n15766) );
  XOR U19864 ( .A(n15767), .B(n15768), .Z(n15765) );
  ANDN U19865 ( .B(n15769), .A(n9032), .Z(n15767) );
  XNOR U19866 ( .A(b[205]), .B(n15768), .Z(n15769) );
  XOR U19867 ( .A(n15770), .B(n15771), .Z(n15768) );
  ANDN U19868 ( .B(n15772), .A(n9073), .Z(n15770) );
  XNOR U19869 ( .A(b[204]), .B(n15771), .Z(n15772) );
  XOR U19870 ( .A(n15773), .B(n15774), .Z(n15771) );
  ANDN U19871 ( .B(n15775), .A(n9114), .Z(n15773) );
  XNOR U19872 ( .A(b[203]), .B(n15774), .Z(n15775) );
  XOR U19873 ( .A(n15776), .B(n15777), .Z(n15774) );
  ANDN U19874 ( .B(n15778), .A(n9155), .Z(n15776) );
  XNOR U19875 ( .A(b[202]), .B(n15777), .Z(n15778) );
  XOR U19876 ( .A(n15779), .B(n15780), .Z(n15777) );
  ANDN U19877 ( .B(n15781), .A(n9196), .Z(n15779) );
  XNOR U19878 ( .A(b[201]), .B(n15780), .Z(n15781) );
  XOR U19879 ( .A(n15782), .B(n15783), .Z(n15780) );
  ANDN U19880 ( .B(n15784), .A(n9237), .Z(n15782) );
  XNOR U19881 ( .A(b[200]), .B(n15783), .Z(n15784) );
  XOR U19882 ( .A(n15785), .B(n15786), .Z(n15783) );
  ANDN U19883 ( .B(n15787), .A(n9280), .Z(n15785) );
  XNOR U19884 ( .A(b[199]), .B(n15786), .Z(n15787) );
  XOR U19885 ( .A(n15788), .B(n15789), .Z(n15786) );
  ANDN U19886 ( .B(n15790), .A(n9321), .Z(n15788) );
  XNOR U19887 ( .A(b[198]), .B(n15789), .Z(n15790) );
  XOR U19888 ( .A(n15791), .B(n15792), .Z(n15789) );
  ANDN U19889 ( .B(n15793), .A(n9362), .Z(n15791) );
  XNOR U19890 ( .A(b[197]), .B(n15792), .Z(n15793) );
  XOR U19891 ( .A(n15794), .B(n15795), .Z(n15792) );
  ANDN U19892 ( .B(n15796), .A(n9403), .Z(n15794) );
  XNOR U19893 ( .A(b[196]), .B(n15795), .Z(n15796) );
  XOR U19894 ( .A(n15797), .B(n15798), .Z(n15795) );
  ANDN U19895 ( .B(n15799), .A(n9444), .Z(n15797) );
  XNOR U19896 ( .A(b[195]), .B(n15798), .Z(n15799) );
  XOR U19897 ( .A(n15800), .B(n15801), .Z(n15798) );
  ANDN U19898 ( .B(n15802), .A(n9485), .Z(n15800) );
  XNOR U19899 ( .A(b[194]), .B(n15801), .Z(n15802) );
  XOR U19900 ( .A(n15803), .B(n15804), .Z(n15801) );
  ANDN U19901 ( .B(n15805), .A(n9526), .Z(n15803) );
  XNOR U19902 ( .A(b[193]), .B(n15804), .Z(n15805) );
  XOR U19903 ( .A(n15806), .B(n15807), .Z(n15804) );
  ANDN U19904 ( .B(n15808), .A(n9567), .Z(n15806) );
  XNOR U19905 ( .A(b[192]), .B(n15807), .Z(n15808) );
  XOR U19906 ( .A(n15809), .B(n15810), .Z(n15807) );
  ANDN U19907 ( .B(n15811), .A(n9608), .Z(n15809) );
  XNOR U19908 ( .A(b[191]), .B(n15810), .Z(n15811) );
  XOR U19909 ( .A(n15812), .B(n15813), .Z(n15810) );
  ANDN U19910 ( .B(n15814), .A(n9649), .Z(n15812) );
  XNOR U19911 ( .A(b[190]), .B(n15813), .Z(n15814) );
  XOR U19912 ( .A(n15815), .B(n15816), .Z(n15813) );
  ANDN U19913 ( .B(n15817), .A(n9691), .Z(n15815) );
  XNOR U19914 ( .A(b[189]), .B(n15816), .Z(n15817) );
  XOR U19915 ( .A(n15818), .B(n15819), .Z(n15816) );
  ANDN U19916 ( .B(n15820), .A(n9732), .Z(n15818) );
  XNOR U19917 ( .A(b[188]), .B(n15819), .Z(n15820) );
  XOR U19918 ( .A(n15821), .B(n15822), .Z(n15819) );
  ANDN U19919 ( .B(n15823), .A(n9773), .Z(n15821) );
  XNOR U19920 ( .A(b[187]), .B(n15822), .Z(n15823) );
  XOR U19921 ( .A(n15824), .B(n15825), .Z(n15822) );
  ANDN U19922 ( .B(n15826), .A(n9814), .Z(n15824) );
  XNOR U19923 ( .A(b[186]), .B(n15825), .Z(n15826) );
  XOR U19924 ( .A(n15827), .B(n15828), .Z(n15825) );
  ANDN U19925 ( .B(n15829), .A(n9855), .Z(n15827) );
  XNOR U19926 ( .A(b[185]), .B(n15828), .Z(n15829) );
  XOR U19927 ( .A(n15830), .B(n15831), .Z(n15828) );
  ANDN U19928 ( .B(n15832), .A(n9896), .Z(n15830) );
  XNOR U19929 ( .A(b[184]), .B(n15831), .Z(n15832) );
  XOR U19930 ( .A(n15833), .B(n15834), .Z(n15831) );
  ANDN U19931 ( .B(n15835), .A(n9937), .Z(n15833) );
  XNOR U19932 ( .A(b[183]), .B(n15834), .Z(n15835) );
  XOR U19933 ( .A(n15836), .B(n15837), .Z(n15834) );
  ANDN U19934 ( .B(n15838), .A(n9978), .Z(n15836) );
  XNOR U19935 ( .A(b[182]), .B(n15837), .Z(n15838) );
  XOR U19936 ( .A(n15839), .B(n15840), .Z(n15837) );
  ANDN U19937 ( .B(n15841), .A(n10019), .Z(n15839) );
  XNOR U19938 ( .A(b[181]), .B(n15840), .Z(n15841) );
  XOR U19939 ( .A(n15842), .B(n15843), .Z(n15840) );
  ANDN U19940 ( .B(n15844), .A(n10060), .Z(n15842) );
  XNOR U19941 ( .A(b[180]), .B(n15843), .Z(n15844) );
  XOR U19942 ( .A(n15845), .B(n15846), .Z(n15843) );
  ANDN U19943 ( .B(n15847), .A(n10102), .Z(n15845) );
  XNOR U19944 ( .A(b[179]), .B(n15846), .Z(n15847) );
  XOR U19945 ( .A(n15848), .B(n15849), .Z(n15846) );
  ANDN U19946 ( .B(n15850), .A(n10143), .Z(n15848) );
  XNOR U19947 ( .A(b[178]), .B(n15849), .Z(n15850) );
  XOR U19948 ( .A(n15851), .B(n15852), .Z(n15849) );
  ANDN U19949 ( .B(n15853), .A(n10184), .Z(n15851) );
  XNOR U19950 ( .A(b[177]), .B(n15852), .Z(n15853) );
  XOR U19951 ( .A(n15854), .B(n15855), .Z(n15852) );
  ANDN U19952 ( .B(n15856), .A(n10225), .Z(n15854) );
  XNOR U19953 ( .A(b[176]), .B(n15855), .Z(n15856) );
  XOR U19954 ( .A(n15857), .B(n15858), .Z(n15855) );
  ANDN U19955 ( .B(n15859), .A(n10266), .Z(n15857) );
  XNOR U19956 ( .A(b[175]), .B(n15858), .Z(n15859) );
  XOR U19957 ( .A(n15860), .B(n15861), .Z(n15858) );
  ANDN U19958 ( .B(n15862), .A(n10307), .Z(n15860) );
  XNOR U19959 ( .A(b[174]), .B(n15861), .Z(n15862) );
  XOR U19960 ( .A(n15863), .B(n15864), .Z(n15861) );
  ANDN U19961 ( .B(n15865), .A(n10348), .Z(n15863) );
  XNOR U19962 ( .A(b[173]), .B(n15864), .Z(n15865) );
  XOR U19963 ( .A(n15866), .B(n15867), .Z(n15864) );
  ANDN U19964 ( .B(n15868), .A(n10389), .Z(n15866) );
  XNOR U19965 ( .A(b[172]), .B(n15867), .Z(n15868) );
  XOR U19966 ( .A(n15869), .B(n15870), .Z(n15867) );
  ANDN U19967 ( .B(n15871), .A(n10430), .Z(n15869) );
  XNOR U19968 ( .A(b[171]), .B(n15870), .Z(n15871) );
  XOR U19969 ( .A(n15872), .B(n15873), .Z(n15870) );
  ANDN U19970 ( .B(n15874), .A(n10471), .Z(n15872) );
  XNOR U19971 ( .A(b[170]), .B(n15873), .Z(n15874) );
  XOR U19972 ( .A(n15875), .B(n15876), .Z(n15873) );
  ANDN U19973 ( .B(n15877), .A(n10513), .Z(n15875) );
  XNOR U19974 ( .A(b[169]), .B(n15876), .Z(n15877) );
  XOR U19975 ( .A(n15878), .B(n15879), .Z(n15876) );
  ANDN U19976 ( .B(n15880), .A(n10554), .Z(n15878) );
  XNOR U19977 ( .A(b[168]), .B(n15879), .Z(n15880) );
  XOR U19978 ( .A(n15881), .B(n15882), .Z(n15879) );
  ANDN U19979 ( .B(n15883), .A(n10595), .Z(n15881) );
  XNOR U19980 ( .A(b[167]), .B(n15882), .Z(n15883) );
  XOR U19981 ( .A(n15884), .B(n15885), .Z(n15882) );
  ANDN U19982 ( .B(n15886), .A(n10636), .Z(n15884) );
  XNOR U19983 ( .A(b[166]), .B(n15885), .Z(n15886) );
  XOR U19984 ( .A(n15887), .B(n15888), .Z(n15885) );
  ANDN U19985 ( .B(n15889), .A(n10677), .Z(n15887) );
  XNOR U19986 ( .A(b[165]), .B(n15888), .Z(n15889) );
  XOR U19987 ( .A(n15890), .B(n15891), .Z(n15888) );
  ANDN U19988 ( .B(n15892), .A(n10718), .Z(n15890) );
  XNOR U19989 ( .A(b[164]), .B(n15891), .Z(n15892) );
  XOR U19990 ( .A(n15893), .B(n15894), .Z(n15891) );
  ANDN U19991 ( .B(n15895), .A(n10759), .Z(n15893) );
  XNOR U19992 ( .A(b[163]), .B(n15894), .Z(n15895) );
  XOR U19993 ( .A(n15896), .B(n15897), .Z(n15894) );
  ANDN U19994 ( .B(n15898), .A(n10800), .Z(n15896) );
  XNOR U19995 ( .A(b[162]), .B(n15897), .Z(n15898) );
  XOR U19996 ( .A(n15899), .B(n15900), .Z(n15897) );
  ANDN U19997 ( .B(n15901), .A(n10841), .Z(n15899) );
  XNOR U19998 ( .A(b[161]), .B(n15900), .Z(n15901) );
  XOR U19999 ( .A(n15902), .B(n15903), .Z(n15900) );
  ANDN U20000 ( .B(n15904), .A(n10882), .Z(n15902) );
  XNOR U20001 ( .A(b[160]), .B(n15903), .Z(n15904) );
  XOR U20002 ( .A(n15905), .B(n15906), .Z(n15903) );
  ANDN U20003 ( .B(n15907), .A(n10924), .Z(n15905) );
  XNOR U20004 ( .A(b[159]), .B(n15906), .Z(n15907) );
  XOR U20005 ( .A(n15908), .B(n15909), .Z(n15906) );
  ANDN U20006 ( .B(n15910), .A(n10965), .Z(n15908) );
  XNOR U20007 ( .A(b[158]), .B(n15909), .Z(n15910) );
  XOR U20008 ( .A(n15911), .B(n15912), .Z(n15909) );
  ANDN U20009 ( .B(n15913), .A(n11006), .Z(n15911) );
  XNOR U20010 ( .A(b[157]), .B(n15912), .Z(n15913) );
  XOR U20011 ( .A(n15914), .B(n15915), .Z(n15912) );
  ANDN U20012 ( .B(n15916), .A(n11047), .Z(n15914) );
  XNOR U20013 ( .A(b[156]), .B(n15915), .Z(n15916) );
  XOR U20014 ( .A(n15917), .B(n15918), .Z(n15915) );
  ANDN U20015 ( .B(n15919), .A(n11088), .Z(n15917) );
  XNOR U20016 ( .A(b[155]), .B(n15918), .Z(n15919) );
  XOR U20017 ( .A(n15920), .B(n15921), .Z(n15918) );
  ANDN U20018 ( .B(n15922), .A(n11129), .Z(n15920) );
  XNOR U20019 ( .A(b[154]), .B(n15921), .Z(n15922) );
  XOR U20020 ( .A(n15923), .B(n15924), .Z(n15921) );
  ANDN U20021 ( .B(n15925), .A(n11170), .Z(n15923) );
  XNOR U20022 ( .A(b[153]), .B(n15924), .Z(n15925) );
  XOR U20023 ( .A(n15926), .B(n15927), .Z(n15924) );
  ANDN U20024 ( .B(n15928), .A(n11211), .Z(n15926) );
  XNOR U20025 ( .A(b[152]), .B(n15927), .Z(n15928) );
  XOR U20026 ( .A(n15929), .B(n15930), .Z(n15927) );
  ANDN U20027 ( .B(n15931), .A(n11252), .Z(n15929) );
  XNOR U20028 ( .A(b[151]), .B(n15930), .Z(n15931) );
  XOR U20029 ( .A(n15932), .B(n15933), .Z(n15930) );
  ANDN U20030 ( .B(n15934), .A(n11293), .Z(n15932) );
  XNOR U20031 ( .A(b[150]), .B(n15933), .Z(n15934) );
  XOR U20032 ( .A(n15935), .B(n15936), .Z(n15933) );
  ANDN U20033 ( .B(n15937), .A(n11335), .Z(n15935) );
  XNOR U20034 ( .A(b[149]), .B(n15936), .Z(n15937) );
  XOR U20035 ( .A(n15938), .B(n15939), .Z(n15936) );
  ANDN U20036 ( .B(n15940), .A(n11376), .Z(n15938) );
  XNOR U20037 ( .A(b[148]), .B(n15939), .Z(n15940) );
  XOR U20038 ( .A(n15941), .B(n15942), .Z(n15939) );
  ANDN U20039 ( .B(n15943), .A(n11417), .Z(n15941) );
  XNOR U20040 ( .A(b[147]), .B(n15942), .Z(n15943) );
  XOR U20041 ( .A(n15944), .B(n15945), .Z(n15942) );
  ANDN U20042 ( .B(n15946), .A(n11458), .Z(n15944) );
  XNOR U20043 ( .A(b[146]), .B(n15945), .Z(n15946) );
  XOR U20044 ( .A(n15947), .B(n15948), .Z(n15945) );
  ANDN U20045 ( .B(n15949), .A(n11499), .Z(n15947) );
  XNOR U20046 ( .A(b[145]), .B(n15948), .Z(n15949) );
  XOR U20047 ( .A(n15950), .B(n15951), .Z(n15948) );
  ANDN U20048 ( .B(n15952), .A(n11540), .Z(n15950) );
  XNOR U20049 ( .A(b[144]), .B(n15951), .Z(n15952) );
  XOR U20050 ( .A(n15953), .B(n15954), .Z(n15951) );
  ANDN U20051 ( .B(n15955), .A(n11581), .Z(n15953) );
  XNOR U20052 ( .A(b[143]), .B(n15954), .Z(n15955) );
  XOR U20053 ( .A(n15956), .B(n15957), .Z(n15954) );
  ANDN U20054 ( .B(n15958), .A(n11622), .Z(n15956) );
  XNOR U20055 ( .A(b[142]), .B(n15957), .Z(n15958) );
  XOR U20056 ( .A(n15959), .B(n15960), .Z(n15957) );
  ANDN U20057 ( .B(n15961), .A(n11663), .Z(n15959) );
  XNOR U20058 ( .A(b[141]), .B(n15960), .Z(n15961) );
  XOR U20059 ( .A(n15962), .B(n15963), .Z(n15960) );
  ANDN U20060 ( .B(n15964), .A(n11704), .Z(n15962) );
  XNOR U20061 ( .A(b[140]), .B(n15963), .Z(n15964) );
  XOR U20062 ( .A(n15965), .B(n15966), .Z(n15963) );
  ANDN U20063 ( .B(n15967), .A(n11746), .Z(n15965) );
  XNOR U20064 ( .A(b[139]), .B(n15966), .Z(n15967) );
  XOR U20065 ( .A(n15968), .B(n15969), .Z(n15966) );
  ANDN U20066 ( .B(n15970), .A(n11787), .Z(n15968) );
  XNOR U20067 ( .A(b[138]), .B(n15969), .Z(n15970) );
  XOR U20068 ( .A(n15971), .B(n15972), .Z(n15969) );
  ANDN U20069 ( .B(n15973), .A(n11828), .Z(n15971) );
  XNOR U20070 ( .A(b[137]), .B(n15972), .Z(n15973) );
  XOR U20071 ( .A(n15974), .B(n15975), .Z(n15972) );
  ANDN U20072 ( .B(n15976), .A(n11869), .Z(n15974) );
  XNOR U20073 ( .A(b[136]), .B(n15975), .Z(n15976) );
  XOR U20074 ( .A(n15977), .B(n15978), .Z(n15975) );
  ANDN U20075 ( .B(n15979), .A(n11910), .Z(n15977) );
  XNOR U20076 ( .A(b[135]), .B(n15978), .Z(n15979) );
  XOR U20077 ( .A(n15980), .B(n15981), .Z(n15978) );
  ANDN U20078 ( .B(n15982), .A(n11951), .Z(n15980) );
  XNOR U20079 ( .A(b[134]), .B(n15981), .Z(n15982) );
  XOR U20080 ( .A(n15983), .B(n15984), .Z(n15981) );
  ANDN U20081 ( .B(n15985), .A(n11992), .Z(n15983) );
  XNOR U20082 ( .A(b[133]), .B(n15984), .Z(n15985) );
  XOR U20083 ( .A(n15986), .B(n15987), .Z(n15984) );
  ANDN U20084 ( .B(n15988), .A(n12033), .Z(n15986) );
  XNOR U20085 ( .A(b[132]), .B(n15987), .Z(n15988) );
  XOR U20086 ( .A(n15989), .B(n15990), .Z(n15987) );
  ANDN U20087 ( .B(n15991), .A(n12074), .Z(n15989) );
  XNOR U20088 ( .A(b[131]), .B(n15990), .Z(n15991) );
  XOR U20089 ( .A(n15992), .B(n15993), .Z(n15990) );
  ANDN U20090 ( .B(n15994), .A(n12115), .Z(n15992) );
  XNOR U20091 ( .A(b[130]), .B(n15993), .Z(n15994) );
  XOR U20092 ( .A(n15995), .B(n15996), .Z(n15993) );
  ANDN U20093 ( .B(n15997), .A(n12157), .Z(n15995) );
  XNOR U20094 ( .A(b[129]), .B(n15996), .Z(n15997) );
  XOR U20095 ( .A(n15998), .B(n15999), .Z(n15996) );
  ANDN U20096 ( .B(n16000), .A(n12198), .Z(n15998) );
  XNOR U20097 ( .A(b[128]), .B(n15999), .Z(n16000) );
  XOR U20098 ( .A(n16001), .B(n16002), .Z(n15999) );
  ANDN U20099 ( .B(n16003), .A(n12239), .Z(n16001) );
  XNOR U20100 ( .A(b[127]), .B(n16002), .Z(n16003) );
  XOR U20101 ( .A(n16004), .B(n16005), .Z(n16002) );
  ANDN U20102 ( .B(n16006), .A(n12280), .Z(n16004) );
  XNOR U20103 ( .A(b[126]), .B(n16005), .Z(n16006) );
  XOR U20104 ( .A(n16007), .B(n16008), .Z(n16005) );
  ANDN U20105 ( .B(n16009), .A(n12321), .Z(n16007) );
  XNOR U20106 ( .A(b[125]), .B(n16008), .Z(n16009) );
  XOR U20107 ( .A(n16010), .B(n16011), .Z(n16008) );
  ANDN U20108 ( .B(n16012), .A(n12362), .Z(n16010) );
  XNOR U20109 ( .A(b[124]), .B(n16011), .Z(n16012) );
  XOR U20110 ( .A(n16013), .B(n16014), .Z(n16011) );
  ANDN U20111 ( .B(n16015), .A(n12403), .Z(n16013) );
  XNOR U20112 ( .A(b[123]), .B(n16014), .Z(n16015) );
  XOR U20113 ( .A(n16016), .B(n16017), .Z(n16014) );
  ANDN U20114 ( .B(n16018), .A(n12444), .Z(n16016) );
  XNOR U20115 ( .A(b[122]), .B(n16017), .Z(n16018) );
  XOR U20116 ( .A(n16019), .B(n16020), .Z(n16017) );
  ANDN U20117 ( .B(n16021), .A(n12485), .Z(n16019) );
  XNOR U20118 ( .A(b[121]), .B(n16020), .Z(n16021) );
  XOR U20119 ( .A(n16022), .B(n16023), .Z(n16020) );
  ANDN U20120 ( .B(n16024), .A(n12526), .Z(n16022) );
  XNOR U20121 ( .A(b[120]), .B(n16023), .Z(n16024) );
  XOR U20122 ( .A(n16025), .B(n16026), .Z(n16023) );
  ANDN U20123 ( .B(n16027), .A(n12568), .Z(n16025) );
  XNOR U20124 ( .A(b[119]), .B(n16026), .Z(n16027) );
  XOR U20125 ( .A(n16028), .B(n16029), .Z(n16026) );
  ANDN U20126 ( .B(n16030), .A(n12609), .Z(n16028) );
  XNOR U20127 ( .A(b[118]), .B(n16029), .Z(n16030) );
  XOR U20128 ( .A(n16031), .B(n16032), .Z(n16029) );
  ANDN U20129 ( .B(n16033), .A(n12650), .Z(n16031) );
  XNOR U20130 ( .A(b[117]), .B(n16032), .Z(n16033) );
  XOR U20131 ( .A(n16034), .B(n16035), .Z(n16032) );
  ANDN U20132 ( .B(n16036), .A(n12691), .Z(n16034) );
  XNOR U20133 ( .A(b[116]), .B(n16035), .Z(n16036) );
  XOR U20134 ( .A(n16037), .B(n16038), .Z(n16035) );
  ANDN U20135 ( .B(n16039), .A(n12732), .Z(n16037) );
  XNOR U20136 ( .A(b[115]), .B(n16038), .Z(n16039) );
  XOR U20137 ( .A(n16040), .B(n16041), .Z(n16038) );
  ANDN U20138 ( .B(n16042), .A(n12773), .Z(n16040) );
  XNOR U20139 ( .A(b[114]), .B(n16041), .Z(n16042) );
  XOR U20140 ( .A(n16043), .B(n16044), .Z(n16041) );
  ANDN U20141 ( .B(n16045), .A(n12814), .Z(n16043) );
  XNOR U20142 ( .A(b[113]), .B(n16044), .Z(n16045) );
  XOR U20143 ( .A(n16046), .B(n16047), .Z(n16044) );
  ANDN U20144 ( .B(n16048), .A(n12855), .Z(n16046) );
  XNOR U20145 ( .A(b[112]), .B(n16047), .Z(n16048) );
  XOR U20146 ( .A(n16049), .B(n16050), .Z(n16047) );
  ANDN U20147 ( .B(n16051), .A(n12896), .Z(n16049) );
  XNOR U20148 ( .A(b[111]), .B(n16050), .Z(n16051) );
  XOR U20149 ( .A(n16052), .B(n16053), .Z(n16050) );
  ANDN U20150 ( .B(n16054), .A(n12937), .Z(n16052) );
  XNOR U20151 ( .A(b[110]), .B(n16053), .Z(n16054) );
  XOR U20152 ( .A(n16055), .B(n16056), .Z(n16053) );
  ANDN U20153 ( .B(n16057), .A(n12979), .Z(n16055) );
  XNOR U20154 ( .A(b[109]), .B(n16056), .Z(n16057) );
  XOR U20155 ( .A(n16058), .B(n16059), .Z(n16056) );
  ANDN U20156 ( .B(n16060), .A(n13020), .Z(n16058) );
  XNOR U20157 ( .A(b[108]), .B(n16059), .Z(n16060) );
  XOR U20158 ( .A(n16061), .B(n16062), .Z(n16059) );
  ANDN U20159 ( .B(n16063), .A(n13061), .Z(n16061) );
  XNOR U20160 ( .A(b[107]), .B(n16062), .Z(n16063) );
  XOR U20161 ( .A(n16064), .B(n16065), .Z(n16062) );
  ANDN U20162 ( .B(n16066), .A(n13102), .Z(n16064) );
  XNOR U20163 ( .A(b[106]), .B(n16065), .Z(n16066) );
  XOR U20164 ( .A(n16067), .B(n16068), .Z(n16065) );
  ANDN U20165 ( .B(n16069), .A(n13143), .Z(n16067) );
  XNOR U20166 ( .A(b[105]), .B(n16068), .Z(n16069) );
  XOR U20167 ( .A(n16070), .B(n16071), .Z(n16068) );
  ANDN U20168 ( .B(n16072), .A(n13184), .Z(n16070) );
  XNOR U20169 ( .A(b[104]), .B(n16071), .Z(n16072) );
  XOR U20170 ( .A(n16073), .B(n16074), .Z(n16071) );
  ANDN U20171 ( .B(n16075), .A(n13225), .Z(n16073) );
  XNOR U20172 ( .A(b[103]), .B(n16074), .Z(n16075) );
  XOR U20173 ( .A(n16076), .B(n16077), .Z(n16074) );
  ANDN U20174 ( .B(n16078), .A(n13266), .Z(n16076) );
  XNOR U20175 ( .A(b[102]), .B(n16077), .Z(n16078) );
  XOR U20176 ( .A(n16079), .B(n16080), .Z(n16077) );
  ANDN U20177 ( .B(n16081), .A(n13307), .Z(n16079) );
  XNOR U20178 ( .A(b[101]), .B(n16080), .Z(n16081) );
  XOR U20179 ( .A(n16082), .B(n16083), .Z(n16080) );
  ANDN U20180 ( .B(n16084), .A(n13348), .Z(n16082) );
  XNOR U20181 ( .A(b[100]), .B(n16083), .Z(n16084) );
  XOR U20182 ( .A(n16085), .B(n16086), .Z(n16083) );
  ANDN U20183 ( .B(n16087), .A(n7), .Z(n16085) );
  XNOR U20184 ( .A(b[99]), .B(n16086), .Z(n16087) );
  XOR U20185 ( .A(n16088), .B(n16089), .Z(n16086) );
  ANDN U20186 ( .B(n16090), .A(n18), .Z(n16088) );
  XNOR U20187 ( .A(b[98]), .B(n16089), .Z(n16090) );
  XOR U20188 ( .A(n16091), .B(n16092), .Z(n16089) );
  ANDN U20189 ( .B(n16093), .A(n29), .Z(n16091) );
  XNOR U20190 ( .A(b[97]), .B(n16092), .Z(n16093) );
  XOR U20191 ( .A(n16094), .B(n16095), .Z(n16092) );
  ANDN U20192 ( .B(n16096), .A(n40), .Z(n16094) );
  XNOR U20193 ( .A(b[96]), .B(n16095), .Z(n16096) );
  XOR U20194 ( .A(n16097), .B(n16098), .Z(n16095) );
  ANDN U20195 ( .B(n16099), .A(n51), .Z(n16097) );
  XNOR U20196 ( .A(b[95]), .B(n16098), .Z(n16099) );
  XOR U20197 ( .A(n16100), .B(n16101), .Z(n16098) );
  ANDN U20198 ( .B(n16102), .A(n62), .Z(n16100) );
  XNOR U20199 ( .A(b[94]), .B(n16101), .Z(n16102) );
  XOR U20200 ( .A(n16103), .B(n16104), .Z(n16101) );
  ANDN U20201 ( .B(n16105), .A(n73), .Z(n16103) );
  XNOR U20202 ( .A(b[93]), .B(n16104), .Z(n16105) );
  XOR U20203 ( .A(n16106), .B(n16107), .Z(n16104) );
  ANDN U20204 ( .B(n16108), .A(n84), .Z(n16106) );
  XNOR U20205 ( .A(b[92]), .B(n16107), .Z(n16108) );
  XOR U20206 ( .A(n16109), .B(n16110), .Z(n16107) );
  ANDN U20207 ( .B(n16111), .A(n95), .Z(n16109) );
  XNOR U20208 ( .A(b[91]), .B(n16110), .Z(n16111) );
  XOR U20209 ( .A(n16112), .B(n16113), .Z(n16110) );
  ANDN U20210 ( .B(n16114), .A(n106), .Z(n16112) );
  XNOR U20211 ( .A(b[90]), .B(n16113), .Z(n16114) );
  XOR U20212 ( .A(n16115), .B(n16116), .Z(n16113) );
  ANDN U20213 ( .B(n16117), .A(n118), .Z(n16115) );
  XNOR U20214 ( .A(b[89]), .B(n16116), .Z(n16117) );
  XOR U20215 ( .A(n16118), .B(n16119), .Z(n16116) );
  ANDN U20216 ( .B(n16120), .A(n129), .Z(n16118) );
  XNOR U20217 ( .A(b[88]), .B(n16119), .Z(n16120) );
  XOR U20218 ( .A(n16121), .B(n16122), .Z(n16119) );
  ANDN U20219 ( .B(n16123), .A(n140), .Z(n16121) );
  XNOR U20220 ( .A(b[87]), .B(n16122), .Z(n16123) );
  XOR U20221 ( .A(n16124), .B(n16125), .Z(n16122) );
  ANDN U20222 ( .B(n16126), .A(n151), .Z(n16124) );
  XNOR U20223 ( .A(b[86]), .B(n16125), .Z(n16126) );
  XOR U20224 ( .A(n16127), .B(n16128), .Z(n16125) );
  ANDN U20225 ( .B(n16129), .A(n162), .Z(n16127) );
  XNOR U20226 ( .A(b[85]), .B(n16128), .Z(n16129) );
  XOR U20227 ( .A(n16130), .B(n16131), .Z(n16128) );
  ANDN U20228 ( .B(n16132), .A(n173), .Z(n16130) );
  XNOR U20229 ( .A(b[84]), .B(n16131), .Z(n16132) );
  XOR U20230 ( .A(n16133), .B(n16134), .Z(n16131) );
  ANDN U20231 ( .B(n16135), .A(n184), .Z(n16133) );
  XNOR U20232 ( .A(b[83]), .B(n16134), .Z(n16135) );
  XOR U20233 ( .A(n16136), .B(n16137), .Z(n16134) );
  ANDN U20234 ( .B(n16138), .A(n195), .Z(n16136) );
  XNOR U20235 ( .A(b[82]), .B(n16137), .Z(n16138) );
  XOR U20236 ( .A(n16139), .B(n16140), .Z(n16137) );
  ANDN U20237 ( .B(n16141), .A(n206), .Z(n16139) );
  XNOR U20238 ( .A(b[81]), .B(n16140), .Z(n16141) );
  XOR U20239 ( .A(n16142), .B(n16143), .Z(n16140) );
  ANDN U20240 ( .B(n16144), .A(n217), .Z(n16142) );
  XNOR U20241 ( .A(b[80]), .B(n16143), .Z(n16144) );
  XOR U20242 ( .A(n16145), .B(n16146), .Z(n16143) );
  ANDN U20243 ( .B(n16147), .A(n229), .Z(n16145) );
  XNOR U20244 ( .A(b[79]), .B(n16146), .Z(n16147) );
  XOR U20245 ( .A(n16148), .B(n16149), .Z(n16146) );
  ANDN U20246 ( .B(n16150), .A(n240), .Z(n16148) );
  XNOR U20247 ( .A(b[78]), .B(n16149), .Z(n16150) );
  XOR U20248 ( .A(n16151), .B(n16152), .Z(n16149) );
  ANDN U20249 ( .B(n16153), .A(n251), .Z(n16151) );
  XNOR U20250 ( .A(b[77]), .B(n16152), .Z(n16153) );
  XOR U20251 ( .A(n16154), .B(n16155), .Z(n16152) );
  ANDN U20252 ( .B(n16156), .A(n262), .Z(n16154) );
  XNOR U20253 ( .A(b[76]), .B(n16155), .Z(n16156) );
  XOR U20254 ( .A(n16157), .B(n16158), .Z(n16155) );
  ANDN U20255 ( .B(n16159), .A(n273), .Z(n16157) );
  XNOR U20256 ( .A(b[75]), .B(n16158), .Z(n16159) );
  XOR U20257 ( .A(n16160), .B(n16161), .Z(n16158) );
  ANDN U20258 ( .B(n16162), .A(n284), .Z(n16160) );
  XNOR U20259 ( .A(b[74]), .B(n16161), .Z(n16162) );
  XOR U20260 ( .A(n16163), .B(n16164), .Z(n16161) );
  ANDN U20261 ( .B(n16165), .A(n295), .Z(n16163) );
  XNOR U20262 ( .A(b[73]), .B(n16164), .Z(n16165) );
  XOR U20263 ( .A(n16166), .B(n16167), .Z(n16164) );
  ANDN U20264 ( .B(n16168), .A(n306), .Z(n16166) );
  XNOR U20265 ( .A(b[72]), .B(n16167), .Z(n16168) );
  XOR U20266 ( .A(n16169), .B(n16170), .Z(n16167) );
  ANDN U20267 ( .B(n16171), .A(n317), .Z(n16169) );
  XNOR U20268 ( .A(b[71]), .B(n16170), .Z(n16171) );
  XOR U20269 ( .A(n16172), .B(n16173), .Z(n16170) );
  ANDN U20270 ( .B(n16174), .A(n328), .Z(n16172) );
  XNOR U20271 ( .A(b[70]), .B(n16173), .Z(n16174) );
  XOR U20272 ( .A(n16175), .B(n16176), .Z(n16173) );
  ANDN U20273 ( .B(n16177), .A(n340), .Z(n16175) );
  XNOR U20274 ( .A(b[69]), .B(n16176), .Z(n16177) );
  XOR U20275 ( .A(n16178), .B(n16179), .Z(n16176) );
  ANDN U20276 ( .B(n16180), .A(n351), .Z(n16178) );
  XNOR U20277 ( .A(b[68]), .B(n16179), .Z(n16180) );
  XOR U20278 ( .A(n16181), .B(n16182), .Z(n16179) );
  ANDN U20279 ( .B(n16183), .A(n362), .Z(n16181) );
  XNOR U20280 ( .A(b[67]), .B(n16182), .Z(n16183) );
  XOR U20281 ( .A(n16184), .B(n16185), .Z(n16182) );
  ANDN U20282 ( .B(n16186), .A(n373), .Z(n16184) );
  XNOR U20283 ( .A(b[66]), .B(n16185), .Z(n16186) );
  XOR U20284 ( .A(n16187), .B(n16188), .Z(n16185) );
  ANDN U20285 ( .B(n16189), .A(n384), .Z(n16187) );
  XNOR U20286 ( .A(b[65]), .B(n16188), .Z(n16189) );
  XOR U20287 ( .A(n16190), .B(n16191), .Z(n16188) );
  ANDN U20288 ( .B(n16192), .A(n395), .Z(n16190) );
  XNOR U20289 ( .A(b[64]), .B(n16191), .Z(n16192) );
  XOR U20290 ( .A(n16193), .B(n16194), .Z(n16191) );
  ANDN U20291 ( .B(n16195), .A(n406), .Z(n16193) );
  XNOR U20292 ( .A(b[63]), .B(n16194), .Z(n16195) );
  XOR U20293 ( .A(n16196), .B(n16197), .Z(n16194) );
  ANDN U20294 ( .B(n16198), .A(n417), .Z(n16196) );
  XNOR U20295 ( .A(b[62]), .B(n16197), .Z(n16198) );
  XOR U20296 ( .A(n16199), .B(n16200), .Z(n16197) );
  ANDN U20297 ( .B(n16201), .A(n428), .Z(n16199) );
  XNOR U20298 ( .A(b[61]), .B(n16200), .Z(n16201) );
  XOR U20299 ( .A(n16202), .B(n16203), .Z(n16200) );
  ANDN U20300 ( .B(n16204), .A(n439), .Z(n16202) );
  XNOR U20301 ( .A(b[60]), .B(n16203), .Z(n16204) );
  XOR U20302 ( .A(n16205), .B(n16206), .Z(n16203) );
  ANDN U20303 ( .B(n16207), .A(n451), .Z(n16205) );
  XNOR U20304 ( .A(b[59]), .B(n16206), .Z(n16207) );
  XOR U20305 ( .A(n16208), .B(n16209), .Z(n16206) );
  ANDN U20306 ( .B(n16210), .A(n462), .Z(n16208) );
  XNOR U20307 ( .A(b[58]), .B(n16209), .Z(n16210) );
  XOR U20308 ( .A(n16211), .B(n16212), .Z(n16209) );
  ANDN U20309 ( .B(n16213), .A(n473), .Z(n16211) );
  XNOR U20310 ( .A(b[57]), .B(n16212), .Z(n16213) );
  XOR U20311 ( .A(n16214), .B(n16215), .Z(n16212) );
  ANDN U20312 ( .B(n16216), .A(n484), .Z(n16214) );
  XNOR U20313 ( .A(b[56]), .B(n16215), .Z(n16216) );
  XOR U20314 ( .A(n16217), .B(n16218), .Z(n16215) );
  ANDN U20315 ( .B(n16219), .A(n495), .Z(n16217) );
  XNOR U20316 ( .A(b[55]), .B(n16218), .Z(n16219) );
  XOR U20317 ( .A(n16220), .B(n16221), .Z(n16218) );
  ANDN U20318 ( .B(n16222), .A(n506), .Z(n16220) );
  XNOR U20319 ( .A(b[54]), .B(n16221), .Z(n16222) );
  XOR U20320 ( .A(n16223), .B(n16224), .Z(n16221) );
  ANDN U20321 ( .B(n16225), .A(n517), .Z(n16223) );
  XNOR U20322 ( .A(b[53]), .B(n16224), .Z(n16225) );
  XOR U20323 ( .A(n16226), .B(n16227), .Z(n16224) );
  ANDN U20324 ( .B(n16228), .A(n528), .Z(n16226) );
  XNOR U20325 ( .A(b[52]), .B(n16227), .Z(n16228) );
  XOR U20326 ( .A(n16229), .B(n16230), .Z(n16227) );
  ANDN U20327 ( .B(n16231), .A(n539), .Z(n16229) );
  XNOR U20328 ( .A(b[51]), .B(n16230), .Z(n16231) );
  XOR U20329 ( .A(n16232), .B(n16233), .Z(n16230) );
  ANDN U20330 ( .B(n16234), .A(n550), .Z(n16232) );
  XNOR U20331 ( .A(b[50]), .B(n16233), .Z(n16234) );
  XOR U20332 ( .A(n16235), .B(n16236), .Z(n16233) );
  ANDN U20333 ( .B(n16237), .A(n562), .Z(n16235) );
  XNOR U20334 ( .A(b[49]), .B(n16236), .Z(n16237) );
  XOR U20335 ( .A(n16238), .B(n16239), .Z(n16236) );
  ANDN U20336 ( .B(n16240), .A(n573), .Z(n16238) );
  XNOR U20337 ( .A(b[48]), .B(n16239), .Z(n16240) );
  XOR U20338 ( .A(n16241), .B(n16242), .Z(n16239) );
  ANDN U20339 ( .B(n16243), .A(n584), .Z(n16241) );
  XNOR U20340 ( .A(b[47]), .B(n16242), .Z(n16243) );
  XOR U20341 ( .A(n16244), .B(n16245), .Z(n16242) );
  ANDN U20342 ( .B(n16246), .A(n595), .Z(n16244) );
  XNOR U20343 ( .A(b[46]), .B(n16245), .Z(n16246) );
  XOR U20344 ( .A(n16247), .B(n16248), .Z(n16245) );
  ANDN U20345 ( .B(n16249), .A(n606), .Z(n16247) );
  XNOR U20346 ( .A(b[45]), .B(n16248), .Z(n16249) );
  XOR U20347 ( .A(n16250), .B(n16251), .Z(n16248) );
  ANDN U20348 ( .B(n16252), .A(n617), .Z(n16250) );
  XNOR U20349 ( .A(b[44]), .B(n16251), .Z(n16252) );
  XOR U20350 ( .A(n16253), .B(n16254), .Z(n16251) );
  ANDN U20351 ( .B(n16255), .A(n628), .Z(n16253) );
  XNOR U20352 ( .A(b[43]), .B(n16254), .Z(n16255) );
  XOR U20353 ( .A(n16256), .B(n16257), .Z(n16254) );
  ANDN U20354 ( .B(n16258), .A(n639), .Z(n16256) );
  XNOR U20355 ( .A(b[42]), .B(n16257), .Z(n16258) );
  XOR U20356 ( .A(n16259), .B(n16260), .Z(n16257) );
  ANDN U20357 ( .B(n16261), .A(n650), .Z(n16259) );
  XNOR U20358 ( .A(b[41]), .B(n16260), .Z(n16261) );
  XOR U20359 ( .A(n16262), .B(n16263), .Z(n16260) );
  ANDN U20360 ( .B(n16264), .A(n661), .Z(n16262) );
  XNOR U20361 ( .A(b[40]), .B(n16263), .Z(n16264) );
  XOR U20362 ( .A(n16265), .B(n16266), .Z(n16263) );
  ANDN U20363 ( .B(n16267), .A(n1057), .Z(n16265) );
  XNOR U20364 ( .A(b[39]), .B(n16266), .Z(n16267) );
  XOR U20365 ( .A(n16268), .B(n16269), .Z(n16266) );
  ANDN U20366 ( .B(n16270), .A(n1468), .Z(n16268) );
  XNOR U20367 ( .A(b[38]), .B(n16269), .Z(n16270) );
  XOR U20368 ( .A(n16271), .B(n16272), .Z(n16269) );
  ANDN U20369 ( .B(n16273), .A(n1879), .Z(n16271) );
  XNOR U20370 ( .A(b[37]), .B(n16272), .Z(n16273) );
  XOR U20371 ( .A(n16274), .B(n16275), .Z(n16272) );
  ANDN U20372 ( .B(n16276), .A(n2290), .Z(n16274) );
  XNOR U20373 ( .A(b[36]), .B(n16275), .Z(n16276) );
  XOR U20374 ( .A(n16277), .B(n16278), .Z(n16275) );
  ANDN U20375 ( .B(n16279), .A(n2701), .Z(n16277) );
  XNOR U20376 ( .A(b[35]), .B(n16278), .Z(n16279) );
  XOR U20377 ( .A(n16280), .B(n16281), .Z(n16278) );
  ANDN U20378 ( .B(n16282), .A(n3112), .Z(n16280) );
  XNOR U20379 ( .A(b[34]), .B(n16281), .Z(n16282) );
  XOR U20380 ( .A(n16283), .B(n16284), .Z(n16281) );
  ANDN U20381 ( .B(n16285), .A(n3523), .Z(n16283) );
  XNOR U20382 ( .A(b[33]), .B(n16284), .Z(n16285) );
  XOR U20383 ( .A(n16286), .B(n16287), .Z(n16284) );
  ANDN U20384 ( .B(n16288), .A(n3934), .Z(n16286) );
  XNOR U20385 ( .A(b[32]), .B(n16287), .Z(n16288) );
  XOR U20386 ( .A(n16289), .B(n16290), .Z(n16287) );
  ANDN U20387 ( .B(n16291), .A(n4345), .Z(n16289) );
  XNOR U20388 ( .A(b[31]), .B(n16290), .Z(n16291) );
  XOR U20389 ( .A(n16292), .B(n16293), .Z(n16290) );
  ANDN U20390 ( .B(n16294), .A(n4756), .Z(n16292) );
  XNOR U20391 ( .A(b[30]), .B(n16293), .Z(n16294) );
  XOR U20392 ( .A(n16295), .B(n16296), .Z(n16293) );
  ANDN U20393 ( .B(n16297), .A(n5168), .Z(n16295) );
  XNOR U20394 ( .A(b[29]), .B(n16296), .Z(n16297) );
  XOR U20395 ( .A(n16298), .B(n16299), .Z(n16296) );
  ANDN U20396 ( .B(n16300), .A(n5579), .Z(n16298) );
  XNOR U20397 ( .A(b[28]), .B(n16299), .Z(n16300) );
  XOR U20398 ( .A(n16301), .B(n16302), .Z(n16299) );
  ANDN U20399 ( .B(n16303), .A(n5990), .Z(n16301) );
  XNOR U20400 ( .A(b[27]), .B(n16302), .Z(n16303) );
  XOR U20401 ( .A(n16304), .B(n16305), .Z(n16302) );
  ANDN U20402 ( .B(n16306), .A(n6401), .Z(n16304) );
  XNOR U20403 ( .A(b[26]), .B(n16305), .Z(n16306) );
  XOR U20404 ( .A(n16307), .B(n16308), .Z(n16305) );
  ANDN U20405 ( .B(n16309), .A(n6812), .Z(n16307) );
  XNOR U20406 ( .A(b[25]), .B(n16308), .Z(n16309) );
  XOR U20407 ( .A(n16310), .B(n16311), .Z(n16308) );
  ANDN U20408 ( .B(n16312), .A(n7223), .Z(n16310) );
  XNOR U20409 ( .A(b[24]), .B(n16311), .Z(n16312) );
  XOR U20410 ( .A(n16313), .B(n16314), .Z(n16311) );
  ANDN U20411 ( .B(n16315), .A(n7634), .Z(n16313) );
  XNOR U20412 ( .A(b[23]), .B(n16314), .Z(n16315) );
  XOR U20413 ( .A(n16316), .B(n16317), .Z(n16314) );
  ANDN U20414 ( .B(n16318), .A(n8045), .Z(n16316) );
  XNOR U20415 ( .A(b[22]), .B(n16317), .Z(n16318) );
  XOR U20416 ( .A(n16319), .B(n16320), .Z(n16317) );
  ANDN U20417 ( .B(n16321), .A(n8456), .Z(n16319) );
  XNOR U20418 ( .A(b[21]), .B(n16320), .Z(n16321) );
  XOR U20419 ( .A(n16322), .B(n16323), .Z(n16320) );
  ANDN U20420 ( .B(n16324), .A(n8867), .Z(n16322) );
  XNOR U20421 ( .A(b[20]), .B(n16323), .Z(n16324) );
  XOR U20422 ( .A(n16325), .B(n16326), .Z(n16323) );
  ANDN U20423 ( .B(n16327), .A(n9279), .Z(n16325) );
  XNOR U20424 ( .A(b[19]), .B(n16326), .Z(n16327) );
  XOR U20425 ( .A(n16328), .B(n16329), .Z(n16326) );
  ANDN U20426 ( .B(n16330), .A(n9690), .Z(n16328) );
  XNOR U20427 ( .A(b[18]), .B(n16329), .Z(n16330) );
  XOR U20428 ( .A(n16331), .B(n16332), .Z(n16329) );
  ANDN U20429 ( .B(n16333), .A(n10101), .Z(n16331) );
  XNOR U20430 ( .A(b[17]), .B(n16332), .Z(n16333) );
  XOR U20431 ( .A(n16334), .B(n16335), .Z(n16332) );
  ANDN U20432 ( .B(n16336), .A(n10512), .Z(n16334) );
  XNOR U20433 ( .A(b[16]), .B(n16335), .Z(n16336) );
  XOR U20434 ( .A(n16337), .B(n16338), .Z(n16335) );
  ANDN U20435 ( .B(n16339), .A(n10923), .Z(n16337) );
  XNOR U20436 ( .A(b[15]), .B(n16338), .Z(n16339) );
  XOR U20437 ( .A(n16340), .B(n16341), .Z(n16338) );
  ANDN U20438 ( .B(n16342), .A(n11334), .Z(n16340) );
  XNOR U20439 ( .A(b[14]), .B(n16341), .Z(n16342) );
  XOR U20440 ( .A(n16343), .B(n16344), .Z(n16341) );
  ANDN U20441 ( .B(n16345), .A(n11745), .Z(n16343) );
  XNOR U20442 ( .A(b[13]), .B(n16344), .Z(n16345) );
  XOR U20443 ( .A(n16346), .B(n16347), .Z(n16344) );
  ANDN U20444 ( .B(n16348), .A(n12156), .Z(n16346) );
  XNOR U20445 ( .A(b[12]), .B(n16347), .Z(n16348) );
  XOR U20446 ( .A(n16349), .B(n16350), .Z(n16347) );
  ANDN U20447 ( .B(n16351), .A(n12567), .Z(n16349) );
  XNOR U20448 ( .A(b[11]), .B(n16350), .Z(n16351) );
  XOR U20449 ( .A(n16352), .B(n16353), .Z(n16350) );
  ANDN U20450 ( .B(n16354), .A(n12978), .Z(n16352) );
  XNOR U20451 ( .A(b[10]), .B(n16353), .Z(n16354) );
  XOR U20452 ( .A(n16355), .B(n16356), .Z(n16353) );
  ANDN U20453 ( .B(n16357), .A(n6), .Z(n16355) );
  XNOR U20454 ( .A(b[9]), .B(n16356), .Z(n16357) );
  XOR U20455 ( .A(n16358), .B(n16359), .Z(n16356) );
  ANDN U20456 ( .B(n16360), .A(n117), .Z(n16358) );
  XNOR U20457 ( .A(b[8]), .B(n16359), .Z(n16360) );
  XOR U20458 ( .A(n16361), .B(n16362), .Z(n16359) );
  ANDN U20459 ( .B(n16363), .A(n228), .Z(n16361) );
  XNOR U20460 ( .A(b[7]), .B(n16362), .Z(n16363) );
  XOR U20461 ( .A(n16364), .B(n16365), .Z(n16362) );
  ANDN U20462 ( .B(n16366), .A(n339), .Z(n16364) );
  XNOR U20463 ( .A(b[6]), .B(n16365), .Z(n16366) );
  XOR U20464 ( .A(n16367), .B(n16368), .Z(n16365) );
  ANDN U20465 ( .B(n16369), .A(n450), .Z(n16367) );
  XNOR U20466 ( .A(b[5]), .B(n16368), .Z(n16369) );
  XOR U20467 ( .A(n16370), .B(n16371), .Z(n16368) );
  ANDN U20468 ( .B(n16372), .A(n561), .Z(n16370) );
  XNOR U20469 ( .A(b[4]), .B(n16371), .Z(n16372) );
  XOR U20470 ( .A(n16373), .B(n16374), .Z(n16371) );
  ANDN U20471 ( .B(n16375), .A(n1056), .Z(n16373) );
  XNOR U20472 ( .A(b[3]), .B(n16374), .Z(n16375) );
  XOR U20473 ( .A(n16376), .B(n16377), .Z(n16374) );
  ANDN U20474 ( .B(n16378), .A(n5167), .Z(n16376) );
  XNOR U20475 ( .A(b[2]), .B(n16377), .Z(n16378) );
  XOR U20476 ( .A(n16379), .B(n16380), .Z(n16377) );
  ANDN U20477 ( .B(n16381), .A(n9278), .Z(n16379) );
  XNOR U20478 ( .A(b[1]), .B(n16380), .Z(n16381) );
  XOR U20479 ( .A(carry_on), .B(n16382), .Z(n16380) );
  NANDN U20480 ( .A(n16383), .B(n16384), .Z(n16382) );
  XOR U20481 ( .A(carry_on), .B(b[0]), .Z(n16384) );
  XNOR U20482 ( .A(b[0]), .B(n16383), .Z(c[0]) );
  XNOR U20483 ( .A(a[0]), .B(carry_on), .Z(n16383) );
endmodule

